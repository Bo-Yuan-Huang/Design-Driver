
module oc8051_gm_top(clk, rst, word_in, xram_data_in, RD_IRAM_0_ABSTR_ADDR, RD_IRAM_1_ABSTR_ADDR, RD_ROM_1_ABSTR_ADDR, RD_ROM_2_ABSTR_ADDR, ACC_abstr, P2_abstr, P0_abstr, P1_abstr, P3_abstr, SP_abstr, PC_abstr, B_abstr, DPL_abstr, PSW_abstr, DPH_abstr, XRAM_DATA_OUT_abstr, XRAM_ADDR_abstr, WR_COND_ABSTR_IRAM_0, WR_ADDR_ABSTR_IRAM_0, WR_DATA_ABSTR_IRAM_0, WR_COND_ABSTR_IRAM_1, WR_ADDR_ABSTR_IRAM_1, WR_DATA_ABSTR_IRAM_1, p0_in, p1_in, p2_in, p3_in, property_invalid_pc, property_invalid_acc, property_invalid_b_reg, property_invalid_dpl, property_invalid_dph, property_invalid_iram, property_invalid_p0, property_invalid_p1, property_invalid_p2, property_invalid_p3, property_invalid_psw, property_invalid_xram_addr, property_invalid_xram_data_out);
  wire _00000_;
  wire _00001_;
  wire _00002_;
  wire _00003_;
  wire [7:0] _00004_;
  wire [7:0] _00005_;
  wire [7:0] _00006_;
  wire [7:0] _00007_;
  wire _00008_;
  wire _00009_;
  wire [7:0] _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  wire _08001_;
  wire _08002_;
  wire _08003_;
  wire _08004_;
  wire _08005_;
  wire _08006_;
  wire _08007_;
  wire _08008_;
  wire _08009_;
  wire _08010_;
  wire _08011_;
  wire _08012_;
  wire _08013_;
  wire _08014_;
  wire _08015_;
  wire _08016_;
  wire _08017_;
  wire _08018_;
  wire _08019_;
  wire _08020_;
  wire _08021_;
  wire _08022_;
  wire _08023_;
  wire _08024_;
  wire _08025_;
  wire _08026_;
  wire _08027_;
  wire _08028_;
  wire _08029_;
  wire _08030_;
  wire _08031_;
  wire _08032_;
  wire _08033_;
  wire _08034_;
  wire _08035_;
  wire _08036_;
  wire _08037_;
  wire _08038_;
  wire _08039_;
  wire _08040_;
  wire _08041_;
  wire _08042_;
  wire _08043_;
  wire _08044_;
  wire _08045_;
  wire _08046_;
  wire _08047_;
  wire _08048_;
  wire _08049_;
  wire _08050_;
  wire _08051_;
  wire _08052_;
  wire _08053_;
  wire _08054_;
  wire _08055_;
  wire _08056_;
  wire _08057_;
  wire _08058_;
  wire _08059_;
  wire _08060_;
  wire _08061_;
  wire _08062_;
  wire _08063_;
  wire _08064_;
  wire _08065_;
  wire _08066_;
  wire _08067_;
  wire _08068_;
  wire _08069_;
  wire _08070_;
  wire _08071_;
  wire _08072_;
  wire _08073_;
  wire _08074_;
  wire _08075_;
  wire _08076_;
  wire _08077_;
  wire _08078_;
  wire _08079_;
  wire _08080_;
  wire _08081_;
  wire _08082_;
  wire _08083_;
  wire _08084_;
  wire _08085_;
  wire _08086_;
  wire _08087_;
  wire _08088_;
  wire _08089_;
  wire _08090_;
  wire _08091_;
  wire _08092_;
  wire _08093_;
  wire _08094_;
  wire _08095_;
  wire _08096_;
  wire _08097_;
  wire _08098_;
  wire _08099_;
  wire _08100_;
  wire _08101_;
  wire _08102_;
  wire _08103_;
  wire _08104_;
  wire _08105_;
  wire _08106_;
  wire _08107_;
  wire _08108_;
  wire _08109_;
  wire _08110_;
  wire _08111_;
  wire _08112_;
  wire _08113_;
  wire _08114_;
  wire _08115_;
  wire _08116_;
  wire _08117_;
  wire _08118_;
  wire _08119_;
  wire _08120_;
  wire _08121_;
  wire _08122_;
  wire _08123_;
  wire _08124_;
  wire _08125_;
  wire _08126_;
  wire _08127_;
  wire _08128_;
  wire _08129_;
  wire _08130_;
  wire _08131_;
  wire _08132_;
  wire _08133_;
  wire _08134_;
  wire _08135_;
  wire _08136_;
  wire _08137_;
  wire _08138_;
  wire _08139_;
  wire _08140_;
  wire _08141_;
  wire _08142_;
  wire _08143_;
  wire _08144_;
  wire _08145_;
  wire _08146_;
  wire _08147_;
  wire _08148_;
  wire _08149_;
  wire _08150_;
  wire _08151_;
  wire _08152_;
  wire _08153_;
  wire _08154_;
  wire _08155_;
  wire _08156_;
  wire _08157_;
  wire _08158_;
  wire _08159_;
  wire _08160_;
  wire _08161_;
  wire _08162_;
  wire _08163_;
  wire _08164_;
  wire _08165_;
  wire _08166_;
  wire _08167_;
  wire _08168_;
  wire _08169_;
  wire _08170_;
  wire _08171_;
  wire _08172_;
  wire _08173_;
  wire _08174_;
  wire _08175_;
  wire _08176_;
  wire _08177_;
  wire _08178_;
  wire _08179_;
  wire _08180_;
  wire _08181_;
  wire _08182_;
  wire _08183_;
  wire _08184_;
  wire _08185_;
  wire _08186_;
  wire _08187_;
  wire _08188_;
  wire _08189_;
  wire _08190_;
  wire _08191_;
  wire _08192_;
  wire _08193_;
  wire _08194_;
  wire _08195_;
  wire _08196_;
  wire _08197_;
  wire _08198_;
  wire _08199_;
  wire _08200_;
  wire _08201_;
  wire _08202_;
  wire _08203_;
  wire _08204_;
  wire _08205_;
  wire _08206_;
  wire _08207_;
  wire _08208_;
  wire _08209_;
  wire _08210_;
  wire _08211_;
  wire _08212_;
  wire _08213_;
  wire _08214_;
  wire _08215_;
  wire _08216_;
  wire _08217_;
  wire _08218_;
  wire _08219_;
  wire _08220_;
  wire _08221_;
  wire _08222_;
  wire _08223_;
  wire _08224_;
  wire _08225_;
  wire _08226_;
  wire _08227_;
  wire _08228_;
  wire _08229_;
  wire _08230_;
  wire _08231_;
  wire _08232_;
  wire _08233_;
  wire _08234_;
  wire _08235_;
  wire _08236_;
  wire _08237_;
  wire _08238_;
  wire _08239_;
  wire _08240_;
  wire _08241_;
  wire _08242_;
  wire _08243_;
  wire _08244_;
  wire _08245_;
  wire _08246_;
  wire _08247_;
  wire _08248_;
  wire _08249_;
  wire _08250_;
  wire _08251_;
  wire _08252_;
  wire _08253_;
  wire _08254_;
  wire _08255_;
  wire _08256_;
  wire _08257_;
  wire _08258_;
  wire _08259_;
  wire _08260_;
  wire _08261_;
  wire _08262_;
  wire _08263_;
  wire _08264_;
  wire _08265_;
  wire _08266_;
  wire _08267_;
  wire _08268_;
  wire _08269_;
  wire _08270_;
  wire _08271_;
  wire _08272_;
  wire _08273_;
  wire _08274_;
  wire _08275_;
  wire _08276_;
  wire _08277_;
  wire _08278_;
  wire _08279_;
  wire _08280_;
  wire _08281_;
  wire _08282_;
  wire _08283_;
  wire _08284_;
  wire _08285_;
  wire _08286_;
  wire _08287_;
  wire _08288_;
  wire _08289_;
  wire _08290_;
  wire _08291_;
  wire _08292_;
  wire _08293_;
  wire _08294_;
  wire _08295_;
  wire _08296_;
  wire _08297_;
  wire _08298_;
  wire _08299_;
  wire _08300_;
  wire _08301_;
  wire _08302_;
  wire _08303_;
  wire _08304_;
  wire _08305_;
  wire _08306_;
  wire _08307_;
  wire _08308_;
  wire _08309_;
  wire _08310_;
  wire _08311_;
  wire _08312_;
  wire _08313_;
  wire _08314_;
  wire _08315_;
  wire _08316_;
  wire _08317_;
  wire _08318_;
  wire _08319_;
  wire _08320_;
  wire _08321_;
  wire _08322_;
  wire _08323_;
  wire _08324_;
  wire _08325_;
  wire _08326_;
  wire _08327_;
  wire _08328_;
  wire _08329_;
  wire _08330_;
  wire _08331_;
  wire _08332_;
  wire _08333_;
  wire _08334_;
  wire _08335_;
  wire _08336_;
  wire _08337_;
  wire _08338_;
  wire _08339_;
  wire _08340_;
  wire _08341_;
  wire _08342_;
  wire _08343_;
  wire _08344_;
  wire _08345_;
  wire _08346_;
  wire _08347_;
  wire _08348_;
  wire _08349_;
  wire _08350_;
  wire _08351_;
  wire _08352_;
  wire _08353_;
  wire _08354_;
  wire _08355_;
  wire _08356_;
  wire _08357_;
  wire _08358_;
  wire _08359_;
  wire _08360_;
  wire _08361_;
  wire _08362_;
  wire _08363_;
  wire _08364_;
  wire _08365_;
  wire _08366_;
  wire _08367_;
  wire _08368_;
  wire _08369_;
  wire _08370_;
  wire _08371_;
  wire _08372_;
  wire _08373_;
  wire _08374_;
  wire _08375_;
  wire _08376_;
  wire _08377_;
  wire _08378_;
  wire _08379_;
  wire _08380_;
  wire _08381_;
  wire _08382_;
  wire _08383_;
  wire _08384_;
  wire _08385_;
  wire _08386_;
  wire _08387_;
  wire _08388_;
  wire _08389_;
  wire _08390_;
  wire _08391_;
  wire _08392_;
  wire _08393_;
  wire _08394_;
  wire _08395_;
  wire _08396_;
  wire _08397_;
  wire _08398_;
  wire _08399_;
  wire _08400_;
  wire _08401_;
  wire _08402_;
  wire _08403_;
  wire _08404_;
  wire _08405_;
  wire _08406_;
  wire _08407_;
  wire _08408_;
  wire _08409_;
  wire _08410_;
  wire _08411_;
  wire _08412_;
  wire _08413_;
  wire _08414_;
  wire _08415_;
  wire _08416_;
  wire _08417_;
  wire _08418_;
  wire _08419_;
  wire _08420_;
  wire _08421_;
  wire _08422_;
  wire _08423_;
  wire _08424_;
  wire _08425_;
  wire _08426_;
  wire _08427_;
  wire _08428_;
  wire _08429_;
  wire _08430_;
  wire _08431_;
  wire _08432_;
  wire _08433_;
  wire _08434_;
  wire _08435_;
  wire _08436_;
  wire _08437_;
  wire _08438_;
  wire _08439_;
  wire _08440_;
  wire _08441_;
  wire _08442_;
  wire _08443_;
  wire _08444_;
  wire _08445_;
  wire _08446_;
  wire _08447_;
  wire _08448_;
  wire _08449_;
  wire _08450_;
  wire _08451_;
  wire _08452_;
  wire _08453_;
  wire _08454_;
  wire _08455_;
  wire _08456_;
  wire _08457_;
  wire _08458_;
  wire _08459_;
  wire _08460_;
  wire _08461_;
  wire _08462_;
  wire _08463_;
  wire _08464_;
  wire _08465_;
  wire _08466_;
  wire _08467_;
  wire _08468_;
  wire _08469_;
  wire _08470_;
  wire _08471_;
  wire _08472_;
  wire _08473_;
  wire _08474_;
  wire _08475_;
  wire _08476_;
  wire _08477_;
  wire _08478_;
  wire _08479_;
  wire _08480_;
  wire _08481_;
  wire _08482_;
  wire _08483_;
  wire _08484_;
  wire _08485_;
  wire _08486_;
  wire _08487_;
  wire _08488_;
  wire _08489_;
  wire _08490_;
  wire _08491_;
  wire _08492_;
  wire _08493_;
  wire _08494_;
  wire _08495_;
  wire _08496_;
  wire _08497_;
  wire _08498_;
  wire _08499_;
  wire _08500_;
  wire _08501_;
  wire _08502_;
  wire _08503_;
  wire _08504_;
  wire _08505_;
  wire _08506_;
  wire _08507_;
  wire _08508_;
  wire _08509_;
  wire _08510_;
  wire _08511_;
  wire _08512_;
  wire _08513_;
  wire _08514_;
  wire _08515_;
  wire _08516_;
  wire _08517_;
  wire _08518_;
  wire _08519_;
  wire _08520_;
  wire _08521_;
  wire _08522_;
  wire _08523_;
  wire _08524_;
  wire _08525_;
  wire _08526_;
  wire _08527_;
  wire _08528_;
  wire _08529_;
  wire _08530_;
  wire _08531_;
  wire _08532_;
  wire _08533_;
  wire _08534_;
  wire _08535_;
  wire _08536_;
  wire _08537_;
  wire _08538_;
  wire _08539_;
  wire _08540_;
  wire _08541_;
  wire _08542_;
  wire _08543_;
  wire _08544_;
  wire _08545_;
  wire _08546_;
  wire _08547_;
  wire _08548_;
  wire _08549_;
  wire _08550_;
  wire _08551_;
  wire _08552_;
  wire _08553_;
  wire _08554_;
  wire _08555_;
  wire _08556_;
  wire _08557_;
  wire _08558_;
  wire _08559_;
  wire _08560_;
  wire _08561_;
  wire _08562_;
  wire _08563_;
  wire _08564_;
  wire _08565_;
  wire _08566_;
  wire _08567_;
  wire _08568_;
  wire _08569_;
  wire _08570_;
  wire _08571_;
  wire _08572_;
  wire _08573_;
  wire _08574_;
  wire _08575_;
  wire _08576_;
  wire _08577_;
  wire _08578_;
  wire _08579_;
  wire _08580_;
  wire _08581_;
  wire _08582_;
  wire _08583_;
  wire _08584_;
  wire _08585_;
  wire _08586_;
  wire _08587_;
  wire _08588_;
  wire _08589_;
  wire _08590_;
  wire _08591_;
  wire _08592_;
  wire _08593_;
  wire _08594_;
  wire _08595_;
  wire _08596_;
  wire _08597_;
  wire _08598_;
  wire _08599_;
  wire _08600_;
  wire _08601_;
  wire _08602_;
  wire _08603_;
  wire _08604_;
  wire _08605_;
  wire _08606_;
  wire _08607_;
  wire _08608_;
  wire _08609_;
  wire _08610_;
  wire _08611_;
  wire _08612_;
  wire _08613_;
  wire _08614_;
  wire _08615_;
  wire _08616_;
  wire _08617_;
  wire _08618_;
  wire _08619_;
  wire _08620_;
  wire _08621_;
  wire _08622_;
  wire _08623_;
  wire _08624_;
  wire _08625_;
  wire _08626_;
  wire _08627_;
  wire _08628_;
  wire _08629_;
  wire _08630_;
  wire _08631_;
  wire _08632_;
  wire _08633_;
  wire _08634_;
  wire _08635_;
  wire _08636_;
  wire _08637_;
  wire _08638_;
  wire _08639_;
  wire _08640_;
  wire _08641_;
  wire _08642_;
  wire _08643_;
  wire _08644_;
  wire _08645_;
  wire _08646_;
  wire _08647_;
  wire _08648_;
  wire _08649_;
  wire _08650_;
  wire _08651_;
  wire _08652_;
  wire _08653_;
  wire _08654_;
  wire _08655_;
  wire _08656_;
  wire _08657_;
  wire _08658_;
  wire _08659_;
  wire _08660_;
  wire _08661_;
  wire _08662_;
  wire _08663_;
  wire _08664_;
  wire _08665_;
  wire _08666_;
  wire _08667_;
  wire _08668_;
  wire _08669_;
  wire _08670_;
  wire _08671_;
  wire _08672_;
  wire _08673_;
  wire _08674_;
  wire _08675_;
  wire _08676_;
  wire _08677_;
  wire _08678_;
  wire _08679_;
  wire _08680_;
  wire _08681_;
  wire _08682_;
  wire _08683_;
  wire _08684_;
  wire _08685_;
  wire _08686_;
  wire _08687_;
  wire _08688_;
  wire _08689_;
  wire _08690_;
  wire _08691_;
  wire _08692_;
  wire _08693_;
  wire _08694_;
  wire _08695_;
  wire _08696_;
  wire _08697_;
  wire _08698_;
  wire _08699_;
  wire _08700_;
  wire _08701_;
  wire _08702_;
  wire _08703_;
  wire _08704_;
  wire _08705_;
  wire _08706_;
  wire _08707_;
  wire _08708_;
  wire _08709_;
  wire _08710_;
  wire _08711_;
  wire _08712_;
  wire _08713_;
  wire _08714_;
  wire _08715_;
  wire _08716_;
  wire _08717_;
  wire _08718_;
  wire _08719_;
  wire _08720_;
  wire _08721_;
  wire _08722_;
  wire _08723_;
  wire _08724_;
  wire _08725_;
  wire _08726_;
  wire _08727_;
  wire _08728_;
  wire _08729_;
  wire _08730_;
  wire _08731_;
  wire _08732_;
  wire _08733_;
  wire _08734_;
  wire _08735_;
  wire _08736_;
  wire _08737_;
  wire _08738_;
  wire _08739_;
  wire _08740_;
  wire _08741_;
  wire _08742_;
  wire _08743_;
  wire _08744_;
  wire _08745_;
  wire _08746_;
  wire _08747_;
  wire _08748_;
  wire _08749_;
  wire _08750_;
  wire _08751_;
  wire _08752_;
  wire _08753_;
  wire _08754_;
  wire _08755_;
  wire _08756_;
  wire _08757_;
  wire _08758_;
  wire _08759_;
  wire _08760_;
  wire _08761_;
  wire _08762_;
  wire _08763_;
  wire _08764_;
  wire _08765_;
  wire _08766_;
  wire _08767_;
  wire _08768_;
  wire _08769_;
  wire _08770_;
  wire _08771_;
  wire _08772_;
  wire _08773_;
  wire _08774_;
  wire _08775_;
  wire _08776_;
  wire _08777_;
  wire _08778_;
  wire _08779_;
  wire _08780_;
  wire _08781_;
  wire _08782_;
  wire _08783_;
  wire _08784_;
  wire _08785_;
  wire _08786_;
  wire _08787_;
  wire _08788_;
  wire _08789_;
  wire _08790_;
  wire _08791_;
  wire _08792_;
  wire _08793_;
  wire _08794_;
  wire _08795_;
  wire _08796_;
  wire _08797_;
  wire _08798_;
  wire _08799_;
  wire _08800_;
  wire _08801_;
  wire _08802_;
  wire _08803_;
  wire _08804_;
  wire _08805_;
  wire _08806_;
  wire _08807_;
  wire _08808_;
  wire _08809_;
  wire _08810_;
  wire _08811_;
  wire _08812_;
  wire _08813_;
  wire _08814_;
  wire _08815_;
  wire _08816_;
  wire _08817_;
  wire _08818_;
  wire _08819_;
  wire _08820_;
  wire _08821_;
  wire _08822_;
  wire _08823_;
  wire _08824_;
  wire _08825_;
  wire _08826_;
  wire _08827_;
  wire _08828_;
  wire _08829_;
  wire _08830_;
  wire _08831_;
  wire _08832_;
  wire _08833_;
  wire _08834_;
  wire _08835_;
  wire _08836_;
  wire _08837_;
  wire _08838_;
  wire _08839_;
  wire _08840_;
  wire _08841_;
  wire _08842_;
  wire _08843_;
  wire _08844_;
  wire _08845_;
  wire _08846_;
  wire _08847_;
  wire _08848_;
  wire _08849_;
  wire _08850_;
  wire _08851_;
  wire _08852_;
  wire _08853_;
  wire _08854_;
  wire _08855_;
  wire _08856_;
  wire _08857_;
  wire _08858_;
  wire _08859_;
  wire _08860_;
  wire _08861_;
  wire _08862_;
  wire _08863_;
  wire _08864_;
  wire _08865_;
  wire _08866_;
  wire _08867_;
  wire _08868_;
  wire _08869_;
  wire _08870_;
  wire _08871_;
  wire _08872_;
  wire _08873_;
  wire _08874_;
  wire _08875_;
  wire _08876_;
  wire _08877_;
  wire _08878_;
  wire _08879_;
  wire _08880_;
  wire _08881_;
  wire _08882_;
  wire _08883_;
  wire _08884_;
  wire _08885_;
  wire _08886_;
  wire _08887_;
  wire _08888_;
  wire _08889_;
  wire _08890_;
  wire _08891_;
  wire _08892_;
  wire _08893_;
  wire _08894_;
  wire _08895_;
  wire _08896_;
  wire _08897_;
  wire _08898_;
  wire _08899_;
  wire _08900_;
  wire _08901_;
  wire _08902_;
  wire _08903_;
  wire _08904_;
  wire _08905_;
  wire _08906_;
  wire _08907_;
  wire _08908_;
  wire _08909_;
  wire _08910_;
  wire _08911_;
  wire _08912_;
  wire _08913_;
  wire _08914_;
  wire _08915_;
  wire _08916_;
  wire _08917_;
  wire _08918_;
  wire _08919_;
  wire _08920_;
  wire _08921_;
  wire _08922_;
  wire _08923_;
  wire _08924_;
  wire _08925_;
  wire _08926_;
  wire _08927_;
  wire _08928_;
  wire _08929_;
  wire _08930_;
  wire _08931_;
  wire _08932_;
  wire _08933_;
  wire _08934_;
  wire _08935_;
  wire _08936_;
  wire _08937_;
  wire _08938_;
  wire _08939_;
  wire _08940_;
  wire _08941_;
  wire _08942_;
  wire _08943_;
  wire _08944_;
  wire _08945_;
  wire _08946_;
  wire _08947_;
  wire _08948_;
  wire _08949_;
  wire _08950_;
  wire _08951_;
  wire _08952_;
  wire _08953_;
  wire _08954_;
  wire _08955_;
  wire _08956_;
  wire _08957_;
  wire _08958_;
  wire _08959_;
  wire _08960_;
  wire _08961_;
  wire _08962_;
  wire _08963_;
  wire _08964_;
  wire _08965_;
  wire _08966_;
  wire _08967_;
  wire _08968_;
  wire _08969_;
  wire _08970_;
  wire _08971_;
  wire _08972_;
  wire _08973_;
  wire _08974_;
  wire _08975_;
  wire _08976_;
  wire _08977_;
  wire _08978_;
  wire _08979_;
  wire _08980_;
  wire _08981_;
  wire _08982_;
  wire _08983_;
  wire _08984_;
  wire _08985_;
  wire _08986_;
  wire _08987_;
  wire _08988_;
  wire _08989_;
  wire _08990_;
  wire _08991_;
  wire _08992_;
  wire _08993_;
  wire _08994_;
  wire _08995_;
  wire _08996_;
  wire _08997_;
  wire _08998_;
  wire _08999_;
  wire _09000_;
  wire _09001_;
  wire _09002_;
  wire _09003_;
  wire _09004_;
  wire _09005_;
  wire _09006_;
  wire _09007_;
  wire _09008_;
  wire _09009_;
  wire _09010_;
  wire _09011_;
  wire _09012_;
  wire _09013_;
  wire _09014_;
  wire _09015_;
  wire _09016_;
  wire _09017_;
  wire _09018_;
  wire _09019_;
  wire _09020_;
  wire _09021_;
  wire _09022_;
  wire _09023_;
  wire _09024_;
  wire _09025_;
  wire _09026_;
  wire _09027_;
  wire _09028_;
  wire _09029_;
  wire _09030_;
  wire _09031_;
  wire _09032_;
  wire _09033_;
  wire _09034_;
  wire _09035_;
  wire _09036_;
  wire _09037_;
  wire _09038_;
  wire _09039_;
  wire _09040_;
  wire _09041_;
  wire _09042_;
  wire _09043_;
  wire _09044_;
  wire _09045_;
  wire _09046_;
  wire _09047_;
  wire _09048_;
  wire _09049_;
  wire _09050_;
  wire _09051_;
  wire _09052_;
  wire _09053_;
  wire _09054_;
  wire _09055_;
  wire _09056_;
  wire _09057_;
  wire _09058_;
  wire _09059_;
  wire _09060_;
  wire _09061_;
  wire _09062_;
  wire _09063_;
  wire _09064_;
  wire _09065_;
  wire _09066_;
  wire _09067_;
  wire _09068_;
  wire _09069_;
  wire _09070_;
  wire _09071_;
  wire _09072_;
  wire _09073_;
  wire _09074_;
  wire _09075_;
  wire _09076_;
  wire _09077_;
  wire _09078_;
  wire _09079_;
  wire _09080_;
  wire _09081_;
  wire _09082_;
  wire _09083_;
  wire _09084_;
  wire _09085_;
  wire _09086_;
  wire _09087_;
  wire _09088_;
  wire _09089_;
  wire _09090_;
  wire _09091_;
  wire _09092_;
  wire _09093_;
  wire _09094_;
  wire _09095_;
  wire _09096_;
  wire _09097_;
  wire _09098_;
  wire _09099_;
  wire _09100_;
  wire _09101_;
  wire _09102_;
  wire _09103_;
  wire _09104_;
  wire _09105_;
  wire _09106_;
  wire _09107_;
  wire _09108_;
  wire _09109_;
  wire _09110_;
  wire _09111_;
  wire _09112_;
  wire _09113_;
  wire _09114_;
  wire _09115_;
  wire _09116_;
  wire _09117_;
  wire _09118_;
  wire _09119_;
  wire _09120_;
  wire _09121_;
  wire _09122_;
  wire _09123_;
  wire _09124_;
  wire _09125_;
  wire _09126_;
  wire _09127_;
  wire _09128_;
  wire _09129_;
  wire _09130_;
  wire _09131_;
  wire _09132_;
  wire _09133_;
  wire _09134_;
  wire _09135_;
  wire _09136_;
  wire _09137_;
  wire _09138_;
  wire _09139_;
  wire _09140_;
  wire _09141_;
  wire _09142_;
  wire _09143_;
  wire _09144_;
  wire _09145_;
  wire _09146_;
  wire _09147_;
  wire _09148_;
  wire _09149_;
  wire _09150_;
  wire _09151_;
  wire _09152_;
  wire _09153_;
  wire _09154_;
  wire _09155_;
  wire _09156_;
  wire _09157_;
  wire _09158_;
  wire _09159_;
  wire _09160_;
  wire _09161_;
  wire _09162_;
  wire _09163_;
  wire _09164_;
  wire _09165_;
  wire _09166_;
  wire _09167_;
  wire _09168_;
  wire _09169_;
  wire _09170_;
  wire _09171_;
  wire _09172_;
  wire _09173_;
  wire _09174_;
  wire _09175_;
  wire _09176_;
  wire _09177_;
  wire _09178_;
  wire _09179_;
  wire _09180_;
  wire _09181_;
  wire _09182_;
  wire _09183_;
  wire _09184_;
  wire _09185_;
  wire _09186_;
  wire _09187_;
  wire _09188_;
  wire _09189_;
  wire _09190_;
  wire _09191_;
  wire _09192_;
  wire _09193_;
  wire _09194_;
  wire _09195_;
  wire _09196_;
  wire _09197_;
  wire _09198_;
  wire _09199_;
  wire _09200_;
  wire _09201_;
  wire _09202_;
  wire _09203_;
  wire _09204_;
  wire _09205_;
  wire _09206_;
  wire _09207_;
  wire _09208_;
  wire _09209_;
  wire _09210_;
  wire _09211_;
  wire _09212_;
  wire _09213_;
  wire _09214_;
  wire _09215_;
  wire _09216_;
  wire _09217_;
  wire _09218_;
  wire _09219_;
  wire _09220_;
  wire _09221_;
  wire _09222_;
  wire _09223_;
  wire _09224_;
  wire _09225_;
  wire _09226_;
  wire _09227_;
  wire _09228_;
  wire _09229_;
  wire _09230_;
  wire _09231_;
  wire _09232_;
  wire _09233_;
  wire _09234_;
  wire _09235_;
  wire _09236_;
  wire _09237_;
  wire _09238_;
  wire _09239_;
  wire _09240_;
  wire _09241_;
  wire _09242_;
  wire _09243_;
  wire _09244_;
  wire _09245_;
  wire _09246_;
  wire _09247_;
  wire _09248_;
  wire _09249_;
  wire _09250_;
  wire _09251_;
  wire _09252_;
  wire _09253_;
  wire _09254_;
  wire _09255_;
  wire _09256_;
  wire _09257_;
  wire _09258_;
  wire _09259_;
  wire _09260_;
  wire _09261_;
  wire _09262_;
  wire _09263_;
  wire _09264_;
  wire _09265_;
  wire _09266_;
  wire _09267_;
  wire _09268_;
  wire _09269_;
  wire _09270_;
  wire _09271_;
  wire _09272_;
  wire _09273_;
  wire _09274_;
  wire _09275_;
  wire _09276_;
  wire _09277_;
  wire _09278_;
  wire _09279_;
  wire _09280_;
  wire _09281_;
  wire _09282_;
  wire _09283_;
  wire _09284_;
  wire _09285_;
  wire _09286_;
  wire _09287_;
  wire _09288_;
  wire _09289_;
  wire _09290_;
  wire _09291_;
  wire _09292_;
  wire _09293_;
  wire _09294_;
  wire _09295_;
  wire _09296_;
  wire _09297_;
  wire _09298_;
  wire _09299_;
  wire _09300_;
  wire _09301_;
  wire _09302_;
  wire _09303_;
  wire _09304_;
  wire _09305_;
  wire _09306_;
  wire _09307_;
  wire _09308_;
  wire _09309_;
  wire _09310_;
  wire _09311_;
  wire _09312_;
  wire _09313_;
  wire _09314_;
  wire _09315_;
  wire _09316_;
  wire _09317_;
  wire _09318_;
  wire _09319_;
  wire _09320_;
  wire _09321_;
  wire _09322_;
  wire _09323_;
  wire _09324_;
  wire _09325_;
  wire _09326_;
  wire _09327_;
  wire _09328_;
  wire _09329_;
  wire _09330_;
  wire _09331_;
  wire _09332_;
  wire _09333_;
  wire _09334_;
  wire _09335_;
  wire _09336_;
  wire _09337_;
  wire _09338_;
  wire _09339_;
  wire _09340_;
  wire _09341_;
  wire _09342_;
  wire _09343_;
  wire _09344_;
  wire _09345_;
  wire _09346_;
  wire _09347_;
  wire _09348_;
  wire _09349_;
  wire _09350_;
  wire _09351_;
  wire _09352_;
  wire _09353_;
  wire _09354_;
  wire _09355_;
  wire _09356_;
  wire _09357_;
  wire _09358_;
  wire _09359_;
  wire _09360_;
  wire _09361_;
  wire _09362_;
  wire _09363_;
  wire _09364_;
  wire _09365_;
  wire _09366_;
  wire _09367_;
  wire _09368_;
  wire _09369_;
  wire _09370_;
  wire _09371_;
  wire _09372_;
  wire _09373_;
  wire _09374_;
  wire _09375_;
  wire _09376_;
  wire _09377_;
  wire _09378_;
  wire _09379_;
  wire _09380_;
  wire _09381_;
  wire _09382_;
  wire _09383_;
  wire _09384_;
  wire _09385_;
  wire _09386_;
  wire _09387_;
  wire _09388_;
  wire _09389_;
  wire _09390_;
  wire _09391_;
  wire _09392_;
  wire _09393_;
  wire _09394_;
  wire _09395_;
  wire _09396_;
  wire _09397_;
  wire _09398_;
  wire _09399_;
  wire _09400_;
  wire _09401_;
  wire _09402_;
  wire _09403_;
  wire _09404_;
  wire _09405_;
  wire _09406_;
  wire _09407_;
  wire _09408_;
  wire _09409_;
  wire _09410_;
  wire _09411_;
  wire _09412_;
  wire _09413_;
  wire _09414_;
  wire _09415_;
  wire _09416_;
  wire _09417_;
  wire _09418_;
  wire _09419_;
  wire _09420_;
  wire _09421_;
  wire _09422_;
  wire _09423_;
  wire _09424_;
  wire _09425_;
  wire _09426_;
  wire _09427_;
  wire _09428_;
  wire _09429_;
  wire _09430_;
  wire _09431_;
  wire _09432_;
  wire _09433_;
  wire _09434_;
  wire _09435_;
  wire _09436_;
  wire _09437_;
  wire _09438_;
  wire _09439_;
  wire _09440_;
  wire _09441_;
  wire _09442_;
  wire _09443_;
  wire _09444_;
  wire _09445_;
  wire _09446_;
  wire _09447_;
  wire _09448_;
  wire _09449_;
  wire _09450_;
  wire _09451_;
  wire _09452_;
  wire _09453_;
  wire _09454_;
  wire _09455_;
  wire _09456_;
  wire _09457_;
  wire _09458_;
  wire _09459_;
  wire _09460_;
  wire _09461_;
  wire _09462_;
  wire _09463_;
  wire _09464_;
  wire _09465_;
  wire _09466_;
  wire _09467_;
  wire _09468_;
  wire _09469_;
  wire _09470_;
  wire _09471_;
  wire _09472_;
  wire _09473_;
  wire _09474_;
  wire _09475_;
  wire _09476_;
  wire _09477_;
  wire _09478_;
  wire _09479_;
  wire _09480_;
  wire _09481_;
  wire _09482_;
  wire _09483_;
  wire _09484_;
  wire _09485_;
  wire _09486_;
  wire _09487_;
  wire _09488_;
  wire _09489_;
  wire _09490_;
  wire _09491_;
  wire _09492_;
  wire _09493_;
  wire _09494_;
  wire _09495_;
  wire _09496_;
  wire _09497_;
  wire _09498_;
  wire _09499_;
  wire _09500_;
  wire _09501_;
  wire _09502_;
  wire _09503_;
  wire _09504_;
  wire _09505_;
  wire _09506_;
  wire _09507_;
  wire _09508_;
  wire _09509_;
  wire _09510_;
  wire _09511_;
  wire _09512_;
  wire _09513_;
  wire _09514_;
  wire _09515_;
  wire _09516_;
  wire _09517_;
  wire _09518_;
  wire _09519_;
  wire _09520_;
  wire _09521_;
  wire _09522_;
  wire _09523_;
  wire _09524_;
  wire _09525_;
  wire _09526_;
  wire _09527_;
  wire _09528_;
  wire _09529_;
  wire _09530_;
  wire _09531_;
  wire _09532_;
  wire _09533_;
  wire _09534_;
  wire _09535_;
  wire _09536_;
  wire _09537_;
  wire _09538_;
  wire _09539_;
  wire _09540_;
  wire _09541_;
  wire _09542_;
  wire _09543_;
  wire _09544_;
  wire _09545_;
  wire _09546_;
  wire _09547_;
  wire _09548_;
  wire _09549_;
  wire _09550_;
  wire _09551_;
  wire _09552_;
  wire _09553_;
  wire _09554_;
  wire _09555_;
  wire _09556_;
  wire _09557_;
  wire _09558_;
  wire _09559_;
  wire _09560_;
  wire _09561_;
  wire _09562_;
  wire _09563_;
  wire _09564_;
  wire _09565_;
  wire _09566_;
  wire _09567_;
  wire _09568_;
  wire _09569_;
  wire _09570_;
  wire _09571_;
  wire _09572_;
  wire _09573_;
  wire _09574_;
  wire _09575_;
  wire _09576_;
  wire _09577_;
  wire _09578_;
  wire _09579_;
  wire _09580_;
  wire _09581_;
  wire _09582_;
  wire _09583_;
  wire _09584_;
  wire _09585_;
  wire _09586_;
  wire _09587_;
  wire _09588_;
  wire _09589_;
  wire _09590_;
  wire _09591_;
  wire _09592_;
  wire _09593_;
  wire _09594_;
  wire _09595_;
  wire _09596_;
  wire _09597_;
  wire _09598_;
  wire _09599_;
  wire _09600_;
  wire _09601_;
  wire _09602_;
  wire _09603_;
  wire _09604_;
  wire _09605_;
  wire _09606_;
  wire _09607_;
  wire _09608_;
  wire _09609_;
  wire _09610_;
  wire _09611_;
  wire _09612_;
  wire _09613_;
  wire _09614_;
  wire _09615_;
  wire _09616_;
  wire _09617_;
  wire _09618_;
  wire _09619_;
  wire _09620_;
  wire _09621_;
  wire _09622_;
  wire _09623_;
  wire _09624_;
  wire _09625_;
  wire _09626_;
  wire _09627_;
  wire _09628_;
  wire _09629_;
  wire _09630_;
  wire _09631_;
  wire _09632_;
  wire _09633_;
  wire _09634_;
  wire _09635_;
  wire _09636_;
  wire _09637_;
  wire _09638_;
  wire _09639_;
  wire _09640_;
  wire _09641_;
  wire _09642_;
  wire _09643_;
  wire _09644_;
  wire _09645_;
  wire _09646_;
  wire _09647_;
  wire _09648_;
  wire _09649_;
  wire _09650_;
  wire _09651_;
  wire _09652_;
  wire _09653_;
  wire _09654_;
  wire _09655_;
  wire _09656_;
  wire _09657_;
  wire _09658_;
  wire _09659_;
  wire _09660_;
  wire _09661_;
  wire _09662_;
  wire _09663_;
  wire _09664_;
  wire _09665_;
  wire _09666_;
  wire _09667_;
  wire _09668_;
  wire _09669_;
  wire _09670_;
  wire _09671_;
  wire _09672_;
  wire _09673_;
  wire _09674_;
  wire _09675_;
  wire _09676_;
  wire _09677_;
  wire _09678_;
  wire _09679_;
  wire _09680_;
  wire _09681_;
  wire _09682_;
  wire _09683_;
  wire _09684_;
  wire _09685_;
  wire _09686_;
  wire _09687_;
  wire _09688_;
  wire _09689_;
  wire _09690_;
  wire _09691_;
  wire _09692_;
  wire _09693_;
  wire _09694_;
  wire _09695_;
  wire _09696_;
  wire _09697_;
  wire _09698_;
  wire _09699_;
  wire _09700_;
  wire _09701_;
  wire _09702_;
  wire _09703_;
  wire _09704_;
  wire _09705_;
  wire _09706_;
  wire _09707_;
  wire _09708_;
  wire _09709_;
  wire _09710_;
  wire _09711_;
  wire _09712_;
  wire _09713_;
  wire _09714_;
  wire _09715_;
  wire _09716_;
  wire _09717_;
  wire _09718_;
  wire _09719_;
  wire _09720_;
  wire _09721_;
  wire _09722_;
  wire _09723_;
  wire _09724_;
  wire _09725_;
  wire _09726_;
  wire _09727_;
  wire _09728_;
  wire _09729_;
  wire _09730_;
  wire _09731_;
  wire _09732_;
  wire _09733_;
  wire _09734_;
  wire _09735_;
  wire _09736_;
  wire _09737_;
  wire _09738_;
  wire _09739_;
  wire _09740_;
  wire _09741_;
  wire _09742_;
  wire _09743_;
  wire _09744_;
  wire _09745_;
  wire _09746_;
  wire _09747_;
  wire _09748_;
  wire _09749_;
  wire _09750_;
  wire _09751_;
  wire _09752_;
  wire _09753_;
  wire _09754_;
  wire _09755_;
  wire _09756_;
  wire _09757_;
  wire _09758_;
  wire _09759_;
  wire _09760_;
  wire _09761_;
  wire _09762_;
  wire _09763_;
  wire _09764_;
  wire _09765_;
  wire _09766_;
  wire _09767_;
  wire _09768_;
  wire _09769_;
  wire _09770_;
  wire _09771_;
  wire _09772_;
  wire _09773_;
  wire _09774_;
  wire _09775_;
  wire _09776_;
  wire _09777_;
  wire _09778_;
  wire _09779_;
  wire _09780_;
  wire _09781_;
  wire _09782_;
  wire _09783_;
  wire _09784_;
  wire _09785_;
  wire _09786_;
  wire _09787_;
  wire _09788_;
  wire _09789_;
  wire _09790_;
  wire _09791_;
  wire _09792_;
  wire _09793_;
  wire _09794_;
  wire _09795_;
  wire _09796_;
  wire _09797_;
  wire _09798_;
  wire _09799_;
  wire _09800_;
  wire _09801_;
  wire _09802_;
  wire _09803_;
  wire _09804_;
  wire _09805_;
  wire _09806_;
  wire _09807_;
  wire _09808_;
  wire _09809_;
  wire _09810_;
  wire _09811_;
  wire _09812_;
  wire _09813_;
  wire _09814_;
  wire _09815_;
  wire _09816_;
  wire _09817_;
  wire _09818_;
  wire _09819_;
  wire _09820_;
  wire _09821_;
  wire _09822_;
  wire _09823_;
  wire _09824_;
  wire _09825_;
  wire _09826_;
  wire _09827_;
  wire _09828_;
  wire _09829_;
  wire _09830_;
  wire _09831_;
  wire _09832_;
  wire _09833_;
  wire _09834_;
  wire _09835_;
  wire _09836_;
  wire _09837_;
  wire _09838_;
  wire _09839_;
  wire _09840_;
  wire _09841_;
  wire _09842_;
  wire _09843_;
  wire _09844_;
  wire _09845_;
  wire _09846_;
  wire _09847_;
  wire _09848_;
  wire _09849_;
  wire _09850_;
  wire _09851_;
  wire _09852_;
  wire _09853_;
  wire _09854_;
  wire _09855_;
  wire _09856_;
  wire _09857_;
  wire _09858_;
  wire _09859_;
  wire _09860_;
  wire _09861_;
  wire _09862_;
  wire _09863_;
  wire _09864_;
  wire _09865_;
  wire _09866_;
  wire _09867_;
  wire _09868_;
  wire _09869_;
  wire _09870_;
  wire _09871_;
  wire _09872_;
  wire _09873_;
  wire _09874_;
  wire _09875_;
  wire _09876_;
  wire _09877_;
  wire _09878_;
  wire _09879_;
  wire _09880_;
  wire _09881_;
  wire _09882_;
  wire _09883_;
  wire _09884_;
  wire _09885_;
  wire _09886_;
  wire _09887_;
  wire _09888_;
  wire _09889_;
  wire _09890_;
  wire _09891_;
  wire _09892_;
  wire _09893_;
  wire _09894_;
  wire _09895_;
  wire _09896_;
  wire _09897_;
  wire _09898_;
  wire _09899_;
  wire _09900_;
  wire _09901_;
  wire _09902_;
  wire _09903_;
  wire _09904_;
  wire _09905_;
  wire _09906_;
  wire _09907_;
  wire _09908_;
  wire _09909_;
  wire _09910_;
  wire _09911_;
  wire _09912_;
  wire _09913_;
  wire _09914_;
  wire _09915_;
  wire _09916_;
  wire _09917_;
  wire _09918_;
  wire _09919_;
  wire _09920_;
  wire _09921_;
  wire _09922_;
  wire _09923_;
  wire _09924_;
  wire _09925_;
  wire _09926_;
  wire _09927_;
  wire _09928_;
  wire _09929_;
  wire _09930_;
  wire _09931_;
  wire _09932_;
  wire _09933_;
  wire _09934_;
  wire _09935_;
  wire _09936_;
  wire _09937_;
  wire _09938_;
  wire _09939_;
  wire _09940_;
  wire _09941_;
  wire _09942_;
  wire _09943_;
  wire _09944_;
  wire _09945_;
  wire _09946_;
  wire _09947_;
  wire _09948_;
  wire _09949_;
  wire _09950_;
  wire _09951_;
  wire _09952_;
  wire _09953_;
  wire _09954_;
  wire _09955_;
  wire _09956_;
  wire _09957_;
  wire _09958_;
  wire _09959_;
  wire _09960_;
  wire _09961_;
  wire _09962_;
  wire _09963_;
  wire _09964_;
  wire _09965_;
  wire _09966_;
  wire _09967_;
  wire _09968_;
  wire _09969_;
  wire _09970_;
  wire _09971_;
  wire _09972_;
  wire _09973_;
  wire _09974_;
  wire _09975_;
  wire _09976_;
  wire _09977_;
  wire _09978_;
  wire _09979_;
  wire _09980_;
  wire _09981_;
  wire _09982_;
  wire _09983_;
  wire _09984_;
  wire _09985_;
  wire _09986_;
  wire _09987_;
  wire _09988_;
  wire _09989_;
  wire _09990_;
  wire _09991_;
  wire _09992_;
  wire _09993_;
  wire _09994_;
  wire _09995_;
  wire _09996_;
  wire _09997_;
  wire _09998_;
  wire _09999_;
  wire _10000_;
  wire _10001_;
  wire _10002_;
  wire _10003_;
  wire _10004_;
  wire _10005_;
  wire _10006_;
  wire _10007_;
  wire _10008_;
  wire _10009_;
  wire _10010_;
  wire _10011_;
  wire _10012_;
  wire _10013_;
  wire _10014_;
  wire _10015_;
  wire _10016_;
  wire _10017_;
  wire _10018_;
  wire _10019_;
  wire _10020_;
  wire _10021_;
  wire _10022_;
  wire _10023_;
  wire _10024_;
  wire _10025_;
  wire _10026_;
  wire _10027_;
  wire _10028_;
  wire _10029_;
  wire _10030_;
  wire _10031_;
  wire _10032_;
  wire _10033_;
  wire _10034_;
  wire _10035_;
  wire _10036_;
  wire _10037_;
  wire _10038_;
  wire _10039_;
  wire _10040_;
  wire _10041_;
  wire _10042_;
  wire _10043_;
  wire _10044_;
  wire _10045_;
  wire _10046_;
  wire _10047_;
  wire _10048_;
  wire _10049_;
  wire _10050_;
  wire _10051_;
  wire _10052_;
  wire _10053_;
  wire _10054_;
  wire _10055_;
  wire _10056_;
  wire _10057_;
  wire _10058_;
  wire _10059_;
  wire _10060_;
  wire _10061_;
  wire _10062_;
  wire _10063_;
  wire _10064_;
  wire _10065_;
  wire _10066_;
  wire _10067_;
  wire _10068_;
  wire _10069_;
  wire _10070_;
  wire _10071_;
  wire _10072_;
  wire _10073_;
  wire _10074_;
  wire _10075_;
  wire _10076_;
  wire _10077_;
  wire _10078_;
  wire _10079_;
  wire _10080_;
  wire _10081_;
  wire _10082_;
  wire _10083_;
  wire _10084_;
  wire _10085_;
  wire _10086_;
  wire _10087_;
  wire _10088_;
  wire _10089_;
  wire _10090_;
  wire _10091_;
  wire _10092_;
  wire _10093_;
  wire _10094_;
  wire _10095_;
  wire _10096_;
  wire _10097_;
  wire _10098_;
  wire _10099_;
  wire _10100_;
  wire _10101_;
  wire _10102_;
  wire _10103_;
  wire _10104_;
  wire _10105_;
  wire _10106_;
  wire _10107_;
  wire _10108_;
  wire _10109_;
  wire _10110_;
  wire _10111_;
  wire _10112_;
  wire _10113_;
  wire _10114_;
  wire _10115_;
  wire _10116_;
  wire _10117_;
  wire _10118_;
  wire _10119_;
  wire _10120_;
  wire _10121_;
  wire _10122_;
  wire _10123_;
  wire _10124_;
  wire _10125_;
  wire _10126_;
  wire _10127_;
  wire _10128_;
  wire _10129_;
  wire _10130_;
  wire _10131_;
  wire _10132_;
  wire _10133_;
  wire _10134_;
  wire _10135_;
  wire _10136_;
  wire _10137_;
  wire _10138_;
  wire _10139_;
  wire _10140_;
  wire _10141_;
  wire _10142_;
  wire _10143_;
  wire _10144_;
  wire _10145_;
  wire _10146_;
  wire _10147_;
  wire _10148_;
  wire _10149_;
  wire _10150_;
  wire _10151_;
  wire _10152_;
  wire _10153_;
  wire _10154_;
  wire _10155_;
  wire _10156_;
  wire _10157_;
  wire _10158_;
  wire _10159_;
  wire _10160_;
  wire _10161_;
  wire _10162_;
  wire _10163_;
  wire _10164_;
  wire _10165_;
  wire _10166_;
  wire _10167_;
  wire _10168_;
  wire _10169_;
  wire _10170_;
  wire _10171_;
  wire _10172_;
  wire _10173_;
  wire _10174_;
  wire _10175_;
  wire _10176_;
  wire _10177_;
  wire _10178_;
  wire _10179_;
  wire _10180_;
  wire _10181_;
  wire _10182_;
  wire _10183_;
  wire _10184_;
  wire _10185_;
  wire _10186_;
  wire _10187_;
  wire _10188_;
  wire _10189_;
  wire _10190_;
  wire _10191_;
  wire _10192_;
  wire _10193_;
  wire _10194_;
  wire _10195_;
  wire _10196_;
  wire _10197_;
  wire _10198_;
  wire _10199_;
  wire _10200_;
  wire _10201_;
  wire _10202_;
  wire _10203_;
  wire _10204_;
  wire _10205_;
  wire _10206_;
  wire _10207_;
  wire _10208_;
  wire _10209_;
  wire _10210_;
  wire _10211_;
  wire _10212_;
  wire _10213_;
  wire _10214_;
  wire _10215_;
  wire _10216_;
  wire _10217_;
  wire _10218_;
  wire _10219_;
  wire _10220_;
  wire _10221_;
  wire _10222_;
  wire _10223_;
  wire _10224_;
  wire _10225_;
  wire _10226_;
  wire _10227_;
  wire _10228_;
  wire _10229_;
  wire _10230_;
  wire _10231_;
  wire _10232_;
  wire _10233_;
  wire _10234_;
  wire _10235_;
  wire _10236_;
  wire _10237_;
  wire _10238_;
  wire _10239_;
  wire _10240_;
  wire _10241_;
  wire _10242_;
  wire _10243_;
  wire _10244_;
  wire _10245_;
  wire _10246_;
  wire _10247_;
  wire _10248_;
  wire _10249_;
  wire _10250_;
  wire _10251_;
  wire _10252_;
  wire _10253_;
  wire _10254_;
  wire _10255_;
  wire _10256_;
  wire _10257_;
  wire _10258_;
  wire _10259_;
  wire _10260_;
  wire _10261_;
  wire _10262_;
  wire _10263_;
  wire _10264_;
  wire _10265_;
  wire _10266_;
  wire _10267_;
  wire _10268_;
  wire _10269_;
  wire _10270_;
  wire _10271_;
  wire _10272_;
  wire _10273_;
  wire _10274_;
  wire _10275_;
  wire _10276_;
  wire _10277_;
  wire _10278_;
  wire _10279_;
  wire _10280_;
  wire _10281_;
  wire _10282_;
  wire _10283_;
  wire _10284_;
  wire _10285_;
  wire _10286_;
  wire _10287_;
  wire _10288_;
  wire _10289_;
  wire _10290_;
  wire _10291_;
  wire _10292_;
  wire _10293_;
  wire _10294_;
  wire _10295_;
  wire _10296_;
  wire _10297_;
  wire _10298_;
  wire _10299_;
  wire _10300_;
  wire _10301_;
  wire _10302_;
  wire _10303_;
  wire _10304_;
  wire _10305_;
  wire _10306_;
  wire _10307_;
  wire _10308_;
  wire _10309_;
  wire _10310_;
  wire _10311_;
  wire _10312_;
  wire _10313_;
  wire _10314_;
  wire _10315_;
  wire _10316_;
  wire _10317_;
  wire _10318_;
  wire _10319_;
  wire _10320_;
  wire _10321_;
  wire _10322_;
  wire _10323_;
  wire _10324_;
  wire _10325_;
  wire _10326_;
  wire _10327_;
  wire _10328_;
  wire _10329_;
  wire _10330_;
  wire _10331_;
  wire _10332_;
  wire _10333_;
  wire _10334_;
  wire _10335_;
  wire _10336_;
  wire _10337_;
  wire _10338_;
  wire _10339_;
  wire _10340_;
  wire _10341_;
  wire _10342_;
  wire _10343_;
  wire _10344_;
  wire _10345_;
  wire _10346_;
  wire _10347_;
  wire _10348_;
  wire _10349_;
  wire _10350_;
  wire _10351_;
  wire _10352_;
  wire _10353_;
  wire _10354_;
  wire _10355_;
  wire _10356_;
  wire _10357_;
  wire _10358_;
  wire _10359_;
  wire _10360_;
  wire _10361_;
  wire _10362_;
  wire _10363_;
  wire _10364_;
  wire _10365_;
  wire _10366_;
  wire _10367_;
  wire _10368_;
  wire _10369_;
  wire _10370_;
  wire _10371_;
  wire _10372_;
  wire _10373_;
  wire _10374_;
  wire _10375_;
  wire _10376_;
  wire _10377_;
  wire _10378_;
  wire _10379_;
  wire _10380_;
  wire _10381_;
  wire _10382_;
  wire _10383_;
  wire _10384_;
  wire _10385_;
  wire _10386_;
  wire _10387_;
  wire _10388_;
  wire _10389_;
  wire _10390_;
  wire _10391_;
  wire _10392_;
  wire _10393_;
  wire _10394_;
  wire _10395_;
  wire _10396_;
  wire _10397_;
  wire _10398_;
  wire _10399_;
  wire _10400_;
  wire _10401_;
  wire _10402_;
  wire _10403_;
  wire _10404_;
  wire _10405_;
  wire _10406_;
  wire _10407_;
  wire _10408_;
  wire _10409_;
  wire _10410_;
  wire _10411_;
  wire _10412_;
  wire _10413_;
  wire _10414_;
  wire _10415_;
  wire _10416_;
  wire _10417_;
  wire _10418_;
  wire _10419_;
  wire _10420_;
  wire _10421_;
  wire _10422_;
  wire _10423_;
  wire _10424_;
  wire _10425_;
  wire _10426_;
  wire _10427_;
  wire _10428_;
  wire _10429_;
  wire _10430_;
  wire _10431_;
  wire _10432_;
  wire _10433_;
  wire _10434_;
  wire _10435_;
  wire _10436_;
  wire _10437_;
  wire _10438_;
  wire _10439_;
  wire _10440_;
  wire _10441_;
  wire _10442_;
  wire _10443_;
  wire _10444_;
  wire _10445_;
  wire _10446_;
  wire _10447_;
  wire _10448_;
  wire _10449_;
  wire _10450_;
  wire _10451_;
  wire _10452_;
  wire _10453_;
  wire _10454_;
  wire _10455_;
  wire _10456_;
  wire _10457_;
  wire _10458_;
  wire _10459_;
  wire _10460_;
  wire _10461_;
  wire _10462_;
  wire _10463_;
  wire _10464_;
  wire _10465_;
  wire _10466_;
  wire _10467_;
  wire _10468_;
  wire _10469_;
  wire _10470_;
  wire _10471_;
  wire _10472_;
  wire _10473_;
  wire _10474_;
  wire _10475_;
  wire _10476_;
  wire _10477_;
  wire _10478_;
  wire _10479_;
  wire _10480_;
  wire _10481_;
  wire _10482_;
  wire _10483_;
  wire _10484_;
  wire _10485_;
  wire _10486_;
  wire _10487_;
  wire _10488_;
  wire _10489_;
  wire _10490_;
  wire _10491_;
  wire _10492_;
  wire _10493_;
  wire _10494_;
  wire _10495_;
  wire _10496_;
  wire _10497_;
  wire _10498_;
  wire _10499_;
  wire _10500_;
  wire _10501_;
  wire _10502_;
  wire _10503_;
  wire _10504_;
  wire _10505_;
  wire _10506_;
  wire _10507_;
  wire _10508_;
  wire _10509_;
  wire _10510_;
  wire _10511_;
  wire _10512_;
  wire _10513_;
  wire _10514_;
  wire _10515_;
  wire _10516_;
  wire _10517_;
  wire _10518_;
  wire _10519_;
  wire _10520_;
  wire _10521_;
  wire _10522_;
  wire _10523_;
  wire _10524_;
  wire _10525_;
  wire _10526_;
  wire _10527_;
  wire _10528_;
  wire _10529_;
  wire _10530_;
  wire _10531_;
  wire _10532_;
  wire _10533_;
  wire _10534_;
  wire _10535_;
  wire _10536_;
  wire _10537_;
  wire _10538_;
  wire _10539_;
  wire _10540_;
  wire _10541_;
  wire _10542_;
  wire _10543_;
  wire _10544_;
  wire _10545_;
  wire _10546_;
  wire _10547_;
  wire _10548_;
  wire _10549_;
  wire _10550_;
  wire _10551_;
  wire _10552_;
  wire _10553_;
  wire _10554_;
  wire _10555_;
  wire _10556_;
  wire _10557_;
  wire _10558_;
  wire _10559_;
  wire _10560_;
  wire _10561_;
  wire _10562_;
  wire _10563_;
  wire _10564_;
  wire _10565_;
  wire _10566_;
  wire _10567_;
  wire _10568_;
  wire _10569_;
  wire _10570_;
  wire _10571_;
  wire _10572_;
  wire _10573_;
  wire _10574_;
  wire _10575_;
  wire _10576_;
  wire _10577_;
  wire _10578_;
  wire _10579_;
  wire _10580_;
  wire _10581_;
  wire _10582_;
  wire _10583_;
  wire _10584_;
  wire _10585_;
  wire _10586_;
  wire _10587_;
  wire _10588_;
  wire _10589_;
  wire _10590_;
  wire _10591_;
  wire _10592_;
  wire _10593_;
  wire _10594_;
  wire _10595_;
  wire _10596_;
  wire _10597_;
  wire _10598_;
  wire _10599_;
  wire _10600_;
  wire _10601_;
  wire _10602_;
  wire _10603_;
  wire _10604_;
  wire _10605_;
  wire _10606_;
  wire _10607_;
  wire _10608_;
  wire _10609_;
  wire _10610_;
  wire _10611_;
  wire _10612_;
  wire _10613_;
  wire _10614_;
  wire _10615_;
  wire _10616_;
  wire _10617_;
  wire _10618_;
  wire _10619_;
  wire _10620_;
  wire _10621_;
  wire _10622_;
  wire _10623_;
  wire _10624_;
  wire _10625_;
  wire _10626_;
  wire _10627_;
  wire _10628_;
  wire _10629_;
  wire _10630_;
  wire _10631_;
  wire _10632_;
  wire _10633_;
  wire _10634_;
  wire _10635_;
  wire _10636_;
  wire _10637_;
  wire _10638_;
  wire _10639_;
  wire _10640_;
  wire _10641_;
  wire _10642_;
  wire _10643_;
  wire _10644_;
  wire _10645_;
  wire _10646_;
  wire _10647_;
  wire _10648_;
  wire _10649_;
  wire _10650_;
  wire _10651_;
  wire _10652_;
  wire _10653_;
  wire _10654_;
  wire _10655_;
  wire _10656_;
  wire _10657_;
  wire _10658_;
  wire _10659_;
  wire _10660_;
  wire _10661_;
  wire _10662_;
  wire _10663_;
  wire _10664_;
  wire _10665_;
  wire _10666_;
  wire _10667_;
  wire _10668_;
  wire _10669_;
  wire _10670_;
  wire _10671_;
  wire _10672_;
  wire _10673_;
  wire _10674_;
  wire _10675_;
  wire _10676_;
  wire _10677_;
  wire _10678_;
  wire _10679_;
  wire _10680_;
  wire _10681_;
  wire _10682_;
  wire _10683_;
  wire _10684_;
  wire _10685_;
  wire _10686_;
  wire _10687_;
  wire _10688_;
  wire _10689_;
  wire _10690_;
  wire _10691_;
  wire _10692_;
  wire _10693_;
  wire _10694_;
  wire _10695_;
  wire _10696_;
  wire _10697_;
  wire _10698_;
  wire _10699_;
  wire _10700_;
  wire _10701_;
  wire _10702_;
  wire _10703_;
  wire _10704_;
  wire _10705_;
  wire _10706_;
  wire _10707_;
  wire _10708_;
  wire _10709_;
  wire _10710_;
  wire _10711_;
  wire _10712_;
  wire _10713_;
  wire _10714_;
  wire _10715_;
  wire _10716_;
  wire _10717_;
  wire _10718_;
  wire _10719_;
  wire _10720_;
  wire _10721_;
  wire _10722_;
  wire _10723_;
  wire _10724_;
  wire _10725_;
  wire _10726_;
  wire _10727_;
  wire _10728_;
  wire _10729_;
  wire _10730_;
  wire _10731_;
  wire _10732_;
  wire _10733_;
  wire _10734_;
  wire _10735_;
  wire _10736_;
  wire _10737_;
  wire _10738_;
  wire _10739_;
  wire _10740_;
  wire _10741_;
  wire _10742_;
  wire _10743_;
  wire _10744_;
  wire _10745_;
  wire _10746_;
  wire _10747_;
  wire _10748_;
  wire _10749_;
  wire _10750_;
  wire _10751_;
  wire _10752_;
  wire _10753_;
  wire _10754_;
  wire _10755_;
  wire _10756_;
  wire _10757_;
  wire _10758_;
  wire _10759_;
  wire _10760_;
  wire _10761_;
  wire _10762_;
  wire _10763_;
  wire _10764_;
  wire _10765_;
  wire _10766_;
  wire _10767_;
  wire _10768_;
  wire _10769_;
  wire _10770_;
  wire _10771_;
  wire _10772_;
  wire _10773_;
  wire _10774_;
  wire _10775_;
  wire _10776_;
  wire _10777_;
  wire _10778_;
  wire _10779_;
  wire _10780_;
  wire _10781_;
  wire _10782_;
  wire _10783_;
  wire _10784_;
  wire _10785_;
  wire _10786_;
  wire _10787_;
  wire _10788_;
  wire _10789_;
  wire _10790_;
  wire _10791_;
  wire _10792_;
  wire _10793_;
  wire _10794_;
  wire _10795_;
  wire _10796_;
  wire _10797_;
  wire _10798_;
  wire _10799_;
  wire _10800_;
  wire _10801_;
  wire _10802_;
  wire _10803_;
  wire _10804_;
  wire _10805_;
  wire _10806_;
  wire _10807_;
  wire _10808_;
  wire _10809_;
  wire _10810_;
  wire _10811_;
  wire _10812_;
  wire _10813_;
  wire _10814_;
  wire _10815_;
  wire _10816_;
  wire _10817_;
  wire _10818_;
  wire _10819_;
  wire _10820_;
  wire _10821_;
  wire _10822_;
  wire _10823_;
  wire _10824_;
  wire _10825_;
  wire _10826_;
  wire _10827_;
  wire _10828_;
  wire _10829_;
  wire _10830_;
  wire _10831_;
  wire _10832_;
  wire _10833_;
  wire _10834_;
  wire _10835_;
  wire _10836_;
  wire _10837_;
  wire _10838_;
  wire _10839_;
  wire _10840_;
  wire _10841_;
  wire _10842_;
  wire _10843_;
  wire _10844_;
  wire _10845_;
  wire _10846_;
  wire _10847_;
  wire _10848_;
  wire _10849_;
  wire _10850_;
  wire _10851_;
  wire _10852_;
  wire _10853_;
  wire _10854_;
  wire _10855_;
  wire _10856_;
  wire _10857_;
  wire _10858_;
  wire _10859_;
  wire _10860_;
  wire _10861_;
  wire _10862_;
  wire _10863_;
  wire _10864_;
  wire _10865_;
  wire _10866_;
  wire _10867_;
  wire _10868_;
  wire _10869_;
  wire _10870_;
  wire _10871_;
  wire _10872_;
  wire _10873_;
  wire _10874_;
  wire _10875_;
  wire _10876_;
  wire _10877_;
  wire _10878_;
  wire _10879_;
  wire _10880_;
  wire _10881_;
  wire _10882_;
  wire _10883_;
  wire _10884_;
  wire _10885_;
  wire _10886_;
  wire _10887_;
  wire _10888_;
  wire _10889_;
  wire _10890_;
  wire _10891_;
  wire _10892_;
  wire _10893_;
  wire _10894_;
  wire _10895_;
  wire _10896_;
  wire _10897_;
  wire _10898_;
  wire _10899_;
  wire _10900_;
  wire _10901_;
  wire _10902_;
  wire _10903_;
  wire _10904_;
  wire _10905_;
  wire _10906_;
  wire _10907_;
  wire _10908_;
  wire _10909_;
  wire _10910_;
  wire _10911_;
  wire _10912_;
  wire _10913_;
  wire _10914_;
  wire _10915_;
  wire _10916_;
  wire _10917_;
  wire _10918_;
  wire _10919_;
  wire _10920_;
  wire _10921_;
  wire _10922_;
  wire _10923_;
  wire _10924_;
  wire _10925_;
  wire _10926_;
  wire _10927_;
  wire _10928_;
  wire _10929_;
  wire _10930_;
  wire _10931_;
  wire _10932_;
  wire _10933_;
  wire _10934_;
  wire _10935_;
  wire _10936_;
  wire _10937_;
  wire _10938_;
  wire _10939_;
  wire _10940_;
  wire _10941_;
  wire _10942_;
  wire _10943_;
  wire _10944_;
  wire _10945_;
  wire _10946_;
  wire _10947_;
  wire _10948_;
  wire _10949_;
  wire _10950_;
  wire _10951_;
  wire _10952_;
  wire _10953_;
  wire _10954_;
  wire _10955_;
  wire _10956_;
  wire _10957_;
  wire _10958_;
  wire _10959_;
  wire _10960_;
  wire _10961_;
  wire _10962_;
  wire _10963_;
  wire _10964_;
  wire _10965_;
  wire _10966_;
  wire _10967_;
  wire _10968_;
  wire _10969_;
  wire _10970_;
  wire _10971_;
  wire _10972_;
  wire _10973_;
  wire _10974_;
  wire _10975_;
  wire _10976_;
  wire _10977_;
  wire _10978_;
  wire _10979_;
  wire _10980_;
  wire _10981_;
  wire _10982_;
  wire _10983_;
  wire _10984_;
  wire _10985_;
  wire _10986_;
  wire _10987_;
  wire _10988_;
  wire _10989_;
  wire _10990_;
  wire _10991_;
  wire _10992_;
  wire _10993_;
  wire _10994_;
  wire _10995_;
  wire _10996_;
  wire _10997_;
  wire _10998_;
  wire _10999_;
  wire _11000_;
  wire _11001_;
  wire _11002_;
  wire _11003_;
  wire _11004_;
  wire _11005_;
  wire _11006_;
  wire _11007_;
  wire _11008_;
  wire _11009_;
  wire _11010_;
  wire _11011_;
  wire _11012_;
  wire _11013_;
  wire _11014_;
  wire _11015_;
  wire _11016_;
  wire _11017_;
  wire _11018_;
  wire _11019_;
  wire _11020_;
  wire _11021_;
  wire _11022_;
  wire _11023_;
  wire _11024_;
  wire _11025_;
  wire _11026_;
  wire _11027_;
  wire _11028_;
  wire _11029_;
  wire _11030_;
  wire _11031_;
  wire _11032_;
  wire _11033_;
  wire _11034_;
  wire _11035_;
  wire _11036_;
  wire _11037_;
  wire _11038_;
  wire _11039_;
  wire _11040_;
  wire _11041_;
  wire _11042_;
  wire _11043_;
  wire _11044_;
  wire _11045_;
  wire _11046_;
  wire _11047_;
  wire _11048_;
  wire _11049_;
  wire _11050_;
  wire _11051_;
  wire _11052_;
  wire _11053_;
  wire _11054_;
  wire _11055_;
  wire _11056_;
  wire _11057_;
  wire _11058_;
  wire _11059_;
  wire _11060_;
  wire _11061_;
  wire _11062_;
  wire _11063_;
  wire _11064_;
  wire _11065_;
  wire _11066_;
  wire _11067_;
  wire _11068_;
  wire _11069_;
  wire _11070_;
  wire _11071_;
  wire _11072_;
  wire _11073_;
  wire _11074_;
  wire _11075_;
  wire _11076_;
  wire _11077_;
  wire _11078_;
  wire _11079_;
  wire _11080_;
  wire _11081_;
  wire _11082_;
  wire _11083_;
  wire _11084_;
  wire _11085_;
  wire _11086_;
  wire _11087_;
  wire _11088_;
  wire _11089_;
  wire _11090_;
  wire _11091_;
  wire _11092_;
  wire _11093_;
  wire _11094_;
  wire _11095_;
  wire _11096_;
  wire _11097_;
  wire _11098_;
  wire _11099_;
  wire _11100_;
  wire _11101_;
  wire _11102_;
  wire _11103_;
  wire _11104_;
  wire _11105_;
  wire _11106_;
  wire _11107_;
  wire _11108_;
  wire _11109_;
  wire _11110_;
  wire _11111_;
  wire _11112_;
  wire _11113_;
  wire _11114_;
  wire _11115_;
  wire _11116_;
  wire _11117_;
  wire _11118_;
  wire _11119_;
  wire _11120_;
  wire _11121_;
  wire _11122_;
  wire _11123_;
  wire _11124_;
  wire _11125_;
  wire _11126_;
  wire _11127_;
  wire _11128_;
  wire _11129_;
  wire _11130_;
  wire _11131_;
  wire _11132_;
  wire _11133_;
  wire _11134_;
  wire _11135_;
  wire _11136_;
  wire _11137_;
  wire _11138_;
  wire _11139_;
  wire _11140_;
  wire _11141_;
  wire _11142_;
  wire _11143_;
  wire _11144_;
  wire _11145_;
  wire _11146_;
  wire _11147_;
  wire _11148_;
  wire _11149_;
  wire _11150_;
  wire _11151_;
  wire _11152_;
  wire _11153_;
  wire _11154_;
  wire _11155_;
  wire _11156_;
  wire _11157_;
  wire _11158_;
  wire _11159_;
  wire _11160_;
  wire _11161_;
  wire _11162_;
  wire _11163_;
  wire _11164_;
  wire _11165_;
  wire _11166_;
  wire _11167_;
  wire _11168_;
  wire _11169_;
  wire _11170_;
  wire _11171_;
  wire _11172_;
  wire _11173_;
  wire _11174_;
  wire _11175_;
  wire _11176_;
  wire _11177_;
  wire _11178_;
  wire _11179_;
  wire _11180_;
  wire _11181_;
  wire _11182_;
  wire _11183_;
  wire _11184_;
  wire _11185_;
  wire _11186_;
  wire _11187_;
  wire _11188_;
  wire _11189_;
  wire _11190_;
  wire _11191_;
  wire _11192_;
  wire _11193_;
  wire _11194_;
  wire _11195_;
  wire _11196_;
  wire _11197_;
  wire _11198_;
  wire _11199_;
  wire _11200_;
  wire _11201_;
  wire _11202_;
  wire _11203_;
  wire _11204_;
  wire _11205_;
  wire _11206_;
  wire _11207_;
  wire _11208_;
  wire _11209_;
  wire _11210_;
  wire _11211_;
  wire _11212_;
  wire _11213_;
  wire _11214_;
  wire _11215_;
  wire _11216_;
  wire _11217_;
  wire _11218_;
  wire _11219_;
  wire _11220_;
  wire _11221_;
  wire _11222_;
  wire _11223_;
  wire _11224_;
  wire _11225_;
  wire _11226_;
  wire _11227_;
  wire _11228_;
  wire _11229_;
  wire _11230_;
  wire _11231_;
  wire _11232_;
  wire _11233_;
  wire _11234_;
  wire _11235_;
  wire _11236_;
  wire _11237_;
  wire _11238_;
  wire _11239_;
  wire _11240_;
  wire _11241_;
  wire _11242_;
  wire _11243_;
  wire _11244_;
  wire _11245_;
  wire _11246_;
  wire _11247_;
  wire _11248_;
  wire _11249_;
  wire _11250_;
  wire _11251_;
  wire _11252_;
  wire _11253_;
  wire _11254_;
  wire _11255_;
  wire _11256_;
  wire _11257_;
  wire _11258_;
  wire _11259_;
  wire _11260_;
  wire _11261_;
  wire _11262_;
  wire _11263_;
  wire _11264_;
  wire _11265_;
  wire _11266_;
  wire _11267_;
  wire _11268_;
  wire _11269_;
  wire _11270_;
  wire _11271_;
  wire _11272_;
  wire _11273_;
  wire _11274_;
  wire _11275_;
  wire _11276_;
  wire _11277_;
  wire _11278_;
  wire _11279_;
  wire _11280_;
  wire _11281_;
  wire _11282_;
  wire _11283_;
  wire _11284_;
  wire _11285_;
  wire _11286_;
  wire _11287_;
  wire _11288_;
  wire _11289_;
  wire _11290_;
  wire _11291_;
  wire _11292_;
  wire _11293_;
  wire _11294_;
  wire _11295_;
  wire _11296_;
  wire _11297_;
  wire _11298_;
  wire _11299_;
  wire _11300_;
  wire _11301_;
  wire _11302_;
  wire _11303_;
  wire _11304_;
  wire _11305_;
  wire _11306_;
  wire _11307_;
  wire _11308_;
  wire _11309_;
  wire _11310_;
  wire _11311_;
  wire _11312_;
  wire _11313_;
  wire _11314_;
  wire _11315_;
  wire _11316_;
  wire _11317_;
  wire _11318_;
  wire _11319_;
  wire _11320_;
  wire _11321_;
  wire _11322_;
  wire _11323_;
  wire _11324_;
  wire _11325_;
  wire _11326_;
  wire _11327_;
  wire _11328_;
  wire _11329_;
  wire _11330_;
  wire _11331_;
  wire _11332_;
  wire _11333_;
  wire _11334_;
  wire _11335_;
  wire _11336_;
  wire _11337_;
  wire _11338_;
  wire _11339_;
  wire _11340_;
  wire _11341_;
  wire _11342_;
  wire _11343_;
  wire _11344_;
  wire _11345_;
  wire _11346_;
  wire _11347_;
  wire _11348_;
  wire _11349_;
  wire _11350_;
  wire _11351_;
  wire _11352_;
  wire _11353_;
  wire _11354_;
  wire _11355_;
  wire _11356_;
  wire _11357_;
  wire _11358_;
  wire _11359_;
  wire _11360_;
  wire _11361_;
  wire _11362_;
  wire _11363_;
  wire _11364_;
  wire _11365_;
  wire _11366_;
  wire _11367_;
  wire _11368_;
  wire _11369_;
  wire _11370_;
  wire _11371_;
  wire _11372_;
  wire _11373_;
  wire _11374_;
  wire _11375_;
  wire _11376_;
  wire _11377_;
  wire _11378_;
  wire _11379_;
  wire _11380_;
  wire _11381_;
  wire _11382_;
  wire _11383_;
  wire _11384_;
  wire _11385_;
  wire _11386_;
  wire _11387_;
  wire _11388_;
  wire _11389_;
  wire _11390_;
  wire _11391_;
  wire _11392_;
  wire _11393_;
  wire _11394_;
  wire _11395_;
  wire _11396_;
  wire _11397_;
  wire _11398_;
  wire _11399_;
  wire _11400_;
  wire _11401_;
  wire _11402_;
  wire _11403_;
  wire _11404_;
  wire _11405_;
  wire _11406_;
  wire _11407_;
  wire _11408_;
  wire _11409_;
  wire _11410_;
  wire _11411_;
  wire _11412_;
  wire _11413_;
  wire _11414_;
  wire _11415_;
  wire _11416_;
  wire _11417_;
  wire _11418_;
  wire _11419_;
  wire _11420_;
  wire _11421_;
  wire _11422_;
  wire _11423_;
  wire _11424_;
  wire _11425_;
  wire _11426_;
  wire _11427_;
  wire _11428_;
  wire _11429_;
  wire _11430_;
  wire _11431_;
  wire _11432_;
  wire _11433_;
  wire _11434_;
  wire _11435_;
  wire _11436_;
  wire _11437_;
  wire _11438_;
  wire _11439_;
  wire _11440_;
  wire _11441_;
  wire _11442_;
  wire _11443_;
  wire _11444_;
  wire _11445_;
  wire _11446_;
  wire _11447_;
  wire _11448_;
  wire _11449_;
  wire _11450_;
  wire _11451_;
  wire _11452_;
  wire _11453_;
  wire _11454_;
  wire _11455_;
  wire _11456_;
  wire _11457_;
  wire _11458_;
  wire _11459_;
  wire _11460_;
  wire _11461_;
  wire _11462_;
  wire _11463_;
  wire _11464_;
  wire _11465_;
  wire _11466_;
  wire _11467_;
  wire _11468_;
  wire _11469_;
  wire _11470_;
  wire _11471_;
  wire _11472_;
  wire _11473_;
  wire _11474_;
  wire _11475_;
  wire _11476_;
  wire _11477_;
  wire _11478_;
  wire _11479_;
  wire _11480_;
  wire _11481_;
  wire _11482_;
  wire _11483_;
  wire _11484_;
  wire _11485_;
  wire _11486_;
  wire _11487_;
  wire _11488_;
  wire _11489_;
  wire _11490_;
  wire _11491_;
  wire _11492_;
  wire _11493_;
  wire _11494_;
  wire _11495_;
  wire _11496_;
  wire _11497_;
  wire _11498_;
  wire _11499_;
  wire _11500_;
  wire _11501_;
  wire _11502_;
  wire _11503_;
  wire _11504_;
  wire _11505_;
  wire _11506_;
  wire _11507_;
  wire _11508_;
  wire _11509_;
  wire _11510_;
  wire _11511_;
  wire _11512_;
  wire _11513_;
  wire _11514_;
  wire _11515_;
  wire _11516_;
  wire _11517_;
  wire _11518_;
  wire _11519_;
  wire _11520_;
  wire _11521_;
  wire _11522_;
  wire _11523_;
  wire _11524_;
  wire _11525_;
  wire _11526_;
  wire _11527_;
  wire _11528_;
  wire _11529_;
  wire _11530_;
  wire _11531_;
  wire _11532_;
  wire _11533_;
  wire _11534_;
  wire _11535_;
  wire _11536_;
  wire _11537_;
  wire _11538_;
  wire _11539_;
  wire _11540_;
  wire _11541_;
  wire _11542_;
  wire _11543_;
  wire _11544_;
  wire _11545_;
  wire _11546_;
  wire _11547_;
  wire _11548_;
  wire _11549_;
  wire _11550_;
  wire _11551_;
  wire _11552_;
  wire _11553_;
  wire _11554_;
  wire _11555_;
  wire _11556_;
  wire _11557_;
  wire _11558_;
  wire _11559_;
  wire _11560_;
  wire _11561_;
  wire _11562_;
  wire _11563_;
  wire _11564_;
  wire _11565_;
  wire _11566_;
  wire _11567_;
  wire _11568_;
  wire _11569_;
  wire _11570_;
  wire _11571_;
  wire _11572_;
  wire _11573_;
  wire _11574_;
  wire _11575_;
  wire _11576_;
  wire _11577_;
  wire _11578_;
  wire _11579_;
  wire _11580_;
  wire _11581_;
  wire _11582_;
  wire _11583_;
  wire _11584_;
  wire _11585_;
  wire _11586_;
  wire _11587_;
  wire _11588_;
  wire _11589_;
  wire _11590_;
  wire _11591_;
  wire _11592_;
  wire _11593_;
  wire _11594_;
  wire _11595_;
  wire _11596_;
  wire _11597_;
  wire _11598_;
  wire _11599_;
  wire _11600_;
  wire _11601_;
  wire _11602_;
  wire _11603_;
  wire _11604_;
  wire _11605_;
  wire _11606_;
  wire _11607_;
  wire _11608_;
  wire _11609_;
  wire _11610_;
  wire _11611_;
  wire _11612_;
  wire _11613_;
  wire _11614_;
  wire _11615_;
  wire _11616_;
  wire _11617_;
  wire _11618_;
  wire _11619_;
  wire _11620_;
  wire _11621_;
  wire _11622_;
  wire _11623_;
  wire _11624_;
  wire _11625_;
  wire _11626_;
  wire _11627_;
  wire _11628_;
  wire _11629_;
  wire _11630_;
  wire _11631_;
  wire _11632_;
  wire _11633_;
  wire _11634_;
  wire _11635_;
  wire _11636_;
  wire _11637_;
  wire _11638_;
  wire _11639_;
  wire _11640_;
  wire _11641_;
  wire _11642_;
  wire _11643_;
  wire _11644_;
  wire _11645_;
  wire _11646_;
  wire _11647_;
  wire _11648_;
  wire _11649_;
  wire _11650_;
  wire _11651_;
  wire _11652_;
  wire _11653_;
  wire _11654_;
  wire _11655_;
  wire _11656_;
  wire _11657_;
  wire _11658_;
  wire _11659_;
  wire _11660_;
  wire _11661_;
  wire _11662_;
  wire _11663_;
  wire _11664_;
  wire _11665_;
  wire _11666_;
  wire _11667_;
  wire _11668_;
  wire _11669_;
  wire _11670_;
  wire _11671_;
  wire _11672_;
  wire _11673_;
  wire _11674_;
  wire _11675_;
  wire _11676_;
  wire _11677_;
  wire _11678_;
  wire _11679_;
  wire _11680_;
  wire _11681_;
  wire _11682_;
  wire _11683_;
  wire _11684_;
  wire _11685_;
  wire _11686_;
  wire _11687_;
  wire _11688_;
  wire _11689_;
  wire _11690_;
  wire _11691_;
  wire _11692_;
  wire _11693_;
  wire _11694_;
  wire _11695_;
  wire _11696_;
  wire _11697_;
  wire _11698_;
  wire _11699_;
  wire _11700_;
  wire _11701_;
  wire _11702_;
  wire _11703_;
  wire _11704_;
  wire _11705_;
  wire _11706_;
  wire _11707_;
  wire _11708_;
  wire _11709_;
  wire _11710_;
  wire _11711_;
  wire _11712_;
  wire _11713_;
  wire _11714_;
  wire _11715_;
  wire _11716_;
  wire _11717_;
  wire _11718_;
  wire _11719_;
  wire _11720_;
  wire _11721_;
  wire _11722_;
  wire _11723_;
  wire _11724_;
  wire _11725_;
  wire _11726_;
  wire _11727_;
  wire _11728_;
  wire _11729_;
  wire _11730_;
  wire _11731_;
  wire _11732_;
  wire _11733_;
  wire _11734_;
  wire _11735_;
  wire _11736_;
  wire _11737_;
  wire _11738_;
  wire _11739_;
  wire _11740_;
  wire _11741_;
  wire _11742_;
  wire _11743_;
  wire _11744_;
  wire _11745_;
  wire _11746_;
  wire _11747_;
  wire _11748_;
  wire _11749_;
  wire _11750_;
  wire _11751_;
  wire _11752_;
  wire _11753_;
  wire _11754_;
  wire _11755_;
  wire _11756_;
  wire _11757_;
  wire _11758_;
  wire _11759_;
  wire _11760_;
  wire _11761_;
  wire _11762_;
  wire _11763_;
  wire _11764_;
  wire _11765_;
  wire _11766_;
  wire _11767_;
  wire _11768_;
  wire _11769_;
  wire _11770_;
  wire _11771_;
  wire _11772_;
  wire _11773_;
  wire _11774_;
  wire _11775_;
  wire _11776_;
  wire _11777_;
  wire _11778_;
  wire _11779_;
  wire _11780_;
  wire _11781_;
  wire _11782_;
  wire _11783_;
  wire _11784_;
  wire _11785_;
  wire _11786_;
  wire _11787_;
  wire _11788_;
  wire _11789_;
  wire _11790_;
  wire _11791_;
  wire _11792_;
  wire _11793_;
  wire _11794_;
  wire _11795_;
  wire _11796_;
  wire _11797_;
  wire _11798_;
  wire _11799_;
  wire _11800_;
  wire _11801_;
  wire _11802_;
  wire _11803_;
  wire _11804_;
  wire _11805_;
  wire _11806_;
  wire _11807_;
  wire _11808_;
  wire _11809_;
  wire _11810_;
  wire _11811_;
  wire _11812_;
  wire _11813_;
  wire _11814_;
  wire _11815_;
  wire _11816_;
  wire _11817_;
  wire _11818_;
  wire _11819_;
  wire _11820_;
  wire _11821_;
  wire _11822_;
  wire _11823_;
  wire _11824_;
  wire _11825_;
  wire _11826_;
  wire _11827_;
  wire _11828_;
  wire _11829_;
  wire _11830_;
  wire _11831_;
  wire _11832_;
  wire _11833_;
  wire _11834_;
  wire _11835_;
  wire _11836_;
  wire _11837_;
  wire _11838_;
  wire _11839_;
  wire _11840_;
  wire _11841_;
  wire _11842_;
  wire _11843_;
  wire _11844_;
  wire _11845_;
  wire _11846_;
  wire _11847_;
  wire _11848_;
  wire _11849_;
  wire _11850_;
  wire _11851_;
  wire _11852_;
  wire _11853_;
  wire _11854_;
  wire _11855_;
  wire _11856_;
  wire _11857_;
  wire _11858_;
  wire _11859_;
  wire _11860_;
  wire _11861_;
  wire _11862_;
  wire _11863_;
  wire _11864_;
  wire _11865_;
  wire _11866_;
  wire _11867_;
  wire _11868_;
  wire _11869_;
  wire _11870_;
  wire _11871_;
  wire _11872_;
  wire _11873_;
  wire _11874_;
  wire _11875_;
  wire _11876_;
  wire _11877_;
  wire _11878_;
  wire _11879_;
  wire _11880_;
  wire _11881_;
  wire _11882_;
  wire _11883_;
  wire _11884_;
  wire _11885_;
  wire _11886_;
  wire _11887_;
  wire _11888_;
  wire _11889_;
  wire _11890_;
  wire _11891_;
  wire _11892_;
  wire _11893_;
  wire _11894_;
  wire _11895_;
  wire _11896_;
  wire _11897_;
  wire _11898_;
  wire _11899_;
  wire _11900_;
  wire _11901_;
  wire _11902_;
  wire _11903_;
  wire _11904_;
  wire _11905_;
  wire _11906_;
  wire _11907_;
  wire _11908_;
  wire _11909_;
  wire _11910_;
  wire _11911_;
  wire _11912_;
  wire _11913_;
  wire _11914_;
  wire _11915_;
  wire _11916_;
  wire _11917_;
  wire _11918_;
  wire _11919_;
  wire _11920_;
  wire _11921_;
  wire _11922_;
  wire _11923_;
  wire _11924_;
  wire _11925_;
  wire _11926_;
  wire _11927_;
  wire _11928_;
  wire _11929_;
  wire _11930_;
  wire _11931_;
  wire _11932_;
  wire _11933_;
  wire _11934_;
  wire _11935_;
  wire _11936_;
  wire _11937_;
  wire _11938_;
  wire _11939_;
  wire _11940_;
  wire _11941_;
  wire _11942_;
  wire _11943_;
  wire _11944_;
  wire _11945_;
  wire _11946_;
  wire _11947_;
  wire _11948_;
  wire _11949_;
  wire _11950_;
  wire _11951_;
  wire _11952_;
  wire _11953_;
  wire _11954_;
  wire _11955_;
  wire _11956_;
  wire _11957_;
  wire _11958_;
  wire _11959_;
  wire _11960_;
  wire _11961_;
  wire _11962_;
  wire _11963_;
  wire _11964_;
  wire _11965_;
  wire _11966_;
  wire _11967_;
  wire _11968_;
  wire _11969_;
  wire _11970_;
  wire _11971_;
  wire _11972_;
  wire _11973_;
  wire _11974_;
  wire _11975_;
  wire _11976_;
  wire _11977_;
  wire _11978_;
  wire _11979_;
  wire _11980_;
  wire _11981_;
  wire _11982_;
  wire _11983_;
  wire _11984_;
  wire _11985_;
  wire _11986_;
  wire _11987_;
  wire _11988_;
  wire _11989_;
  wire _11990_;
  wire _11991_;
  wire _11992_;
  wire _11993_;
  wire _11994_;
  wire _11995_;
  wire _11996_;
  wire _11997_;
  wire _11998_;
  wire _11999_;
  wire _12000_;
  wire _12001_;
  wire _12002_;
  wire _12003_;
  wire _12004_;
  wire _12005_;
  wire _12006_;
  wire _12007_;
  wire _12008_;
  wire _12009_;
  wire _12010_;
  wire _12011_;
  wire _12012_;
  wire _12013_;
  wire _12014_;
  wire _12015_;
  wire _12016_;
  wire _12017_;
  wire _12018_;
  wire _12019_;
  wire _12020_;
  wire _12021_;
  wire _12022_;
  wire _12023_;
  wire _12024_;
  wire _12025_;
  wire _12026_;
  wire _12027_;
  wire _12028_;
  wire _12029_;
  wire _12030_;
  wire _12031_;
  wire _12032_;
  wire _12033_;
  wire _12034_;
  wire _12035_;
  wire _12036_;
  wire _12037_;
  wire _12038_;
  wire _12039_;
  wire _12040_;
  wire _12041_;
  wire _12042_;
  wire _12043_;
  wire _12044_;
  wire _12045_;
  wire _12046_;
  wire _12047_;
  wire _12048_;
  wire _12049_;
  wire _12050_;
  wire _12051_;
  wire _12052_;
  wire _12053_;
  wire _12054_;
  wire _12055_;
  wire _12056_;
  wire _12057_;
  wire _12058_;
  wire _12059_;
  wire _12060_;
  wire _12061_;
  wire _12062_;
  wire _12063_;
  wire _12064_;
  wire _12065_;
  wire _12066_;
  wire _12067_;
  wire _12068_;
  wire _12069_;
  wire _12070_;
  wire _12071_;
  wire _12072_;
  wire _12073_;
  wire _12074_;
  wire _12075_;
  wire _12076_;
  wire _12077_;
  wire _12078_;
  wire _12079_;
  wire _12080_;
  wire _12081_;
  wire _12082_;
  wire _12083_;
  wire _12084_;
  wire _12085_;
  wire _12086_;
  wire _12087_;
  wire _12088_;
  wire _12089_;
  wire _12090_;
  wire _12091_;
  wire _12092_;
  wire _12093_;
  wire _12094_;
  wire _12095_;
  wire _12096_;
  wire _12097_;
  wire _12098_;
  wire _12099_;
  wire _12100_;
  wire _12101_;
  wire _12102_;
  wire _12103_;
  wire _12104_;
  wire _12105_;
  wire _12106_;
  wire _12107_;
  wire _12108_;
  wire _12109_;
  wire _12110_;
  wire _12111_;
  wire _12112_;
  wire _12113_;
  wire _12114_;
  wire _12115_;
  wire _12116_;
  wire _12117_;
  wire _12118_;
  wire _12119_;
  wire _12120_;
  wire _12121_;
  wire _12122_;
  wire _12123_;
  wire _12124_;
  wire _12125_;
  wire _12126_;
  wire _12127_;
  wire _12128_;
  wire _12129_;
  wire _12130_;
  wire _12131_;
  wire _12132_;
  wire _12133_;
  wire _12134_;
  wire _12135_;
  wire _12136_;
  wire _12137_;
  wire _12138_;
  wire _12139_;
  wire _12140_;
  wire _12141_;
  wire _12142_;
  wire _12143_;
  wire _12144_;
  wire _12145_;
  wire _12146_;
  wire _12147_;
  wire _12148_;
  wire _12149_;
  wire _12150_;
  wire _12151_;
  wire _12152_;
  wire _12153_;
  wire _12154_;
  wire _12155_;
  wire _12156_;
  wire _12157_;
  wire _12158_;
  wire _12159_;
  wire _12160_;
  wire _12161_;
  wire _12162_;
  wire _12163_;
  wire _12164_;
  wire _12165_;
  wire _12166_;
  wire _12167_;
  wire _12168_;
  wire _12169_;
  wire _12170_;
  wire _12171_;
  wire _12172_;
  wire _12173_;
  wire _12174_;
  wire _12175_;
  wire _12176_;
  wire _12177_;
  wire _12178_;
  wire _12179_;
  wire _12180_;
  wire _12181_;
  wire _12182_;
  wire _12183_;
  wire _12184_;
  wire _12185_;
  wire _12186_;
  wire _12187_;
  wire _12188_;
  wire _12189_;
  wire _12190_;
  wire _12191_;
  wire _12192_;
  wire _12193_;
  wire _12194_;
  wire _12195_;
  wire _12196_;
  wire _12197_;
  wire _12198_;
  wire _12199_;
  wire _12200_;
  wire _12201_;
  wire _12202_;
  wire _12203_;
  wire _12204_;
  wire _12205_;
  wire _12206_;
  wire _12207_;
  wire _12208_;
  wire _12209_;
  wire _12210_;
  wire _12211_;
  wire _12212_;
  wire _12213_;
  wire _12214_;
  wire _12215_;
  wire _12216_;
  wire _12217_;
  wire _12218_;
  wire _12219_;
  wire _12220_;
  wire _12221_;
  wire _12222_;
  wire _12223_;
  wire _12224_;
  wire _12225_;
  wire _12226_;
  wire _12227_;
  wire _12228_;
  wire _12229_;
  wire _12230_;
  wire _12231_;
  wire _12232_;
  wire _12233_;
  wire _12234_;
  wire _12235_;
  wire _12236_;
  wire _12237_;
  wire _12238_;
  wire _12239_;
  wire _12240_;
  wire _12241_;
  wire _12242_;
  wire _12243_;
  wire _12244_;
  wire _12245_;
  wire _12246_;
  wire _12247_;
  wire _12248_;
  wire _12249_;
  wire _12250_;
  wire _12251_;
  wire _12252_;
  wire _12253_;
  wire _12254_;
  wire _12255_;
  wire _12256_;
  wire _12257_;
  wire _12258_;
  wire _12259_;
  wire _12260_;
  wire _12261_;
  wire _12262_;
  wire _12263_;
  wire _12264_;
  wire _12265_;
  wire _12266_;
  wire _12267_;
  wire _12268_;
  wire _12269_;
  wire _12270_;
  wire _12271_;
  wire _12272_;
  wire _12273_;
  wire _12274_;
  wire _12275_;
  wire _12276_;
  wire _12277_;
  wire _12278_;
  wire _12279_;
  wire _12280_;
  wire _12281_;
  wire _12282_;
  wire _12283_;
  wire _12284_;
  wire _12285_;
  wire _12286_;
  wire _12287_;
  wire _12288_;
  wire _12289_;
  wire _12290_;
  wire _12291_;
  wire _12292_;
  wire _12293_;
  wire _12294_;
  wire _12295_;
  wire _12296_;
  wire _12297_;
  wire _12298_;
  wire _12299_;
  wire _12300_;
  wire _12301_;
  wire _12302_;
  wire _12303_;
  wire _12304_;
  wire _12305_;
  wire _12306_;
  wire _12307_;
  wire _12308_;
  wire _12309_;
  wire _12310_;
  wire _12311_;
  wire _12312_;
  wire _12313_;
  wire _12314_;
  wire _12315_;
  wire _12316_;
  wire _12317_;
  wire _12318_;
  wire _12319_;
  wire _12320_;
  wire _12321_;
  wire _12322_;
  wire _12323_;
  wire _12324_;
  wire _12325_;
  wire _12326_;
  wire _12327_;
  wire _12328_;
  wire _12329_;
  wire _12330_;
  wire _12331_;
  wire _12332_;
  wire _12333_;
  wire _12334_;
  wire _12335_;
  wire _12336_;
  wire _12337_;
  wire _12338_;
  wire _12339_;
  wire _12340_;
  wire _12341_;
  wire _12342_;
  wire _12343_;
  wire _12344_;
  wire _12345_;
  wire _12346_;
  wire _12347_;
  wire _12348_;
  wire _12349_;
  wire _12350_;
  wire _12351_;
  wire _12352_;
  wire _12353_;
  wire _12354_;
  wire _12355_;
  wire _12356_;
  wire _12357_;
  wire _12358_;
  wire _12359_;
  wire _12360_;
  wire _12361_;
  wire _12362_;
  wire _12363_;
  wire _12364_;
  wire _12365_;
  wire _12366_;
  wire _12367_;
  wire _12368_;
  wire _12369_;
  wire _12370_;
  wire _12371_;
  wire _12372_;
  wire _12373_;
  wire _12374_;
  wire _12375_;
  wire _12376_;
  wire _12377_;
  wire _12378_;
  wire _12379_;
  wire _12380_;
  wire _12381_;
  wire _12382_;
  wire _12383_;
  wire _12384_;
  wire _12385_;
  wire _12386_;
  wire _12387_;
  wire _12388_;
  wire _12389_;
  wire _12390_;
  wire _12391_;
  wire _12392_;
  wire _12393_;
  wire _12394_;
  wire _12395_;
  wire _12396_;
  wire _12397_;
  wire _12398_;
  wire _12399_;
  wire _12400_;
  wire _12401_;
  wire _12402_;
  wire _12403_;
  wire _12404_;
  wire _12405_;
  wire _12406_;
  wire _12407_;
  wire _12408_;
  wire _12409_;
  wire _12410_;
  wire _12411_;
  wire _12412_;
  wire _12413_;
  wire _12414_;
  wire _12415_;
  wire _12416_;
  wire _12417_;
  wire _12418_;
  wire _12419_;
  wire _12420_;
  wire _12421_;
  wire _12422_;
  wire _12423_;
  wire _12424_;
  wire _12425_;
  wire _12426_;
  wire _12427_;
  wire _12428_;
  wire _12429_;
  wire _12430_;
  wire _12431_;
  wire _12432_;
  wire _12433_;
  wire _12434_;
  wire _12435_;
  wire _12436_;
  wire _12437_;
  wire _12438_;
  wire _12439_;
  wire _12440_;
  wire _12441_;
  wire _12442_;
  wire _12443_;
  wire _12444_;
  wire _12445_;
  wire _12446_;
  wire _12447_;
  wire _12448_;
  wire _12449_;
  wire _12450_;
  wire _12451_;
  wire _12452_;
  wire _12453_;
  wire _12454_;
  wire _12455_;
  wire _12456_;
  wire _12457_;
  wire _12458_;
  wire _12459_;
  wire _12460_;
  wire _12461_;
  wire _12462_;
  wire _12463_;
  wire _12464_;
  wire _12465_;
  wire _12466_;
  wire _12467_;
  wire _12468_;
  wire _12469_;
  wire _12470_;
  wire _12471_;
  wire _12472_;
  wire _12473_;
  wire _12474_;
  wire _12475_;
  wire _12476_;
  wire _12477_;
  wire _12478_;
  wire _12479_;
  wire _12480_;
  wire _12481_;
  wire _12482_;
  wire _12483_;
  wire _12484_;
  wire _12485_;
  wire _12486_;
  wire _12487_;
  wire _12488_;
  wire _12489_;
  wire _12490_;
  wire _12491_;
  wire _12492_;
  wire _12493_;
  wire _12494_;
  wire _12495_;
  wire _12496_;
  wire _12497_;
  wire _12498_;
  wire _12499_;
  wire _12500_;
  wire _12501_;
  wire _12502_;
  wire _12503_;
  wire _12504_;
  wire _12505_;
  wire _12506_;
  wire _12507_;
  wire _12508_;
  wire _12509_;
  wire _12510_;
  wire _12511_;
  wire _12512_;
  wire _12513_;
  wire _12514_;
  wire _12515_;
  wire _12516_;
  wire _12517_;
  wire _12518_;
  wire _12519_;
  wire _12520_;
  wire _12521_;
  wire _12522_;
  wire _12523_;
  wire _12524_;
  wire _12525_;
  wire _12526_;
  wire _12527_;
  wire _12528_;
  wire _12529_;
  wire _12530_;
  wire _12531_;
  wire _12532_;
  wire _12533_;
  wire _12534_;
  wire _12535_;
  wire _12536_;
  wire _12537_;
  wire _12538_;
  wire _12539_;
  wire _12540_;
  wire _12541_;
  wire _12542_;
  wire _12543_;
  wire _12544_;
  wire _12545_;
  wire _12546_;
  wire _12547_;
  wire _12548_;
  wire _12549_;
  wire _12550_;
  wire _12551_;
  wire _12552_;
  wire _12553_;
  wire _12554_;
  wire _12555_;
  wire _12556_;
  wire _12557_;
  wire _12558_;
  wire _12559_;
  wire _12560_;
  wire _12561_;
  wire _12562_;
  wire _12563_;
  wire _12564_;
  wire _12565_;
  wire _12566_;
  wire _12567_;
  wire _12568_;
  wire _12569_;
  wire _12570_;
  wire _12571_;
  wire _12572_;
  wire _12573_;
  wire _12574_;
  wire _12575_;
  wire _12576_;
  wire _12577_;
  wire _12578_;
  wire _12579_;
  wire _12580_;
  wire _12581_;
  wire _12582_;
  wire _12583_;
  wire _12584_;
  wire _12585_;
  wire _12586_;
  wire _12587_;
  wire _12588_;
  wire _12589_;
  wire _12590_;
  wire _12591_;
  wire _12592_;
  wire _12593_;
  wire _12594_;
  wire _12595_;
  wire _12596_;
  wire _12597_;
  wire _12598_;
  wire _12599_;
  wire _12600_;
  wire _12601_;
  wire _12602_;
  wire _12603_;
  wire _12604_;
  wire _12605_;
  wire _12606_;
  wire _12607_;
  wire _12608_;
  wire _12609_;
  wire _12610_;
  wire _12611_;
  wire _12612_;
  wire _12613_;
  wire _12614_;
  wire _12615_;
  wire _12616_;
  wire _12617_;
  wire _12618_;
  wire _12619_;
  wire _12620_;
  wire _12621_;
  wire _12622_;
  wire _12623_;
  wire _12624_;
  wire _12625_;
  wire _12626_;
  wire _12627_;
  wire _12628_;
  wire _12629_;
  wire _12630_;
  wire _12631_;
  wire _12632_;
  wire _12633_;
  wire _12634_;
  wire _12635_;
  wire _12636_;
  wire _12637_;
  wire _12638_;
  wire _12639_;
  wire _12640_;
  wire _12641_;
  wire _12642_;
  wire _12643_;
  wire _12644_;
  wire _12645_;
  wire _12646_;
  wire _12647_;
  wire _12648_;
  wire _12649_;
  wire _12650_;
  wire _12651_;
  wire _12652_;
  wire _12653_;
  wire _12654_;
  wire _12655_;
  wire _12656_;
  wire _12657_;
  wire _12658_;
  wire _12659_;
  wire _12660_;
  wire _12661_;
  wire _12662_;
  wire _12663_;
  wire _12664_;
  wire _12665_;
  wire _12666_;
  wire _12667_;
  wire _12668_;
  wire _12669_;
  wire _12670_;
  wire _12671_;
  wire _12672_;
  wire _12673_;
  wire _12674_;
  wire _12675_;
  wire _12676_;
  wire _12677_;
  wire _12678_;
  wire _12679_;
  wire _12680_;
  wire _12681_;
  wire _12682_;
  wire _12683_;
  wire _12684_;
  wire _12685_;
  wire _12686_;
  wire _12687_;
  wire _12688_;
  wire _12689_;
  wire _12690_;
  wire _12691_;
  wire _12692_;
  wire _12693_;
  wire _12694_;
  wire _12695_;
  wire _12696_;
  wire _12697_;
  wire _12698_;
  wire _12699_;
  wire _12700_;
  wire _12701_;
  wire _12702_;
  wire _12703_;
  wire _12704_;
  wire _12705_;
  wire _12706_;
  wire _12707_;
  wire _12708_;
  wire _12709_;
  wire _12710_;
  wire _12711_;
  wire _12712_;
  wire _12713_;
  wire _12714_;
  wire _12715_;
  wire _12716_;
  wire _12717_;
  wire _12718_;
  wire _12719_;
  wire _12720_;
  wire _12721_;
  wire _12722_;
  wire _12723_;
  wire _12724_;
  wire _12725_;
  wire _12726_;
  wire _12727_;
  wire _12728_;
  wire _12729_;
  wire _12730_;
  wire _12731_;
  wire _12732_;
  wire _12733_;
  wire _12734_;
  wire _12735_;
  wire _12736_;
  wire _12737_;
  wire _12738_;
  wire _12739_;
  wire _12740_;
  wire _12741_;
  wire _12742_;
  wire _12743_;
  wire _12744_;
  wire _12745_;
  wire _12746_;
  wire _12747_;
  wire _12748_;
  wire _12749_;
  wire _12750_;
  wire _12751_;
  wire _12752_;
  wire _12753_;
  wire _12754_;
  wire _12755_;
  wire _12756_;
  wire _12757_;
  wire _12758_;
  wire _12759_;
  wire _12760_;
  wire _12761_;
  wire _12762_;
  wire _12763_;
  wire _12764_;
  wire _12765_;
  wire _12766_;
  wire _12767_;
  wire _12768_;
  wire _12769_;
  wire _12770_;
  wire _12771_;
  wire _12772_;
  wire _12773_;
  wire _12774_;
  wire _12775_;
  wire _12776_;
  wire _12777_;
  wire _12778_;
  wire _12779_;
  wire _12780_;
  wire _12781_;
  wire _12782_;
  wire _12783_;
  wire _12784_;
  wire _12785_;
  wire _12786_;
  wire _12787_;
  wire _12788_;
  wire _12789_;
  wire _12790_;
  wire _12791_;
  wire _12792_;
  wire _12793_;
  wire _12794_;
  wire _12795_;
  wire _12796_;
  wire _12797_;
  wire _12798_;
  wire _12799_;
  wire _12800_;
  wire _12801_;
  wire _12802_;
  wire _12803_;
  wire _12804_;
  wire _12805_;
  wire _12806_;
  wire _12807_;
  wire _12808_;
  wire _12809_;
  wire _12810_;
  wire _12811_;
  wire _12812_;
  wire _12813_;
  wire _12814_;
  wire _12815_;
  wire _12816_;
  wire _12817_;
  wire _12818_;
  wire _12819_;
  wire _12820_;
  wire _12821_;
  wire _12822_;
  wire _12823_;
  wire _12824_;
  wire _12825_;
  wire _12826_;
  wire _12827_;
  wire _12828_;
  wire _12829_;
  wire _12830_;
  wire _12831_;
  wire _12832_;
  wire _12833_;
  wire _12834_;
  wire _12835_;
  wire _12836_;
  wire _12837_;
  wire _12838_;
  wire _12839_;
  wire _12840_;
  wire _12841_;
  wire _12842_;
  wire _12843_;
  wire _12844_;
  wire _12845_;
  wire _12846_;
  wire _12847_;
  wire _12848_;
  wire _12849_;
  wire _12850_;
  wire _12851_;
  wire _12852_;
  wire _12853_;
  wire _12854_;
  wire _12855_;
  wire _12856_;
  wire _12857_;
  wire _12858_;
  wire _12859_;
  wire _12860_;
  wire _12861_;
  wire _12862_;
  wire _12863_;
  wire _12864_;
  wire _12865_;
  wire _12866_;
  wire _12867_;
  wire _12868_;
  wire _12869_;
  wire _12870_;
  wire _12871_;
  wire _12872_;
  wire _12873_;
  wire _12874_;
  wire _12875_;
  wire _12876_;
  wire _12877_;
  wire _12878_;
  wire _12879_;
  wire _12880_;
  wire _12881_;
  wire _12882_;
  wire _12883_;
  wire _12884_;
  wire _12885_;
  wire _12886_;
  wire _12887_;
  wire _12888_;
  wire _12889_;
  wire _12890_;
  wire _12891_;
  wire _12892_;
  wire _12893_;
  wire _12894_;
  wire _12895_;
  wire _12896_;
  wire _12897_;
  wire _12898_;
  wire _12899_;
  wire _12900_;
  wire _12901_;
  wire _12902_;
  wire _12903_;
  wire _12904_;
  wire _12905_;
  wire _12906_;
  wire _12907_;
  wire _12908_;
  wire _12909_;
  wire _12910_;
  wire _12911_;
  wire _12912_;
  wire _12913_;
  wire _12914_;
  wire _12915_;
  wire _12916_;
  wire _12917_;
  wire _12918_;
  wire _12919_;
  wire _12920_;
  wire _12921_;
  wire _12922_;
  wire _12923_;
  wire _12924_;
  wire _12925_;
  wire _12926_;
  wire _12927_;
  wire _12928_;
  wire _12929_;
  wire _12930_;
  wire _12931_;
  wire _12932_;
  wire _12933_;
  wire _12934_;
  wire _12935_;
  wire _12936_;
  wire _12937_;
  wire _12938_;
  wire _12939_;
  wire _12940_;
  wire _12941_;
  wire _12942_;
  wire _12943_;
  wire _12944_;
  wire _12945_;
  wire _12946_;
  wire _12947_;
  wire _12948_;
  wire _12949_;
  wire _12950_;
  wire _12951_;
  wire _12952_;
  wire _12953_;
  wire _12954_;
  wire _12955_;
  wire _12956_;
  wire _12957_;
  wire _12958_;
  wire _12959_;
  wire _12960_;
  wire _12961_;
  wire _12962_;
  wire _12963_;
  wire _12964_;
  wire _12965_;
  wire _12966_;
  wire _12967_;
  wire _12968_;
  wire _12969_;
  wire _12970_;
  wire _12971_;
  wire _12972_;
  wire _12973_;
  wire _12974_;
  wire _12975_;
  wire _12976_;
  wire _12977_;
  wire _12978_;
  wire _12979_;
  wire _12980_;
  wire _12981_;
  wire _12982_;
  wire _12983_;
  wire _12984_;
  wire _12985_;
  wire _12986_;
  wire _12987_;
  wire _12988_;
  wire _12989_;
  wire _12990_;
  wire _12991_;
  wire _12992_;
  wire _12993_;
  wire _12994_;
  wire _12995_;
  wire _12996_;
  wire _12997_;
  wire _12998_;
  wire _12999_;
  wire _13000_;
  wire _13001_;
  wire _13002_;
  wire _13003_;
  wire _13004_;
  wire _13005_;
  wire _13006_;
  wire _13007_;
  wire _13008_;
  wire _13009_;
  wire _13010_;
  wire _13011_;
  wire _13012_;
  wire _13013_;
  wire _13014_;
  wire _13015_;
  wire _13016_;
  wire _13017_;
  wire _13018_;
  wire _13019_;
  wire _13020_;
  wire _13021_;
  wire _13022_;
  wire _13023_;
  wire _13024_;
  wire _13025_;
  wire _13026_;
  wire _13027_;
  wire _13028_;
  wire _13029_;
  wire _13030_;
  wire _13031_;
  wire _13032_;
  wire _13033_;
  wire _13034_;
  wire _13035_;
  wire _13036_;
  wire _13037_;
  wire _13038_;
  wire _13039_;
  wire _13040_;
  wire _13041_;
  wire _13042_;
  wire _13043_;
  wire _13044_;
  wire _13045_;
  wire _13046_;
  wire _13047_;
  wire _13048_;
  wire _13049_;
  wire _13050_;
  wire _13051_;
  wire _13052_;
  wire _13053_;
  wire _13054_;
  wire _13055_;
  wire _13056_;
  wire _13057_;
  wire _13058_;
  wire _13059_;
  wire _13060_;
  wire _13061_;
  wire _13062_;
  wire _13063_;
  wire _13064_;
  wire _13065_;
  wire _13066_;
  wire _13067_;
  wire _13068_;
  wire _13069_;
  wire _13070_;
  wire _13071_;
  wire _13072_;
  wire _13073_;
  wire _13074_;
  wire _13075_;
  wire _13076_;
  wire _13077_;
  wire _13078_;
  wire _13079_;
  wire _13080_;
  wire _13081_;
  wire _13082_;
  wire _13083_;
  wire _13084_;
  wire _13085_;
  wire _13086_;
  wire _13087_;
  wire _13088_;
  wire _13089_;
  wire _13090_;
  wire _13091_;
  wire _13092_;
  wire _13093_;
  wire _13094_;
  wire _13095_;
  wire _13096_;
  wire _13097_;
  wire _13098_;
  wire _13099_;
  wire _13100_;
  wire _13101_;
  wire _13102_;
  wire _13103_;
  wire _13104_;
  wire _13105_;
  wire _13106_;
  wire _13107_;
  wire _13108_;
  wire _13109_;
  wire _13110_;
  wire _13111_;
  wire _13112_;
  wire _13113_;
  wire _13114_;
  wire _13115_;
  wire _13116_;
  wire _13117_;
  wire _13118_;
  wire _13119_;
  wire _13120_;
  wire _13121_;
  wire _13122_;
  wire _13123_;
  wire _13124_;
  wire _13125_;
  wire _13126_;
  wire _13127_;
  wire _13128_;
  wire _13129_;
  wire _13130_;
  wire _13131_;
  wire _13132_;
  wire _13133_;
  wire _13134_;
  wire _13135_;
  wire _13136_;
  wire _13137_;
  wire _13138_;
  wire _13139_;
  wire _13140_;
  wire _13141_;
  wire _13142_;
  wire _13143_;
  wire _13144_;
  wire _13145_;
  wire _13146_;
  wire _13147_;
  wire _13148_;
  wire _13149_;
  wire _13150_;
  wire _13151_;
  wire _13152_;
  wire _13153_;
  wire _13154_;
  wire _13155_;
  wire _13156_;
  wire _13157_;
  wire _13158_;
  wire _13159_;
  wire _13160_;
  wire _13161_;
  wire _13162_;
  wire _13163_;
  wire _13164_;
  wire _13165_;
  wire _13166_;
  wire _13167_;
  wire _13168_;
  wire _13169_;
  wire _13170_;
  wire _13171_;
  wire _13172_;
  wire _13173_;
  wire _13174_;
  wire _13175_;
  wire _13176_;
  wire _13177_;
  wire _13178_;
  wire _13179_;
  wire _13180_;
  wire _13181_;
  wire _13182_;
  wire _13183_;
  wire _13184_;
  wire _13185_;
  wire _13186_;
  wire _13187_;
  wire _13188_;
  wire _13189_;
  wire _13190_;
  wire _13191_;
  wire _13192_;
  wire _13193_;
  wire _13194_;
  wire _13195_;
  wire _13196_;
  wire _13197_;
  wire _13198_;
  wire _13199_;
  wire _13200_;
  wire _13201_;
  wire _13202_;
  wire _13203_;
  wire _13204_;
  wire _13205_;
  wire _13206_;
  wire _13207_;
  wire _13208_;
  wire _13209_;
  wire _13210_;
  wire _13211_;
  wire _13212_;
  wire _13213_;
  wire _13214_;
  wire _13215_;
  wire _13216_;
  wire _13217_;
  wire _13218_;
  wire _13219_;
  wire _13220_;
  wire _13221_;
  wire _13222_;
  wire _13223_;
  wire _13224_;
  wire _13225_;
  wire _13226_;
  wire _13227_;
  wire _13228_;
  wire _13229_;
  wire _13230_;
  wire _13231_;
  wire _13232_;
  wire _13233_;
  wire _13234_;
  wire _13235_;
  wire _13236_;
  wire _13237_;
  wire _13238_;
  wire _13239_;
  wire _13240_;
  wire _13241_;
  wire _13242_;
  wire _13243_;
  wire _13244_;
  wire _13245_;
  wire _13246_;
  wire _13247_;
  wire _13248_;
  wire _13249_;
  wire _13250_;
  wire _13251_;
  wire _13252_;
  wire _13253_;
  wire _13254_;
  wire _13255_;
  wire _13256_;
  wire _13257_;
  wire _13258_;
  wire _13259_;
  wire _13260_;
  wire _13261_;
  wire _13262_;
  wire _13263_;
  wire _13264_;
  wire _13265_;
  wire _13266_;
  wire _13267_;
  wire _13268_;
  wire _13269_;
  wire _13270_;
  wire _13271_;
  wire _13272_;
  wire _13273_;
  wire _13274_;
  wire _13275_;
  wire _13276_;
  wire _13277_;
  wire _13278_;
  wire _13279_;
  wire _13280_;
  wire _13281_;
  wire _13282_;
  wire _13283_;
  wire _13284_;
  wire _13285_;
  wire _13286_;
  wire _13287_;
  wire _13288_;
  wire _13289_;
  wire _13290_;
  wire _13291_;
  wire _13292_;
  wire _13293_;
  wire _13294_;
  wire _13295_;
  wire _13296_;
  wire _13297_;
  wire _13298_;
  wire _13299_;
  wire _13300_;
  wire _13301_;
  wire _13302_;
  wire _13303_;
  wire _13304_;
  wire _13305_;
  wire _13306_;
  wire _13307_;
  wire _13308_;
  wire _13309_;
  wire _13310_;
  wire _13311_;
  wire _13312_;
  wire _13313_;
  wire _13314_;
  wire _13315_;
  wire _13316_;
  wire _13317_;
  wire _13318_;
  wire _13319_;
  wire _13320_;
  wire _13321_;
  wire _13322_;
  wire _13323_;
  wire _13324_;
  wire _13325_;
  wire _13326_;
  wire _13327_;
  wire _13328_;
  wire _13329_;
  wire _13330_;
  wire _13331_;
  wire _13332_;
  wire _13333_;
  wire _13334_;
  wire _13335_;
  wire _13336_;
  wire _13337_;
  wire _13338_;
  wire _13339_;
  wire _13340_;
  wire _13341_;
  wire _13342_;
  wire _13343_;
  wire _13344_;
  wire _13345_;
  wire _13346_;
  wire _13347_;
  wire _13348_;
  wire _13349_;
  wire _13350_;
  wire _13351_;
  wire _13352_;
  wire _13353_;
  wire _13354_;
  wire _13355_;
  wire _13356_;
  wire _13357_;
  wire _13358_;
  wire _13359_;
  wire _13360_;
  wire _13361_;
  wire _13362_;
  wire _13363_;
  wire _13364_;
  wire _13365_;
  wire _13366_;
  wire _13367_;
  wire _13368_;
  wire _13369_;
  wire _13370_;
  wire _13371_;
  wire _13372_;
  wire _13373_;
  wire _13374_;
  wire _13375_;
  wire _13376_;
  wire _13377_;
  wire _13378_;
  wire _13379_;
  wire _13380_;
  wire _13381_;
  wire _13382_;
  wire _13383_;
  wire _13384_;
  wire _13385_;
  wire _13386_;
  wire _13387_;
  wire _13388_;
  wire _13389_;
  wire _13390_;
  wire _13391_;
  wire _13392_;
  wire _13393_;
  wire _13394_;
  wire _13395_;
  wire _13396_;
  wire _13397_;
  wire _13398_;
  wire _13399_;
  wire _13400_;
  wire _13401_;
  wire _13402_;
  wire _13403_;
  wire _13404_;
  wire _13405_;
  wire _13406_;
  wire _13407_;
  wire _13408_;
  wire _13409_;
  wire _13410_;
  wire _13411_;
  wire _13412_;
  wire _13413_;
  wire _13414_;
  wire _13415_;
  wire _13416_;
  wire _13417_;
  wire _13418_;
  wire _13419_;
  wire _13420_;
  wire _13421_;
  wire _13422_;
  wire _13423_;
  wire _13424_;
  wire _13425_;
  wire _13426_;
  wire _13427_;
  wire _13428_;
  wire _13429_;
  wire _13430_;
  wire _13431_;
  wire _13432_;
  wire _13433_;
  wire _13434_;
  wire _13435_;
  wire _13436_;
  wire _13437_;
  wire _13438_;
  wire _13439_;
  wire _13440_;
  wire _13441_;
  wire _13442_;
  wire _13443_;
  wire _13444_;
  wire _13445_;
  wire _13446_;
  wire _13447_;
  wire _13448_;
  wire _13449_;
  wire _13450_;
  wire _13451_;
  wire _13452_;
  wire _13453_;
  wire _13454_;
  wire _13455_;
  wire _13456_;
  wire _13457_;
  wire _13458_;
  wire _13459_;
  wire _13460_;
  wire _13461_;
  wire _13462_;
  wire _13463_;
  wire _13464_;
  wire _13465_;
  wire _13466_;
  wire _13467_;
  wire _13468_;
  wire _13469_;
  wire _13470_;
  wire _13471_;
  wire _13472_;
  wire _13473_;
  wire _13474_;
  wire _13475_;
  wire _13476_;
  wire _13477_;
  wire _13478_;
  wire _13479_;
  wire _13480_;
  wire _13481_;
  wire _13482_;
  wire _13483_;
  wire _13484_;
  wire _13485_;
  wire _13486_;
  wire _13487_;
  wire _13488_;
  wire _13489_;
  wire _13490_;
  wire _13491_;
  wire _13492_;
  wire _13493_;
  wire _13494_;
  wire _13495_;
  wire _13496_;
  wire _13497_;
  wire _13498_;
  wire _13499_;
  wire _13500_;
  wire _13501_;
  wire _13502_;
  wire _13503_;
  wire _13504_;
  wire _13505_;
  wire _13506_;
  wire _13507_;
  wire _13508_;
  wire _13509_;
  wire _13510_;
  wire _13511_;
  wire _13512_;
  wire _13513_;
  wire _13514_;
  wire _13515_;
  wire _13516_;
  wire _13517_;
  wire _13518_;
  wire _13519_;
  wire _13520_;
  wire _13521_;
  wire _13522_;
  wire _13523_;
  wire _13524_;
  wire _13525_;
  wire _13526_;
  wire _13527_;
  wire _13528_;
  wire _13529_;
  wire _13530_;
  wire _13531_;
  wire _13532_;
  wire _13533_;
  wire _13534_;
  wire _13535_;
  wire _13536_;
  wire _13537_;
  wire _13538_;
  wire _13539_;
  wire _13540_;
  wire _13541_;
  wire _13542_;
  wire _13543_;
  wire _13544_;
  wire _13545_;
  wire _13546_;
  wire _13547_;
  wire _13548_;
  wire _13549_;
  wire _13550_;
  wire _13551_;
  wire _13552_;
  wire _13553_;
  wire _13554_;
  wire _13555_;
  wire _13556_;
  wire _13557_;
  wire _13558_;
  wire _13559_;
  wire _13560_;
  wire _13561_;
  wire _13562_;
  wire _13563_;
  wire _13564_;
  wire _13565_;
  wire _13566_;
  wire _13567_;
  wire _13568_;
  wire _13569_;
  wire _13570_;
  wire _13571_;
  wire _13572_;
  wire _13573_;
  wire _13574_;
  wire _13575_;
  wire _13576_;
  wire _13577_;
  wire _13578_;
  wire _13579_;
  wire _13580_;
  wire _13581_;
  wire _13582_;
  wire _13583_;
  wire _13584_;
  wire _13585_;
  wire _13586_;
  wire _13587_;
  wire _13588_;
  wire _13589_;
  wire _13590_;
  wire _13591_;
  wire _13592_;
  wire _13593_;
  wire _13594_;
  wire _13595_;
  wire _13596_;
  wire _13597_;
  wire _13598_;
  wire _13599_;
  wire _13600_;
  wire _13601_;
  wire _13602_;
  wire _13603_;
  wire _13604_;
  wire _13605_;
  wire _13606_;
  wire _13607_;
  wire _13608_;
  wire _13609_;
  wire _13610_;
  wire _13611_;
  wire _13612_;
  wire _13613_;
  wire _13614_;
  wire _13615_;
  wire _13616_;
  wire _13617_;
  wire _13618_;
  wire _13619_;
  wire _13620_;
  wire _13621_;
  wire _13622_;
  wire _13623_;
  wire _13624_;
  wire _13625_;
  wire _13626_;
  wire _13627_;
  wire _13628_;
  wire _13629_;
  wire _13630_;
  wire _13631_;
  wire _13632_;
  wire _13633_;
  wire _13634_;
  wire _13635_;
  wire _13636_;
  wire _13637_;
  wire _13638_;
  wire _13639_;
  wire _13640_;
  wire _13641_;
  wire _13642_;
  wire _13643_;
  wire _13644_;
  wire _13645_;
  wire _13646_;
  wire _13647_;
  wire _13648_;
  wire _13649_;
  wire _13650_;
  wire _13651_;
  wire _13652_;
  wire _13653_;
  wire _13654_;
  wire _13655_;
  wire _13656_;
  wire _13657_;
  wire _13658_;
  wire _13659_;
  wire _13660_;
  wire _13661_;
  wire _13662_;
  wire _13663_;
  wire _13664_;
  wire _13665_;
  wire _13666_;
  wire _13667_;
  wire _13668_;
  wire _13669_;
  wire _13670_;
  wire _13671_;
  wire _13672_;
  wire _13673_;
  wire _13674_;
  wire _13675_;
  wire _13676_;
  wire _13677_;
  wire _13678_;
  wire _13679_;
  wire _13680_;
  wire _13681_;
  wire _13682_;
  wire _13683_;
  wire _13684_;
  wire _13685_;
  wire _13686_;
  wire _13687_;
  wire _13688_;
  wire _13689_;
  wire _13690_;
  wire _13691_;
  wire _13692_;
  wire _13693_;
  wire _13694_;
  wire _13695_;
  wire _13696_;
  wire _13697_;
  wire _13698_;
  wire _13699_;
  wire _13700_;
  wire _13701_;
  wire _13702_;
  wire _13703_;
  wire _13704_;
  wire _13705_;
  wire _13706_;
  wire _13707_;
  wire _13708_;
  wire _13709_;
  wire _13710_;
  wire _13711_;
  wire _13712_;
  wire _13713_;
  wire _13714_;
  wire _13715_;
  wire _13716_;
  wire _13717_;
  wire _13718_;
  wire _13719_;
  wire _13720_;
  wire _13721_;
  wire _13722_;
  wire _13723_;
  wire _13724_;
  wire _13725_;
  wire _13726_;
  wire _13727_;
  wire _13728_;
  wire _13729_;
  wire _13730_;
  wire _13731_;
  wire _13732_;
  wire _13733_;
  wire _13734_;
  wire _13735_;
  wire _13736_;
  wire _13737_;
  wire _13738_;
  wire _13739_;
  wire _13740_;
  wire _13741_;
  wire _13742_;
  wire _13743_;
  wire _13744_;
  wire _13745_;
  wire _13746_;
  wire _13747_;
  wire _13748_;
  wire _13749_;
  wire _13750_;
  wire _13751_;
  wire _13752_;
  wire _13753_;
  wire _13754_;
  wire _13755_;
  wire _13756_;
  wire _13757_;
  wire _13758_;
  wire _13759_;
  wire _13760_;
  wire _13761_;
  wire _13762_;
  wire _13763_;
  wire _13764_;
  wire _13765_;
  wire _13766_;
  wire _13767_;
  wire _13768_;
  wire _13769_;
  wire _13770_;
  wire _13771_;
  wire _13772_;
  wire _13773_;
  wire _13774_;
  wire _13775_;
  wire _13776_;
  wire _13777_;
  wire _13778_;
  wire _13779_;
  wire _13780_;
  wire _13781_;
  wire _13782_;
  wire _13783_;
  wire _13784_;
  wire _13785_;
  wire _13786_;
  wire _13787_;
  wire _13788_;
  wire _13789_;
  wire _13790_;
  wire _13791_;
  wire _13792_;
  wire _13793_;
  wire _13794_;
  wire _13795_;
  wire _13796_;
  wire _13797_;
  wire _13798_;
  wire _13799_;
  wire _13800_;
  wire _13801_;
  wire _13802_;
  wire _13803_;
  wire _13804_;
  wire _13805_;
  wire _13806_;
  wire _13807_;
  wire _13808_;
  wire _13809_;
  wire _13810_;
  wire _13811_;
  wire _13812_;
  wire _13813_;
  wire _13814_;
  wire _13815_;
  wire _13816_;
  wire _13817_;
  wire _13818_;
  wire _13819_;
  wire _13820_;
  wire _13821_;
  wire _13822_;
  wire _13823_;
  wire _13824_;
  wire [7:0] _13825_;
  wire [7:0] _13826_;
  wire _13827_;
  wire [7:0] _13828_;
  wire [7:0] _13829_;
  wire [7:0] _13830_;
  wire [7:0] _13831_;
  wire [7:0] _13832_;
  wire [7:0] _13833_;
  wire [7:0] _13834_;
  wire [7:0] _13835_;
  wire [7:0] _13836_;
  wire [7:0] _13837_;
  wire [7:0] _13838_;
  wire [15:0] _13839_;
  wire [7:0] _13840_;
  wire [7:0] _13841_;
  wire [7:0] _13842_;
  wire [7:0] _13843_;
  wire [7:0] _13844_;
  wire [7:0] _13845_;
  wire [7:0] _13846_;
  wire [7:0] _13847_;
  wire [7:0] _13848_;
  wire [7:0] _13849_;
  wire [15:0] _13850_;
  wire [7:0] _13851_;
  wire _13852_;
  wire _13853_;
  wire _13854_;
  wire _13855_;
  wire _13856_;
  wire _13857_;
  wire _13858_;
  wire _13859_;
  wire _13860_;
  wire _13861_;
  wire _13862_;
  wire _13863_;
  wire _13864_;
  wire _13865_;
  wire _13866_;
  wire _13867_;
  wire _13868_;
  wire _13869_;
  wire _13870_;
  wire _13871_;
  wire _13872_;
  wire _13873_;
  wire _13874_;
  wire _13875_;
  wire _13876_;
  wire _13877_;
  wire _13878_;
  wire _13879_;
  wire _13880_;
  wire _13881_;
  wire _13882_;
  wire _13883_;
  wire _13884_;
  wire _13885_;
  wire _13886_;
  wire _13887_;
  wire _13888_;
  wire _13889_;
  wire _13890_;
  wire _13891_;
  wire _13892_;
  wire _13893_;
  wire _13894_;
  wire _13895_;
  wire _13896_;
  wire _13897_;
  wire _13898_;
  wire _13899_;
  wire [7:0] _13900_;
  wire [7:0] _13901_;
  wire [7:0] _13902_;
  wire [7:0] _13903_;
  wire [7:0] _13904_;
  wire [7:0] _13905_;
  wire [7:0] _13906_;
  wire [7:0] _13907_;
  wire [7:0] _13908_;
  wire [7:0] _13909_;
  wire [7:0] _13910_;
  wire [7:0] _13911_;
  wire [7:0] _13912_;
  wire [2:0] _13913_;
  wire [2:0] _13914_;
  wire [1:0] _13915_;
  wire [7:0] _13916_;
  wire _13917_;
  wire [1:0] _13918_;
  wire [1:0] _13919_;
  wire [2:0] _13920_;
  wire [2:0] _13921_;
  wire [1:0] _13922_;
  wire [3:0] _13923_;
  wire [1:0] _13924_;
  wire _13925_;
  wire _13926_;
  wire [15:0] _13927_;
  wire [15:0] _13928_;
  wire _13929_;
  wire _13930_;
  wire [4:0] _13931_;
  wire [7:0] _13932_;
  wire [7:0] _13933_;
  wire [7:0] _13934_;
  wire _13935_;
  wire _13936_;
  wire [7:0] _13937_;
  wire [15:0] _13938_;
  wire [15:0] _13939_;
  wire _13940_;
  wire _13941_;
  wire _13942_;
  wire [7:0] _13943_;
  wire [2:0] _13944_;
  wire [7:0] _13945_;
  wire [7:0] _13946_;
  wire _13947_;
  wire [7:0] _13948_;
  wire _13949_;
  wire _13950_;
  wire [3:0] _13951_;
  wire [31:0] _13952_;
  wire [31:0] _13953_;
  wire [7:0] _13954_;
  wire _13955_;
  wire _13956_;
  wire [15:0] _13957_;
  wire _13958_;
  wire _13959_;
  wire _13960_;
  wire [15:0] _13961_;
  wire _13962_;
  wire _13963_;
  wire [7:0] _13964_;
  wire _13965_;
  wire [2:0] _13966_;
  wire _13967_;
  wire _13968_;
  wire [7:0] _13969_;
  wire _13970_;
  input [7:0] ACC_abstr;
  wire [7:0] ACC_gm;
  input [7:0] B_abstr;
  wire [7:0] B_gm;
  input [7:0] DPH_abstr;
  wire [7:0] DPH_gm;
  input [7:0] DPL_abstr;
  wire [7:0] DPL_gm;
  wire [7:0] IE_gm;
  wire [7:0] IE_gm_next;
  wire [7:0] IP_gm;
  wire [7:0] IP_gm_next;
  input [7:0] P0_abstr;
  wire [7:0] P0_gm;
  input [7:0] P1_abstr;
  wire [7:0] P1_gm;
  input [7:0] P2_abstr;
  wire [7:0] P2_gm;
  input [7:0] P3_abstr;
  wire [7:0] P3_gm;
  wire [7:0] PCON_gm;
  wire [7:0] PCON_gm_next;
  input [15:0] PC_abstr;
  input [7:0] PSW_abstr;
  wire [7:0] PSW_gm;
  input [7:0] RD_IRAM_0_ABSTR_ADDR;
  input [7:0] RD_IRAM_1_ABSTR_ADDR;
  input [15:0] RD_ROM_1_ABSTR_ADDR;
  input [15:0] RD_ROM_2_ABSTR_ADDR;
  wire [7:0] SBUF_gm;
  wire [7:0] SBUF_gm_next;
  wire [7:0] SCON_gm;
  wire [7:0] SCON_gm_next;
  input [7:0] SP_abstr;
  wire [7:0] SP_gm;
  wire [7:0] TCON_gm;
  wire [7:0] TCON_gm_next;
  wire [7:0] TH0_gm;
  wire [7:0] TH0_gm_next;
  wire [7:0] TH1_gm;
  wire [7:0] TH1_gm_next;
  wire [7:0] TL0_gm;
  wire [7:0] TL0_gm_next;
  wire [7:0] TL1_gm;
  wire [7:0] TL1_gm_next;
  wire [7:0] TMOD_gm;
  wire [7:0] TMOD_gm_next;
  input [3:0] WR_ADDR_ABSTR_IRAM_0;
  input [3:0] WR_ADDR_ABSTR_IRAM_1;
  input WR_COND_ABSTR_IRAM_0;
  input WR_COND_ABSTR_IRAM_1;
  input [7:0] WR_DATA_ABSTR_IRAM_0;
  input [7:0] WR_DATA_ABSTR_IRAM_1;
  input [15:0] XRAM_ADDR_abstr;
  input [7:0] XRAM_DATA_OUT_abstr;
  wire [7:0] acc_impl;
  wire [7:0] b_reg_impl;
  input clk;
  wire [31:0] cxrom_data_out;
  wire [15:0] dptr_impl;
  wire eq_state_1;
  wire eq_state_2;
  wire inst_finished_r;
  wire \oc8051_gm_cxrom_1.cell0.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell0.data ;
  wire \oc8051_gm_cxrom_1.cell0.rst ;
  wire \oc8051_gm_cxrom_1.cell0.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell0.word ;
  wire \oc8051_gm_cxrom_1.cell1.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell1.data ;
  wire \oc8051_gm_cxrom_1.cell1.rst ;
  wire \oc8051_gm_cxrom_1.cell1.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell1.word ;
  wire \oc8051_gm_cxrom_1.cell10.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell10.data ;
  wire \oc8051_gm_cxrom_1.cell10.rst ;
  wire \oc8051_gm_cxrom_1.cell10.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell10.word ;
  wire \oc8051_gm_cxrom_1.cell11.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell11.data ;
  wire \oc8051_gm_cxrom_1.cell11.rst ;
  wire \oc8051_gm_cxrom_1.cell11.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell11.word ;
  wire \oc8051_gm_cxrom_1.cell12.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell12.data ;
  wire \oc8051_gm_cxrom_1.cell12.rst ;
  wire \oc8051_gm_cxrom_1.cell12.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell12.word ;
  wire \oc8051_gm_cxrom_1.cell13.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell13.data ;
  wire \oc8051_gm_cxrom_1.cell13.rst ;
  wire \oc8051_gm_cxrom_1.cell13.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell13.word ;
  wire \oc8051_gm_cxrom_1.cell14.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell14.data ;
  wire \oc8051_gm_cxrom_1.cell14.rst ;
  wire \oc8051_gm_cxrom_1.cell14.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell14.word ;
  wire \oc8051_gm_cxrom_1.cell15.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell15.data ;
  wire \oc8051_gm_cxrom_1.cell15.rst ;
  wire \oc8051_gm_cxrom_1.cell15.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell15.word ;
  wire \oc8051_gm_cxrom_1.cell2.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell2.data ;
  wire \oc8051_gm_cxrom_1.cell2.rst ;
  wire \oc8051_gm_cxrom_1.cell2.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell2.word ;
  wire \oc8051_gm_cxrom_1.cell3.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell3.data ;
  wire \oc8051_gm_cxrom_1.cell3.rst ;
  wire \oc8051_gm_cxrom_1.cell3.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell3.word ;
  wire \oc8051_gm_cxrom_1.cell4.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell4.data ;
  wire \oc8051_gm_cxrom_1.cell4.rst ;
  wire \oc8051_gm_cxrom_1.cell4.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell4.word ;
  wire \oc8051_gm_cxrom_1.cell5.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell5.data ;
  wire \oc8051_gm_cxrom_1.cell5.rst ;
  wire \oc8051_gm_cxrom_1.cell5.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell5.word ;
  wire \oc8051_gm_cxrom_1.cell6.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell6.data ;
  wire \oc8051_gm_cxrom_1.cell6.rst ;
  wire \oc8051_gm_cxrom_1.cell6.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell6.word ;
  wire \oc8051_gm_cxrom_1.cell7.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell7.data ;
  wire \oc8051_gm_cxrom_1.cell7.rst ;
  wire \oc8051_gm_cxrom_1.cell7.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell7.word ;
  wire \oc8051_gm_cxrom_1.cell8.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell8.data ;
  wire \oc8051_gm_cxrom_1.cell8.rst ;
  wire \oc8051_gm_cxrom_1.cell8.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell8.word ;
  wire \oc8051_gm_cxrom_1.cell9.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell9.data ;
  wire \oc8051_gm_cxrom_1.cell9.rst ;
  wire \oc8051_gm_cxrom_1.cell9.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell9.word ;
  wire \oc8051_gm_cxrom_1.clk ;
  wire [31:0] \oc8051_gm_cxrom_1.cxrom_data_out ;
  wire [15:0] \oc8051_gm_cxrom_1.rd_addr_0 ;
  wire [15:0] \oc8051_gm_cxrom_1.rd_addr_2 ;
  wire \oc8051_gm_cxrom_1.rst ;
  wire [127:0] \oc8051_gm_cxrom_1.word_in ;
  wire [7:0] \oc8051_golden_model_1.ACC ;
  wire [7:0] \oc8051_golden_model_1.ACC_abstr ;
  wire [7:0] \oc8051_golden_model_1.B ;
  wire [7:0] \oc8051_golden_model_1.B_abstr ;
  wire [7:0] \oc8051_golden_model_1.DPH ;
  wire [7:0] \oc8051_golden_model_1.DPH_abstr ;
  wire [7:0] \oc8051_golden_model_1.DPL ;
  wire [7:0] \oc8051_golden_model_1.DPL_abstr ;
  wire [7:0] \oc8051_golden_model_1.IE ;
  wire [7:0] \oc8051_golden_model_1.IE_next ;
  wire [7:0] \oc8051_golden_model_1.IP ;
  wire [7:0] \oc8051_golden_model_1.IP_next ;
  wire [7:0] \oc8051_golden_model_1.IRAM[0] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[10] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[11] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[12] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[13] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[14] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[15] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[1] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[2] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[3] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[4] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[5] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[6] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[7] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[8] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[9] ;
  wire [7:0] \oc8051_golden_model_1.P0 ;
  wire [7:0] \oc8051_golden_model_1.P0_abstr ;
  wire [7:0] \oc8051_golden_model_1.P1 ;
  wire [7:0] \oc8051_golden_model_1.P1_abstr ;
  wire [7:0] \oc8051_golden_model_1.P2 ;
  wire [7:0] \oc8051_golden_model_1.P2_abstr ;
  wire [7:0] \oc8051_golden_model_1.P3 ;
  wire [7:0] \oc8051_golden_model_1.P3_abstr ;
  wire [15:0] \oc8051_golden_model_1.PC ;
  wire [7:0] \oc8051_golden_model_1.PCON ;
  wire [7:0] \oc8051_golden_model_1.PCON_next ;
  wire [15:0] \oc8051_golden_model_1.PC_abstr ;
  wire [7:0] \oc8051_golden_model_1.PSW ;
  wire [7:0] \oc8051_golden_model_1.PSW_abstr ;
  wire [7:0] \oc8051_golden_model_1.RD_IRAM_0_ABSTR_ADDR ;
  wire [7:0] \oc8051_golden_model_1.RD_IRAM_1 ;
  wire [7:0] \oc8051_golden_model_1.RD_IRAM_1_ABSTR_ADDR ;
  wire [7:0] \oc8051_golden_model_1.RD_IRAM_1_ADDR ;
  wire [15:0] \oc8051_golden_model_1.RD_ROM_0_ADDR ;
  wire [15:0] \oc8051_golden_model_1.RD_ROM_1_ABSTR_ADDR ;
  wire [15:0] \oc8051_golden_model_1.RD_ROM_2_ABSTR_ADDR ;
  wire [15:0] \oc8051_golden_model_1.RD_ROM_2_ADDR ;
  wire [7:0] \oc8051_golden_model_1.SBUF ;
  wire [7:0] \oc8051_golden_model_1.SBUF_next ;
  wire [7:0] \oc8051_golden_model_1.SCON ;
  wire [7:0] \oc8051_golden_model_1.SCON_next ;
  wire [7:0] \oc8051_golden_model_1.SP ;
  wire [7:0] \oc8051_golden_model_1.SP_abstr ;
  wire [7:0] \oc8051_golden_model_1.TCON ;
  wire [7:0] \oc8051_golden_model_1.TCON_next ;
  wire [7:0] \oc8051_golden_model_1.TH0 ;
  wire [7:0] \oc8051_golden_model_1.TH0_next ;
  wire [7:0] \oc8051_golden_model_1.TH1 ;
  wire [7:0] \oc8051_golden_model_1.TH1_next ;
  wire [7:0] \oc8051_golden_model_1.TL0 ;
  wire [7:0] \oc8051_golden_model_1.TL0_next ;
  wire [7:0] \oc8051_golden_model_1.TL1 ;
  wire [7:0] \oc8051_golden_model_1.TL1_next ;
  wire [7:0] \oc8051_golden_model_1.TMOD ;
  wire [7:0] \oc8051_golden_model_1.TMOD_next ;
  wire [3:0] \oc8051_golden_model_1.WR_ADDR_1_IRAM ;
  wire [3:0] \oc8051_golden_model_1.WR_ADDR_ABSTR_IRAM_0 ;
  wire [3:0] \oc8051_golden_model_1.WR_ADDR_ABSTR_IRAM_1 ;
  wire \oc8051_golden_model_1.WR_COND_ABSTR_IRAM_0 ;
  wire \oc8051_golden_model_1.WR_COND_ABSTR_IRAM_1 ;
  wire [7:0] \oc8051_golden_model_1.WR_DATA_1_IRAM ;
  wire [7:0] \oc8051_golden_model_1.WR_DATA_ABSTR_IRAM_0 ;
  wire [7:0] \oc8051_golden_model_1.WR_DATA_ABSTR_IRAM_1 ;
  wire [15:0] \oc8051_golden_model_1.XRAM_ADDR ;
  wire [15:0] \oc8051_golden_model_1.XRAM_ADDR_abstr ;
  wire [7:0] \oc8051_golden_model_1.XRAM_DATA_IN ;
  wire [7:0] \oc8051_golden_model_1.XRAM_DATA_OUT ;
  wire [7:0] \oc8051_golden_model_1.XRAM_DATA_OUT_abstr ;
  wire \oc8051_golden_model_1.clk ;
  wire [3:0] \oc8051_golden_model_1.n0006 ;
  wire [1:0] \oc8051_golden_model_1.n0115 ;
  wire [7:0] \oc8051_golden_model_1.n0116 ;
  wire [3:0] \oc8051_golden_model_1.n0117 ;
  wire [7:0] \oc8051_golden_model_1.n0120 ;
  wire [3:0] \oc8051_golden_model_1.n0121 ;
  wire [7:0] \oc8051_golden_model_1.n0123 ;
  wire [3:0] \oc8051_golden_model_1.n0124 ;
  wire [7:0] \oc8051_golden_model_1.n0126 ;
  wire [3:0] \oc8051_golden_model_1.n0127 ;
  wire [7:0] \oc8051_golden_model_1.n0129 ;
  wire [3:0] \oc8051_golden_model_1.n0130 ;
  wire [7:0] \oc8051_golden_model_1.n0132 ;
  wire [3:0] \oc8051_golden_model_1.n0133 ;
  wire [7:0] \oc8051_golden_model_1.n0135 ;
  wire [3:0] \oc8051_golden_model_1.n0136 ;
  wire [7:0] \oc8051_golden_model_1.n0138 ;
  wire [3:0] \oc8051_golden_model_1.n0139 ;
  wire \oc8051_golden_model_1.n0246 ;
  wire [7:0] \oc8051_golden_model_1.n0247 ;
  wire [3:0] \oc8051_golden_model_1.n0288 ;
  wire [7:0] \oc8051_golden_model_1.n0289 ;
  wire \oc8051_golden_model_1.rst ;
  wire [7:0] \oc8051_top_1.acc ;
  wire [7:0] \oc8051_top_1.b_reg ;
  wire [31:0] \oc8051_top_1.cxrom_data_out ;
  wire \oc8051_top_1.cy ;
  wire [1:0] \oc8051_top_1.cy_sel ;
  wire [15:0] \oc8051_top_1.dptr ;
  wire [7:0] \oc8051_top_1.dptr_hi ;
  wire [7:0] \oc8051_top_1.dptr_lo ;
  wire \oc8051_top_1.ea_int ;
  wire [31:0] \oc8051_top_1.idat_onchip ;
  wire \oc8051_top_1.int_ack ;
  wire \oc8051_top_1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.mem_act ;
  wire \oc8051_top_1.oc8051_alu1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.divsrc2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.des2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div0 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.div_out ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.rst ;
  wire [5:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.rst ;
  wire [15:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul ;
  wire \oc8051_top_1.oc8051_alu1.rst ;
  wire \oc8051_top_1.oc8051_alu1.srcAc ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.acc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.clk ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.dptr ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op1_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op2_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op3_r ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.pc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_alu_src_sel1.sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_alu_src_sel1.sel2 ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.sel3 ;
  wire [7:0] \oc8051_top_1.oc8051_comp1.acc ;
  wire \oc8051_top_1.oc8051_comp1.cy ;
  wire \oc8051_top_1.oc8051_cy_select1.cy_in ;
  wire [1:0] \oc8051_top_1.oc8051_cy_select1.cy_sel ;
  wire [3:0] \oc8051_top_1.oc8051_decoder1.alu_op ;
  wire \oc8051_top_1.oc8051_decoder1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.cy_sel ;
  wire \oc8051_top_1.oc8051_decoder1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_decoder1.op ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.psw_set ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_wr_sel ;
  wire \oc8051_top_1.oc8051_decoder1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.src_sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.src_sel2 ;
  wire \oc8051_top_1.oc8051_decoder1.src_sel3 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.state ;
  wire \oc8051_top_1.oc8051_decoder1.wait_data ;
  wire \oc8051_top_1.oc8051_decoder1.wr ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.wr_sfr ;
  wire \oc8051_top_1.oc8051_indi_addr1.clk ;
  wire \oc8051_top_1.oc8051_indi_addr1.rst ;
  wire \oc8051_top_1.oc8051_indi_addr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.cdata ;
  wire \oc8051_top_1.oc8051_memory_interface1.cdone ;
  wire \oc8051_top_1.oc8051_memory_interface1.clk ;
  wire \oc8051_top_1.oc8051_memory_interface1.dack_i ;
  wire \oc8051_top_1.oc8051_memory_interface1.dack_ir ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dadr_o ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dadr_ot ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_i ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_ir ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.dmem_wait ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dptr ;
  wire \oc8051_top_1.oc8051_memory_interface1.dstb_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.dwe_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.ea_int ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.iadr_t ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_cur ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_old ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_onchip ;
  wire \oc8051_top_1.oc8051_memory_interface1.imem_wait ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm2_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_t ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_vec_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.istb_t ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op2_buff ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op3_buff ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.op_pos ;
  wire \oc8051_top_1.oc8051_memory_interface1.out_of_rst ;
  wire [3:0] \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_buf ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log_prev ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_addr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_ind ;
  wire \oc8051_top_1.oc8051_memory_interface1.reti ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ri_r ;
  wire [4:0] \oc8051_top_1.oc8051_memory_interface1.rn_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.sfr ;
  wire \oc8051_top_1.oc8051_memory_interface1.sfr_bit ;
  wire \oc8051_top_1.oc8051_ram_top1.bit_addr_r ;
  wire [2:0] \oc8051_top_1.oc8051_ram_top1.bit_select ;
  wire \oc8051_top_1.oc8051_ram_top1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.rd_data_m ;
  wire \oc8051_top_1.oc8051_ram_top1.rd_en_r ;
  wire \oc8051_top_1.oc8051_ram_top1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.wr_data_r ;
  wire \oc8051_top_1.oc8051_rom1.clk ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.cxrom_data_out ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.data_o ;
  wire \oc8051_top_1.oc8051_rom1.ea_int ;
  wire \oc8051_top_1.oc8051_rom1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.b_reg ;
  wire \oc8051_top_1.oc8051_sfr1.bit_out ;
  wire \oc8051_top_1.oc8051_sfr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.cy ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_lo ;
  wire \oc8051_top_1.oc8051_sfr1.int_ack ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.p ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ack ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.set ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.p ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw_next ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.psw_set ;
  wire \oc8051_top_1.oc8051_sfr1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.srcAc ;
  wire \oc8051_top_1.oc8051_sfr1.wait_data ;
  wire \oc8051_top_1.oc8051_sfr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.p0_o ;
  wire [7:0] \oc8051_top_1.p1_o ;
  wire [7:0] \oc8051_top_1.p2_o ;
  wire [7:0] \oc8051_top_1.p3_o ;
  wire [15:0] \oc8051_top_1.pc ;
  wire [15:0] \oc8051_top_1.pc_log ;
  wire [15:0] \oc8051_top_1.pc_log_prev ;
  wire [7:0] \oc8051_top_1.psw ;
  wire [1:0] \oc8051_top_1.psw_set ;
  wire \oc8051_top_1.rd_ind ;
  wire \oc8051_top_1.reti ;
  wire \oc8051_top_1.sfr_bit ;
  wire [7:0] \oc8051_top_1.sfr_out ;
  wire \oc8051_top_1.srcAc ;
  wire [2:0] \oc8051_top_1.src_sel1 ;
  wire [1:0] \oc8051_top_1.src_sel2 ;
  wire \oc8051_top_1.src_sel3 ;
  wire \oc8051_top_1.wait_data ;
  wire \oc8051_top_1.wb_clk_i ;
  wire \oc8051_top_1.wb_rst_i ;
  wire \oc8051_top_1.wbd_ack_i ;
  wire [15:0] \oc8051_top_1.wbd_adr_o ;
  wire \oc8051_top_1.wbd_cyc_o ;
  wire [7:0] \oc8051_top_1.wbd_dat_i ;
  wire [7:0] \oc8051_top_1.wbd_dat_o ;
  wire \oc8051_top_1.wbd_stb_o ;
  wire \oc8051_top_1.wbd_we_o ;
  wire op0_cnst;
  input [7:0] p0_in;
  wire [7:0] p0_out;
  wire [7:0] p0in_reg;
  input [7:0] p1_in;
  wire [7:0] p1_out;
  wire [7:0] p1in_reg;
  input [7:0] p2_in;
  wire [7:0] p2_out;
  wire [7:0] p2in_reg;
  input [7:0] p3_in;
  wire [7:0] p3_out;
  wire [7:0] p3in_reg;
  wire [15:0] pc1;
  wire [15:0] pc2;
  output property_invalid_acc;
  output property_invalid_b_reg;
  output property_invalid_dph;
  output property_invalid_dpl;
  output property_invalid_iram;
  output property_invalid_p0;
  output property_invalid_p1;
  output property_invalid_p2;
  output property_invalid_p3;
  output property_invalid_pc;
  output property_invalid_psw;
  output property_invalid_xram_addr;
  output property_invalid_xram_data_out;
  wire property_valid_psw_1_r;
  wire [7:0] psw_impl;
  wire [15:0] rd_rom_0_addr;
  wire [15:0] rd_rom_2_addr;
  input rst;
  wire this_op_cnst_r;
  wire wbd_ack_i;
  wire [15:0] wbd_adr_o;
  wire wbd_cyc_o;
  wire [7:0] wbd_dat_i;
  wire [7:0] wbd_dat_o;
  wire wbd_stb_o;
  wire wbd_we_o;
  input [127:0] word_in;
  input [7:0] xram_data_in;
  wire [7:0] xram_data_in_model;
  wire [7:0] xram_data_in_reg;
  not (_13707_, rst);
  not (_06840_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  not (_06841_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_06842_, \oc8051_top_1.oc8051_decoder1.alu_op [1], _06841_);
  and (_06843_, _06842_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_06844_, \oc8051_top_1.oc8051_decoder1.alu_op [2], _06841_);
  and (_06845_, \oc8051_top_1.oc8051_decoder1.alu_op [3], _06841_);
  nor (_06846_, _06845_, _06844_);
  and (_06847_, _06846_, _06843_);
  nor (_06848_, _06847_, _06840_);
  and (_06849_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], _06840_);
  not (_06850_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  and (_06851_, _06850_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  or (_06852_, _06851_, _06849_);
  and (_06853_, _06852_, _06847_);
  or (_06854_, _06853_, _06848_);
  and (_07572_, _06854_, _13707_);
  nor (_06855_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  not (_06856_, _06855_);
  and (_06857_, _06856_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12]);
  and (_06858_, _06856_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7]);
  not (_06859_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  not (_06860_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  not (_06861_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  nand (_06862_, _06861_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  or (_06863_, _06862_, _06860_);
  or (_06864_, _06863_, _06859_);
  not (_06865_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  or (_06866_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  or (_06867_, _06866_, _06860_);
  or (_06868_, _06867_, _06865_);
  and (_06869_, _06868_, _06864_);
  nor (_06870_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_06871_, _06870_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  nand (_06872_, _06871_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  not (_06873_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  or (_06874_, _06862_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  or (_06875_, _06874_, _06873_);
  and (_06876_, _06875_, _06872_);
  and (_06877_, _06876_, _06869_);
  not (_06878_, \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  and (_06879_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _06878_);
  or (_06880_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  not (_06881_, \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  or (_06882_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _06881_);
  and (_06883_, _06882_, _06880_);
  or (_06884_, _06883_, _06879_);
  nand (_06885_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _06878_);
  or (_06886_, _06885_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  nand (_06887_, _06886_, _06884_);
  or (_06888_, _06866_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  or (_06889_, _06888_, _06887_);
  and (_06890_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and (_06891_, _06890_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  nand (_06892_, _06891_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [4]);
  not (_06893_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nand (_06894_, _06890_, _06860_);
  or (_06895_, _06894_, _06893_);
  and (_06896_, _06895_, _06892_);
  and (_06897_, _06896_, _06889_);
  and (_06898_, _06897_, _06877_);
  not (_06899_, _06898_);
  not (_06900_, _06851_);
  or (_06901_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  or (_06902_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  or (_06903_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _06881_);
  and (_06904_, _06903_, _06902_);
  or (_06905_, _06904_, _06879_);
  or (_06906_, _06885_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  nand (_06907_, _06906_, _06905_);
  or (_06908_, _06907_, _06901_);
  not (_06909_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  nand (_06910_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  or (_06911_, _06910_, _06909_);
  not (_06912_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  not (_06913_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  nand (_06914_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], _06913_);
  or (_06915_, _06914_, _06912_);
  and (_06916_, _06915_, _06911_);
  and (_06917_, _06916_, _06908_);
  or (_06918_, _06917_, _06900_);
  not (_06919_, _06849_);
  or (_06920_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  or (_06921_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _06881_);
  and (_06922_, _06921_, _06920_);
  or (_06923_, _06922_, _06879_);
  or (_06924_, _06885_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  nand (_06925_, _06924_, _06923_);
  or (_06926_, _06925_, _06901_);
  not (_06927_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  or (_06928_, _06910_, _06927_);
  not (_06929_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or (_06930_, _06914_, _06929_);
  and (_06931_, _06930_, _06928_);
  and (_06932_, _06931_, _06926_);
  or (_06933_, _06932_, _06919_);
  and (_06934_, _06933_, _06918_);
  or (_06935_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  or (_06936_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _06881_);
  and (_06937_, _06936_, _06935_);
  or (_06938_, _06937_, _06879_);
  or (_06939_, _06885_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  nand (_06940_, _06939_, _06938_);
  or (_06941_, _06940_, _06901_);
  not (_06942_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  or (_06943_, _06910_, _06942_);
  not (_06944_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_06945_, _06914_, _06944_);
  and (_06946_, _06945_, _06943_);
  and (_06947_, _06946_, _06941_);
  or (_06948_, _06947_, _06852_);
  and (_06949_, _06948_, _06856_);
  nand (_06950_, _06949_, _06934_);
  or (_06951_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  or (_06952_, _06881_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [7]);
  and (_06953_, _06952_, _06951_);
  or (_06954_, _06953_, _06879_);
  or (_06955_, _06885_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  nand (_06956_, _06955_, _06954_);
  or (_06957_, _06956_, _06901_);
  not (_06958_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  nor (_06959_, _06910_, _06958_);
  not (_06960_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor (_06961_, _06914_, _06960_);
  nor (_06962_, _06961_, _06959_);
  and (_06963_, _06962_, _06957_);
  nand (_06964_, _06963_, _06855_);
  and (_06965_, _06964_, _06950_);
  and (_06966_, _06965_, _06899_);
  or (_06967_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  or (_06968_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _06881_);
  and (_06969_, _06968_, _06967_);
  or (_06970_, _06969_, _06879_);
  or (_06971_, _06885_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  nand (_06972_, _06971_, _06970_);
  or (_06973_, _06972_, _06901_);
  not (_06974_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  or (_06975_, _06910_, _06974_);
  not (_06976_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_06977_, _06914_, _06976_);
  and (_06978_, _06977_, _06975_);
  and (_06979_, _06978_, _06973_);
  or (_06980_, _06979_, _06900_);
  or (_06981_, _06887_, _06901_);
  or (_06982_, _06910_, _06873_);
  or (_06983_, _06914_, _06893_);
  and (_06984_, _06983_, _06982_);
  and (_06985_, _06984_, _06981_);
  or (_06986_, _06985_, _06919_);
  and (_06987_, _06986_, _06980_);
  or (_06988_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  or (_06989_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _06881_);
  and (_06990_, _06989_, _06988_);
  or (_06991_, _06990_, _06879_);
  or (_06992_, _06885_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  nand (_06993_, _06992_, _06991_);
  or (_06994_, _06993_, _06901_);
  not (_06995_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  or (_06996_, _06910_, _06995_);
  not (_06997_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_06998_, _06914_, _06997_);
  and (_06999_, _06998_, _06996_);
  and (_07000_, _06999_, _06994_);
  or (_07001_, _07000_, _06852_);
  and (_07002_, _07001_, _06856_);
  nand (_07003_, _07002_, _06987_);
  or (_07004_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  or (_07005_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _06881_);
  and (_07006_, _07005_, _07004_);
  or (_07007_, _07006_, _06879_);
  or (_07008_, _06885_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  nand (_07009_, _07008_, _07007_);
  or (_07010_, _07009_, _06901_);
  not (_07011_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  or (_07012_, _06910_, _07011_);
  not (_07013_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_07014_, _06914_, _07013_);
  and (_07015_, _07014_, _07012_);
  nand (_07016_, _07015_, _07010_);
  or (_07017_, _07016_, _06856_);
  and (_07018_, _07017_, _07003_);
  not (_07019_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  or (_07020_, _06863_, _07019_);
  not (_07021_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  or (_07022_, _06867_, _07021_);
  and (_07023_, _07022_, _07020_);
  nand (_07024_, _06871_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  or (_07025_, _06874_, _06909_);
  and (_07026_, _07025_, _07024_);
  and (_07027_, _07026_, _07023_);
  or (_07028_, _06907_, _06888_);
  nand (_07029_, _06891_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [3]);
  or (_07030_, _06894_, _06912_);
  and (_07031_, _07030_, _07029_);
  and (_07032_, _07031_, _07028_);
  and (_07033_, _07032_, _07027_);
  not (_07034_, _07033_);
  and (_07035_, _07034_, _07018_);
  and (_07036_, _07035_, _06966_);
  and (_07037_, _06899_, _07018_);
  not (_07038_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  or (_07039_, _06863_, _07038_);
  not (_07040_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  or (_07041_, _06867_, _07040_);
  and (_07042_, _07041_, _07039_);
  nand (_07043_, _06871_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  or (_07044_, _06874_, _06927_);
  and (_07045_, _07044_, _07043_);
  and (_07046_, _07045_, _07042_);
  or (_07047_, _06925_, _06888_);
  nand (_07048_, _06891_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [5]);
  or (_07049_, _06894_, _06929_);
  and (_07050_, _07049_, _07048_);
  and (_07051_, _07050_, _07047_);
  nand (_07052_, _07051_, _07046_);
  and (_07053_, _07052_, _06965_);
  nand (_07054_, _07053_, _07037_);
  and (_07055_, _07052_, _07018_);
  or (_07056_, _07055_, _06966_);
  and (_07057_, _07056_, _07054_);
  and (_07058_, _07057_, _07036_);
  and (_07059_, _07053_, _07037_);
  not (_07060_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  or (_07061_, _06863_, _07060_);
  not (_07062_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  or (_07063_, _06867_, _07062_);
  and (_07064_, _07063_, _07061_);
  nand (_07065_, _06871_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  or (_07066_, _06874_, _07011_);
  and (_07067_, _07066_, _07065_);
  and (_07068_, _07067_, _07064_);
  or (_07069_, _06888_, _07009_);
  nand (_07070_, _06891_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [6]);
  or (_07071_, _06894_, _07013_);
  and (_07072_, _07071_, _07070_);
  and (_07073_, _07072_, _07069_);
  and (_07074_, _07073_, _07068_);
  not (_07075_, _07074_);
  and (_07076_, _07075_, _07018_);
  or (_07077_, _07076_, _07059_);
  or (_07078_, _07074_, _07054_);
  and (_07079_, _07078_, _07077_);
  nand (_07080_, _07079_, _07053_);
  or (_07081_, _07076_, _07053_);
  and (_07082_, _07081_, _07080_);
  nand (_07083_, _07082_, _07058_);
  not (_07084_, _07083_);
  not (_07085_, _07078_);
  nand (_07086_, _06964_, _06950_);
  or (_07087_, _07074_, _07086_);
  nand (_07088_, _07017_, _07003_);
  or (_07089_, _06874_, _06958_);
  nand (_07090_, _06871_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  and (_07091_, _07090_, _07089_);
  not (_07092_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  or (_07093_, _06867_, _07092_);
  not (_07094_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  or (_07095_, _06863_, _07094_);
  and (_07096_, _07095_, _07093_);
  and (_07097_, _07096_, _07091_);
  or (_07098_, _06956_, _06888_);
  nand (_07099_, _06891_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [7]);
  or (_07100_, _06894_, _06960_);
  and (_07101_, _07100_, _07099_);
  and (_07102_, _07101_, _07098_);
  and (_07103_, _07102_, _07097_);
  or (_07104_, _07103_, _07088_);
  or (_07105_, _07104_, _07087_);
  nand (_07106_, _07104_, _07087_);
  and (_07107_, _07106_, _07105_);
  and (_07108_, _07107_, _07085_);
  not (_07109_, _07108_);
  and (_07110_, _07079_, _07053_);
  nand (_07111_, _07107_, _07110_);
  or (_07112_, _07107_, _07110_);
  nand (_07113_, _07112_, _07111_);
  nand (_07114_, _07113_, _07078_);
  and (_07115_, _07114_, _07109_);
  nand (_07116_, _07115_, _07084_);
  or (_07117_, _07115_, _07084_);
  nand (_07118_, _07117_, _07116_);
  not (_07119_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  or (_07120_, _06863_, _07119_);
  not (_07121_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  or (_07122_, _06867_, _07121_);
  and (_07123_, _07122_, _07120_);
  nand (_07124_, _06871_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  or (_07125_, _06874_, _06942_);
  and (_07126_, _07125_, _07124_);
  and (_07127_, _07126_, _07123_);
  or (_07128_, _06940_, _06888_);
  nand (_07129_, _06891_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [1]);
  or (_07130_, _06894_, _06944_);
  and (_07131_, _07130_, _07129_);
  and (_07132_, _07131_, _07128_);
  nand (_07133_, _07132_, _07127_);
  and (_07134_, _07133_, _06965_);
  nand (_07135_, _06891_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [2]);
  or (_07136_, _06894_, _06976_);
  and (_07137_, _07136_, _07135_);
  not (_07138_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  or (_07139_, _06863_, _07138_);
  not (_07140_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  or (_07141_, _06867_, _07140_);
  and (_07142_, _07141_, _07139_);
  and (_07143_, _07142_, _07137_);
  or (_07144_, _06888_, _06972_);
  or (_07145_, _06874_, _06974_);
  nand (_07146_, _06871_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  and (_07147_, _07146_, _07145_);
  and (_07148_, _07147_, _07144_);
  nand (_07149_, _07148_, _07143_);
  and (_07150_, _07149_, _07018_);
  and (_07151_, _07150_, _07134_);
  not (_07152_, _07151_);
  and (_07153_, _07133_, _07018_);
  not (_07154_, _07153_);
  and (_07155_, _07149_, _06965_);
  and (_07156_, _07155_, _07154_);
  nand (_07157_, _07156_, _07035_);
  nand (_07158_, _07157_, _07152_);
  not (_07159_, _07036_);
  and (_07160_, _07034_, _06965_);
  or (_07161_, _07160_, _07037_);
  and (_07162_, _07161_, _07159_);
  and (_07163_, _07162_, _07158_);
  not (_07164_, _07058_);
  or (_07165_, _07057_, _07036_);
  and (_07166_, _07165_, _07164_);
  and (_07167_, _07166_, _07163_);
  or (_07168_, _07082_, _07058_);
  and (_07169_, _07168_, _07083_);
  nand (_07170_, _07169_, _07167_);
  not (_07171_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor (_07172_, _06863_, _07171_);
  not (_07173_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor (_07174_, _06867_, _07173_);
  nor (_07175_, _07174_, _07172_);
  and (_07176_, _06871_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  nor (_07177_, _06874_, _06995_);
  nor (_07178_, _07177_, _07176_);
  and (_07179_, _07178_, _07175_);
  or (_07180_, _06888_, _06993_);
  nor (_07181_, _06894_, _06997_);
  and (_07182_, _06891_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [0]);
  nor (_07183_, _07182_, _07181_);
  and (_07184_, _07183_, _07180_);
  and (_07185_, _07184_, _07179_);
  not (_07186_, _07185_);
  and (_07187_, _07186_, _06965_);
  and (_07188_, _07187_, _07153_);
  or (_07189_, _07150_, _07134_);
  and (_07190_, _07189_, _07152_);
  and (_07191_, _07190_, _07188_);
  or (_07192_, _07156_, _07035_);
  and (_07193_, _07192_, _07157_);
  nand (_07194_, _07193_, _07191_);
  not (_07195_, _07194_);
  nand (_07196_, _07162_, _07158_);
  or (_07197_, _07162_, _07158_);
  and (_07198_, _07197_, _07196_);
  nand (_07199_, _07198_, _07195_);
  nand (_07200_, _07166_, _07163_);
  or (_07201_, _07166_, _07163_);
  nand (_07202_, _07201_, _07200_);
  or (_07203_, _07202_, _07199_);
  or (_07204_, _07169_, _07167_);
  nand (_07205_, _07204_, _07170_);
  or (_07206_, _07205_, _07203_);
  and (_07207_, _07206_, _07170_);
  or (_07208_, _07207_, _07118_);
  nand (_07209_, _07208_, _07116_);
  not (_07210_, _07103_);
  and (_07211_, _07210_, _06965_);
  and (_07212_, _07105_, _07211_);
  not (_07213_, _07212_);
  and (_07214_, _07109_, _07111_);
  nor (_07215_, _07214_, _07213_);
  and (_07216_, _07214_, _07213_);
  nor (_07217_, _07216_, _07215_);
  nand (_07218_, _07217_, _07209_);
  not (_07219_, _07215_);
  and (_07220_, _07219_, _07105_);
  nand (_07221_, _07220_, _07218_);
  nand (_07222_, _07221_, _06858_);
  or (_07223_, _07221_, _06858_);
  nand (_07224_, _07223_, _07222_);
  and (_07225_, _06856_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6]);
  or (_07226_, _07217_, _07209_);
  and (_07227_, _07226_, _07218_);
  nand (_07228_, _07227_, _07225_);
  or (_07229_, _07228_, _07224_);
  nand (_07230_, _07229_, _07222_);
  and (_07231_, _06856_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8]);
  and (_07232_, _06856_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  and (_07233_, _07232_, _07231_);
  and (_07234_, _07233_, _07230_);
  and (_07235_, _06856_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5]);
  nand (_07236_, _07207_, _07118_);
  and (_07237_, _07236_, _07208_);
  nand (_07238_, _07237_, _07235_);
  or (_07239_, _07237_, _07235_);
  nand (_07240_, _07239_, _07238_);
  and (_07241_, _06856_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4]);
  nand (_07242_, _07205_, _07203_);
  and (_07243_, _07242_, _07206_);
  nand (_07244_, _07243_, _07241_);
  or (_07245_, _07243_, _07241_);
  nand (_07246_, _07245_, _07244_);
  and (_07247_, _06856_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3]);
  nand (_07248_, _07202_, _07199_);
  and (_07249_, _07248_, _07203_);
  nand (_07250_, _07249_, _07247_);
  or (_07251_, _07249_, _07247_);
  nand (_07252_, _07251_, _07250_);
  and (_07253_, _06856_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2]);
  or (_07254_, _07198_, _07195_);
  and (_07255_, _07254_, _07199_);
  nand (_07256_, _07255_, _07253_);
  and (_07257_, _06856_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1]);
  or (_07258_, _07193_, _07191_);
  and (_07259_, _07258_, _07194_);
  nand (_07260_, _07259_, _07257_);
  and (_07261_, _06856_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0]);
  nand (_07262_, _07190_, _07188_);
  or (_07263_, _07190_, _07188_);
  and (_07264_, _07263_, _07262_);
  and (_07265_, _07264_, _07261_);
  not (_07266_, _07265_);
  or (_07267_, _07259_, _07257_);
  nand (_07268_, _07267_, _07260_);
  or (_07269_, _07268_, _07266_);
  and (_07270_, _07269_, _07260_);
  or (_07271_, _07255_, _07253_);
  nand (_07272_, _07271_, _07256_);
  or (_07273_, _07272_, _07270_);
  and (_07274_, _07273_, _07256_);
  or (_07275_, _07274_, _07252_);
  and (_07276_, _07275_, _07250_);
  or (_07277_, _07276_, _07246_);
  and (_07278_, _07277_, _07244_);
  or (_07279_, _07278_, _07240_);
  nand (_07280_, _07279_, _07238_);
  and (_07281_, _07223_, _07222_);
  or (_07282_, _07227_, _07225_);
  and (_07283_, _07282_, _07228_);
  and (_07284_, _07283_, _07281_);
  and (_07285_, _07233_, _07284_);
  and (_07286_, _07285_, _07280_);
  or (_07287_, _07286_, _07234_);
  and (_07288_, _06856_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10]);
  and (_07289_, _06856_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  and (_07291_, _07289_, _07288_);
  and (_07293_, _07291_, _07287_);
  nand (_07295_, _07293_, _06857_);
  nor (_07297_, _07295_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  not (_07299_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  nor (_07301_, _06855_, _07299_);
  and (_07302_, _07301_, _07295_);
  or (_07303_, _07302_, _07297_);
  and (_07759_, _07303_, _13707_);
  nor (_07304_, _06847_, _06850_);
  and (_07305_, _06847_, _06850_);
  or (_07306_, _07305_, _07304_);
  and (_02746_, _07306_, _13707_);
  and (_07307_, _07186_, _07018_);
  and (_02947_, _07307_, _13707_);
  nor (_07308_, _07187_, _07153_);
  nor (_07309_, _07308_, _07188_);
  and (_03159_, _07309_, _13707_);
  nor (_07310_, _07264_, _07261_);
  nor (_07311_, _07310_, _07265_);
  and (_03362_, _07311_, _13707_);
  and (_07312_, _07268_, _07266_);
  not (_07313_, _07312_);
  and (_07314_, _07313_, _07269_);
  and (_03563_, _07314_, _13707_);
  and (_07315_, _07272_, _07270_);
  not (_07316_, _07315_);
  and (_07317_, _07316_, _07273_);
  and (_03764_, _07317_, _13707_);
  and (_07318_, _07274_, _07252_);
  not (_07319_, _07318_);
  and (_07320_, _07319_, _07275_);
  and (_03957_, _07320_, _13707_);
  and (_07321_, _07276_, _07246_);
  not (_07322_, _07321_);
  and (_07323_, _07322_, _07277_);
  and (_04143_, _07323_, _13707_);
  and (_07324_, _07278_, _07240_);
  not (_07325_, _07324_);
  and (_07326_, _07325_, _07279_);
  and (_04316_, _07326_, _13707_);
  nand (_07327_, _07283_, _07280_);
  or (_07328_, _07283_, _07280_);
  and (_07329_, _07328_, _07327_);
  and (_04402_, _07329_, _13707_);
  and (_07330_, _07327_, _07228_);
  or (_07331_, _07330_, _07224_);
  nand (_07332_, _07330_, _07224_);
  and (_07333_, _07332_, _07331_);
  and (_04488_, _07333_, _13707_);
  nand (_07334_, _07331_, _07222_);
  nand (_07335_, _07334_, _07231_);
  or (_07336_, _07334_, _07231_);
  and (_07337_, _07336_, _07335_);
  and (_04574_, _07337_, _13707_);
  not (_07338_, _07232_);
  and (_07339_, _07338_, _07335_);
  nor (_07340_, _07339_, _07287_);
  and (_04659_, _07340_, _13707_);
  nand (_07341_, _07288_, _07287_);
  or (_07342_, _07288_, _07287_);
  and (_07343_, _07342_, _07341_);
  and (_04745_, _07343_, _13707_);
  not (_07344_, _07289_);
  and (_07345_, _07344_, _07341_);
  nor (_07346_, _07345_, _07293_);
  and (_04830_, _07346_, _13707_);
  or (_07347_, _07293_, _06857_);
  and (_07348_, _07347_, _07295_);
  and (_04921_, _07348_, _13707_);
  and (_07349_, \oc8051_top_1.oc8051_decoder1.alu_op [0], _06841_);
  nor (_07350_, _07349_, _06842_);
  not (_07351_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and (_07352_, _06844_, _07351_);
  and (_07353_, _07352_, _07350_);
  and (_07354_, _07353_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand (_07356_, _07354_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_07357_, _07354_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_07358_, _07357_, _07356_);
  and (_01017_, _07358_, _13707_);
  and (_01048_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _13707_);
  nor (_07359_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nand (_07360_, _07359_, _07103_);
  nor (_07361_, _07359_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7]);
  not (_07362_, _07361_);
  and (_07363_, _07362_, _07360_);
  nand (_07364_, _06946_, _06941_);
  or (_07365_, _07364_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  not (_07366_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand (_07367_, _06916_, _06908_);
  or (_07368_, _07367_, _07366_);
  and (_07369_, _07368_, _07365_);
  nor (_07370_, _07369_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nand (_07371_, _06931_, _06926_);
  or (_07372_, _07371_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand (_07373_, _06963_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand (_07374_, _07373_, _07372_);
  and (_07375_, _07374_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nor (_07376_, _07375_, _07370_);
  not (_07377_, _07376_);
  not (_07378_, _07016_);
  and (_07379_, _06963_, _07378_);
  nor (_07380_, _07379_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  not (_07381_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nand (_07382_, _06984_, _06981_);
  or (_07383_, _07382_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_07384_, _07016_, _07366_);
  and (_07385_, _07384_, _07383_);
  or (_07386_, _07367_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_07387_, _07371_, _07366_);
  and (_07388_, _07387_, _07386_);
  nor (_07389_, _07388_, _07385_);
  nand (_07390_, _06978_, _06973_);
  or (_07391_, _07390_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_07392_, _07382_, _07366_);
  and (_07393_, _07392_, _07391_);
  not (_07394_, _07393_);
  and (_07395_, _07374_, _07394_);
  nand (_07396_, _07395_, _07389_);
  and (_07397_, _07396_, _07381_);
  nor (_07398_, _07397_, _07380_);
  and (_07399_, _07398_, _07377_);
  nand (_07400_, _06999_, _06994_);
  or (_07401_, _07400_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_07402_, _07390_, _07366_);
  and (_07403_, _07402_, _07401_);
  or (_07404_, _07403_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_07405_, _07385_, _07381_);
  nand (_07406_, _07405_, _07404_);
  nand (_07407_, _07406_, _07363_);
  nor (_07408_, _07359_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6]);
  not (_07409_, _07408_);
  nand (_07410_, _07359_, _07074_);
  and (_07411_, _07410_, _07409_);
  and (_07412_, _07364_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_07413_, _07412_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_07414_, _07388_, _07381_);
  nand (_07415_, _07414_, _07413_);
  nand (_07416_, _07415_, _07411_);
  or (_07417_, _07406_, _07363_);
  nand (_07418_, _07417_, _07407_);
  or (_07419_, _07418_, _07416_);
  and (_07420_, _07419_, _07407_);
  not (_07421_, _07359_);
  or (_07422_, _07421_, _07052_);
  nor (_07423_, _07359_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5]);
  not (_07424_, _07423_);
  nand (_07425_, _07424_, _07422_);
  and (_07426_, _07400_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_07427_, _07426_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_07428_, _07393_, _07381_);
  and (_07429_, _07428_, _07427_);
  nor (_07430_, _07429_, _07425_);
  and (_07431_, _07369_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nand (_07432_, _07359_, _06898_);
  nor (_07433_, _07359_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4]);
  not (_07434_, _07433_);
  and (_07435_, _07434_, _07432_);
  not (_07436_, _07435_);
  or (_07437_, _07436_, _07431_);
  not (_07438_, _07437_);
  and (_07439_, _07429_, _07425_);
  nor (_07440_, _07439_, _07430_);
  and (_07441_, _07440_, _07438_);
  or (_07442_, _07441_, _07430_);
  or (_07443_, _07415_, _07411_);
  nand (_07444_, _07443_, _07416_);
  nor (_07445_, _07418_, _07444_);
  nand (_07446_, _07445_, _07442_);
  and (_07447_, _07446_, _07420_);
  and (_07448_, _07403_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nor (_07449_, _07359_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3]);
  not (_07450_, _07449_);
  nand (_07451_, _07359_, _07033_);
  and (_07452_, _07451_, _07450_);
  not (_07453_, _07452_);
  or (_07454_, _07453_, _07448_);
  not (_07455_, _07448_);
  or (_07456_, _07452_, _07455_);
  nand (_07457_, _07456_, _07454_);
  nand (_07458_, _07412_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nor (_07459_, _07359_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2]);
  not (_07460_, _07459_);
  or (_07461_, _07421_, _07149_);
  and (_07462_, _07461_, _07460_);
  nand (_07463_, _07462_, _07458_);
  and (_07464_, _07426_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_07465_, _07421_, _07133_);
  nor (_07466_, _07359_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1]);
  not (_07467_, _07466_);
  nand (_07468_, _07467_, _07465_);
  and (_07469_, _07468_, _07464_);
  or (_07470_, _07462_, _07458_);
  nand (_07471_, _07470_, _07463_);
  or (_07472_, _07471_, _07469_);
  and (_07473_, _07472_, _07463_);
  or (_07474_, _07473_, _07457_);
  nand (_07475_, _07474_, _07454_);
  not (_07476_, _07431_);
  or (_07477_, _07435_, _07476_);
  and (_07478_, _07477_, _07437_);
  and (_07479_, _07440_, _07478_);
  and (_07480_, _07445_, _07479_);
  nand (_07481_, _07480_, _07475_);
  nand (_07482_, _07481_, _07447_);
  nand (_07483_, _07482_, _07399_);
  and (_07484_, _07483_, _07363_);
  not (_07485_, _07416_);
  and (_07486_, _07478_, _07475_);
  nor (_07487_, _07486_, _07438_);
  nor (_07488_, _07487_, _07439_);
  nor (_07489_, _07488_, _07430_);
  nor (_07490_, _07489_, _07444_);
  nor (_07491_, _07490_, _07485_);
  not (_07492_, _07407_);
  and (_07493_, _07399_, _07492_);
  not (_07494_, _07493_);
  nor (_07495_, _07494_, _07491_);
  or (_07496_, _07495_, _07484_);
  nand (_07497_, _07496_, _07377_);
  or (_07498_, _07496_, _07377_);
  and (_07499_, _07489_, _07444_);
  nor (_07500_, _07499_, _07490_);
  nor (_07501_, _07500_, _07483_);
  and (_07502_, _07482_, _07399_);
  nor (_07503_, _07502_, _07411_);
  nor (_07504_, _07503_, _07501_);
  and (_07505_, _07504_, _07406_);
  nand (_07506_, _07505_, _07498_);
  and (_07507_, _07506_, _07497_);
  and (_07508_, _07498_, _07497_);
  nor (_07509_, _07504_, _07406_);
  nor (_07510_, _07509_, _07505_);
  and (_07511_, _07510_, _07508_);
  nor (_07512_, _07440_, _07487_);
  and (_07513_, _07440_, _07487_);
  or (_07514_, _07513_, _07512_);
  nor (_07515_, _07514_, _07483_);
  and (_07516_, _07483_, _07425_);
  nor (_07517_, _07516_, _07515_);
  and (_07518_, _07517_, _07415_);
  nand (_07519_, _07428_, _07427_);
  nor (_07520_, _07478_, _07475_);
  nor (_07521_, _07520_, _07486_);
  nor (_07522_, _07521_, _07483_);
  and (_07523_, _07483_, _07436_);
  nor (_07524_, _07523_, _07522_);
  and (_07526_, _07524_, _07519_);
  nor (_07528_, _07517_, _07415_);
  or (_07530_, _07528_, _07518_);
  not (_07532_, _07530_);
  and (_07534_, _07532_, _07526_);
  nor (_07536_, _07534_, _07518_);
  and (_07538_, _07473_, _07457_);
  not (_07539_, _07538_);
  and (_07540_, _07539_, _07474_);
  nor (_07541_, _07540_, _07483_);
  and (_07542_, _07483_, _07453_);
  nor (_07543_, _07542_, _07541_);
  and (_07544_, _07543_, _07476_);
  nor (_07545_, _07543_, _07476_);
  nor (_07546_, _07545_, _07544_);
  and (_07547_, _07471_, _07469_);
  not (_07548_, _07547_);
  and (_07549_, _07548_, _07472_);
  or (_07550_, _07549_, _07483_);
  or (_07551_, _07502_, _07462_);
  and (_07552_, _07551_, _07550_);
  nand (_07553_, _07552_, _07455_);
  not (_07554_, _07464_);
  or (_07555_, _07483_, _07554_);
  nand (_07556_, _07555_, _07468_);
  or (_07557_, _07555_, _07468_);
  and (_07558_, _07557_, _07556_);
  nand (_07559_, _07558_, _07458_);
  or (_07560_, _07558_, _07458_);
  and (_07561_, _07560_, _07559_);
  and (_07562_, _07359_, _07185_);
  nor (_07563_, _07359_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0]);
  nor (_07564_, _07563_, _07562_);
  nor (_07565_, _07564_, _07554_);
  not (_07566_, _07565_);
  nand (_07567_, _07566_, _07561_);
  and (_07568_, _07567_, _07559_);
  or (_07569_, _07552_, _07455_);
  nand (_07570_, _07569_, _07553_);
  or (_07571_, _07570_, _07568_);
  nand (_07573_, _07571_, _07553_);
  and (_07574_, _07573_, _07546_);
  or (_07575_, _07574_, _07544_);
  nor (_07576_, _07524_, _07519_);
  nor (_07577_, _07576_, _07526_);
  and (_07578_, _07532_, _07577_);
  nand (_07579_, _07578_, _07575_);
  nand (_07580_, _07579_, _07536_);
  nand (_07581_, _07580_, _07511_);
  nand (_07582_, _07581_, _07507_);
  and (_07583_, _07582_, _07398_);
  or (_07584_, _07583_, _07496_);
  not (_07585_, _07505_);
  nand (_07586_, _07580_, _07510_);
  and (_07587_, _07586_, _07585_);
  or (_07588_, _07587_, _07508_);
  nand (_07589_, _07587_, _07508_);
  and (_07590_, _07589_, _07588_);
  nand (_07591_, _07590_, _07583_);
  and (_07592_, _07591_, _07584_);
  and (_01069_, _07592_, _13707_);
  and (_03008_, _07583_, _13707_);
  and (_03019_, _07502_, _13707_);
  and (_03040_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _13707_);
  and (_03061_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _13707_);
  and (_03082_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _13707_);
  or (_07593_, _07353_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_07594_, _07354_, rst);
  and (_03093_, _07594_, _07593_);
  not (_07595_, _07564_);
  and (_07596_, _07583_, _07464_);
  nor (_07597_, _07596_, _07595_);
  and (_07598_, _07596_, _07595_);
  or (_07599_, _07598_, _07597_);
  and (_03104_, _07599_, _13707_);
  nand (_07600_, _07582_, _07398_);
  or (_07601_, _07566_, _07561_);
  and (_07602_, _07601_, _07567_);
  or (_07603_, _07602_, _07600_);
  or (_07604_, _07583_, _07558_);
  and (_07605_, _07604_, _07603_);
  and (_03115_, _07605_, _13707_);
  and (_07606_, _07570_, _07568_);
  not (_07607_, _07606_);
  and (_07608_, _07607_, _07571_);
  or (_07609_, _07608_, _07600_);
  or (_07610_, _07583_, _07552_);
  and (_07611_, _07610_, _07609_);
  and (_03126_, _07611_, _13707_);
  nor (_07612_, _07573_, _07546_);
  nor (_07613_, _07612_, _07574_);
  or (_07614_, _07613_, _07600_);
  or (_07615_, _07583_, _07543_);
  and (_07616_, _07615_, _07614_);
  and (_03137_, _07616_, _13707_);
  and (_07617_, _07577_, _07575_);
  nor (_07618_, _07577_, _07575_);
  or (_07619_, _07618_, _07617_);
  nand (_07620_, _07619_, _07583_);
  or (_07621_, _07583_, _07524_);
  and (_07622_, _07621_, _07620_);
  and (_03148_, _07622_, _13707_);
  nor (_07623_, _07617_, _07526_);
  nand (_07624_, _07530_, _07623_);
  or (_07625_, _07530_, _07623_);
  nand (_07626_, _07625_, _07624_);
  nand (_07627_, _07626_, _07583_);
  or (_07628_, _07583_, _07517_);
  and (_07629_, _07628_, _07627_);
  and (_03160_, _07629_, _13707_);
  or (_07630_, _07580_, _07510_);
  nand (_07631_, _07630_, _07586_);
  nand (_07632_, _07631_, _07583_);
  or (_07633_, _07583_, _07504_);
  and (_07634_, _07633_, _07632_);
  and (_03171_, _07634_, _13707_);
  and (_07635_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and (_07636_, _07635_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  and (_07637_, _07636_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  and (_07638_, _07637_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  and (_07639_, _07638_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  and (_07640_, _07639_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  not (_07641_, _07640_);
  not (_07642_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_07643_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _06841_);
  and (_07644_, _07643_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  and (_07645_, _07644_, _07642_);
  not (_07646_, _07645_);
  nor (_07647_, _07639_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor (_07648_, _07647_, _07646_);
  and (_07649_, _07648_, _07641_);
  not (_07650_, _07649_);
  and (_07651_, _07644_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  not (_07652_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  and (_07653_, _07643_, _07652_);
  and (_07654_, _07653_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_07655_, _07654_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [6]);
  nor (_07656_, _07655_, _07651_);
  not (_07657_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  and (_07658_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _06841_);
  and (_07659_, _07658_, _07642_);
  and (_07660_, _07659_, _07657_);
  and (_07661_, _07660_, \oc8051_top_1.oc8051_memory_interface1.ri_r [6]);
  and (_07662_, _07653_, _07642_);
  and (_07663_, _07662_, \oc8051_top_1.oc8051_memory_interface1.imm_r [6]);
  nor (_07664_, _07663_, _07661_);
  and (_07665_, _07664_, _07656_);
  and (_07666_, _07665_, _07650_);
  nor (_07667_, _07638_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  not (_07668_, _07667_);
  nor (_07669_, _07646_, _07639_);
  and (_07670_, _07669_, _07668_);
  not (_07671_, _07670_);
  and (_07672_, _07662_, \oc8051_top_1.oc8051_memory_interface1.imm_r [5]);
  nor (_07673_, _07672_, _07651_);
  and (_07674_, _07660_, \oc8051_top_1.oc8051_memory_interface1.ri_r [5]);
  and (_07675_, _07654_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [5]);
  nor (_07676_, _07675_, _07674_);
  and (_07677_, _07676_, _07673_);
  and (_07678_, _07677_, _07671_);
  nor (_07679_, _07678_, _07666_);
  not (_07680_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  nor (_07681_, _07640_, _07680_);
  and (_07682_, _07640_, _07680_);
  nor (_07683_, _07682_, _07681_);
  nor (_07684_, _07683_, _07646_);
  not (_07685_, _07684_);
  and (_07686_, _07660_, \oc8051_top_1.oc8051_memory_interface1.ri_r [7]);
  not (_07687_, _07686_);
  not (_07688_, _07651_);
  and (_07689_, _07662_, \oc8051_top_1.oc8051_memory_interface1.imm_r [7]);
  and (_07690_, _07654_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [7]);
  nor (_07691_, _07690_, _07689_);
  and (_07692_, _07691_, _07688_);
  and (_07693_, _07692_, _07687_);
  and (_07694_, _07693_, _07685_);
  not (_07695_, _07694_);
  and (_07696_, _07654_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [3]);
  and (_07697_, _07662_, \oc8051_top_1.oc8051_memory_interface1.imm_r [3]);
  nor (_07698_, _07697_, _07696_);
  not (_07699_, _07637_);
  nor (_07700_, _07636_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor (_07701_, _07700_, _07646_);
  and (_07702_, _07701_, _07699_);
  or (_07703_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_07704_, _07703_, _06841_);
  nor (_07705_, _07704_, _07643_);
  and (_07706_, _07705_, \oc8051_top_1.oc8051_memory_interface1.rn_r [3]);
  and (_07707_, _07660_, \oc8051_top_1.oc8051_memory_interface1.ri_r [3]);
  nor (_07708_, _07707_, _07706_);
  not (_07709_, _07708_);
  nor (_07710_, _07709_, _07702_);
  and (_07711_, _07710_, _07698_);
  nor (_07712_, _07637_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  or (_07713_, _07712_, _07646_);
  nor (_07714_, _07713_, _07638_);
  and (_07715_, _07654_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [4]);
  nor (_07716_, _07715_, _07714_);
  and (_07717_, _07705_, \oc8051_top_1.oc8051_memory_interface1.rn_r [4]);
  and (_07718_, _07662_, \oc8051_top_1.oc8051_memory_interface1.imm_r [4]);
  nor (_07719_, _07718_, _07717_);
  and (_07720_, _07660_, \oc8051_top_1.oc8051_memory_interface1.ri_r [4]);
  nor (_07721_, _07720_, _07651_);
  and (_07722_, _07721_, _07719_);
  and (_07723_, _07722_, _07716_);
  not (_07724_, _07723_);
  and (_07725_, _07724_, _07711_);
  and (_07726_, _07725_, _07695_);
  and (_07727_, _07726_, _07679_);
  and (_07728_, _07654_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [0]);
  and (_07729_, _07662_, \oc8051_top_1.oc8051_memory_interface1.imm_r [0]);
  nor (_07730_, _07729_, _07728_);
  and (_07731_, _07660_, \oc8051_top_1.oc8051_memory_interface1.ri_r [0]);
  not (_07732_, _07731_);
  not (_07733_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and (_07734_, _07645_, _07733_);
  and (_07735_, _07705_, \oc8051_top_1.oc8051_memory_interface1.rn_r [0]);
  nor (_07736_, _07735_, _07734_);
  and (_07737_, _07736_, _07732_);
  and (_07738_, _07737_, _07730_);
  nor (_07739_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  nor (_07740_, _07739_, _07635_);
  and (_07741_, _07740_, _07645_);
  and (_07742_, _07660_, \oc8051_top_1.oc8051_memory_interface1.ri_r [1]);
  nor (_07743_, _07742_, _07741_);
  and (_07744_, _07654_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [1]);
  and (_07745_, _07662_, \oc8051_top_1.oc8051_memory_interface1.imm_r [1]);
  and (_07746_, _07705_, \oc8051_top_1.oc8051_memory_interface1.rn_r [1]);
  or (_07747_, _07746_, _07745_);
  nor (_07748_, _07747_, _07744_);
  and (_07749_, _07748_, _07743_);
  nor (_07750_, _07635_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_07751_, _07750_, _07636_);
  and (_07752_, _07751_, _07645_);
  and (_07753_, _07660_, \oc8051_top_1.oc8051_memory_interface1.ri_r [2]);
  nor (_07754_, _07753_, _07752_);
  and (_07755_, _07654_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [2]);
  and (_07756_, _07662_, \oc8051_top_1.oc8051_memory_interface1.imm_r [2]);
  and (_07757_, _07705_, \oc8051_top_1.oc8051_memory_interface1.rn_r [2]);
  or (_07758_, _07757_, _07756_);
  nor (_07760_, _07758_, _07755_);
  and (_07761_, _07760_, _07754_);
  and (_07762_, _07761_, _07749_);
  and (_07763_, _07762_, _07738_);
  nand (_07764_, _07763_, _07727_);
  nand (_07765_, _07592_, _07353_);
  nand (_07766_, _07303_, _06847_);
  not (_07767_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_07768_, _06842_, _07767_);
  and (_07769_, _07768_, _06846_);
  not (_07770_, _07769_);
  nor (_07771_, _07103_, _06963_);
  and (_07772_, _07103_, _06963_);
  nor (_07773_, _07772_, _07771_);
  nor (_07774_, _07074_, _07016_);
  nor (_07775_, _07074_, _07378_);
  and (_07776_, _07074_, _07378_);
  nor (_07777_, _07776_, _07775_);
  and (_07778_, _07052_, _06932_);
  and (_07779_, _07052_, _07371_);
  nor (_07780_, _07052_, _07371_);
  nor (_07781_, _07780_, _07779_);
  and (_07782_, _06898_, _07382_);
  nor (_07783_, _07782_, _07781_);
  nor (_07784_, _07783_, _07778_);
  nor (_07785_, _07784_, _07777_);
  nor (_07786_, _07785_, _07774_);
  and (_07787_, _07784_, _07777_);
  nor (_07788_, _07787_, _07785_);
  not (_07789_, _07788_);
  and (_07790_, _07782_, _07781_);
  nor (_07791_, _07790_, _07783_);
  not (_07792_, _07791_);
  nor (_07793_, _06898_, _06985_);
  and (_07794_, _06898_, _06985_);
  nor (_07795_, _07794_, _07793_);
  not (_07796_, _07795_);
  and (_07797_, _07033_, _06917_);
  nor (_07798_, _07033_, _06917_);
  nor (_07799_, _07798_, _07797_);
  and (_07800_, _07149_, _07390_);
  nor (_07801_, _07149_, _07390_);
  nor (_07802_, _07801_, _07800_);
  and (_07803_, _07133_, _07364_);
  nor (_07804_, _07133_, _07364_);
  nor (_07805_, _07804_, _07803_);
  and (_07806_, _07185_, _07400_);
  nor (_07807_, _07806_, _07805_);
  and (_07808_, _07133_, _06947_);
  nor (_07809_, _07808_, _07807_);
  nor (_07810_, _07809_, _07802_);
  and (_07811_, _07149_, _06979_);
  nor (_07812_, _07811_, _07810_);
  nor (_07813_, _07812_, _07799_);
  and (_07814_, _07812_, _07799_);
  nor (_07815_, _07814_, _07813_);
  not (_07816_, _07815_);
  and (_07817_, _07809_, _07802_);
  nor (_07818_, _07817_, _07810_);
  not (_07819_, _07818_);
  and (_07820_, _07806_, _07805_);
  nor (_07821_, _07820_, _07807_);
  not (_07822_, _07821_);
  nor (_07823_, _07185_, _07000_);
  and (_07824_, _07185_, _07000_);
  nor (_07825_, _07824_, _07823_);
  nor (_07826_, _06885_, \oc8051_top_1.oc8051_sfr1.bit_out );
  not (_07827_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_07828_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_07829_, _07828_, _06953_);
  nor (_07830_, _07829_, _07827_);
  nor (_07831_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_07832_, _07831_, _06883_);
  not (_07833_, _07832_);
  not (_07834_, \oc8051_top_1.oc8051_ram_top1.bit_select [0]);
  and (_07835_, _07834_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_07836_, _07835_, _07006_);
  not (_07837_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_07838_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], _07837_);
  and (_07839_, _07838_, _06922_);
  nor (_07840_, _07839_, _07836_);
  and (_07841_, _07840_, _07833_);
  and (_07842_, _07841_, _07830_);
  and (_07843_, _07828_, _06904_);
  nor (_07844_, _07843_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_07845_, _07838_, _06937_);
  not (_07846_, _07845_);
  and (_07847_, _07835_, _06969_);
  and (_07848_, _07831_, _06990_);
  nor (_07849_, _07848_, _07847_);
  and (_07850_, _07849_, _07846_);
  and (_07851_, _07850_, _07844_);
  nor (_07852_, _07851_, _07842_);
  nor (_07853_, _07852_, _06879_);
  nor (_07854_, _07853_, _07826_);
  and (_07855_, \oc8051_top_1.oc8051_decoder1.cy_sel [0], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_07856_, _07855_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  not (_07857_, _07856_);
  and (_07858_, _07857_, _07854_);
  and (_07859_, _07857_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  nor (_07860_, _07859_, _07858_);
  nor (_07861_, _07860_, _07825_);
  and (_07862_, _07861_, _07822_);
  and (_07863_, _07862_, _07819_);
  and (_07864_, _07863_, _07816_);
  or (_07865_, _07033_, _07367_);
  and (_07866_, _07033_, _07367_);
  or (_07867_, _07812_, _07866_);
  and (_07868_, _07867_, _07865_);
  or (_07869_, _07868_, _07864_);
  and (_07870_, _07869_, _07796_);
  and (_07871_, _07870_, _07792_);
  and (_07872_, _07871_, _07789_);
  nor (_07873_, _07872_, _07786_);
  nor (_07874_, _07873_, _07773_);
  and (_07875_, _07873_, _07773_);
  nor (_07876_, _07875_, _07874_);
  nor (_07877_, _07876_, _07770_);
  not (_07878_, _07877_);
  not (_07879_, _07773_);
  not (_07880_, _07802_);
  and (_07881_, _07823_, _07805_);
  nor (_07882_, _07881_, _07803_);
  nor (_07883_, _07882_, _07880_);
  nor (_07884_, _07883_, _07800_);
  nor (_07885_, _07884_, _07799_);
  and (_07886_, _07884_, _07799_);
  nor (_07887_, _07886_, _07885_);
  not (_07888_, _07825_);
  nor (_07889_, _07860_, _07888_);
  and (_07890_, _07889_, _07805_);
  and (_07891_, _07882_, _07880_);
  nor (_07892_, _07891_, _07883_);
  and (_07893_, _07892_, _07890_);
  not (_07894_, _07893_);
  nor (_07895_, _07894_, _07887_);
  nor (_07896_, _07884_, _07797_);
  or (_07897_, _07896_, _07798_);
  or (_07898_, _07897_, _07895_);
  and (_07899_, _07898_, _07795_);
  and (_07900_, _07899_, _07781_);
  not (_07901_, _07777_);
  and (_07902_, _07793_, _07781_);
  nor (_07903_, _07902_, _07779_);
  nor (_07904_, _07903_, _07901_);
  and (_07905_, _07903_, _07901_);
  nor (_07906_, _07905_, _07904_);
  and (_07907_, _07906_, _07900_);
  nor (_07908_, _07904_, _07775_);
  not (_07909_, _07908_);
  nor (_07910_, _07909_, _07907_);
  and (_07911_, _07910_, _07879_);
  nor (_07912_, _07910_, _07879_);
  not (_07913_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  and (_07914_, _07349_, _07913_);
  and (_07915_, _07914_, _06846_);
  not (_07916_, _07915_);
  or (_07917_, _07916_, _07912_);
  nor (_07918_, _07917_, _07911_);
  not (_07919_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and (_07920_, _06845_, _07919_);
  and (_07921_, _07920_, _07914_);
  not (_07922_, _07921_);
  nor (_07923_, _07922_, _07772_);
  and (_07924_, _07920_, _07350_);
  and (_07925_, _07924_, _07773_);
  nor (_07926_, _07925_, _07923_);
  and (_07927_, _06845_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and (_07928_, _07927_, _07350_);
  and (_07929_, _07928_, _07186_);
  and (_07930_, _07920_, _06842_);
  and (_07931_, _07930_, _07075_);
  nor (_07932_, _07931_, _07929_);
  not (_07933_, _07860_);
  and (_07934_, _07927_, _07914_);
  and (_07935_, _07934_, _07933_);
  and (_07936_, _07352_, _06843_);
  and (_07937_, _07936_, _07771_);
  and (_07938_, _07768_, _07352_);
  and (_07939_, _07938_, _07103_);
  nor (_07940_, _07939_, _07937_);
  and (_07941_, _07350_, _06846_);
  not (_07942_, _07941_);
  nor (_07943_, _07942_, _07103_);
  not (_07944_, _07943_);
  nand (_07945_, _07944_, _07940_);
  nor (_07946_, _07945_, _07935_);
  and (_07947_, _07946_, _07932_);
  and (_07948_, _07927_, _07768_);
  and (_07949_, _07186_, _07133_);
  and (_07950_, _07949_, _07149_);
  and (_07951_, _07950_, _07034_);
  and (_07952_, _07951_, _06899_);
  and (_07953_, _07952_, _07052_);
  and (_07954_, _07953_, _07075_);
  and (_07955_, _07954_, _07860_);
  not (_07956_, _07052_);
  and (_07957_, _07074_, _07956_);
  nor (_07958_, _07149_, _07133_);
  and (_07959_, _07958_, _07185_);
  and (_07960_, _07959_, _07033_);
  and (_07961_, _07960_, _06898_);
  and (_07962_, _07961_, _07957_);
  and (_07963_, _07962_, _07933_);
  nor (_07964_, _07963_, _07955_);
  and (_07965_, _07964_, _07103_);
  nor (_07966_, _07964_, _07103_);
  nor (_07967_, _07966_, _07965_);
  and (_07968_, _07967_, _07948_);
  not (_07969_, _06963_);
  nor (_07970_, _07860_, _07969_);
  not (_07971_, _07970_);
  and (_07972_, _07860_, _07103_);
  and (_07973_, _07927_, _06843_);
  not (_07974_, _07973_);
  nor (_07975_, _07974_, _07972_);
  and (_07976_, _07975_, _07971_);
  nor (_07977_, _07976_, _07968_);
  and (_07978_, _07914_, _07352_);
  not (_07979_, _07978_);
  not (_07980_, _07957_);
  nor (_07981_, _07958_, _07033_);
  and (_07982_, _07981_, _07978_);
  and (_07983_, _07982_, _06899_);
  nor (_07984_, _07983_, _07980_);
  nor (_07985_, _07957_, _07103_);
  nor (_07986_, _07985_, _07982_);
  and (_07987_, _07986_, _07860_);
  nor (_07988_, _07987_, _07984_);
  and (_07989_, _07988_, _07103_);
  nor (_07990_, _07988_, _07103_);
  nor (_07991_, _07990_, _07989_);
  nor (_07992_, _07991_, _07979_);
  not (_07993_, _07992_);
  and (_07994_, _07993_, _07977_);
  and (_07995_, _07994_, _07947_);
  and (_07996_, _07995_, _07926_);
  not (_07997_, _07996_);
  nor (_07998_, _07997_, _07918_);
  and (_07999_, _07998_, _07878_);
  and (_08000_, _07999_, _07766_);
  and (_08001_, _08000_, _07765_);
  not (_08002_, _08001_);
  or (_08003_, _08002_, _07764_);
  not (_08004_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_08005_, \oc8051_top_1.oc8051_decoder1.wr , _06841_);
  not (_08006_, _08005_);
  nor (_08007_, _08006_, _07659_);
  and (_08008_, _08007_, _08004_);
  not (_08009_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  nand (_08010_, _07764_, _08009_);
  and (_08011_, _08010_, _08008_);
  and (_08012_, _08011_, _08003_);
  nor (_08013_, _08007_, _08009_);
  nor (_08014_, _07912_, _07771_);
  nor (_08015_, _08014_, _07916_);
  not (_08016_, _08015_);
  and (_08017_, _07103_, _07969_);
  nor (_08018_, _08017_, _07874_);
  nor (_08019_, _08018_, _07770_);
  and (_08020_, _07984_, _07860_);
  nor (_08021_, _08020_, _07972_);
  not (_08022_, _07984_);
  nor (_08023_, _07860_, _07103_);
  and (_08024_, _08023_, _08022_);
  nor (_08025_, _08024_, _07979_);
  and (_08026_, _08025_, _08021_);
  not (_08027_, _08026_);
  nor (_08028_, _07942_, _07860_);
  not (_08029_, _08028_);
  and (_08030_, _07920_, _06843_);
  not (_08031_, _08030_);
  nor (_08032_, _08031_, _07103_);
  not (_08033_, _08032_);
  and (_08034_, _07934_, _07186_);
  nor (_08035_, _08034_, _07982_);
  and (_08036_, _08035_, _08033_);
  and (_08037_, _08036_, _08029_);
  nor (_08038_, _07859_, _07854_);
  not (_08039_, _07924_);
  nor (_08040_, _08039_, _07858_);
  nor (_08041_, _08040_, _07921_);
  or (_08042_, _08041_, _08038_);
  and (_08043_, _07856_, _07854_);
  and (_08044_, _07920_, _07768_);
  and (_08045_, _07936_, _07854_);
  nor (_08046_, _08045_, _08044_);
  nor (_08047_, _08046_, _08043_);
  and (_08048_, _07938_, _07860_);
  not (_08049_, _07928_);
  nor (_08050_, _08049_, _07854_);
  and (_08051_, _08050_, _07933_);
  or (_08052_, _08051_, _08048_);
  nor (_08053_, _08052_, _08047_);
  and (_08054_, _08053_, _08042_);
  and (_08055_, _08054_, _08037_);
  and (_08056_, _08055_, _08027_);
  not (_08057_, _08056_);
  nor (_08058_, _08057_, _08019_);
  and (_08059_, _08058_, _08016_);
  not (_08060_, _07738_);
  nor (_08061_, _07761_, _07749_);
  and (_08062_, _08061_, _08060_);
  and (_08063_, _08062_, _07727_);
  nand (_08064_, _08063_, _08059_);
  and (_08065_, _08007_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  or (_08066_, _08063_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_08067_, _08066_, _08065_);
  and (_08068_, _08067_, _08064_);
  or (_08069_, _08068_, _08013_);
  or (_08070_, _08069_, _08012_);
  and (_06303_, _08070_, _13707_);
  nand (_08071_, _07599_, _07353_);
  and (_08072_, _07329_, _06847_);
  and (_08073_, _07860_, _07888_);
  nor (_08074_, _08073_, _07889_);
  nor (_08075_, _07915_, _07769_);
  not (_08076_, _08075_);
  and (_08077_, _08076_, _08074_);
  not (_08078_, _08077_);
  nor (_08079_, _08031_, _07860_);
  not (_08080_, _08079_);
  nor (_08081_, _08039_, _07823_);
  nor (_08082_, _08081_, _07921_);
  or (_08083_, _08082_, _07824_);
  and (_08084_, _07936_, _07823_);
  and (_08085_, _07938_, _07185_);
  nor (_08086_, _08085_, _08084_);
  and (_08087_, _07973_, _07400_);
  and (_08088_, _07948_, _07185_);
  nor (_08089_, _08088_, _08087_);
  and (_08090_, _07927_, _07913_);
  and (_08091_, _08090_, _07133_);
  and (_08092_, _08044_, _07210_);
  nor (_08093_, _08092_, _08091_);
  or (_08094_, _07941_, _07978_);
  and (_08095_, _08094_, _07186_);
  not (_08096_, _08095_);
  and (_08097_, _08096_, _08093_);
  and (_08098_, _08097_, _08089_);
  and (_08099_, _08098_, _08086_);
  and (_08100_, _08099_, _08083_);
  and (_08101_, _08100_, _08080_);
  and (_08102_, _08101_, _08078_);
  not (_08103_, _08102_);
  nor (_08104_, _08103_, _08072_);
  and (_08105_, _08104_, _08071_);
  not (_08106_, _08105_);
  or (_08107_, _08106_, _07764_);
  not (_08108_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nand (_08109_, _07764_, _08108_);
  and (_08110_, _08109_, _08008_);
  and (_08111_, _08110_, _08107_);
  nor (_08112_, _08007_, _08108_);
  not (_08113_, _08059_);
  or (_08114_, _08113_, _07764_);
  and (_08115_, _08109_, _08065_);
  and (_08116_, _08115_, _08114_);
  or (_08117_, _08116_, _08112_);
  or (_08118_, _08117_, _08111_);
  and (_06807_, _08118_, _13707_);
  nand (_08119_, _07605_, _07353_);
  nand (_08120_, _07333_, _06847_);
  nor (_08121_, _07823_, _07805_);
  or (_08122_, _08121_, _07881_);
  and (_08123_, _08122_, _07889_);
  nor (_08124_, _08122_, _07889_);
  or (_08125_, _08124_, _08123_);
  and (_08126_, _08125_, _07915_);
  nor (_08127_, _07861_, _07822_);
  nor (_08128_, _08127_, _07862_);
  nor (_08129_, _08128_, _07770_);
  nor (_08130_, _08129_, _08126_);
  and (_08131_, _07973_, _07364_);
  not (_08132_, _07133_);
  and (_08133_, _07185_, _08132_);
  nor (_08134_, _08133_, _07949_);
  not (_08135_, _08134_);
  nor (_08136_, _08135_, _07860_);
  and (_08137_, _08135_, _07860_);
  nor (_08138_, _08137_, _08136_);
  and (_08139_, _08138_, _07948_);
  nor (_08140_, _08139_, _08131_);
  nor (_08141_, _07981_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_08142_, _08141_, _07133_);
  nor (_08143_, _08141_, _07133_);
  nor (_08144_, _08143_, _08142_);
  nor (_08145_, _08144_, _07979_);
  not (_08146_, _08145_);
  and (_08147_, _07924_, _07805_);
  nor (_08148_, _07922_, _07804_);
  not (_08149_, _08148_);
  and (_08150_, _07936_, _07803_);
  and (_08151_, _07938_, _08132_);
  nor (_08152_, _08151_, _08150_);
  nand (_08153_, _08152_, _08149_);
  nor (_08154_, _08153_, _08147_);
  and (_08155_, _07941_, _07133_);
  not (_08156_, _08155_);
  and (_08157_, _08090_, _07149_);
  and (_08158_, _07930_, _07186_);
  nor (_08159_, _08158_, _08157_);
  and (_08160_, _08159_, _08156_);
  and (_08161_, _08160_, _08154_);
  and (_08162_, _08161_, _08146_);
  and (_08163_, _08162_, _08140_);
  and (_08164_, _08163_, _08130_);
  and (_08165_, _08164_, _08120_);
  nand (_08166_, _08165_, _08119_);
  or (_08167_, _08166_, _07764_);
  not (_08168_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  nand (_08169_, _07764_, _08168_);
  and (_08170_, _08169_, _08008_);
  and (_08171_, _08170_, _08167_);
  nor (_08172_, _08007_, _08168_);
  and (_08173_, _07762_, _08060_);
  and (_08174_, _08173_, _07727_);
  or (_08175_, _08174_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_08176_, _08175_, _08065_);
  nand (_08177_, _08174_, _08059_);
  and (_08178_, _08177_, _08176_);
  or (_08179_, _08178_, _08172_);
  or (_08180_, _08179_, _08171_);
  and (_06808_, _08180_, _13707_);
  nand (_08181_, _07337_, _06847_);
  nand (_08182_, _07611_, _07353_);
  and (_08183_, _07973_, _07390_);
  not (_08184_, _07149_);
  and (_08185_, _08133_, _07933_);
  and (_08186_, _07949_, _07860_);
  nor (_08187_, _08186_, _08185_);
  nor (_08188_, _08187_, _08184_);
  not (_08189_, _07948_);
  and (_08190_, _08187_, _08184_);
  or (_08191_, _08190_, _08189_);
  nor (_08192_, _08191_, _08188_);
  nor (_08193_, _08192_, _08183_);
  nor (_08194_, _07862_, _07819_);
  nor (_08195_, _08194_, _07863_);
  nor (_08196_, _08195_, _07770_);
  not (_08197_, _08196_);
  and (_08198_, _08090_, _07034_);
  and (_08199_, _07936_, _07800_);
  and (_08200_, _07938_, _08184_);
  nor (_08201_, _08200_, _08199_);
  nor (_08202_, _07922_, _07801_);
  and (_08203_, _07924_, _07802_);
  nor (_08204_, _08203_, _08202_);
  and (_08205_, _07930_, _07133_);
  and (_08206_, _07941_, _07149_);
  nor (_08207_, _08206_, _08205_);
  and (_08208_, _08207_, _08204_);
  nand (_08209_, _08208_, _08201_);
  nor (_08210_, _08209_, _08198_);
  and (_08211_, _08210_, _08197_);
  nor (_08212_, _07892_, _07890_);
  nor (_08213_, _08212_, _07916_);
  and (_08214_, _08213_, _07894_);
  nor (_08215_, _08143_, _08184_);
  and (_08216_, _07958_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_08217_, _08216_, _08215_);
  nor (_08218_, _08217_, _07979_);
  nor (_08219_, _08218_, _08214_);
  and (_08220_, _08219_, _08211_);
  and (_08221_, _08220_, _08193_);
  and (_08222_, _08221_, _08182_);
  and (_08223_, _08222_, _08181_);
  not (_08224_, _08223_);
  or (_08225_, _08224_, _07764_);
  not (_08226_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  nand (_08227_, _07764_, _08226_);
  and (_08228_, _08227_, _08008_);
  and (_08229_, _08228_, _08225_);
  nor (_08230_, _08007_, _08226_);
  nand (_08231_, _07761_, _07727_);
  nor (_08232_, _07749_, _07738_);
  or (_08233_, _08232_, _08231_);
  and (_08234_, _08233_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  not (_08235_, _07749_);
  and (_08236_, _07761_, _08235_);
  and (_08237_, _08236_, _07738_);
  and (_08238_, _08237_, _08113_);
  and (_08239_, _07762_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or (_08240_, _08239_, _08238_);
  and (_08241_, _08240_, _07727_);
  or (_08242_, _08241_, _08234_);
  and (_08243_, _08242_, _08065_);
  or (_08244_, _08243_, _08230_);
  or (_08245_, _08244_, _08229_);
  and (_06809_, _08245_, _13707_);
  nand (_08246_, _07340_, _06847_);
  nand (_08247_, _07616_, _07353_);
  nor (_08248_, _07863_, _07816_);
  nor (_08249_, _08248_, _07864_);
  nor (_08250_, _08249_, _07770_);
  not (_08251_, _08250_);
  and (_08252_, _07936_, _07798_);
  and (_08253_, _07938_, _07033_);
  nor (_08254_, _08253_, _08252_);
  and (_08255_, _08090_, _06899_);
  and (_08256_, _07930_, _07149_);
  nor (_08257_, _07942_, _07033_);
  or (_08258_, _08257_, _08256_);
  nor (_08259_, _08258_, _08255_);
  and (_08260_, _08259_, _08254_);
  and (_08261_, _07894_, _07887_);
  or (_08262_, _08261_, _07916_);
  nor (_08263_, _08262_, _07895_);
  and (_08264_, _07973_, _07367_);
  nor (_08265_, _07959_, _07860_);
  nor (_08266_, _07950_, _07933_);
  nor (_08267_, _08266_, _08265_);
  and (_08268_, _08267_, _07034_);
  nor (_08269_, _08267_, _07034_);
  or (_08270_, _08269_, _08189_);
  nor (_08271_, _08270_, _08268_);
  nor (_08272_, _08271_, _08264_);
  not (_08273_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_08274_, _07958_, _08273_);
  nor (_08275_, _08274_, _07034_);
  or (_08276_, _08275_, _07979_);
  nor (_08277_, _08276_, _07981_);
  not (_08278_, _08277_);
  nor (_08279_, _07922_, _07797_);
  and (_08280_, _07924_, _07799_);
  nor (_08281_, _08280_, _08279_);
  and (_08282_, _08281_, _08278_);
  nand (_08283_, _08282_, _08272_);
  nor (_08284_, _08283_, _08263_);
  and (_08285_, _08284_, _08260_);
  and (_08286_, _08285_, _08251_);
  and (_08287_, _08286_, _08247_);
  nand (_08288_, _08287_, _08246_);
  or (_08289_, _08288_, _07764_);
  not (_08290_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nand (_08291_, _07764_, _08290_);
  and (_08292_, _08291_, _08008_);
  and (_08293_, _08292_, _08289_);
  nor (_08294_, _08007_, _08290_);
  and (_08295_, _08231_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_08296_, _08232_, _07761_);
  not (_08297_, _08296_);
  nor (_08298_, _08297_, _08059_);
  not (_08299_, _07761_);
  or (_08300_, _08232_, _08299_);
  nor (_08301_, _08300_, _08290_);
  or (_08302_, _08301_, _08298_);
  and (_08303_, _08302_, _07727_);
  or (_08304_, _08303_, _08295_);
  and (_08305_, _08304_, _08065_);
  or (_08306_, _08305_, _08294_);
  or (_08307_, _08306_, _08293_);
  and (_06810_, _08307_, _13707_);
  nand (_08308_, _07622_, _07353_);
  nand (_08309_, _07343_, _06847_);
  nor (_08310_, _07869_, _07795_);
  and (_08311_, _07869_, _07795_);
  nor (_08312_, _08311_, _08310_);
  and (_08313_, _08312_, _07769_);
  not (_08314_, _08313_);
  nor (_08315_, _07898_, _07795_);
  nor (_08316_, _08315_, _07899_);
  and (_08317_, _08316_, _07915_);
  and (_08318_, _07860_, _06899_);
  nor (_08319_, _07860_, _06985_);
  or (_08320_, _08319_, _08318_);
  and (_08321_, _08320_, _07973_);
  and (_08322_, _07951_, _07860_);
  and (_08323_, _07960_, _07933_);
  nor (_08324_, _08323_, _08322_);
  nor (_08325_, _08324_, _06898_);
  not (_08326_, _08325_);
  and (_08327_, _08324_, _06898_);
  nor (_08328_, _08327_, _08189_);
  and (_08329_, _08328_, _08326_);
  nor (_08330_, _08329_, _08321_);
  nor (_08331_, _07982_, _06899_);
  nor (_08332_, _08331_, _07983_);
  and (_08333_, _08332_, _07978_);
  not (_08334_, _08333_);
  and (_08335_, _07924_, _07795_);
  and (_08336_, _07936_, _07793_);
  nor (_08337_, _07922_, _07794_);
  and (_08338_, _07938_, _06898_);
  or (_08339_, _08338_, _08337_);
  or (_08340_, _08339_, _08336_);
  nor (_08341_, _08340_, _08335_);
  and (_08342_, _08090_, _07052_);
  and (_08343_, _07930_, _07034_);
  nor (_08344_, _07942_, _06898_);
  or (_08345_, _08344_, _08343_);
  nor (_08346_, _08345_, _08342_);
  and (_08347_, _08346_, _08341_);
  and (_08348_, _08347_, _08334_);
  and (_08349_, _08348_, _08330_);
  not (_08350_, _08349_);
  nor (_08351_, _08350_, _08317_);
  and (_08352_, _08351_, _08314_);
  and (_08353_, _08352_, _08309_);
  nand (_08354_, _08353_, _08308_);
  or (_08355_, _08354_, _07764_);
  not (_08356_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nand (_08357_, _07764_, _08356_);
  and (_08358_, _08357_, _08008_);
  and (_08359_, _08358_, _08355_);
  nor (_08360_, _08007_, _08356_);
  not (_08361_, _07727_);
  and (_08362_, _07749_, _07738_);
  and (_08363_, _08362_, _08299_);
  nor (_08364_, _08362_, _08299_);
  nor (_08365_, _08364_, _08363_);
  or (_08366_, _08365_, _08361_);
  and (_08367_, _08366_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  not (_08368_, _08363_);
  nor (_08369_, _08368_, _08059_);
  and (_08370_, _08364_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  or (_08371_, _08370_, _08369_);
  and (_08372_, _08371_, _07727_);
  or (_08373_, _08372_, _08367_);
  and (_08374_, _08373_, _08065_);
  or (_08375_, _08374_, _08360_);
  or (_08376_, _08375_, _08359_);
  and (_06811_, _08376_, _13707_);
  nand (_08377_, _07629_, _07353_);
  nand (_08378_, _07346_, _06847_);
  nor (_08379_, _07870_, _07792_);
  nor (_08380_, _08379_, _07871_);
  nor (_08381_, _08380_, _07770_);
  not (_08382_, _08381_);
  nor (_08383_, _07793_, _07781_);
  nor (_08384_, _08383_, _07902_);
  nor (_08385_, _08384_, _07899_);
  nor (_08386_, _08385_, _07900_);
  and (_08387_, _08386_, _07915_);
  nor (_08388_, _07860_, _06932_);
  and (_08389_, _07860_, _07052_);
  nor (_08390_, _08389_, _08388_);
  nor (_08391_, _08390_, _07974_);
  nor (_08392_, _07952_, _07933_);
  nor (_08393_, _07961_, _07860_);
  nor (_08394_, _08393_, _08392_);
  nor (_08395_, _08394_, _07052_);
  and (_08396_, _08394_, _07052_);
  or (_08397_, _08396_, _08189_);
  nor (_08398_, _08397_, _08395_);
  nor (_08399_, _08398_, _08391_);
  nor (_08400_, _07983_, _07052_);
  not (_08401_, _07987_);
  and (_08402_, _08401_, _08400_);
  nor (_08403_, _07987_, _07983_);
  nor (_08404_, _08403_, _07956_);
  nor (_08405_, _08404_, _08402_);
  nor (_08406_, _08405_, _07979_);
  and (_08407_, _07924_, _07781_);
  and (_08408_, _07936_, _07779_);
  nor (_08409_, _07922_, _07780_);
  and (_08410_, _07938_, _07956_);
  or (_08411_, _08410_, _08409_);
  or (_08412_, _08411_, _08408_);
  nor (_08413_, _08412_, _08407_);
  and (_08414_, _08090_, _07075_);
  not (_08415_, _08414_);
  and (_08416_, _07941_, _07052_);
  and (_08417_, _07930_, _06899_);
  nor (_08418_, _08417_, _08416_);
  and (_08419_, _08418_, _08415_);
  and (_08420_, _08419_, _08413_);
  not (_08421_, _08420_);
  nor (_08422_, _08421_, _08406_);
  and (_08423_, _08422_, _08399_);
  not (_08424_, _08423_);
  nor (_08425_, _08424_, _08387_);
  and (_08426_, _08425_, _08382_);
  and (_08427_, _08426_, _08378_);
  nand (_08428_, _08427_, _08377_);
  or (_08429_, _08428_, _07764_);
  not (_08430_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nand (_08431_, _07764_, _08430_);
  and (_08432_, _08431_, _08008_);
  and (_08433_, _08432_, _08429_);
  nor (_08434_, _08007_, _08430_);
  and (_08435_, _08299_, _07749_);
  nor (_08436_, _08435_, _08236_);
  or (_08437_, _08436_, _08361_);
  and (_08438_, _08437_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_08439_, _07749_, _08060_);
  and (_08440_, _08439_, _08299_);
  not (_08441_, _08440_);
  nor (_08442_, _08441_, _08059_);
  or (_08443_, _08363_, _08236_);
  and (_08444_, _08443_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  or (_08445_, _08444_, _08442_);
  and (_08446_, _08445_, _07727_);
  or (_08447_, _08446_, _08438_);
  and (_08448_, _08447_, _08065_);
  or (_08449_, _08448_, _08434_);
  or (_08450_, _08449_, _08433_);
  and (_06812_, _08450_, _13707_);
  nand (_08451_, _07634_, _07353_);
  nand (_08452_, _07348_, _06847_);
  nor (_08453_, _07906_, _07900_);
  not (_08454_, _08453_);
  nor (_08455_, _07916_, _07907_);
  and (_08456_, _08455_, _08454_);
  not (_08457_, _08456_);
  nor (_08458_, _07871_, _07789_);
  nor (_08459_, _08458_, _07872_);
  nor (_08460_, _08459_, _07770_);
  and (_08461_, _07860_, _07075_);
  nor (_08462_, _07860_, _07378_);
  or (_08463_, _08462_, _08461_);
  and (_08464_, _08463_, _07973_);
  nor (_08465_, _07860_, _07052_);
  nand (_08466_, _08465_, _07961_);
  nand (_08467_, _07953_, _07860_);
  and (_08468_, _08467_, _08466_);
  and (_08469_, _08468_, _07074_);
  nor (_08470_, _08468_, _07074_);
  or (_08471_, _08470_, _08189_);
  nor (_08472_, _08471_, _08469_);
  nor (_08473_, _08472_, _08464_);
  nor (_08474_, _08402_, _07074_);
  and (_08475_, _08402_, _07074_);
  nor (_08476_, _08475_, _08474_);
  nor (_08477_, _08476_, _07979_);
  and (_08478_, _07924_, _07777_);
  and (_08479_, _07936_, _07775_);
  nor (_08480_, _07922_, _07776_);
  and (_08481_, _07938_, _07074_);
  or (_08482_, _08481_, _08480_);
  or (_08483_, _08482_, _08479_);
  nor (_08484_, _08483_, _08478_);
  nor (_08485_, _07942_, _07074_);
  not (_08486_, _08485_);
  and (_08487_, _08090_, _07210_);
  and (_08488_, _07930_, _07052_);
  nor (_08489_, _08488_, _08487_);
  and (_08490_, _08489_, _08486_);
  and (_08491_, _08490_, _08484_);
  not (_08492_, _08491_);
  nor (_08493_, _08492_, _08477_);
  and (_08494_, _08493_, _08473_);
  not (_08495_, _08494_);
  nor (_08496_, _08495_, _08460_);
  and (_08497_, _08496_, _08457_);
  and (_08498_, _08497_, _08452_);
  and (_08499_, _08498_, _08451_);
  not (_08500_, _08499_);
  or (_08501_, _08500_, _07764_);
  not (_08502_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  nand (_08503_, _07764_, _08502_);
  and (_08504_, _08503_, _08008_);
  and (_08505_, _08504_, _08501_);
  nor (_08506_, _08007_, _08502_);
  not (_08507_, _08062_);
  nand (_08508_, _08507_, _07727_);
  and (_08509_, _08508_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_08510_, _08061_, _07738_);
  not (_08511_, _08510_);
  nor (_08512_, _08511_, _08059_);
  nor (_08513_, _08061_, _08502_);
  or (_08514_, _08513_, _08512_);
  and (_08515_, _08514_, _07727_);
  or (_08516_, _08515_, _08509_);
  and (_08517_, _08516_, _08065_);
  or (_08518_, _08517_, _08506_);
  or (_08519_, _08518_, _08505_);
  and (_06813_, _08519_, _13707_);
  and (_08520_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_08521_, \oc8051_top_1.oc8051_decoder1.state [0], \oc8051_top_1.oc8051_decoder1.state [1]);
  nor (_08522_, _08521_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_08523_, _08522_);
  not (_08524_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  nor (_08525_, \oc8051_top_1.oc8051_memory_interface1.imem_wait , \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and (_08526_, _08525_, _08524_);
  and (_08527_, _08521_, _06841_);
  and (_08528_, _08527_, _08526_);
  and (_08529_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  not (_08530_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_08531_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], \oc8051_top_1.oc8051_memory_interface1.cdone );
  not (_08532_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_08533_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  not (_08534_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  not (_08535_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_08536_, _08535_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_08537_, _08536_, _08534_);
  and (_08538_, _08537_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  not (_08539_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_08540_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], _08539_);
  and (_08541_, _08540_, _08534_);
  and (_08542_, _08541_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_08543_, _08542_, _08538_);
  nor (_08544_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_08545_, _08544_, _08534_);
  and (_08546_, _08545_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_08548_, _08544_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_08549_, _08548_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor (_08551_, _08549_, _08546_);
  and (_08552_, _08544_, _08534_);
  and (_08554_, _08552_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  and (_08555_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_08557_, _08555_, _08534_);
  and (_08558_, _08557_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_08559_, _08558_, _08554_);
  and (_08560_, _08559_, _08551_);
  and (_08561_, _08560_, _08543_);
  nor (_08562_, _08561_, _08533_);
  and (_08563_, _08562_, _08532_);
  or (_08564_, _08563_, _08531_);
  and (_08565_, _08564_, _08530_);
  or (_08566_, _08565_, _08529_);
  and (_08567_, _08566_, _08528_);
  not (_08568_, _08528_);
  and (_08569_, _08526_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and (_08570_, _08569_, _08568_);
  or (_08571_, _08570_, _08567_);
  and (_08572_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  not (_08573_, _08572_);
  nand (_08574_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_08575_, _08541_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  and (_08576_, _08537_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor (_08577_, _08576_, _08575_);
  and (_08578_, _08545_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_08579_, _08548_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor (_08580_, _08579_, _08578_);
  and (_08581_, _08552_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  and (_08582_, _08557_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_08583_, _08582_, _08581_);
  and (_08584_, _08583_, _08580_);
  and (_08585_, _08584_, _08577_);
  nor (_08586_, _08585_, _08533_);
  nand (_08587_, _08586_, _08532_);
  and (_08588_, _08587_, _08574_);
  or (_08589_, _08588_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_08590_, _08589_, _08573_);
  or (_08591_, _08590_, _08568_);
  and (_08592_, _08526_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and (_08593_, _08592_, _08568_);
  not (_08594_, _08593_);
  and (_08595_, _08594_, _08591_);
  and (_08596_, _08595_, _08571_);
  and (_08597_, _08545_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_08598_, _08552_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  and (_08599_, _08548_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_08600_, _08557_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_08601_, _08600_, _08599_);
  and (_08602_, _08541_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  and (_08603_, _08537_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor (_08604_, _08603_, _08602_);
  nand (_08605_, _08604_, _08601_);
  or (_08606_, _08605_, _08598_);
  or (_08607_, _08606_, _08597_);
  or (_08608_, _08607_, _08533_);
  or (_08609_, _08608_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor (_08610_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], _08532_);
  nor (_08611_, _08610_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_08612_, _08611_, _08609_);
  and (_08613_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  or (_08614_, _08613_, _08612_);
  nand (_08615_, _08614_, _08528_);
  and (_08616_, _08526_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and (_08617_, _08616_, _08568_);
  not (_08618_, _08617_);
  and (_08619_, _08618_, _08615_);
  and (_08620_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  not (_08621_, _08620_);
  nand (_08622_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_08623_, _08541_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  and (_08624_, _08537_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor (_08625_, _08624_, _08623_);
  and (_08626_, _08545_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_08627_, _08548_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor (_08628_, _08627_, _08626_);
  and (_08629_, _08552_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  and (_08630_, _08557_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_08631_, _08630_, _08629_);
  and (_08632_, _08631_, _08628_);
  and (_08633_, _08632_, _08625_);
  nor (_08634_, _08633_, _08533_);
  nand (_08635_, _08634_, _08532_);
  and (_08636_, _08635_, _08622_);
  or (_08637_, _08636_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_08638_, _08637_, _08621_);
  or (_08639_, _08638_, _08568_);
  and (_08640_, _08526_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and (_08641_, _08640_, _08568_);
  not (_08642_, _08641_);
  and (_08643_, _08642_, _08639_);
  not (_08644_, _08643_);
  and (_08645_, _08644_, _08619_);
  and (_08646_, _08645_, _08596_);
  and (_08647_, _08557_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  and (_08648_, _08548_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor (_08649_, _08648_, _08647_);
  and (_08650_, _08541_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_08651_, _08650_, _08533_);
  and (_08652_, _08651_, _08649_);
  and (_08653_, _08537_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  not (_08654_, _08653_);
  and (_08655_, _08552_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  and (_08656_, _08545_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nor (_08657_, _08656_, _08655_);
  and (_08658_, _08657_, _08654_);
  and (_08659_, _08658_, _08652_);
  and (_08660_, _08659_, _08532_);
  nor (_08661_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], _08532_);
  or (_08662_, _08661_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_08663_, _08662_, _08660_);
  and (_08664_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  or (_08665_, _08664_, _08663_);
  and (_08666_, _08665_, _08528_);
  and (_08667_, _08526_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and (_08668_, _08667_, _08568_);
  nor (_08669_, _08668_, _08666_);
  not (_08670_, _08669_);
  and (_08671_, \oc8051_top_1.oc8051_memory_interface1.dack_ir , \oc8051_top_1.oc8051_memory_interface1.ddat_ir [7]);
  not (_08672_, _08671_);
  and (_08673_, _08548_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_08674_, _08537_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  nor (_08675_, _08674_, _08673_);
  and (_08676_, _08557_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  and (_08677_, _08541_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_08678_, _08677_, _08676_);
  and (_08679_, _08678_, _08675_);
  and (_08680_, _08545_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_08681_, _08552_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  nor (_08682_, _08681_, _08680_);
  and (_08683_, _08682_, _08679_);
  or (_08684_, _08683_, _08533_);
  nand (_08685_, _08684_, _08532_);
  nor (_08686_, _08532_, \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  nor (_08687_, _08686_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nand (_08688_, _08687_, _08685_);
  and (_08689_, _08688_, _08672_);
  or (_08690_, _08689_, _08568_);
  and (_08691_, _08526_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and (_08692_, _08691_, _08568_);
  not (_08693_, _08692_);
  and (_08694_, _08693_, _08690_);
  not (_08695_, _08694_);
  and (_08696_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  not (_08697_, _08696_);
  and (_08698_, _08548_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_08699_, _08537_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor (_08700_, _08699_, _08698_);
  and (_08701_, _08557_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  and (_08702_, _08541_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_08703_, _08702_, _08701_);
  and (_08704_, _08703_, _08700_);
  and (_08705_, _08545_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_08706_, _08552_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  nor (_08707_, _08706_, _08705_);
  and (_08708_, _08707_, _08704_);
  or (_08709_, _08708_, _08533_);
  nand (_08710_, _08709_, _08532_);
  nor (_08711_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], _08532_);
  nor (_08712_, _08711_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nand (_08713_, _08712_, _08710_);
  and (_08714_, _08713_, _08697_);
  or (_08715_, _08714_, _08568_);
  and (_08716_, _08526_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and (_08717_, _08716_, _08568_);
  not (_08718_, _08717_);
  and (_08719_, _08718_, _08715_);
  and (_08720_, _08719_, _08695_);
  and (_08721_, _08720_, _08670_);
  and (_08722_, _08721_, _08646_);
  and (_08723_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  not (_08724_, _08723_);
  nand (_08725_, \oc8051_top_1.oc8051_memory_interface1.cdata [5], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_08726_, _08552_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  and (_08727_, _08541_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_08728_, _08727_, _08726_);
  and (_08729_, _08545_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_08730_, _08548_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor (_08731_, _08730_, _08729_);
  and (_08732_, _08557_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  and (_08733_, _08537_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor (_08734_, _08733_, _08732_);
  and (_08735_, _08734_, _08731_);
  and (_08736_, _08735_, _08728_);
  nor (_08737_, _08736_, _08533_);
  nand (_08738_, _08737_, _08532_);
  and (_08739_, _08738_, _08725_);
  or (_08740_, _08739_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_08741_, _08740_, _08724_);
  or (_08742_, _08741_, _08568_);
  and (_08743_, _08526_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and (_08744_, _08743_, _08568_);
  not (_08745_, _08744_);
  and (_08746_, _08745_, _08742_);
  not (_08747_, _08746_);
  and (_08748_, _08747_, _08720_);
  not (_08749_, _08619_);
  and (_08750_, _08749_, _08596_);
  and (_08751_, _08750_, _08669_);
  and (_08752_, _08751_, _08748_);
  nor (_08753_, _08719_, _08694_);
  and (_08754_, _08753_, _08747_);
  and (_08755_, _08754_, _08669_);
  and (_08756_, _08755_, _08646_);
  or (_08757_, _08756_, _08752_);
  or (_08758_, _08757_, _08722_);
  not (_08759_, _08719_);
  and (_08760_, _08759_, _08694_);
  and (_08761_, _08760_, _08746_);
  and (_08762_, _08761_, _08670_);
  and (_08763_, _08719_, _08694_);
  and (_08764_, _08763_, _08747_);
  or (_08765_, _08764_, _08762_);
  and (_08766_, _08765_, _08646_);
  not (_08767_, _08571_);
  and (_08768_, _08595_, _08767_);
  and (_08769_, _08768_, _08749_);
  and (_08770_, _08769_, _08643_);
  and (_08771_, _08770_, _08764_);
  and (_08772_, _08763_, _08746_);
  and (_08773_, _08772_, _08669_);
  and (_08774_, _08773_, _08646_);
  not (_08775_, _08595_);
  and (_08776_, _08748_, _08669_);
  and (_08777_, _08776_, _08775_);
  or (_08778_, _08777_, _08774_);
  or (_08779_, _08778_, _08771_);
  or (_08780_, _08779_, _08766_);
  and (_08781_, _08753_, _08746_);
  and (_08782_, _08781_, _08670_);
  and (_08783_, _08782_, _08770_);
  and (_08784_, _08776_, _08770_);
  nor (_08785_, _08784_, _08783_);
  not (_08786_, _08785_);
  and (_08787_, _08760_, _08747_);
  and (_08788_, _08787_, _08669_);
  and (_08789_, _08788_, _08646_);
  and (_08790_, _08781_, _08669_);
  and (_08791_, _08790_, _08646_);
  or (_08792_, _08791_, _08789_);
  or (_08793_, _08792_, _08786_);
  or (_08794_, _08793_, _08780_);
  or (_08795_, _08794_, _08758_);
  and (_08796_, _08746_, _08669_);
  and (_08797_, _08796_, _08760_);
  and (_08798_, _08797_, _08769_);
  not (_08799_, _08798_);
  and (_08800_, _08772_, _08670_);
  and (_08801_, _08800_, _08646_);
  and (_08802_, _08748_, _08670_);
  and (_08803_, _08643_, _08619_);
  and (_08804_, _08803_, _08768_);
  and (_08805_, _08804_, _08802_);
  nor (_08806_, _08805_, _08801_);
  and (_08807_, _08806_, _08799_);
  and (_08808_, _08787_, _08670_);
  and (_08809_, _08808_, _08770_);
  and (_08810_, _08782_, _08646_);
  nor (_08811_, _08810_, _08809_);
  and (_08812_, _08811_, _08807_);
  and (_08813_, _08797_, _08646_);
  and (_08814_, _08804_, _08776_);
  nor (_08815_, _08814_, _08813_);
  and (_08816_, _08770_, _08802_);
  and (_08817_, _08790_, _08770_);
  nor (_08818_, _08817_, _08816_);
  and (_08819_, _08818_, _08815_);
  and (_08820_, _08819_, _08812_);
  and (_08821_, _08746_, _08720_);
  and (_08822_, _08821_, _08670_);
  and (_08823_, _08770_, _08822_);
  and (_08824_, _08796_, _08720_);
  and (_08825_, _08824_, _08646_);
  or (_08826_, _08825_, _08823_);
  and (_08827_, _08804_, _08781_);
  and (_08828_, _08788_, _08769_);
  or (_08829_, _08828_, _08827_);
  or (_08830_, _08829_, _08826_);
  and (_08831_, _08824_, _08770_);
  and (_08832_, _08769_, _08762_);
  or (_08833_, _08832_, _08831_);
  and (_08834_, _08804_, _08764_);
  and (_08835_, _08834_, _08669_);
  and (_08836_, _08764_, _08670_);
  or (_08837_, _08800_, _08836_);
  and (_08838_, _08837_, _08804_);
  nor (_08839_, _08838_, _08835_);
  not (_08840_, _08839_);
  or (_08841_, _08840_, _08833_);
  nor (_08842_, _08841_, _08830_);
  nand (_08843_, _08842_, _08820_);
  or (_08844_, _08843_, _08795_);
  and (_08845_, _08844_, _08523_);
  not (_08846_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and (_08847_, _06841_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_08848_, _08847_, _08846_);
  and (_08849_, _08804_, _08800_);
  or (_08850_, _08849_, _08835_);
  and (_08851_, _08850_, _08848_);
  and (_08852_, _08804_, _08760_);
  and (_08853_, _08852_, _08848_);
  nand (_08854_, _08771_, _08847_);
  nor (_08855_, _08854_, _08846_);
  or (_08856_, _08855_, _08853_);
  or (_08857_, _08856_, _08851_);
  nor (_08858_, _08857_, _08845_);
  nor (_08859_, _08858_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_08860_, _08859_, _08520_);
  not (_08861_, _08860_);
  and (_08862_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_08863_, _08761_, _08754_);
  and (_08864_, _08863_, _08751_);
  and (_08865_, _08804_, _08782_);
  and (_08866_, _08788_, _08750_);
  or (_08867_, _08866_, _08865_);
  or (_08868_, _08867_, _08864_);
  and (_08869_, _08765_, _08750_);
  and (_08870_, _08824_, _08750_);
  or (_08871_, _08870_, _08771_);
  and (_08872_, _08781_, _08750_);
  nor (_08873_, _08619_, _08767_);
  and (_08874_, _08670_, _08595_);
  and (_08875_, _08874_, _08873_);
  and (_08876_, _08875_, _08821_);
  or (_08877_, _08876_, _08872_);
  and (_08878_, _08875_, _08748_);
  and (_08879_, _08772_, _08750_);
  or (_08880_, _08879_, _08878_);
  or (_08881_, _08880_, _08877_);
  or (_08882_, _08881_, _08871_);
  or (_08883_, _08882_, _08869_);
  or (_08884_, _08883_, _08868_);
  and (_08885_, _08884_, _08523_);
  and (_08886_, _08769_, _08644_);
  and (_08887_, _08886_, _08776_);
  and (_08888_, _08886_, _08808_);
  and (_08889_, _08886_, _08822_);
  nor (_08890_, _08889_, _08888_);
  not (_08891_, _08890_);
  nor (_08892_, _08891_, _08887_);
  nor (_08893_, _08892_, _08522_);
  and (_08894_, _08848_, _08787_);
  and (_08895_, _08894_, _08804_);
  or (_08896_, _08895_, _08855_);
  or (_08897_, _08896_, _08893_);
  or (_08898_, _08897_, _08885_);
  and (_08899_, _08898_, _06841_);
  or (_08900_, _08899_, _08862_);
  and (_08901_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_08902_, _08803_, _08596_);
  and (_08903_, _08902_, _08824_);
  and (_08904_, _08902_, _08776_);
  nor (_08905_, _08904_, _08903_);
  not (_08906_, _08905_);
  nor (_08907_, _08906_, _08853_);
  not (_08908_, _08907_);
  nor (_08909_, _08908_, _08893_);
  nor (_08910_, _08909_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_08911_, _08910_, _08901_);
  and (_08912_, _08911_, _13707_);
  and (_13962_, _08912_, _08900_);
  and (_06814_, _13962_, _08861_);
  and (_08913_, _08008_, _07711_);
  and (_08914_, _07678_, _07666_);
  nor (_08915_, _07724_, _07694_);
  and (_08916_, _08915_, _08914_);
  and (_08917_, _08916_, _08173_);
  and (_08918_, _08917_, _08913_);
  not (_08919_, _08918_);
  and (_08920_, _08919_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  or (_08921_, _07353_, _06847_);
  and (_08922_, _07914_, _07351_);
  or (_08923_, _07930_, _08922_);
  or (_08924_, _08923_, _07941_);
  or (_08925_, _08924_, _08921_);
  nor (_08926_, _08925_, _08090_);
  nor (_08927_, _08926_, _07074_);
  not (_08928_, _08927_);
  and (_08929_, _08928_, _08484_);
  and (_08930_, _08929_, _08473_);
  nor (_08931_, _08930_, _08919_);
  nor (_08932_, _08931_, _08920_);
  and (_08933_, _08919_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor (_08934_, _08926_, _07956_);
  not (_08935_, _08934_);
  and (_08936_, _08935_, _08413_);
  and (_08937_, _08936_, _08399_);
  nor (_08938_, _08937_, _08919_);
  nor (_08939_, _08938_, _08933_);
  and (_08940_, _08919_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  nor (_08941_, _08926_, _06898_);
  not (_08942_, _08941_);
  and (_08943_, _08942_, _08341_);
  and (_08944_, _08943_, _08330_);
  nor (_08945_, _08944_, _08919_);
  nor (_08946_, _08945_, _08940_);
  and (_08947_, _08919_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor (_08948_, _08926_, _07033_);
  not (_08949_, _08948_);
  and (_08950_, _08949_, _08254_);
  and (_08951_, _08950_, _08281_);
  and (_08952_, _08951_, _08272_);
  nor (_08953_, _08952_, _08919_);
  nor (_08954_, _08953_, _08947_);
  and (_08955_, _08919_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_08956_, _08926_, _08184_);
  not (_08957_, _08956_);
  and (_08958_, _08957_, _08201_);
  and (_08959_, _08958_, _08204_);
  and (_08960_, _08959_, _08193_);
  nor (_08961_, _08960_, _08919_);
  nor (_08962_, _08961_, _08955_);
  and (_08963_, _08919_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  nor (_08964_, _08926_, _08132_);
  not (_08965_, _08964_);
  and (_08966_, _08965_, _08154_);
  and (_08967_, _08966_, _08140_);
  nor (_08968_, _08967_, _08919_);
  nor (_08969_, _08968_, _08963_);
  nor (_08970_, _08918_, _07733_);
  nor (_08971_, _08926_, _07185_);
  not (_08972_, _08971_);
  and (_08973_, _08972_, _08089_);
  and (_08974_, _08973_, _08086_);
  and (_08975_, _08974_, _08083_);
  not (_08976_, _08975_);
  and (_08977_, _08976_, _08918_);
  nor (_08978_, _08977_, _08970_);
  and (_08979_, _08978_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and (_08980_, _08979_, _08969_);
  and (_08981_, _08980_, _08962_);
  and (_08982_, _08981_, _08954_);
  and (_08983_, _08982_, _08946_);
  and (_08984_, _08983_, _08939_);
  and (_08985_, _08984_, _08932_);
  nor (_08986_, _08918_, _07680_);
  nand (_08987_, _08986_, _08985_);
  or (_08988_, _08986_, _08985_);
  and (_08989_, _08988_, _07646_);
  and (_08990_, _08989_, _08987_);
  or (_08991_, _08990_, _07684_);
  and (_08992_, _08991_, _08919_);
  nor (_08993_, _08926_, _07103_);
  not (_08994_, _08993_);
  and (_08995_, _08994_, _07940_);
  and (_08996_, _08995_, _07926_);
  and (_08997_, _08996_, _07977_);
  nor (_08998_, _08997_, _08919_);
  or (_08999_, _08998_, _08992_);
  and (_06815_, _08999_, _13707_);
  not (_09000_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and (_09001_, _08978_, _09000_);
  nor (_09002_, _08978_, _09000_);
  nor (_09003_, _09002_, _09001_);
  and (_09004_, _09003_, _07646_);
  nor (_09005_, _09004_, _07734_);
  nor (_09006_, _09005_, _08918_);
  nor (_09007_, _09006_, _08977_);
  nand (_06816_, _09007_, _13707_);
  nor (_09008_, _08979_, _08969_);
  nor (_09009_, _09008_, _08980_);
  nor (_09010_, _09009_, _07645_);
  nor (_09011_, _09010_, _07741_);
  nor (_09012_, _09011_, _08918_);
  nor (_09013_, _09012_, _08968_);
  nand (_06817_, _09013_, _13707_);
  nor (_09014_, _08980_, _08962_);
  nor (_09015_, _09014_, _08981_);
  nor (_09016_, _09015_, _07645_);
  nor (_09017_, _09016_, _07752_);
  nor (_09018_, _09017_, _08918_);
  nor (_09019_, _09018_, _08961_);
  nand (_06818_, _09019_, _13707_);
  nor (_09020_, _08981_, _08954_);
  nor (_09021_, _09020_, _08982_);
  nor (_09022_, _09021_, _07645_);
  nor (_09023_, _09022_, _07702_);
  nor (_09024_, _09023_, _08918_);
  nor (_09025_, _09024_, _08953_);
  nor (_06819_, _09025_, rst);
  nor (_09026_, _08982_, _08946_);
  nor (_09027_, _09026_, _08983_);
  nor (_09028_, _09027_, _07645_);
  nor (_09029_, _09028_, _07714_);
  nor (_09030_, _09029_, _08918_);
  nor (_09031_, _09030_, _08945_);
  nor (_06820_, _09031_, rst);
  nor (_09032_, _08983_, _08939_);
  nor (_09033_, _09032_, _08984_);
  nor (_09034_, _09033_, _07645_);
  nor (_09035_, _09034_, _07670_);
  nor (_09036_, _09035_, _08918_);
  nor (_09037_, _09036_, _08938_);
  nor (_06821_, _09037_, rst);
  nor (_09038_, _08984_, _08932_);
  nor (_09039_, _09038_, _08985_);
  nor (_09040_, _09039_, _07645_);
  nor (_09041_, _09040_, _07649_);
  nor (_09042_, _09041_, _08918_);
  nor (_09043_, _09042_, _08931_);
  nor (_06822_, _09043_, rst);
  and (_09044_, _08913_, _08296_);
  nand (_09045_, _09044_, _08916_);
  nor (_09046_, _09045_, _08001_);
  and (_09047_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], _06841_);
  and (_09048_, _09047_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_09049_, _09045_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_09050_, _09049_, _09048_);
  or (_09051_, _09050_, _09046_);
  not (_09052_, _09048_);
  nor (_09053_, _07942_, _06963_);
  nor (_09054_, _08031_, _07033_);
  and (_09055_, _07860_, _06932_);
  not (_09056_, _09055_);
  nor (_09057_, _07103_, _07000_);
  and (_09058_, _09057_, _07954_);
  and (_09059_, _09058_, _07364_);
  and (_09060_, _09059_, _07390_);
  and (_09061_, _09060_, _07367_);
  nor (_09062_, _09061_, _07933_);
  and (_09063_, _07860_, _06985_);
  nor (_09064_, _09063_, _09062_);
  and (_09065_, _09064_, _09056_);
  and (_09066_, _07962_, _07103_);
  and (_09067_, _06917_, _06979_);
  and (_09068_, _06947_, _07000_);
  and (_09069_, _09068_, _09067_);
  and (_09070_, _09069_, _09066_);
  and (_09071_, _06932_, _06985_);
  and (_09072_, _09071_, _09070_);
  nor (_09073_, _09072_, _07860_);
  not (_09074_, _09073_);
  and (_09075_, _09074_, _09065_);
  and (_09076_, _07860_, _07378_);
  nor (_09077_, _09076_, _08462_);
  and (_09078_, _09077_, _09075_);
  and (_09079_, _09078_, _07969_);
  nor (_09080_, _09078_, _07969_);
  nor (_09081_, _09080_, _09079_);
  and (_09082_, _09081_, _07948_);
  and (_09083_, _07860_, _07969_);
  nor (_09084_, _09083_, _08023_);
  nor (_09085_, _09084_, _07974_);
  or (_09086_, _09085_, _09082_);
  or (_09087_, _09086_, _09054_);
  and (_09088_, _07353_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  nor (_09089_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  and (_09090_, _07040_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_09091_, _09090_, _09089_);
  nor (_09092_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  and (_09093_, _07021_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_09094_, _09093_, _09092_);
  nor (_09095_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and (_09096_, _07173_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_09097_, _09096_, _09095_);
  not (_09098_, _09097_);
  nor (_09099_, _09098_, _08014_);
  nor (_09100_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  and (_09101_, _07121_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_09102_, _09101_, _09100_);
  and (_09103_, _09102_, _09099_);
  nor (_09104_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  and (_09105_, _07140_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_09106_, _09105_, _09104_);
  and (_09107_, _09106_, _09103_);
  and (_09108_, _09107_, _09094_);
  nor (_09109_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  and (_09110_, _06865_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_09111_, _09110_, _09109_);
  and (_09112_, _09111_, _09108_);
  and (_09113_, _09112_, _09091_);
  nor (_09114_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  and (_09115_, _07062_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_09116_, _09115_, _09114_);
  and (_09117_, _09116_, _09113_);
  nor (_09118_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  and (_09119_, _07092_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_09120_, _09119_, _09118_);
  nor (_09121_, _09120_, _09117_);
  and (_09122_, _09120_, _09117_);
  or (_09123_, _09122_, _09121_);
  nor (_09124_, _09123_, _07916_);
  and (_09125_, _07326_, _06847_);
  or (_09126_, _09125_, _09124_);
  or (_09127_, _09126_, _09088_);
  or (_09128_, _09127_, _09087_);
  or (_09129_, _09128_, _09053_);
  or (_09130_, _09129_, _09052_);
  and (_09131_, _09130_, _13707_);
  and (_06823_, _09131_, _09051_);
  and (_09132_, _08913_, _08237_);
  and (_09133_, _09132_, _08916_);
  nor (_09134_, _09133_, _09048_);
  not (_09135_, _09134_);
  nand (_09136_, _09135_, _08001_);
  not (_09137_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  nand (_09138_, _09134_, _09137_);
  and (_09139_, _09138_, _13707_);
  and (_06824_, _09139_, _09136_);
  nor (_09140_, _09045_, _08105_);
  and (_09141_, _09045_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or (_09142_, _09141_, _09048_);
  or (_09143_, _09142_, _09140_);
  and (_09144_, _09098_, _08014_);
  nor (_09145_, _09144_, _09099_);
  and (_09146_, _09145_, _07915_);
  nand (_09147_, _07583_, _07353_);
  nor (_09148_, _08023_, _07972_);
  not (_09149_, _09148_);
  nor (_09150_, _09149_, _07964_);
  nor (_09151_, _09150_, _07400_);
  and (_09152_, _09150_, _07400_);
  or (_09153_, _09152_, _08189_);
  nor (_09154_, _09153_, _09151_);
  and (_09155_, _07941_, _07400_);
  and (_09156_, _07307_, _06847_);
  nor (_09157_, _08031_, _06898_);
  nor (_09158_, _07974_, _07185_);
  or (_09159_, _09158_, _09157_);
  or (_09160_, _09159_, _09156_);
  nor (_09161_, _09160_, _09155_);
  not (_09162_, _09161_);
  nor (_09163_, _09162_, _09154_);
  nand (_09164_, _09163_, _09147_);
  or (_09165_, _09164_, _09146_);
  or (_09166_, _09165_, _09052_);
  and (_09167_, _09166_, _13707_);
  and (_06825_, _09167_, _09143_);
  not (_09168_, _08166_);
  nor (_09169_, _09045_, _09168_);
  and (_09170_, _09045_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_09171_, _09170_, _09048_);
  or (_09172_, _09171_, _09169_);
  nor (_09173_, _09102_, _09099_);
  not (_09174_, _09173_);
  nor (_09175_, _09103_, _07916_);
  and (_09176_, _09175_, _09174_);
  not (_09177_, _09176_);
  and (_09178_, _07502_, _07353_);
  not (_09179_, _09178_);
  and (_09180_, _07941_, _07364_);
  and (_09181_, _09058_, _07860_);
  and (_09182_, _09066_, _07000_);
  and (_09183_, _09182_, _07933_);
  nor (_09184_, _09183_, _09181_);
  and (_09185_, _09184_, _06947_);
  not (_09186_, _09185_);
  nor (_09187_, _09184_, _06947_);
  nor (_09188_, _09187_, _08189_);
  and (_09189_, _09188_, _09186_);
  and (_09190_, _07309_, _06847_);
  and (_09191_, _08030_, _07052_);
  and (_09192_, _07973_, _07133_);
  or (_09193_, _09192_, _09191_);
  or (_09194_, _09193_, _09190_);
  or (_09195_, _09194_, _09189_);
  nor (_09196_, _09195_, _09180_);
  and (_09197_, _09196_, _09179_);
  and (_09198_, _09197_, _09177_);
  nand (_09199_, _09198_, _09048_);
  and (_09200_, _09199_, _13707_);
  and (_06826_, _09200_, _09172_);
  nor (_09201_, _09045_, _08223_);
  and (_09202_, _09045_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_09203_, _09202_, _09048_);
  or (_09204_, _09203_, _09201_);
  nor (_09205_, _09106_, _09103_);
  nor (_09206_, _09205_, _09107_);
  and (_09207_, _09206_, _07915_);
  not (_09208_, _09207_);
  and (_09209_, _09182_, _06947_);
  and (_09210_, _09209_, _07933_);
  and (_09211_, _09059_, _07860_);
  nor (_09212_, _09211_, _09210_);
  and (_09213_, _09212_, _06979_);
  nor (_09214_, _09212_, _06979_);
  nor (_09215_, _09214_, _09213_);
  and (_09216_, _09215_, _07948_);
  not (_09217_, _09216_);
  and (_09218_, _07973_, _07149_);
  and (_09219_, _07353_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  nor (_09220_, _09219_, _09218_);
  and (_09221_, _07311_, _06847_);
  nor (_09222_, _08031_, _07074_);
  and (_09223_, _07941_, _07390_);
  or (_09224_, _09223_, _09222_);
  nor (_09225_, _09224_, _09221_);
  and (_09226_, _09225_, _09220_);
  and (_09227_, _09226_, _09217_);
  and (_09228_, _09227_, _09208_);
  nand (_09229_, _09228_, _09048_);
  and (_09230_, _09229_, _13707_);
  and (_06827_, _09230_, _09204_);
  not (_09231_, _08288_);
  nor (_09232_, _09045_, _09231_);
  and (_09233_, _09045_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_09234_, _09233_, _09048_);
  or (_09235_, _09234_, _09232_);
  nor (_09236_, _09107_, _09094_);
  nor (_09237_, _09236_, _09108_);
  and (_09238_, _09237_, _07915_);
  not (_09239_, _09238_);
  nor (_09240_, _09060_, _07367_);
  not (_09241_, _09240_);
  and (_09242_, _09241_, _09062_);
  and (_09243_, _09209_, _06979_);
  nor (_09244_, _09243_, _06917_);
  nor (_09245_, _09244_, _09070_);
  nor (_09246_, _09245_, _07860_);
  nor (_09247_, _09246_, _09242_);
  nor (_09248_, _09247_, _08189_);
  and (_09249_, _07941_, _07367_);
  or (_09250_, _09249_, _08032_);
  nor (_09251_, _09250_, _09248_);
  and (_09252_, _07314_, _06847_);
  nor (_09253_, _07974_, _07033_);
  and (_09254_, _07353_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  or (_09255_, _09254_, _09253_);
  nor (_09256_, _09255_, _09252_);
  and (_09257_, _09256_, _09251_);
  and (_09258_, _09257_, _09239_);
  nand (_09259_, _09258_, _09048_);
  and (_09260_, _09259_, _13707_);
  and (_06828_, _09260_, _09235_);
  not (_09261_, _08354_);
  nor (_09262_, _09045_, _09261_);
  and (_09263_, _09045_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or (_09264_, _09263_, _09048_);
  or (_09265_, _09264_, _09262_);
  nor (_09266_, _09111_, _09108_);
  nor (_09267_, _09266_, _09112_);
  and (_09268_, _09267_, _07915_);
  not (_09269_, _09268_);
  and (_09270_, _07317_, _06847_);
  nor (_09271_, _09070_, _07860_);
  nor (_09272_, _09271_, _09062_);
  nor (_09273_, _09272_, _07382_);
  and (_09274_, _09272_, _07382_);
  nor (_09275_, _09274_, _09273_);
  and (_09276_, _09275_, _07948_);
  and (_09277_, _07353_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  nor (_09278_, _07860_, _06899_);
  or (_09279_, _09278_, _07974_);
  nor (_09280_, _09279_, _09063_);
  nor (_09281_, _08031_, _07185_);
  and (_09282_, _07941_, _07382_);
  or (_09283_, _09282_, _09281_);
  or (_09284_, _09283_, _09280_);
  nor (_09285_, _09284_, _09277_);
  not (_09286_, _09285_);
  nor (_09287_, _09286_, _09276_);
  not (_09288_, _09287_);
  nor (_09289_, _09288_, _09270_);
  and (_09290_, _09289_, _09269_);
  nand (_09291_, _09290_, _09048_);
  and (_09292_, _09291_, _13707_);
  and (_06829_, _09292_, _09265_);
  not (_09293_, _08428_);
  nor (_09294_, _09045_, _09293_);
  and (_09295_, _09045_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or (_09296_, _09295_, _09048_);
  or (_09297_, _09296_, _09294_);
  nor (_09298_, _09112_, _09091_);
  not (_09299_, _09298_);
  nor (_09300_, _09113_, _07916_);
  and (_09301_, _09300_, _09299_);
  not (_09302_, _09301_);
  and (_09303_, _07320_, _06847_);
  and (_09304_, _09070_, _06985_);
  nor (_09305_, _09304_, _07860_);
  not (_09306_, _09305_);
  and (_09307_, _09306_, _09064_);
  and (_09308_, _09307_, _06932_);
  nor (_09309_, _09307_, _06932_);
  or (_09310_, _09309_, _09308_);
  and (_09311_, _09310_, _07948_);
  and (_09312_, _07353_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  nor (_09313_, _08465_, _07974_);
  and (_09314_, _09313_, _09056_);
  and (_09315_, _08030_, _07133_);
  and (_09316_, _07941_, _07371_);
  or (_09317_, _09316_, _09315_);
  or (_09318_, _09317_, _09314_);
  nor (_09319_, _09318_, _09312_);
  not (_09320_, _09319_);
  nor (_09321_, _09320_, _09311_);
  not (_09322_, _09321_);
  nor (_09323_, _09322_, _09303_);
  and (_09324_, _09323_, _09302_);
  nand (_09325_, _09324_, _09048_);
  and (_09326_, _09325_, _13707_);
  and (_06830_, _09326_, _09297_);
  nor (_09327_, _09045_, _08499_);
  and (_09328_, _09045_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_09329_, _09328_, _09048_);
  or (_09330_, _09329_, _09327_);
  nor (_09331_, _09116_, _09113_);
  nor (_09332_, _09331_, _09117_);
  and (_09333_, _09332_, _07915_);
  not (_09334_, _09333_);
  and (_09335_, _07323_, _06847_);
  and (_09336_, _09075_, _07378_);
  nor (_09337_, _09075_, _07378_);
  nor (_09338_, _09337_, _09336_);
  nor (_09339_, _09338_, _08189_);
  and (_09340_, _07353_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  nor (_09341_, _07860_, _07075_);
  or (_09342_, _09341_, _07974_);
  nor (_09343_, _09342_, _09076_);
  and (_09344_, _08030_, _07149_);
  and (_09345_, _07941_, _07016_);
  or (_09346_, _09345_, _09344_);
  or (_09347_, _09346_, _09343_);
  nor (_09348_, _09347_, _09340_);
  not (_09349_, _09348_);
  nor (_09350_, _09349_, _09339_);
  not (_09351_, _09350_);
  nor (_09352_, _09351_, _09335_);
  and (_09353_, _09352_, _09334_);
  nand (_09354_, _09353_, _09048_);
  and (_09355_, _09354_, _13707_);
  and (_06831_, _09355_, _09330_);
  nand (_09356_, _09135_, _08105_);
  or (_09357_, _09135_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_09358_, _09357_, _13707_);
  and (_06832_, _09358_, _09356_);
  or (_09359_, _09134_, _08166_);
  or (_09360_, _09135_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_09361_, _09360_, _13707_);
  and (_06833_, _09361_, _09359_);
  nand (_09362_, _09135_, _08223_);
  not (_09363_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  nand (_09364_, _09134_, _09363_);
  and (_09365_, _09364_, _13707_);
  and (_06834_, _09365_, _09362_);
  or (_09366_, _09134_, _08288_);
  or (_09367_, _09135_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_09368_, _09367_, _13707_);
  and (_06835_, _09368_, _09366_);
  or (_09369_, _09134_, _08354_);
  or (_09370_, _09135_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_09371_, _09370_, _13707_);
  and (_06836_, _09371_, _09369_);
  or (_09372_, _09134_, _08428_);
  or (_09373_, _09135_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_09374_, _09373_, _13707_);
  and (_06837_, _09374_, _09372_);
  nand (_09375_, _09135_, _08499_);
  or (_09376_, _09135_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_09377_, _09376_, _13707_);
  and (_06838_, _09377_, _09375_);
  nor (_09378_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  nor (_09379_, _09378_, _08059_);
  nor (_09380_, _07694_, _07666_);
  and (_09381_, _07725_, _07678_);
  and (_09382_, _09381_, _09380_);
  and (_09383_, _09382_, _08065_);
  and (_09384_, _09378_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or (_09385_, _09384_, _09383_);
  or (_09386_, _09385_, _09379_);
  and (_09387_, _08008_, _07763_);
  and (_09388_, _09387_, _09382_);
  not (_09389_, _09388_);
  nor (_09390_, _08507_, _08059_);
  not (_09391_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or (_09392_, _08062_, _09391_);
  nand (_09393_, _09392_, _09383_);
  or (_09394_, _09393_, _09390_);
  and (_09395_, _09394_, _09389_);
  and (_09396_, _09395_, _09386_);
  nor (_09397_, _09389_, _08997_);
  or (_09398_, _09397_, _09396_);
  and (_06839_, _09398_, _13707_);
  nand (_09399_, _09388_, _08967_);
  nand (_09400_, _09383_, _08173_);
  and (_09401_, _09400_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  or (_09402_, _09401_, _09388_);
  nor (_09403_, _09400_, _08059_);
  or (_09404_, _09403_, _09402_);
  and (_09405_, _09404_, _09399_);
  and (_07290_, _09405_, _13707_);
  or (_09406_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_09407_, _07333_, _07329_);
  or (_09408_, _09407_, _07337_);
  or (_09409_, _09408_, _07340_);
  or (_09410_, _07346_, _07343_);
  or (_09411_, _07348_, _07303_);
  or (_09412_, _09411_, _09410_);
  or (_09413_, _09412_, _09409_);
  and (_09414_, _09413_, _06847_);
  or (_09415_, _08018_, _07873_);
  not (_09416_, _08017_);
  nand (_09417_, _09416_, _07873_);
  and (_09418_, _09417_, _07769_);
  and (_09419_, _09418_, _09415_);
  not (_09420_, _07771_);
  nand (_09421_, _07910_, _09420_);
  or (_09422_, _07910_, _07772_);
  and (_09423_, _07915_, _09422_);
  and (_09424_, _09423_, _09421_);
  and (_09425_, _09071_, _07379_);
  and (_09426_, _09069_, _07353_);
  nand (_09427_, _09426_, _09425_);
  nand (_09428_, _09427_, \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or (_09429_, _09428_, _09424_);
  or (_09430_, _09429_, _09419_);
  or (_09431_, _09430_, _09414_);
  and (_09432_, _09431_, _09406_);
  or (_09433_, _09432_, _09383_);
  not (_09434_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_09435_, _08237_, _09434_);
  nand (_09436_, _09435_, _09383_);
  or (_09437_, _09436_, _08238_);
  and (_09438_, _09437_, _09389_);
  and (_09439_, _09438_, _09433_);
  nor (_09440_, _09389_, _08960_);
  or (_09441_, _09440_, _09439_);
  and (_07292_, _09441_, _13707_);
  and (_09442_, _09383_, _08296_);
  nand (_09443_, _09442_, _08059_);
  or (_09444_, _09442_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_09445_, _09444_, _09389_);
  and (_09446_, _09445_, _09443_);
  nor (_09447_, _09389_, _08952_);
  or (_09448_, _09447_, _09446_);
  and (_07294_, _09448_, _13707_);
  and (_09449_, _08364_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  or (_09450_, _09449_, _08369_);
  and (_09451_, _09450_, _09383_);
  nor (_09452_, _09389_, _08944_);
  not (_09453_, _09383_);
  or (_09454_, _09453_, _08365_);
  not (_09455_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  nor (_09456_, _09388_, _09455_);
  and (_09457_, _09456_, _09454_);
  or (_09458_, _09457_, _09452_);
  or (_09459_, _09458_, _09451_);
  and (_07296_, _09459_, _13707_);
  nand (_09460_, _09388_, _08937_);
  and (_09461_, _08443_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  or (_09462_, _09461_, _08442_);
  and (_09463_, _09462_, _09383_);
  or (_09464_, _09453_, _08436_);
  and (_09465_, _09464_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  or (_09466_, _09465_, _09388_);
  or (_09467_, _09466_, _09463_);
  and (_09468_, _09467_, _09460_);
  and (_07298_, _09468_, _13707_);
  or (_09469_, _08510_, _08273_);
  nand (_09470_, _09469_, _09383_);
  or (_09471_, _09470_, _08512_);
  and (_09472_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  and (_09473_, _07915_, _07898_);
  and (_09474_, _07869_, _07769_);
  or (_09475_, _09474_, _09473_);
  and (_09476_, _09475_, _09472_);
  nand (_09477_, _09472_, _07942_);
  and (_09478_, _09477_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  or (_09479_, _09478_, _09383_);
  or (_09480_, _09479_, _09476_);
  and (_09481_, _09480_, _09389_);
  and (_09482_, _09481_, _09471_);
  nor (_09483_, _09389_, _08930_);
  or (_09484_, _09483_, _09482_);
  and (_07300_, _09484_, _13707_);
  not (_09485_, _09047_);
  and (_09486_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], _06841_);
  and (_09487_, _09486_, _09485_);
  not (_09488_, _09487_);
  not (_09489_, _07678_);
  and (_09490_, _07763_, _09489_);
  and (_09491_, _07723_, _07711_);
  and (_09492_, _09491_, _08008_);
  and (_09493_, _09492_, _09490_);
  nand (_09494_, _09493_, _09380_);
  and (_09495_, _09494_, _09488_);
  or (_09496_, _09495_, _08001_);
  not (_09497_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_09498_, _09047_, _09497_);
  and (_09499_, _09491_, _07679_);
  and (_09500_, _08065_, _07695_);
  and (_09501_, _09500_, _09499_);
  and (_09502_, _09501_, _08062_);
  and (_09503_, _09502_, _08059_);
  nor (_09504_, _09502_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  not (_09505_, _09498_);
  and (_09506_, _09505_, _09495_);
  not (_09507_, _09506_);
  nor (_09508_, _09507_, _09504_);
  not (_09509_, _09508_);
  nor (_09510_, _09509_, _09503_);
  nor (_09511_, _09510_, _09498_);
  nand (_09512_, _09511_, _09496_);
  or (_09513_, _09505_, _09129_);
  and (_09514_, _09513_, _09512_);
  and (_07355_, _09514_, _13707_);
  or (_09515_, _09495_, _08105_);
  and (_09516_, _09501_, _07763_);
  and (_09517_, _09516_, _08059_);
  nor (_09518_, _09516_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_09519_, _09518_, _09507_);
  not (_09520_, _09519_);
  nor (_09521_, _09520_, _09517_);
  nor (_09522_, _09521_, _09498_);
  nand (_09523_, _09522_, _09515_);
  or (_09524_, _09505_, _09165_);
  and (_09525_, _09524_, _09523_);
  and (_07525_, _09525_, _13707_);
  nor (_09526_, _09505_, _09198_);
  not (_09527_, _09526_);
  or (_09528_, _09495_, _08166_);
  and (_09529_, _09491_, _07695_);
  and (_09530_, _08065_, _07679_);
  and (_09531_, _09530_, _09529_);
  nor (_09532_, _09531_, _06944_);
  not (_09533_, _09495_);
  not (_09534_, _08173_);
  nor (_09535_, _09534_, _08059_);
  nor (_09536_, _08173_, _06944_);
  nor (_09537_, _09536_, _09535_);
  nand (_09538_, _09506_, _09501_);
  nor (_09539_, _09538_, _09537_);
  or (_09540_, _09539_, _09533_);
  or (_09541_, _09540_, _09532_);
  and (_09542_, _09541_, _09505_);
  nand (_09543_, _09542_, _09528_);
  nand (_09544_, _09543_, _09527_);
  and (_07527_, _09544_, _13707_);
  or (_09545_, _09495_, _08223_);
  and (_09546_, _09501_, _08237_);
  and (_09547_, _09546_, _08059_);
  nor (_09548_, _09546_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor (_09549_, _09548_, _09507_);
  not (_09550_, _09549_);
  nor (_09551_, _09550_, _09547_);
  nor (_09552_, _09551_, _09498_);
  nand (_09553_, _09552_, _09545_);
  and (_09554_, _09498_, _09228_);
  not (_09555_, _09554_);
  and (_09556_, _09555_, _09553_);
  and (_07529_, _09556_, _13707_);
  nor (_09557_, _09505_, _09258_);
  not (_09558_, _09557_);
  or (_09559_, _09495_, _08288_);
  nor (_09560_, _09531_, _06912_);
  nor (_09561_, _09560_, _09533_);
  not (_09562_, _09531_);
  nor (_09563_, _08296_, _06912_);
  nor (_09564_, _09563_, _08298_);
  or (_09565_, _09564_, _09562_);
  and (_09566_, _09565_, _09561_);
  nor (_09567_, _09566_, _09498_);
  nand (_09568_, _09567_, _09559_);
  nand (_09569_, _09568_, _09558_);
  and (_07531_, _09569_, _13707_);
  nor (_09570_, _09505_, _09290_);
  not (_09571_, _09570_);
  or (_09572_, _09495_, _08354_);
  nor (_09573_, _09531_, _06893_);
  nor (_09574_, _09573_, _09533_);
  nor (_09575_, _08363_, _06893_);
  nor (_09576_, _09575_, _08369_);
  or (_09577_, _09576_, _09562_);
  and (_09578_, _09577_, _09574_);
  nor (_09579_, _09578_, _09498_);
  nand (_09580_, _09579_, _09572_);
  nand (_09581_, _09580_, _09571_);
  and (_07533_, _09581_, _13707_);
  nor (_09582_, _09505_, _09324_);
  not (_09583_, _09582_);
  or (_09584_, _09495_, _08428_);
  nor (_09585_, _09531_, _06929_);
  nor (_09586_, _09585_, _09533_);
  nor (_09587_, _08440_, _06929_);
  nor (_09588_, _09587_, _08442_);
  or (_09589_, _09588_, _09562_);
  and (_09590_, _09589_, _09586_);
  nor (_09591_, _09590_, _09498_);
  nand (_09592_, _09591_, _09584_);
  nand (_09593_, _09592_, _09583_);
  and (_07535_, _09593_, _13707_);
  or (_09594_, _09495_, _08499_);
  and (_09595_, _09501_, _08510_);
  and (_09596_, _09595_, _08059_);
  nor (_09597_, _09595_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor (_09598_, _09597_, _09507_);
  not (_09599_, _09598_);
  nor (_09600_, _09599_, _09596_);
  nor (_09601_, _09600_, _09498_);
  nand (_09602_, _09601_, _09594_);
  and (_09603_, _09498_, _09353_);
  not (_09604_, _09603_);
  and (_09605_, _09604_, _09602_);
  and (_07537_, _09605_, _13707_);
  and (_09606_, _09529_, _08914_);
  and (_09607_, _09606_, _08062_);
  nand (_09608_, _09607_, _08059_);
  or (_09609_, _09607_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_09610_, _09609_, _08065_);
  and (_09611_, _09610_, _09608_);
  and (_09612_, _09606_, _07763_);
  nand (_09613_, _09612_, _08997_);
  or (_09614_, _09612_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_09615_, _09614_, _08008_);
  and (_09616_, _09615_, _09613_);
  not (_09617_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  nor (_09618_, _08007_, _09617_);
  or (_09619_, _09618_, rst);
  or (_09620_, _09619_, _09616_);
  or (_08547_, _09620_, _09611_);
  and (_09621_, _08914_, _07726_);
  and (_09622_, _09621_, _08062_);
  nand (_09623_, _09622_, _08059_);
  or (_09624_, _09622_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_09625_, _09624_, _08065_);
  and (_09626_, _09625_, _09623_);
  not (_09627_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_09628_, _09621_, _07763_);
  nor (_09629_, _09628_, _09627_);
  not (_09630_, _09628_);
  nor (_09631_, _09630_, _08997_);
  or (_09632_, _09631_, _09629_);
  and (_09633_, _09632_, _08008_);
  nor (_09634_, _08007_, _09627_);
  or (_09635_, _09634_, rst);
  or (_09636_, _09635_, _09633_);
  or (_08550_, _09636_, _09626_);
  and (_09637_, _09489_, _07666_);
  and (_09638_, _09637_, _09529_);
  and (_09639_, _09638_, _08062_);
  nand (_09640_, _09639_, _08059_);
  or (_09641_, _09639_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_09642_, _09641_, _08065_);
  and (_09643_, _09642_, _09640_);
  and (_09644_, _09638_, _07763_);
  not (_09645_, _09644_);
  nor (_09646_, _09645_, _08997_);
  not (_09647_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  nor (_09648_, _09644_, _09647_);
  or (_09649_, _09648_, _09646_);
  and (_09650_, _09649_, _08008_);
  nor (_09651_, _08007_, _09647_);
  or (_09652_, _09651_, rst);
  or (_09653_, _09652_, _09650_);
  or (_08553_, _09653_, _09643_);
  and (_09654_, _09637_, _07726_);
  not (_09655_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  nor (_09656_, _08062_, _09655_);
  or (_09657_, _09656_, _09390_);
  and (_09658_, _09657_, _09654_);
  nor (_09659_, _09654_, _09655_);
  or (_09660_, _09659_, _09658_);
  and (_09661_, _09660_, _08065_);
  and (_09662_, _07763_, _07725_);
  and (_09663_, _09662_, _07695_);
  and (_09664_, _09637_, _09663_);
  nor (_09665_, _09664_, _09655_);
  not (_09666_, _09664_);
  nor (_09667_, _09666_, _08997_);
  or (_09668_, _09667_, _09665_);
  and (_09669_, _09668_, _08008_);
  nor (_09670_, _08007_, _09655_);
  or (_09671_, _09670_, rst);
  or (_09672_, _09671_, _09669_);
  or (_08556_, _09672_, _09661_);
  or (_09673_, _09612_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  nand (_09674_, _09612_, _08059_);
  and (_09675_, _09674_, _08065_);
  nand (_09676_, _09612_, _08975_);
  and (_09677_, _09676_, _08008_);
  or (_09678_, _09677_, _09675_);
  and (_09679_, _09678_, _09673_);
  not (_09680_, _08007_);
  and (_09681_, _09680_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  or (_09682_, _09681_, rst);
  or (_11189_, _09682_, _09679_);
  and (_09683_, _09606_, _08173_);
  nand (_09684_, _09683_, _08059_);
  or (_09685_, _09683_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_09686_, _09685_, _08065_);
  and (_09687_, _09686_, _09684_);
  nand (_09688_, _09612_, _08967_);
  or (_09689_, _09612_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_09690_, _09689_, _08008_);
  and (_09691_, _09690_, _09688_);
  and (_09692_, _09680_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  or (_09693_, _09692_, rst);
  or (_09694_, _09693_, _09691_);
  or (_11191_, _09694_, _09687_);
  not (_09695_, _08300_);
  nand (_09696_, _09606_, _09695_);
  and (_09697_, _09696_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_09698_, _07762_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or (_09699_, _09698_, _08238_);
  and (_09700_, _09699_, _09606_);
  or (_09701_, _09700_, _09697_);
  and (_09702_, _09701_, _08065_);
  nand (_09703_, _09612_, _08960_);
  or (_09704_, _09612_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_09705_, _09704_, _08008_);
  and (_09706_, _09705_, _09703_);
  not (_09707_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  nor (_09708_, _08007_, _09707_);
  or (_09709_, _09708_, rst);
  or (_09710_, _09709_, _09706_);
  or (_11193_, _09710_, _09702_);
  nand (_09711_, _09606_, _07761_);
  and (_09712_, _09711_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_09713_, _09695_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or (_09714_, _09713_, _08298_);
  and (_09715_, _09714_, _09606_);
  or (_09716_, _09715_, _09712_);
  and (_09717_, _09716_, _08065_);
  nand (_09718_, _09612_, _08952_);
  or (_09719_, _09612_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_09720_, _09719_, _08008_);
  and (_09721_, _09720_, _09718_);
  and (_09722_, _09680_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or (_09723_, _09722_, rst);
  or (_09724_, _09723_, _09721_);
  or (_11195_, _09724_, _09717_);
  and (_09725_, _09606_, _08363_);
  nand (_09726_, _09725_, _08059_);
  or (_09727_, _09725_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_09728_, _09727_, _08065_);
  and (_09729_, _09728_, _09726_);
  nand (_09730_, _09612_, _08944_);
  or (_09731_, _09612_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_09732_, _09731_, _08008_);
  and (_09733_, _09732_, _09730_);
  and (_09734_, _09680_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or (_09735_, _09734_, rst);
  or (_09736_, _09735_, _09733_);
  or (_11197_, _09736_, _09729_);
  and (_09737_, _09606_, _08440_);
  nand (_09738_, _09737_, _08059_);
  or (_09739_, _09737_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_09740_, _09739_, _08065_);
  and (_09741_, _09740_, _09738_);
  nand (_09742_, _09612_, _08937_);
  or (_09743_, _09612_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_09744_, _09743_, _08008_);
  and (_09745_, _09744_, _09742_);
  and (_09746_, _09680_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  or (_09747_, _09746_, rst);
  or (_09748_, _09747_, _09745_);
  or (_11199_, _09748_, _09741_);
  nand (_09749_, _09606_, _08507_);
  and (_09750_, _09749_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  not (_09751_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  nor (_09752_, _08061_, _09751_);
  or (_09753_, _09752_, _08512_);
  and (_09754_, _09753_, _09606_);
  or (_09755_, _09754_, _09750_);
  and (_09756_, _09755_, _08065_);
  nand (_09757_, _09612_, _08930_);
  or (_09758_, _09612_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_09759_, _09758_, _08008_);
  and (_09760_, _09759_, _09757_);
  nor (_09761_, _08007_, _09751_);
  or (_09762_, _09761_, rst);
  or (_09763_, _09762_, _09760_);
  or (_11201_, _09763_, _09756_);
  nand (_09764_, _09628_, _08059_);
  or (_09765_, _09628_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and (_09766_, _09765_, _08065_);
  and (_09767_, _09766_, _09764_);
  and (_09768_, _09630_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and (_09769_, _09628_, _08976_);
  or (_09770_, _09769_, _09768_);
  and (_09771_, _09770_, _08008_);
  and (_09772_, _09680_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  or (_09773_, _09772_, rst);
  or (_09774_, _09773_, _09771_);
  or (_11203_, _09774_, _09767_);
  and (_09775_, _09621_, _08173_);
  nand (_09776_, _09775_, _08059_);
  or (_09777_, _09775_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_09778_, _09777_, _08065_);
  and (_09779_, _09778_, _09776_);
  and (_09780_, _09630_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  nor (_09781_, _09630_, _08967_);
  or (_09782_, _09781_, _09780_);
  and (_09783_, _09782_, _08008_);
  and (_09784_, _09680_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  or (_09785_, _09784_, rst);
  or (_09786_, _09785_, _09783_);
  or (_11205_, _09786_, _09779_);
  and (_09787_, _09621_, _08237_);
  nand (_09788_, _09787_, _08059_);
  or (_09789_, _09787_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_09790_, _09789_, _08065_);
  and (_09791_, _09790_, _09788_);
  not (_09792_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  nor (_09793_, _09628_, _09792_);
  nor (_09794_, _09630_, _08960_);
  or (_09795_, _09794_, _09793_);
  and (_09796_, _09795_, _08008_);
  nor (_09797_, _08007_, _09792_);
  or (_09798_, _09797_, rst);
  or (_09799_, _09798_, _09796_);
  or (_11207_, _09799_, _09791_);
  and (_09800_, _09621_, _08296_);
  nand (_09801_, _09800_, _08059_);
  or (_09802_, _09800_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_09803_, _09802_, _08065_);
  and (_09804_, _09803_, _09801_);
  and (_09805_, _09630_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  nor (_09806_, _09630_, _08952_);
  or (_09807_, _09806_, _09805_);
  and (_09808_, _09807_, _08008_);
  and (_09809_, _09680_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or (_09810_, _09809_, rst);
  or (_09811_, _09810_, _09808_);
  or (_11209_, _09811_, _09804_);
  and (_09812_, _09621_, _08363_);
  nand (_09813_, _09812_, _08059_);
  or (_09814_, _09812_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_09815_, _09814_, _08065_);
  and (_09816_, _09815_, _09813_);
  and (_09817_, _09630_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  nor (_09818_, _09630_, _08944_);
  or (_09819_, _09818_, _09817_);
  and (_09820_, _09819_, _08008_);
  and (_09821_, _09680_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  or (_09822_, _09821_, rst);
  or (_09823_, _09822_, _09820_);
  or (_11211_, _09823_, _09816_);
  and (_09824_, _09621_, _08440_);
  nand (_09825_, _09824_, _08059_);
  or (_09826_, _09824_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_09827_, _09826_, _08065_);
  and (_09828_, _09827_, _09825_);
  and (_09829_, _09630_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  nor (_09830_, _09630_, _08937_);
  or (_09831_, _09830_, _09829_);
  and (_09832_, _09831_, _08008_);
  and (_09833_, _09680_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  or (_09834_, _09833_, rst);
  or (_09835_, _09834_, _09832_);
  or (_11213_, _09835_, _09828_);
  and (_09836_, _09621_, _08510_);
  nand (_09837_, _09836_, _08059_);
  or (_09838_, _09836_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_09839_, _09838_, _08065_);
  and (_09840_, _09839_, _09837_);
  and (_09841_, _09630_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  nor (_09842_, _09630_, _08930_);
  or (_09843_, _09842_, _09841_);
  and (_09844_, _09843_, _08008_);
  and (_09845_, _09680_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  or (_09846_, _09845_, rst);
  or (_09847_, _09846_, _09844_);
  or (_11215_, _09847_, _09840_);
  nand (_09848_, _09644_, _08059_);
  or (_09849_, _09644_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and (_09850_, _09849_, _08065_);
  and (_09851_, _09850_, _09848_);
  and (_09852_, _09644_, _08976_);
  and (_09853_, _09645_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  or (_09854_, _09853_, _09852_);
  and (_09855_, _09854_, _08008_);
  and (_09856_, _09680_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  or (_09857_, _09856_, rst);
  or (_09858_, _09857_, _09855_);
  or (_11217_, _09858_, _09851_);
  and (_09859_, _09638_, _08173_);
  nand (_09860_, _09859_, _08059_);
  or (_09861_, _09859_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_09862_, _09861_, _08065_);
  and (_09863_, _09862_, _09860_);
  nor (_09864_, _09645_, _08967_);
  and (_09865_, _09645_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or (_09866_, _09865_, _09864_);
  and (_09867_, _09866_, _08008_);
  and (_09868_, _09680_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or (_09869_, _09868_, rst);
  or (_09870_, _09869_, _09867_);
  or (_11219_, _09870_, _09863_);
  and (_09871_, _09638_, _08237_);
  nand (_09872_, _09871_, _08059_);
  or (_09873_, _09871_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_09874_, _09873_, _08065_);
  and (_09875_, _09874_, _09872_);
  nor (_09876_, _09645_, _08960_);
  not (_09877_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  nor (_09878_, _09644_, _09877_);
  or (_09879_, _09878_, _09876_);
  and (_09880_, _09879_, _08008_);
  nor (_09881_, _08007_, _09877_);
  or (_09882_, _09881_, rst);
  or (_09883_, _09882_, _09880_);
  or (_11221_, _09883_, _09875_);
  and (_09884_, _09638_, _08296_);
  nand (_09885_, _09884_, _08059_);
  or (_09886_, _09884_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_09887_, _09886_, _08065_);
  and (_09888_, _09887_, _09885_);
  nor (_09889_, _09645_, _08952_);
  and (_09890_, _09645_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_09891_, _09890_, _09889_);
  and (_09892_, _09891_, _08008_);
  and (_09893_, _09680_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_09894_, _09893_, rst);
  or (_09895_, _09894_, _09892_);
  or (_11223_, _09895_, _09888_);
  and (_09896_, _09638_, _08363_);
  nand (_09897_, _09896_, _08059_);
  or (_09898_, _09896_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_09899_, _09898_, _08065_);
  and (_09900_, _09899_, _09897_);
  nor (_09901_, _09645_, _08944_);
  and (_09902_, _09645_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or (_09903_, _09902_, _09901_);
  and (_09904_, _09903_, _08008_);
  and (_09905_, _09680_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or (_09906_, _09905_, rst);
  or (_09907_, _09906_, _09904_);
  or (_11225_, _09907_, _09900_);
  and (_09908_, _09638_, _08440_);
  nand (_09909_, _09908_, _08059_);
  or (_09910_, _09908_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_09911_, _09910_, _08065_);
  and (_09912_, _09911_, _09909_);
  nor (_09913_, _09645_, _08937_);
  and (_09914_, _09645_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or (_09915_, _09914_, _09913_);
  and (_09916_, _09915_, _08008_);
  and (_09917_, _09680_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or (_09918_, _09917_, rst);
  or (_09919_, _09918_, _09916_);
  or (_11227_, _09919_, _09912_);
  and (_09920_, _09638_, _08510_);
  nand (_09921_, _09920_, _08059_);
  or (_09922_, _09920_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_09923_, _09922_, _08065_);
  and (_09924_, _09923_, _09921_);
  nor (_09925_, _09645_, _08930_);
  and (_09926_, _09645_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or (_09927_, _09926_, _09925_);
  and (_09928_, _09927_, _08008_);
  and (_09929_, _09680_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or (_09930_, _09929_, rst);
  or (_09931_, _09930_, _09928_);
  or (_11229_, _09931_, _09924_);
  nand (_09932_, _08059_, _07763_);
  or (_09933_, _07763_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and (_09934_, _09933_, _09654_);
  and (_09935_, _09934_, _09932_);
  not (_09936_, _09654_);
  and (_09937_, _09936_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  or (_09938_, _09937_, _09935_);
  and (_09939_, _09938_, _08065_);
  and (_09940_, _09666_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and (_09941_, _09664_, _08976_);
  or (_09942_, _09941_, _09940_);
  and (_09943_, _09942_, _08008_);
  and (_09944_, _09680_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  or (_09945_, _09944_, rst);
  or (_09946_, _09945_, _09943_);
  or (_11231_, _09946_, _09939_);
  and (_09947_, _09534_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or (_09948_, _09947_, _09535_);
  and (_09949_, _09948_, _09654_);
  and (_09950_, _09936_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or (_09951_, _09950_, _09949_);
  and (_09952_, _09951_, _08065_);
  and (_09953_, _09666_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  nor (_09954_, _09666_, _08967_);
  or (_09955_, _09954_, _09953_);
  and (_09956_, _09955_, _08008_);
  and (_09957_, _09680_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or (_09958_, _09957_, rst);
  or (_09959_, _09958_, _09956_);
  or (_11233_, _09959_, _09952_);
  not (_09960_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  nor (_09961_, _08237_, _09960_);
  or (_09962_, _09961_, _08238_);
  and (_09963_, _09962_, _09654_);
  nor (_09964_, _09654_, _09960_);
  or (_09965_, _09964_, _09963_);
  and (_09966_, _09965_, _08065_);
  nor (_09967_, _09664_, _09960_);
  nor (_09968_, _09666_, _08960_);
  or (_09969_, _09968_, _09967_);
  and (_09970_, _09969_, _08008_);
  nor (_09971_, _08007_, _09960_);
  or (_09972_, _09971_, rst);
  or (_09973_, _09972_, _09970_);
  or (_11235_, _09973_, _09966_);
  and (_09974_, _08297_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_09975_, _09974_, _08298_);
  and (_09976_, _09975_, _09654_);
  and (_09977_, _09936_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_09978_, _09977_, _09976_);
  and (_09979_, _09978_, _08065_);
  and (_09980_, _09666_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  nor (_09981_, _09666_, _08952_);
  or (_09982_, _09981_, _09980_);
  and (_09983_, _09982_, _08008_);
  and (_09984_, _09680_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_09985_, _09984_, rst);
  or (_09986_, _09985_, _09983_);
  or (_11237_, _09986_, _09979_);
  and (_09987_, _08368_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or (_09988_, _09987_, _08369_);
  and (_09989_, _09988_, _09654_);
  and (_09990_, _09936_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or (_09991_, _09990_, _09989_);
  and (_09992_, _09991_, _08065_);
  and (_09993_, _09666_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  nor (_09994_, _09666_, _08944_);
  or (_09995_, _09994_, _09993_);
  and (_09996_, _09995_, _08008_);
  and (_09997_, _09680_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or (_09998_, _09997_, rst);
  or (_09999_, _09998_, _09996_);
  or (_11239_, _09999_, _09992_);
  and (_10000_, _08441_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or (_10001_, _10000_, _08442_);
  and (_10002_, _10001_, _09654_);
  and (_10003_, _09936_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or (_10004_, _10003_, _10002_);
  and (_10005_, _10004_, _08065_);
  and (_10006_, _09666_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  nor (_10007_, _09666_, _08937_);
  or (_10008_, _10007_, _10006_);
  and (_10009_, _10008_, _08008_);
  and (_10010_, _09680_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or (_10011_, _10010_, rst);
  or (_10012_, _10011_, _10009_);
  or (_11241_, _10012_, _10005_);
  and (_10013_, _08511_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or (_10014_, _10013_, _08512_);
  and (_10015_, _10014_, _09654_);
  and (_10016_, _09936_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or (_10017_, _10016_, _10015_);
  and (_10018_, _10017_, _08065_);
  and (_10019_, _09666_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  nor (_10020_, _09666_, _08930_);
  or (_10021_, _10020_, _10019_);
  and (_10022_, _10021_, _08008_);
  and (_10023_, _09680_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or (_10024_, _10023_, rst);
  or (_10025_, _10024_, _10022_);
  or (_11243_, _10025_, _10018_);
  and (_10026_, _07694_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_10027_, _10026_, _09489_);
  nor (_10028_, _07761_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_10029_, _10028_, _10027_);
  not (_10030_, _10029_);
  and (_10031_, _08848_, _08838_);
  not (_10032_, _08823_);
  and (_10033_, _10032_, _08785_);
  nor (_10034_, _08831_, _08805_);
  nor (_10035_, _08814_, _08809_);
  and (_10036_, _10035_, _10034_);
  and (_10037_, _08839_, _08818_);
  and (_10038_, _10037_, _10036_);
  and (_10039_, _10038_, _10033_);
  nor (_10040_, _10039_, _08522_);
  nor (_10041_, _10040_, _10031_);
  not (_10042_, _10041_);
  and (_10043_, _08900_, _08860_);
  and (_10044_, _10043_, _08911_);
  not (_10045_, _07711_);
  and (_10046_, _09389_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  nor (_10047_, _10046_, _09447_);
  nor (_10048_, _10047_, _10045_);
  not (_10049_, _10048_);
  and (_10050_, _10047_, _10045_);
  nor (_10051_, _08643_, _07738_);
  and (_10052_, _08643_, _07738_);
  nor (_10053_, _10052_, _10051_);
  and (_10054_, _08005_, _07692_);
  not (_10055_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and (_10056_, _07762_, _10055_);
  and (_10057_, _10056_, _10054_);
  not (_10058_, _10057_);
  nor (_10059_, _10058_, _10053_);
  not (_10060_, _10059_);
  nor (_10061_, _10060_, _10050_);
  and (_10062_, _10061_, _10049_);
  not (_10063_, _10062_);
  nor (_10064_, _10063_, _08960_);
  nor (_10065_, _10026_, _10045_);
  and (_10066_, _10026_, _07666_);
  nor (_10067_, _10066_, _10065_);
  nor (_10068_, _10067_, _10047_);
  not (_10069_, _10068_);
  and (_10070_, _10067_, _10047_);
  and (_10071_, _10026_, _10045_);
  nor (_10072_, _07738_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_10073_, _10072_, _10071_);
  and (_10074_, _10073_, _08644_);
  nor (_10075_, _10073_, _08644_);
  nor (_10076_, _10075_, _10074_);
  and (_10077_, _10026_, _07724_);
  nor (_10078_, _07749_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_10079_, _10078_, _10077_);
  and (_10080_, _10079_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and (_10081_, _10080_, _10029_);
  and (_10082_, _10081_, _10076_);
  not (_10083_, _10082_);
  nor (_10084_, _10083_, _10070_);
  and (_10085_, _10084_, _10069_);
  not (_10086_, _10085_);
  and (_10087_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , _07827_);
  nand (_10088_, _10087_, _07835_);
  nor (_10089_, _10088_, _08059_);
  nor (_10090_, _08960_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_10091_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_10092_, _10087_, _07828_);
  or (_10093_, _10092_, _10091_);
  and (_10094_, _10087_, _07837_);
  or (_10095_, _10094_, _10093_);
  and (_10096_, _10095_, _06969_);
  or (_10097_, _10096_, _10090_);
  or (_10098_, _10097_, _10089_);
  or (_10099_, _10098_, _10086_);
  nor (_10100_, _10047_, _08643_);
  and (_10101_, _10100_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  and (_10102_, _10047_, _08644_);
  and (_10103_, _10102_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  or (_10104_, _10103_, _10101_);
  and (_10105_, _10047_, _08643_);
  and (_10106_, _10105_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  nor (_10107_, _10047_, _08644_);
  and (_10108_, _10107_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  or (_10109_, _10108_, _10106_);
  or (_10110_, _10109_, _10104_);
  or (_10111_, _10110_, _10085_);
  and (_10112_, _10111_, _10063_);
  and (_10113_, _10112_, _10099_);
  or (_10114_, _10113_, _10064_);
  and (_10115_, _10114_, _10044_);
  not (_10116_, _10115_);
  and (_10117_, _08900_, _08861_);
  and (_10118_, _10117_, _08911_);
  not (_10119_, _09019_);
  and (_10120_, _10119_, _10118_);
  not (_10121_, _10120_);
  not (_10122_, _08911_);
  nor (_10123_, _10122_, _08900_);
  and (_10124_, _10123_, _08860_);
  and (_10125_, _10124_, _08571_);
  nor (_10126_, _08900_, _08860_);
  and (_10127_, _10126_, _08911_);
  not (_10128_, _08527_);
  and (_10129_, _10128_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [2]);
  nor (_10130_, _08533_, _10128_);
  not (_10131_, _10130_);
  and (_10132_, _08545_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_10133_, _08548_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nor (_10134_, _10133_, _10132_);
  and (_10135_, _08552_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  and (_10136_, _08541_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_10137_, _10136_, _10135_);
  and (_10138_, _08557_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_10139_, _08537_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_10140_, _10139_, _10138_);
  and (_10141_, _10140_, _10137_);
  and (_10142_, _10141_, _10134_);
  nor (_10143_, _10142_, _10131_);
  nor (_10144_, _10143_, _10129_);
  not (_10145_, _10144_);
  and (_10146_, _10145_, _10127_);
  nor (_10147_, _10146_, _10125_);
  and (_10148_, _10147_, _10121_);
  and (_10149_, _10148_, _10116_);
  nor (_10150_, _10149_, _10042_);
  nor (_10151_, _10063_, _08937_);
  and (_10152_, _07838_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  not (_10153_, _10152_);
  and (_10154_, _06922_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_10155_, _10154_, _10153_);
  and (_10156_, _10091_, _07838_);
  and (_10157_, _10156_, _08113_);
  nor (_10158_, _08937_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  or (_10159_, _10158_, _10157_);
  nor (_10160_, _10159_, _10155_);
  and (_10161_, _10160_, _10085_);
  and (_10162_, _10107_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  and (_10163_, _10102_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  nor (_10164_, _10163_, _10162_);
  and (_10165_, _10100_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  and (_10166_, _10105_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nor (_10167_, _10166_, _10165_);
  and (_10168_, _10167_, _10164_);
  and (_10169_, _10168_, _10086_);
  nor (_10170_, _10169_, _10062_);
  not (_10171_, _10170_);
  nor (_10172_, _10171_, _10161_);
  or (_10173_, _10172_, _10151_);
  nand (_10174_, _10173_, _10044_);
  not (_10175_, _09037_);
  and (_10176_, _10175_, _10118_);
  not (_10177_, _10176_);
  and (_10178_, _10128_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [5]);
  and (_10179_, _08545_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_10180_, _08548_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  nor (_10181_, _10180_, _10179_);
  and (_10182_, _08557_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_10183_, _08537_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_10184_, _10183_, _10182_);
  and (_10185_, _08552_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  and (_10186_, _08541_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_10187_, _10186_, _10185_);
  and (_10188_, _10187_, _10184_);
  and (_10189_, _10188_, _10181_);
  nor (_10190_, _10189_, _10131_);
  nor (_10191_, _10190_, _10178_);
  not (_10192_, _10191_);
  and (_10193_, _10192_, _10127_);
  not (_10194_, _10126_);
  nor (_10195_, _10043_, _08911_);
  and (_10196_, _10195_, _10194_);
  nor (_10197_, _10196_, _10193_);
  and (_10198_, _10197_, _10177_);
  and (_10199_, _10198_, _10174_);
  not (_10200_, _10199_);
  nand (_10201_, _08804_, _08836_);
  not (_10202_, _08849_);
  and (_10203_, _10202_, _10201_);
  not (_10204_, _08848_);
  nor (_10205_, _10204_, _10203_);
  not (_10206_, _08783_);
  nor (_10207_, _08746_, _08670_);
  and (_10208_, _10207_, _08720_);
  and (_10209_, _10208_, _08804_);
  nor (_10210_, _10209_, _08809_);
  and (_10211_, _10210_, _10206_);
  and (_10212_, _10211_, _10032_);
  and (_10213_, _10208_, _08770_);
  not (_10214_, _10213_);
  and (_10215_, _10214_, _10203_);
  and (_10216_, _10207_, _08763_);
  and (_10217_, _08804_, _10216_);
  not (_10218_, _10217_);
  and (_10219_, _08796_, _08753_);
  and (_10220_, _10219_, _08770_);
  nor (_10221_, _10220_, _08816_);
  and (_10222_, _10221_, _10218_);
  and (_10223_, _10222_, _10215_);
  and (_10224_, _10223_, _10212_);
  and (_10225_, _10224_, _10034_);
  nor (_10226_, _10225_, _08522_);
  nor (_10227_, _10226_, _10205_);
  not (_10228_, _07828_);
  and (_10229_, _10091_, _10228_);
  nor (_10230_, _10229_, _10087_);
  not (_10231_, _10230_);
  and (_10232_, _10231_, _06953_);
  and (_10233_, _10091_, _07828_);
  and (_10234_, _10233_, _08113_);
  nor (_10235_, _08997_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  or (_10236_, _10235_, _10234_);
  or (_10237_, _10236_, _10232_);
  nor (_10238_, _10237_, _10086_);
  and (_10239_, _10102_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  and (_10240_, _10107_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  nor (_10241_, _10240_, _10239_);
  and (_10242_, _10100_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  and (_10243_, _10105_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  nor (_10244_, _10243_, _10242_);
  and (_10245_, _10244_, _10241_);
  and (_10246_, _10245_, _10086_);
  or (_10247_, _10246_, _10238_);
  and (_10248_, _10247_, _10063_);
  and (_10249_, _10062_, _08997_);
  nor (_10250_, _10249_, _10248_);
  nand (_10251_, _10250_, _10044_);
  and (_10252_, _10128_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [7]);
  and (_10253_, _08545_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_10254_, _08548_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nor (_10255_, _10254_, _10253_);
  and (_10256_, _08557_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_10257_, _08537_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_10258_, _10257_, _10256_);
  and (_10259_, _08552_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  and (_10260_, _08541_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor (_10261_, _10260_, _10259_);
  and (_10262_, _10261_, _10258_);
  and (_10263_, _10262_, _10255_);
  nor (_10264_, _10263_, _10131_);
  nor (_10265_, _10264_, _10252_);
  not (_10266_, _10265_);
  and (_10267_, _10266_, _10126_);
  nor (_10268_, _10267_, _10122_);
  nand (_10269_, _08999_, _10117_);
  and (_10270_, _10269_, _10268_);
  and (_10271_, _10270_, _10251_);
  not (_10272_, _10271_);
  nor (_10273_, _10272_, _10227_);
  and (_10274_, _10273_, _10200_);
  nor (_10275_, _10274_, _10150_);
  and (_10276_, _10275_, _10030_);
  not (_10277_, _10073_);
  and (_10278_, _10062_, _08976_);
  and (_10279_, _10087_, _07831_);
  not (_10280_, _10279_);
  nor (_10281_, _10280_, _08059_);
  not (_10282_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand (_10283_, _08975_, _10282_);
  or (_10284_, _06990_, _10282_);
  and (_10285_, _10284_, _10280_);
  and (_10286_, _10285_, _10283_);
  or (_10287_, _10286_, _10281_);
  or (_10288_, _10287_, _10086_);
  and (_10289_, _10105_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  and (_10290_, _10107_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  or (_10291_, _10290_, _10289_);
  and (_10292_, _10100_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  and (_10293_, _10102_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  or (_10294_, _10293_, _10292_);
  or (_10295_, _10294_, _10291_);
  or (_10296_, _10295_, _10085_);
  and (_10297_, _10296_, _10063_);
  and (_10298_, _10297_, _10288_);
  or (_10299_, _10298_, _10278_);
  and (_10300_, _10299_, _10044_);
  not (_10301_, _10300_);
  not (_10302_, _09007_);
  and (_10303_, _10302_, _10118_);
  not (_10304_, _10303_);
  and (_10305_, _10124_, _08644_);
  and (_10306_, _10128_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [0]);
  and (_10307_, _08545_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_10308_, _08548_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nor (_10309_, _10308_, _10307_);
  and (_10310_, _08541_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  and (_10311_, _08537_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_10312_, _10311_, _10310_);
  and (_10313_, _08552_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  and (_10314_, _08557_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor (_10315_, _10314_, _10313_);
  and (_10316_, _10315_, _10312_);
  and (_10317_, _10316_, _10309_);
  nor (_10318_, _10317_, _10131_);
  nor (_10319_, _10318_, _10306_);
  not (_10320_, _10319_);
  and (_10321_, _10320_, _10127_);
  nor (_10322_, _10321_, _10305_);
  and (_10323_, _10322_, _10304_);
  and (_10324_, _10323_, _10301_);
  nor (_10325_, _10324_, _10042_);
  not (_10326_, _08952_);
  and (_10327_, _10062_, _10326_);
  and (_10328_, _10092_, _08113_);
  nor (_10329_, _08952_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_10330_, _10087_, _10228_);
  or (_10331_, _10330_, _10091_);
  and (_10332_, _10331_, _06904_);
  or (_10333_, _10332_, _10329_);
  or (_10334_, _10333_, _10328_);
  or (_10335_, _10334_, _10086_);
  and (_10336_, _10105_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  and (_10337_, _10107_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  or (_10338_, _10337_, _10336_);
  and (_10339_, _10100_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  and (_10340_, _10102_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  or (_10341_, _10340_, _10339_);
  or (_10342_, _10341_, _10338_);
  or (_10343_, _10342_, _10085_);
  and (_10344_, _10343_, _10063_);
  and (_10345_, _10344_, _10335_);
  or (_10346_, _10345_, _10327_);
  and (_10347_, _10346_, _10044_);
  not (_10348_, _10347_);
  not (_10349_, _09025_);
  and (_10350_, _10349_, _10118_);
  not (_10351_, _10350_);
  not (_10352_, _10047_);
  and (_10353_, _10124_, _10352_);
  and (_10354_, _10128_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [3]);
  and (_10355_, _08545_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_10356_, _08548_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nor (_10357_, _10356_, _10355_);
  and (_10358_, _08541_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  and (_10359_, _08537_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_10360_, _10359_, _10358_);
  and (_10361_, _08552_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  and (_10362_, _08557_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor (_10363_, _10362_, _10361_);
  and (_10364_, _10363_, _10360_);
  and (_10365_, _10364_, _10357_);
  nor (_10366_, _10365_, _10131_);
  nor (_10367_, _10366_, _10354_);
  not (_10368_, _10367_);
  and (_10369_, _10368_, _10127_);
  nor (_10370_, _10369_, _10353_);
  and (_10371_, _10370_, _10351_);
  and (_10372_, _10371_, _10348_);
  not (_10373_, _10372_);
  and (_10374_, _10373_, _10273_);
  nor (_10375_, _10374_, _10325_);
  nor (_10376_, _10375_, _10277_);
  nor (_10377_, _10376_, _10276_);
  nor (_10378_, _10275_, _10030_);
  not (_10379_, _10378_);
  not (_10380_, _10067_);
  and (_10381_, _10271_, _10042_);
  nor (_10382_, _10373_, _10381_);
  not (_10383_, _08930_);
  and (_10384_, _10062_, _10383_);
  and (_10385_, _07835_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  not (_10386_, _10385_);
  and (_10387_, _07006_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_10388_, _10387_, _10386_);
  and (_10389_, _10091_, _07835_);
  and (_10390_, _10389_, _08113_);
  nor (_10391_, _08930_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  or (_10392_, _10391_, _10390_);
  nor (_10393_, _10392_, _10388_);
  and (_10394_, _10393_, _10085_);
  and (_10395_, _10105_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  and (_10396_, _10107_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  nor (_10397_, _10396_, _10395_);
  and (_10398_, _10100_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  and (_10399_, _10102_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  nor (_10400_, _10399_, _10398_);
  and (_10401_, _10400_, _10397_);
  and (_10402_, _10401_, _10086_);
  nor (_10403_, _10402_, _10062_);
  not (_10404_, _10403_);
  nor (_10405_, _10404_, _10394_);
  or (_10406_, _10405_, _10384_);
  nand (_10407_, _10406_, _10044_);
  not (_10408_, _09043_);
  and (_10409_, _10408_, _10118_);
  and (_10410_, _10128_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [6]);
  and (_10411_, _08545_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_10412_, _08548_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nor (_10413_, _10412_, _10411_);
  and (_10414_, _08557_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_10415_, _08537_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_10416_, _10415_, _10414_);
  and (_10417_, _08552_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  and (_10418_, _08541_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor (_10419_, _10418_, _10417_);
  and (_10420_, _10419_, _10416_);
  and (_10421_, _10420_, _10413_);
  nor (_10422_, _10421_, _10131_);
  nor (_10423_, _10422_, _10410_);
  not (_10424_, _10423_);
  and (_10425_, _10424_, _10126_);
  nor (_10426_, _10425_, _10195_);
  not (_10427_, _10426_);
  nor (_10428_, _10427_, _10409_);
  and (_10429_, _10428_, _10407_);
  and (_10430_, _10429_, _10381_);
  nor (_10431_, _10430_, _10382_);
  nor (_10432_, _10431_, _10380_);
  and (_10433_, _10431_, _10380_);
  nor (_10434_, _10433_, _10432_);
  and (_10435_, _10434_, _10379_);
  not (_10436_, _08967_);
  and (_10437_, _10062_, _10436_);
  nand (_10438_, _10087_, _07838_);
  nor (_10439_, _10438_, _08059_);
  nor (_10440_, _08967_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_10441_, _10087_, _07834_);
  or (_10442_, _10093_, _10441_);
  and (_10443_, _10442_, _06937_);
  or (_10444_, _10443_, _10440_);
  or (_10445_, _10444_, _10439_);
  or (_10446_, _10445_, _10086_);
  and (_10447_, _10105_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  and (_10448_, _10107_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  or (_10449_, _10448_, _10447_);
  and (_10450_, _10100_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  and (_10451_, _10102_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  or (_10452_, _10451_, _10450_);
  or (_10453_, _10452_, _10449_);
  or (_10454_, _10453_, _10085_);
  and (_10455_, _10454_, _10063_);
  and (_10456_, _10455_, _10446_);
  or (_10457_, _10456_, _10437_);
  and (_10458_, _10457_, _10044_);
  not (_10459_, _10458_);
  not (_10460_, _09013_);
  and (_10461_, _10460_, _10118_);
  not (_10462_, _10461_);
  and (_10463_, _10043_, _10122_);
  not (_10464_, _10463_);
  and (_10465_, _10124_, _08749_);
  and (_10466_, _10128_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [1]);
  and (_10467_, _08545_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_10468_, _08548_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor (_10469_, _10468_, _10467_);
  and (_10470_, _08541_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  and (_10471_, _08537_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_10472_, _10471_, _10470_);
  and (_10473_, _08552_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  and (_10474_, _08557_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nor (_10475_, _10474_, _10473_);
  and (_10476_, _10475_, _10472_);
  and (_10477_, _10476_, _10469_);
  nor (_10478_, _10477_, _10131_);
  nor (_10479_, _10478_, _10466_);
  not (_10480_, _10479_);
  and (_10481_, _10480_, _10127_);
  nor (_10482_, _10481_, _10465_);
  and (_10483_, _10482_, _10464_);
  and (_10484_, _10483_, _10462_);
  and (_10485_, _10484_, _10459_);
  nor (_10486_, _10485_, _10042_);
  not (_10487_, _08944_);
  and (_10488_, _10062_, _10487_);
  and (_10489_, _10102_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  and (_10490_, _10107_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  nor (_10491_, _10490_, _10489_);
  and (_10492_, _10105_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  and (_10493_, _10100_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  nor (_10494_, _10493_, _10492_);
  and (_10495_, _10494_, _10491_);
  and (_10496_, _10495_, _10086_);
  and (_10497_, _07831_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  not (_10498_, _10497_);
  and (_10499_, _06883_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_10500_, _10499_, _10498_);
  and (_10501_, _10091_, _07831_);
  and (_10502_, _10501_, _08113_);
  nor (_10503_, _08944_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  or (_10504_, _10503_, _10502_);
  nor (_10505_, _10504_, _10500_);
  and (_10506_, _10505_, _10085_);
  or (_10507_, _10506_, _10062_);
  nor (_10508_, _10507_, _10496_);
  or (_10509_, _10508_, _10488_);
  nand (_10510_, _10509_, _10044_);
  not (_10511_, _09031_);
  and (_10512_, _10511_, _10118_);
  and (_10513_, _10128_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [4]);
  and (_10514_, _08545_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_10515_, _08548_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nor (_10516_, _10515_, _10514_);
  and (_10517_, _08541_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  and (_10518_, _08537_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_10519_, _10518_, _10517_);
  and (_10520_, _08552_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  and (_10521_, _08557_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor (_10522_, _10521_, _10520_);
  and (_10523_, _10522_, _10519_);
  and (_10524_, _10523_, _10516_);
  nor (_10525_, _10524_, _10131_);
  nor (_10526_, _10525_, _10513_);
  not (_10527_, _10526_);
  and (_10528_, _10527_, _10127_);
  nor (_10529_, _10528_, _10512_);
  nor (_10530_, _08911_, _08900_);
  nor (_10531_, _09456_, _09452_);
  not (_10532_, _10531_);
  and (_10533_, _10532_, _10124_);
  or (_10534_, _10533_, _10530_);
  not (_10535_, _10534_);
  and (_10536_, _10535_, _10529_);
  and (_10537_, _10536_, _10510_);
  not (_10538_, _10537_);
  and (_10539_, _10538_, _10273_);
  nor (_10540_, _10539_, _10486_);
  nand (_10541_, _10540_, _10079_);
  or (_10542_, _10540_, _10079_);
  and (_10543_, _10542_, _10541_);
  not (_10544_, _10543_);
  not (_10545_, _10054_);
  and (_10546_, _10375_, _10277_);
  nor (_10547_, _10546_, _10545_);
  and (_10548_, _10547_, _10544_);
  and (_10549_, _10548_, _10435_);
  and (_10550_, _10549_, _10377_);
  not (_10551_, _10275_);
  and (_10552_, _10375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  not (_10553_, _10375_);
  and (_10554_, _10553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  or (_10555_, _10554_, _10552_);
  and (_10556_, _10555_, _10540_);
  not (_10557_, _10540_);
  not (_10558_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  nor (_10559_, _10375_, _10558_);
  and (_10560_, _10375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  or (_10561_, _10560_, _10559_);
  and (_10562_, _10561_, _10557_);
  or (_10563_, _10562_, _10556_);
  or (_10564_, _10563_, _10551_);
  not (_10565_, _10431_);
  and (_10566_, _10375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  and (_10567_, _10553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  or (_10568_, _10567_, _10566_);
  and (_10569_, _10568_, _10540_);
  not (_10570_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  nor (_10571_, _10375_, _10570_);
  and (_10572_, _10375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  or (_10573_, _10572_, _10571_);
  and (_10574_, _10573_, _10557_);
  or (_10575_, _10574_, _10569_);
  or (_10576_, _10575_, _10275_);
  and (_10577_, _10576_, _10565_);
  and (_10578_, _10577_, _10564_);
  or (_10579_, _10553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  or (_10580_, _10375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  and (_10581_, _10580_, _10579_);
  and (_10582_, _10581_, _10540_);
  or (_10583_, _10375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  not (_10584_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  nand (_10585_, _10375_, _10584_);
  and (_10586_, _10585_, _10583_);
  and (_10587_, _10586_, _10557_);
  or (_10588_, _10587_, _10582_);
  or (_10589_, _10588_, _10551_);
  or (_10590_, _10553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  or (_10591_, _10375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  and (_10592_, _10591_, _10590_);
  and (_10593_, _10592_, _10540_);
  or (_10594_, _10375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  not (_10595_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  nand (_10596_, _10375_, _10595_);
  and (_10597_, _10596_, _10594_);
  and (_10598_, _10597_, _10557_);
  or (_10599_, _10598_, _10593_);
  or (_10600_, _10599_, _10275_);
  and (_10601_, _10600_, _10431_);
  and (_10602_, _10601_, _10589_);
  or (_10603_, _10602_, _10578_);
  or (_10604_, _10603_, _10550_);
  not (_10605_, _10550_);
  or (_10606_, _10605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  and (_10607_, _10606_, _13707_);
  and (_11331_, _10607_, _10604_);
  nor (_10608_, _10073_, _10545_);
  nor (_10609_, _10079_, _10545_);
  and (_10610_, _10609_, _10608_);
  nor (_10611_, _10029_, _10545_);
  and (_10612_, _10067_, _10054_);
  and (_10613_, _10612_, _10611_);
  and (_10614_, _10613_, _10610_);
  and (_10615_, _10237_, _10054_);
  and (_10616_, _10615_, _10614_);
  not (_10617_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  nor (_10618_, _10614_, _10617_);
  or (_11343_, _10618_, _10616_);
  nor (_10619_, _10609_, _10608_);
  nor (_10620_, _10612_, _10611_);
  and (_10621_, _10620_, _10054_);
  and (_10622_, _10621_, _10619_);
  and (_10623_, _10287_, _10054_);
  and (_10624_, _10623_, _10622_);
  not (_10625_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  nor (_10626_, _10622_, _10625_);
  or (_11586_, _10626_, _10624_);
  and (_10627_, _10445_, _10054_);
  and (_10628_, _10627_, _10622_);
  not (_10629_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  nor (_10630_, _10622_, _10629_);
  or (_11591_, _10630_, _10628_);
  and (_10631_, _10098_, _10054_);
  and (_10632_, _10631_, _10622_);
  not (_10633_, _10622_);
  and (_10634_, _10633_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  or (_11596_, _10634_, _10632_);
  and (_10635_, _10334_, _10054_);
  and (_10636_, _10635_, _10622_);
  not (_10637_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  nor (_10638_, _10622_, _10637_);
  or (_11601_, _10638_, _10636_);
  nor (_10639_, _10505_, _10545_);
  and (_10640_, _10639_, _10622_);
  and (_10641_, _10633_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  or (_11606_, _10641_, _10640_);
  nor (_10642_, _10160_, _10545_);
  and (_10643_, _10642_, _10622_);
  and (_10644_, _10633_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  or (_11612_, _10644_, _10643_);
  nor (_10645_, _10393_, _10545_);
  and (_10646_, _10645_, _10622_);
  not (_10647_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  nor (_10648_, _10622_, _10647_);
  or (_11617_, _10648_, _10646_);
  and (_10649_, _10622_, _10615_);
  and (_10650_, _10633_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  or (_11619_, _10650_, _10649_);
  and (_10651_, _10608_, _10079_);
  and (_10652_, _10651_, _10620_);
  and (_10653_, _10652_, _10623_);
  not (_10654_, _10652_);
  and (_10655_, _10654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  or (_11626_, _10655_, _10653_);
  and (_10656_, _10652_, _10627_);
  and (_10657_, _10654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  or (_11630_, _10657_, _10656_);
  and (_10658_, _10652_, _10631_);
  and (_10659_, _10654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  or (_11633_, _10659_, _10658_);
  and (_10660_, _10652_, _10635_);
  and (_10661_, _10654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  or (_11637_, _10661_, _10660_);
  and (_10662_, _10652_, _10639_);
  not (_10663_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  nor (_10664_, _10652_, _10663_);
  or (_11640_, _10664_, _10662_);
  and (_10665_, _10652_, _10642_);
  not (_10666_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  nor (_10667_, _10652_, _10666_);
  or (_11644_, _10667_, _10665_);
  and (_10668_, _10652_, _10645_);
  and (_10669_, _10654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  or (_11647_, _10669_, _10668_);
  and (_10670_, _10652_, _10615_);
  and (_10671_, _10654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  or (_11650_, _10671_, _10670_);
  and (_10672_, _10609_, _10073_);
  and (_10673_, _10672_, _10620_);
  and (_10674_, _10673_, _10623_);
  not (_10675_, _10673_);
  and (_10676_, _10675_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  or (_11657_, _10676_, _10674_);
  and (_10677_, _10673_, _10627_);
  and (_10678_, _10675_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  or (_11660_, _10678_, _10677_);
  and (_10679_, _10673_, _10631_);
  not (_10680_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  nor (_10681_, _10673_, _10680_);
  or (_11664_, _10681_, _10679_);
  and (_10682_, _10673_, _10635_);
  not (_10683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  nor (_10684_, _10673_, _10683_);
  or (_11667_, _10684_, _10682_);
  and (_10685_, _10673_, _10639_);
  not (_10686_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  nor (_10687_, _10673_, _10686_);
  or (_11671_, _10687_, _10685_);
  and (_10688_, _10673_, _10642_);
  not (_10689_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  nor (_10690_, _10673_, _10689_);
  or (_11674_, _10690_, _10688_);
  and (_10691_, _10673_, _10645_);
  and (_10692_, _10675_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  or (_11678_, _10692_, _10691_);
  and (_10693_, _10673_, _10615_);
  not (_10694_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  nor (_10695_, _10673_, _10694_);
  or (_11681_, _10695_, _10693_);
  and (_10696_, _10620_, _10610_);
  and (_10697_, _10696_, _10623_);
  not (_10698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  nor (_10699_, _10696_, _10698_);
  or (_11686_, _10699_, _10697_);
  and (_10700_, _10696_, _10627_);
  not (_10701_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  nor (_10702_, _10696_, _10701_);
  or (_11689_, _10702_, _10700_);
  and (_10703_, _10696_, _10631_);
  not (_10704_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  nor (_10705_, _10696_, _10704_);
  or (_11693_, _10705_, _10703_);
  and (_10706_, _10696_, _10635_);
  not (_10707_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  nor (_10708_, _10696_, _10707_);
  or (_11696_, _10708_, _10706_);
  and (_10709_, _10696_, _10639_);
  not (_10710_, _10696_);
  and (_10711_, _10710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  or (_11700_, _10711_, _10709_);
  and (_10712_, _10696_, _10642_);
  and (_10713_, _10710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  or (_11703_, _10713_, _10712_);
  and (_10714_, _10696_, _10645_);
  not (_10715_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  nor (_10716_, _10696_, _10715_);
  or (_11707_, _10716_, _10714_);
  and (_10717_, _10696_, _10615_);
  nor (_10718_, _10696_, _10558_);
  or (_11710_, _10718_, _10717_);
  and (_10719_, _10611_, _10380_);
  and (_10720_, _10719_, _10619_);
  and (_10721_, _10720_, _10623_);
  not (_10722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  nor (_10723_, _10720_, _10722_);
  or (_11716_, _10723_, _10721_);
  and (_10724_, _10720_, _10627_);
  not (_10725_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  nor (_10726_, _10720_, _10725_);
  or (_11720_, _10726_, _10724_);
  and (_10727_, _10720_, _10631_);
  not (_10728_, _10720_);
  and (_10729_, _10728_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  or (_11723_, _10729_, _10727_);
  and (_10730_, _10720_, _10635_);
  and (_10731_, _10728_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  or (_11727_, _10731_, _10730_);
  and (_10732_, _10720_, _10639_);
  and (_10733_, _10728_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  or (_11730_, _10733_, _10732_);
  and (_10734_, _10720_, _10642_);
  and (_10735_, _10728_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  or (_11734_, _10735_, _10734_);
  and (_10736_, _10720_, _10645_);
  not (_10737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  nor (_10738_, _10720_, _10737_);
  or (_11737_, _10738_, _10736_);
  and (_10739_, _10720_, _10615_);
  and (_10740_, _10728_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  or (_11740_, _10740_, _10739_);
  and (_10741_, _10719_, _10651_);
  and (_10742_, _10741_, _10623_);
  not (_10743_, _10741_);
  and (_10744_, _10743_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  or (_11744_, _10744_, _10742_);
  and (_10745_, _10741_, _10627_);
  and (_10746_, _10743_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  or (_11748_, _10746_, _10745_);
  and (_10747_, _10741_, _10631_);
  and (_10748_, _10743_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  or (_11751_, _10748_, _10747_);
  and (_10749_, _10741_, _10635_);
  not (_10750_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  nor (_10751_, _10741_, _10750_);
  or (_11755_, _10751_, _10749_);
  and (_10752_, _10741_, _10639_);
  not (_10753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  nor (_10754_, _10741_, _10753_);
  or (_11758_, _10754_, _10752_);
  and (_10755_, _10741_, _10642_);
  not (_10756_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  nor (_10757_, _10741_, _10756_);
  or (_11762_, _10757_, _10755_);
  and (_10758_, _10741_, _10645_);
  not (_10759_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  nor (_10760_, _10741_, _10759_);
  or (_11766_, _10760_, _10758_);
  and (_10761_, _10741_, _10615_);
  and (_10762_, _10743_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  or (_11768_, _10762_, _10761_);
  and (_10763_, _10719_, _10672_);
  and (_10764_, _10763_, _10623_);
  not (_10765_, _10763_);
  and (_10766_, _10765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  or (_11773_, _10766_, _10764_);
  and (_10767_, _10763_, _10627_);
  and (_10768_, _10765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  or (_11776_, _10768_, _10767_);
  and (_10769_, _10763_, _10631_);
  not (_10770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  nor (_10771_, _10763_, _10770_);
  or (_11780_, _10771_, _10769_);
  and (_10772_, _10763_, _10635_);
  and (_10773_, _10765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or (_11783_, _10773_, _10772_);
  and (_10774_, _10763_, _10639_);
  not (_10775_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  nor (_10776_, _10763_, _10775_);
  or (_11787_, _10776_, _10774_);
  and (_10777_, _10763_, _10642_);
  not (_10778_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  nor (_10779_, _10763_, _10778_);
  or (_11790_, _10779_, _10777_);
  and (_10780_, _10763_, _10645_);
  not (_10781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  nor (_10782_, _10763_, _10781_);
  or (_11794_, _10782_, _10780_);
  and (_10783_, _10763_, _10615_);
  not (_10784_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  nor (_10785_, _10763_, _10784_);
  or (_11796_, _10785_, _10783_);
  and (_10786_, _10719_, _10610_);
  and (_10787_, _10786_, _10623_);
  not (_10788_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  nor (_10789_, _10786_, _10788_);
  or (_11801_, _10789_, _10787_);
  and (_10790_, _10786_, _10627_);
  not (_10791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  nor (_10792_, _10786_, _10791_);
  or (_11804_, _10792_, _10790_);
  and (_10793_, _10786_, _10631_);
  not (_10794_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  nor (_10795_, _10786_, _10794_);
  or (_11808_, _10795_, _10793_);
  and (_10796_, _10786_, _10635_);
  not (_10797_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  nor (_10798_, _10786_, _10797_);
  or (_11811_, _10798_, _10796_);
  and (_10799_, _10786_, _10639_);
  not (_10800_, _10786_);
  and (_10801_, _10800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  or (_11815_, _10801_, _10799_);
  and (_10802_, _10786_, _10642_);
  and (_10803_, _10800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  or (_11818_, _10803_, _10802_);
  and (_10804_, _10786_, _10645_);
  not (_10805_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  nor (_10806_, _10786_, _10805_);
  or (_11822_, _10806_, _10804_);
  and (_10807_, _10786_, _10615_);
  nor (_10808_, _10786_, _10570_);
  or (_11824_, _10808_, _10807_);
  and (_10809_, _10612_, _10029_);
  and (_10810_, _10809_, _10619_);
  and (_10811_, _10810_, _10623_);
  not (_10812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  nor (_10813_, _10810_, _10812_);
  or (_11831_, _10813_, _10811_);
  and (_10814_, _10810_, _10627_);
  not (_10815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  nor (_10816_, _10810_, _10815_);
  or (_11835_, _10816_, _10814_);
  and (_10817_, _10810_, _10631_);
  not (_10818_, _10810_);
  and (_10819_, _10818_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  or (_11838_, _10819_, _10817_);
  and (_10820_, _10810_, _10635_);
  and (_10821_, _10818_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  or (_11842_, _10821_, _10820_);
  and (_10822_, _10810_, _10639_);
  and (_10823_, _10818_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  or (_11845_, _10823_, _10822_);
  and (_10824_, _10810_, _10642_);
  and (_10825_, _10818_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  or (_11849_, _10825_, _10824_);
  and (_10826_, _10810_, _10645_);
  and (_10827_, _10818_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  or (_11852_, _10827_, _10826_);
  and (_10828_, _10810_, _10615_);
  and (_10829_, _10818_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  or (_11855_, _10829_, _10828_);
  and (_10830_, _10809_, _10651_);
  and (_10831_, _10830_, _10623_);
  not (_10832_, _10830_);
  and (_10833_, _10832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  or (_11859_, _10833_, _10831_);
  and (_10834_, _10830_, _10627_);
  and (_10835_, _10832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  or (_11863_, _10835_, _10834_);
  and (_10836_, _10830_, _10631_);
  and (_10837_, _10832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  or (_11866_, _10837_, _10836_);
  and (_10838_, _10830_, _10635_);
  and (_10839_, _10832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  or (_11870_, _10839_, _10838_);
  and (_10840_, _10830_, _10639_);
  not (_10841_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  nor (_10842_, _10830_, _10841_);
  or (_11873_, _10842_, _10840_);
  and (_10843_, _10830_, _10642_);
  not (_10844_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  nor (_10845_, _10830_, _10844_);
  or (_11877_, _10845_, _10843_);
  and (_10846_, _10830_, _10645_);
  and (_10847_, _10832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  or (_11880_, _10847_, _10846_);
  and (_10848_, _10830_, _10615_);
  and (_10849_, _10832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  or (_11883_, _10849_, _10848_);
  and (_10850_, _10809_, _10672_);
  and (_10851_, _10850_, _10623_);
  not (_10852_, _10850_);
  and (_10853_, _10852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  or (_11887_, _10853_, _10851_);
  and (_10854_, _10850_, _10627_);
  and (_10855_, _10852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  or (_11891_, _10855_, _10854_);
  and (_10856_, _10850_, _10631_);
  not (_10857_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  nor (_10858_, _10850_, _10857_);
  or (_11894_, _10858_, _10856_);
  and (_10859_, _10850_, _10635_);
  not (_10860_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  nor (_10861_, _10850_, _10860_);
  or (_11898_, _10861_, _10859_);
  and (_10862_, _10850_, _10639_);
  not (_10863_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  nor (_10864_, _10850_, _10863_);
  or (_11901_, _10864_, _10862_);
  and (_10865_, _10850_, _10642_);
  not (_10866_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  nor (_10867_, _10850_, _10866_);
  or (_11905_, _10867_, _10865_);
  and (_10868_, _10850_, _10645_);
  and (_10869_, _10852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  or (_11908_, _10869_, _10868_);
  and (_10870_, _10850_, _10615_);
  nor (_10871_, _10850_, _10584_);
  or (_11911_, _10871_, _10870_);
  and (_10872_, _10809_, _10610_);
  and (_10873_, _10872_, _10623_);
  not (_10874_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  nor (_10875_, _10872_, _10874_);
  or (_11915_, _10875_, _10873_);
  and (_10876_, _10872_, _10627_);
  not (_10877_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  nor (_10878_, _10872_, _10877_);
  or (_11919_, _10878_, _10876_);
  and (_10879_, _10872_, _10631_);
  not (_10880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  nor (_10881_, _10872_, _10880_);
  or (_11922_, _10881_, _10879_);
  and (_10882_, _10872_, _10635_);
  not (_10883_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  nor (_10884_, _10872_, _10883_);
  or (_11926_, _10884_, _10882_);
  and (_10885_, _10872_, _10639_);
  not (_10886_, _10872_);
  and (_10887_, _10886_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  or (_11929_, _10887_, _10885_);
  and (_10888_, _10872_, _10642_);
  and (_10889_, _10886_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  or (_11933_, _10889_, _10888_);
  and (_10890_, _10872_, _10645_);
  and (_10891_, _10886_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  or (_11937_, _10891_, _10890_);
  and (_10892_, _10872_, _10615_);
  not (_10893_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  nor (_10894_, _10872_, _10893_);
  or (_11939_, _10894_, _10892_);
  and (_10895_, _10619_, _10613_);
  and (_10896_, _10895_, _10623_);
  not (_10897_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  nor (_10898_, _10895_, _10897_);
  or (_11944_, _10898_, _10896_);
  and (_10899_, _10895_, _10627_);
  not (_10900_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  nor (_10901_, _10895_, _10900_);
  or (_11948_, _10901_, _10899_);
  and (_10902_, _10895_, _10631_);
  not (_10903_, _10895_);
  and (_10904_, _10903_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  or (_11951_, _10904_, _10902_);
  and (_10905_, _10895_, _10635_);
  and (_10906_, _10903_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  or (_11955_, _10906_, _10905_);
  and (_10907_, _10895_, _10639_);
  and (_10908_, _10903_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  or (_11958_, _10908_, _10907_);
  and (_10909_, _10895_, _10642_);
  and (_10910_, _10903_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  or (_11962_, _10910_, _10909_);
  and (_10911_, _10895_, _10645_);
  not (_10912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  nor (_10913_, _10895_, _10912_);
  or (_11965_, _10913_, _10911_);
  and (_10914_, _10895_, _10615_);
  and (_10915_, _10903_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  or (_11968_, _10915_, _10914_);
  and (_10916_, _10651_, _10613_);
  and (_10917_, _10916_, _10623_);
  not (_10918_, _10916_);
  and (_10919_, _10918_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  or (_11972_, _10919_, _10917_);
  and (_10920_, _10916_, _10627_);
  and (_10921_, _10918_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  or (_11976_, _10921_, _10920_);
  and (_10922_, _10916_, _10631_);
  and (_10923_, _10918_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  or (_11979_, _10923_, _10922_);
  and (_10924_, _10916_, _10635_);
  and (_10925_, _10918_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  or (_11983_, _10925_, _10924_);
  and (_10926_, _10916_, _10639_);
  not (_10927_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  nor (_10928_, _10916_, _10927_);
  or (_11986_, _10928_, _10926_);
  and (_10929_, _10916_, _10642_);
  not (_10930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  nor (_10931_, _10916_, _10930_);
  or (_11990_, _10931_, _10929_);
  and (_10932_, _10916_, _10645_);
  not (_10933_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  nor (_10934_, _10916_, _10933_);
  or (_11994_, _10934_, _10932_);
  and (_10935_, _10916_, _10615_);
  and (_10936_, _10918_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  or (_11996_, _10936_, _10935_);
  and (_10937_, _10672_, _10613_);
  and (_10938_, _10937_, _10623_);
  not (_10939_, _10937_);
  and (_10940_, _10939_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  or (_12001_, _10940_, _10938_);
  and (_10941_, _10937_, _10627_);
  and (_10942_, _10939_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  or (_12004_, _10942_, _10941_);
  and (_10943_, _10937_, _10631_);
  not (_10944_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  nor (_10945_, _10937_, _10944_);
  or (_12008_, _10945_, _10943_);
  and (_10946_, _10937_, _10635_);
  and (_10947_, _10939_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  or (_12011_, _10947_, _10946_);
  and (_10948_, _10937_, _10639_);
  not (_10949_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  nor (_10950_, _10937_, _10949_);
  or (_12015_, _10950_, _10948_);
  and (_10951_, _10937_, _10642_);
  not (_10952_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  nor (_10953_, _10937_, _10952_);
  or (_12018_, _10953_, _10951_);
  and (_10954_, _10937_, _10645_);
  not (_10955_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  nor (_10956_, _10937_, _10955_);
  or (_12022_, _10956_, _10954_);
  and (_10957_, _10937_, _10615_);
  nor (_10958_, _10937_, _10595_);
  or (_12024_, _10958_, _10957_);
  and (_10959_, _10623_, _10614_);
  not (_10960_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  nor (_10961_, _10614_, _10960_);
  or (_12029_, _10961_, _10959_);
  and (_10962_, _10627_, _10614_);
  not (_10963_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  nor (_10964_, _10614_, _10963_);
  or (_12032_, _10964_, _10962_);
  and (_10965_, _10631_, _10614_);
  not (_10966_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  nor (_10967_, _10614_, _10966_);
  or (_12036_, _10967_, _10965_);
  and (_10968_, _10635_, _10614_);
  not (_10969_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  nor (_10970_, _10614_, _10969_);
  or (_12039_, _10970_, _10968_);
  and (_10971_, _10639_, _10614_);
  not (_10972_, _10614_);
  and (_10973_, _10972_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  or (_12043_, _10973_, _10971_);
  and (_10974_, _10642_, _10614_);
  and (_10975_, _10972_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  or (_12046_, _10975_, _10974_);
  and (_10976_, _10645_, _10614_);
  not (_10977_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  nor (_10978_, _10614_, _10977_);
  or (_12050_, _10978_, _10976_);
  or (_10979_, _10375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  nand (_10980_, _10375_, _10625_);
  and (_10981_, _10980_, _10540_);
  and (_10982_, _10981_, _10979_);
  nor (_10983_, _10375_, _10698_);
  and (_10984_, _10375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  or (_10985_, _10984_, _10983_);
  and (_10986_, _10985_, _10557_);
  or (_10987_, _10986_, _10982_);
  or (_10988_, _10987_, _10551_);
  or (_10989_, _10375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  nand (_10990_, _10375_, _10722_);
  and (_10991_, _10990_, _10540_);
  and (_10992_, _10991_, _10989_);
  nor (_10993_, _10375_, _10788_);
  and (_10994_, _10375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  or (_10995_, _10994_, _10993_);
  and (_10996_, _10995_, _10557_);
  or (_10997_, _10996_, _10992_);
  or (_10998_, _10997_, _10275_);
  and (_10999_, _10998_, _10565_);
  and (_11000_, _10999_, _10988_);
  nand (_11001_, _10375_, _10812_);
  or (_11002_, _10375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  and (_11003_, _11002_, _11001_);
  and (_11004_, _11003_, _10540_);
  and (_11005_, _10375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  nor (_11006_, _10375_, _10874_);
  or (_11007_, _11006_, _11005_);
  and (_11008_, _11007_, _10557_);
  or (_11009_, _11008_, _11004_);
  or (_11010_, _11009_, _10551_);
  nand (_11011_, _10375_, _10897_);
  or (_11012_, _10375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  and (_11013_, _11012_, _11011_);
  and (_11014_, _11013_, _10540_);
  and (_11015_, _10375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  nor (_11016_, _10375_, _10960_);
  or (_11017_, _11016_, _11015_);
  and (_11018_, _11017_, _10557_);
  or (_11019_, _11018_, _11014_);
  or (_11020_, _11019_, _10275_);
  and (_11021_, _11020_, _10431_);
  and (_11022_, _11021_, _11010_);
  or (_11023_, _11022_, _11000_);
  or (_11024_, _11023_, _10550_);
  or (_11025_, _10605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  and (_11026_, _11025_, _13707_);
  and (_13685_, _11026_, _11024_);
  or (_11027_, _10375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  nand (_11028_, _10375_, _10629_);
  and (_11029_, _11028_, _10540_);
  and (_11030_, _11029_, _11027_);
  nor (_11031_, _10375_, _10701_);
  and (_11032_, _10375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  or (_11033_, _11032_, _11031_);
  and (_11034_, _11033_, _10557_);
  or (_11035_, _11034_, _11030_);
  or (_11036_, _11035_, _10551_);
  or (_11037_, _10375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  nand (_11038_, _10375_, _10725_);
  and (_11039_, _11038_, _10540_);
  and (_11040_, _11039_, _11037_);
  nor (_11041_, _10375_, _10791_);
  and (_11042_, _10375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  or (_11043_, _11042_, _11041_);
  and (_11044_, _11043_, _10557_);
  or (_11045_, _11044_, _11040_);
  or (_11046_, _11045_, _10275_);
  and (_11047_, _11046_, _10565_);
  and (_11048_, _11047_, _11036_);
  nand (_11049_, _10375_, _10815_);
  or (_11050_, _10375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  and (_11051_, _11050_, _11049_);
  and (_11052_, _11051_, _10540_);
  and (_11053_, _10375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  nor (_11054_, _10375_, _10877_);
  or (_11055_, _11054_, _11053_);
  and (_11056_, _11055_, _10557_);
  or (_11057_, _11056_, _11052_);
  or (_11058_, _11057_, _10551_);
  nand (_11059_, _10375_, _10900_);
  or (_11060_, _10375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  and (_11061_, _11060_, _11059_);
  and (_11062_, _11061_, _10540_);
  and (_11063_, _10375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  nor (_11064_, _10375_, _10963_);
  or (_11065_, _11064_, _11063_);
  and (_11066_, _11065_, _10557_);
  or (_11067_, _11066_, _11062_);
  or (_11068_, _11067_, _10275_);
  and (_11069_, _11068_, _10431_);
  and (_11070_, _11069_, _11058_);
  or (_11071_, _11070_, _11048_);
  or (_11072_, _11071_, _10550_);
  or (_11073_, _10605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  and (_11074_, _11073_, _13707_);
  and (_13687_, _11074_, _11072_);
  and (_11075_, _10375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  and (_11076_, _10553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  or (_11077_, _11076_, _11075_);
  and (_11078_, _11077_, _10540_);
  nor (_11079_, _10375_, _10704_);
  and (_11080_, _10375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  or (_11081_, _11080_, _11079_);
  and (_11082_, _11081_, _10557_);
  or (_11083_, _11082_, _11078_);
  or (_11084_, _11083_, _10551_);
  and (_11085_, _10375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  and (_11086_, _10553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  or (_11087_, _11086_, _11085_);
  and (_11088_, _11087_, _10540_);
  nor (_11089_, _10375_, _10794_);
  and (_11090_, _10375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  or (_11091_, _11090_, _11089_);
  and (_11092_, _11091_, _10557_);
  or (_11093_, _11092_, _11088_);
  or (_11094_, _11093_, _10275_);
  and (_11095_, _11094_, _10565_);
  and (_11096_, _11095_, _11084_);
  or (_11097_, _10553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  or (_11098_, _10375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  and (_11099_, _11098_, _11097_);
  and (_11100_, _11099_, _10540_);
  or (_11101_, _10375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  nand (_11102_, _10375_, _10857_);
  and (_11103_, _11102_, _11101_);
  and (_11104_, _11103_, _10557_);
  or (_11105_, _11104_, _11100_);
  or (_11106_, _11105_, _10551_);
  or (_11107_, _10553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  or (_11108_, _10375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  and (_11109_, _11108_, _11107_);
  and (_11110_, _11109_, _10540_);
  or (_11111_, _10375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  nand (_11112_, _10375_, _10944_);
  and (_11113_, _11112_, _11111_);
  and (_11114_, _11113_, _10557_);
  or (_11115_, _11114_, _11110_);
  or (_11116_, _11115_, _10275_);
  and (_11117_, _11116_, _10431_);
  and (_11118_, _11117_, _11106_);
  or (_11119_, _11118_, _11096_);
  or (_11120_, _11119_, _10550_);
  or (_11121_, _10605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  and (_11122_, _11121_, _13707_);
  and (_13688_, _11122_, _11120_);
  or (_11123_, _10375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  nand (_11124_, _10375_, _10637_);
  and (_11125_, _11124_, _10540_);
  and (_11126_, _11125_, _11123_);
  nor (_11127_, _10375_, _10707_);
  and (_11128_, _10375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or (_11129_, _11128_, _11127_);
  and (_11130_, _11129_, _10557_);
  or (_11131_, _11130_, _11126_);
  or (_11132_, _11131_, _10551_);
  and (_11133_, _10375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  nor (_11134_, _10375_, _10750_);
  or (_11135_, _11134_, _11133_);
  and (_11136_, _11135_, _10540_);
  nor (_11137_, _10375_, _10797_);
  and (_11138_, _10375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or (_11139_, _11138_, _11137_);
  and (_11140_, _11139_, _10557_);
  or (_11141_, _11140_, _11136_);
  or (_11142_, _11141_, _10275_);
  and (_11143_, _11142_, _10565_);
  and (_11144_, _11143_, _11132_);
  or (_11145_, _10553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  or (_11146_, _10375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  and (_11147_, _11146_, _11145_);
  and (_11148_, _11147_, _10540_);
  or (_11149_, _10375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  nand (_11150_, _10375_, _10860_);
  and (_11151_, _11150_, _11149_);
  and (_11152_, _11151_, _10557_);
  or (_11153_, _11152_, _11148_);
  or (_11154_, _11153_, _10551_);
  or (_11155_, _10553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  or (_11156_, _10375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  and (_11157_, _11156_, _11155_);
  and (_11158_, _11157_, _10540_);
  and (_11159_, _10375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  nor (_11160_, _10375_, _10969_);
  or (_11161_, _11160_, _11159_);
  and (_11162_, _11161_, _10557_);
  or (_11163_, _11162_, _11158_);
  or (_11164_, _11163_, _10275_);
  and (_11165_, _11164_, _10431_);
  and (_11166_, _11165_, _11154_);
  or (_11167_, _11166_, _11144_);
  or (_11168_, _11167_, _10550_);
  or (_11169_, _10605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  and (_11170_, _11169_, _13707_);
  and (_13690_, _11170_, _11168_);
  and (_11171_, _10375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  nor (_11172_, _10375_, _10663_);
  or (_11173_, _11172_, _11171_);
  and (_11174_, _11173_, _10540_);
  or (_11175_, _10375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  nand (_11176_, _10375_, _10686_);
  and (_11177_, _11176_, _11175_);
  and (_11178_, _11177_, _10557_);
  or (_11179_, _11178_, _11174_);
  or (_11180_, _11179_, _10551_);
  and (_11181_, _10375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  nor (_11182_, _10375_, _10753_);
  or (_11183_, _11182_, _11181_);
  and (_11184_, _11183_, _10540_);
  or (_11185_, _10375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  nand (_11186_, _10375_, _10775_);
  and (_11187_, _11186_, _11185_);
  and (_11188_, _11187_, _10557_);
  or (_11190_, _11188_, _11184_);
  or (_11192_, _11190_, _10275_);
  and (_11194_, _11192_, _10565_);
  and (_11196_, _11194_, _11180_);
  and (_11198_, _10375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  nor (_11200_, _10375_, _10841_);
  or (_11202_, _11200_, _11198_);
  and (_11204_, _11202_, _10540_);
  or (_11206_, _10375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  nand (_11208_, _10375_, _10863_);
  and (_11210_, _11208_, _11206_);
  and (_11212_, _11210_, _10557_);
  or (_11214_, _11212_, _11204_);
  or (_11216_, _11214_, _10551_);
  and (_11218_, _10375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  nor (_11220_, _10375_, _10927_);
  or (_11222_, _11220_, _11218_);
  and (_11224_, _11222_, _10540_);
  or (_11226_, _10375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  nand (_11228_, _10375_, _10949_);
  and (_11230_, _11228_, _11226_);
  and (_11232_, _11230_, _10557_);
  or (_11234_, _11232_, _11224_);
  or (_11236_, _11234_, _10275_);
  and (_11238_, _11236_, _10431_);
  and (_11240_, _11238_, _11216_);
  or (_11242_, _11240_, _11196_);
  or (_11244_, _11242_, _10550_);
  or (_11245_, _10605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  and (_11246_, _11245_, _13707_);
  and (_13692_, _11246_, _11244_);
  and (_11247_, _10375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nor (_11248_, _10375_, _10666_);
  or (_11249_, _11248_, _11247_);
  and (_11250_, _11249_, _10540_);
  or (_11251_, _10375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  nand (_11252_, _10375_, _10689_);
  and (_11253_, _11252_, _11251_);
  and (_11254_, _11253_, _10557_);
  or (_11255_, _11254_, _11250_);
  or (_11256_, _11255_, _10551_);
  and (_11257_, _10375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  nor (_11258_, _10375_, _10756_);
  or (_11259_, _11258_, _11257_);
  and (_11260_, _11259_, _10540_);
  or (_11261_, _10375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  nand (_11262_, _10375_, _10778_);
  and (_11263_, _11262_, _11261_);
  and (_11264_, _11263_, _10557_);
  or (_11265_, _11264_, _11260_);
  or (_11266_, _11265_, _10275_);
  and (_11267_, _11266_, _10565_);
  and (_11268_, _11267_, _11256_);
  and (_11269_, _10375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  nor (_11270_, _10375_, _10844_);
  or (_11271_, _11270_, _11269_);
  and (_11272_, _11271_, _10540_);
  or (_11273_, _10375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  nand (_11274_, _10375_, _10866_);
  and (_11275_, _11274_, _11273_);
  and (_11276_, _11275_, _10557_);
  or (_11277_, _11276_, _11272_);
  or (_11278_, _11277_, _10551_);
  and (_11279_, _10375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  nor (_11280_, _10375_, _10930_);
  or (_11281_, _11280_, _11279_);
  and (_11282_, _11281_, _10540_);
  or (_11283_, _10375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  nand (_11284_, _10375_, _10952_);
  and (_11285_, _11284_, _11283_);
  and (_11286_, _11285_, _10557_);
  or (_11287_, _11286_, _11282_);
  or (_11288_, _11287_, _10275_);
  and (_11289_, _11288_, _10431_);
  and (_11290_, _11289_, _11278_);
  or (_11291_, _11290_, _11268_);
  or (_11292_, _11291_, _10550_);
  or (_11293_, _10605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  and (_11294_, _11293_, _13707_);
  and (_13694_, _11294_, _11292_);
  or (_11295_, _10375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  nand (_11296_, _10375_, _10647_);
  and (_11297_, _11296_, _10540_);
  and (_11298_, _11297_, _11295_);
  nor (_11299_, _10375_, _10715_);
  and (_11300_, _10375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  or (_11301_, _11300_, _11299_);
  and (_11302_, _11301_, _10557_);
  or (_11303_, _11302_, _11298_);
  or (_11304_, _11303_, _10551_);
  and (_11305_, _10375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  nor (_11306_, _10375_, _10759_);
  or (_11307_, _11306_, _11305_);
  and (_11308_, _11307_, _10540_);
  nor (_11309_, _10375_, _10805_);
  and (_11310_, _10375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  or (_11311_, _11310_, _11309_);
  and (_11312_, _11311_, _10557_);
  or (_11313_, _11312_, _11308_);
  or (_11314_, _11313_, _10275_);
  and (_11315_, _11314_, _10565_);
  and (_11316_, _11315_, _11304_);
  or (_11317_, _10553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  or (_11318_, _10375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  and (_11319_, _11318_, _11317_);
  and (_11320_, _11319_, _10540_);
  or (_11321_, _10375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  or (_11322_, _10553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  and (_11323_, _11322_, _11321_);
  and (_11324_, _11323_, _10557_);
  or (_11325_, _11324_, _11320_);
  or (_11326_, _11325_, _10551_);
  nand (_11327_, _10375_, _10912_);
  or (_11328_, _10375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  and (_11329_, _11328_, _11327_);
  and (_11330_, _11329_, _10540_);
  or (_11332_, _10375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  nand (_11333_, _10375_, _10955_);
  and (_11334_, _11333_, _11332_);
  and (_11335_, _11334_, _10557_);
  or (_11336_, _11335_, _11330_);
  or (_11337_, _11336_, _10275_);
  and (_11338_, _11337_, _10431_);
  and (_11339_, _11338_, _11326_);
  or (_11340_, _11339_, _11316_);
  or (_11341_, _11340_, _10550_);
  or (_11342_, _10605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  and (_11344_, _11342_, _13707_);
  and (_13696_, _11344_, _11341_);
  or (_11345_, \oc8051_gm_cxrom_1.cell0.valid , word_in[7]);
  not (_11346_, \oc8051_gm_cxrom_1.cell0.valid );
  or (_11347_, _11346_, \oc8051_gm_cxrom_1.cell0.data [7]);
  and (_11348_, _11347_, _11345_);
  or (_11349_, _11348_, rst);
  or (_11350_, \oc8051_gm_cxrom_1.cell0.data [7], _13707_);
  and (_13704_, _11350_, _11349_);
  or (_11351_, word_in[0], \oc8051_gm_cxrom_1.cell0.valid );
  or (_11352_, \oc8051_gm_cxrom_1.cell0.data [0], _11346_);
  and (_11353_, _11352_, _11351_);
  or (_11354_, _11353_, rst);
  or (_11355_, \oc8051_gm_cxrom_1.cell0.data [0], _13707_);
  and (_13711_, _11355_, _11354_);
  or (_11356_, word_in[1], \oc8051_gm_cxrom_1.cell0.valid );
  or (_11357_, \oc8051_gm_cxrom_1.cell0.data [1], _11346_);
  and (_11358_, _11357_, _11356_);
  or (_11359_, _11358_, rst);
  or (_11360_, \oc8051_gm_cxrom_1.cell0.data [1], _13707_);
  and (_13715_, _11360_, _11359_);
  or (_11361_, word_in[2], \oc8051_gm_cxrom_1.cell0.valid );
  or (_11362_, \oc8051_gm_cxrom_1.cell0.data [2], _11346_);
  and (_11363_, _11362_, _11361_);
  or (_11364_, _11363_, rst);
  or (_11365_, \oc8051_gm_cxrom_1.cell0.data [2], _13707_);
  and (_13718_, _11365_, _11364_);
  or (_11366_, word_in[3], \oc8051_gm_cxrom_1.cell0.valid );
  or (_11367_, \oc8051_gm_cxrom_1.cell0.data [3], _11346_);
  and (_11368_, _11367_, _11366_);
  or (_11369_, _11368_, rst);
  or (_11370_, \oc8051_gm_cxrom_1.cell0.data [3], _13707_);
  and (_13722_, _11370_, _11369_);
  or (_11371_, word_in[4], \oc8051_gm_cxrom_1.cell0.valid );
  or (_11372_, \oc8051_gm_cxrom_1.cell0.data [4], _11346_);
  and (_11373_, _11372_, _11371_);
  or (_11374_, _11373_, rst);
  or (_11375_, \oc8051_gm_cxrom_1.cell0.data [4], _13707_);
  and (_13726_, _11375_, _11374_);
  or (_11376_, word_in[5], \oc8051_gm_cxrom_1.cell0.valid );
  or (_11377_, \oc8051_gm_cxrom_1.cell0.data [5], _11346_);
  and (_11378_, _11377_, _11376_);
  or (_11379_, _11378_, rst);
  or (_11380_, \oc8051_gm_cxrom_1.cell0.data [5], _13707_);
  and (_13730_, _11380_, _11379_);
  or (_11381_, word_in[6], \oc8051_gm_cxrom_1.cell0.valid );
  or (_11382_, \oc8051_gm_cxrom_1.cell0.data [6], _11346_);
  and (_11383_, _11382_, _11381_);
  or (_11384_, _11383_, rst);
  or (_11385_, \oc8051_gm_cxrom_1.cell0.data [6], _13707_);
  and (_13734_, _11385_, _11384_);
  or (_11386_, \oc8051_gm_cxrom_1.cell1.valid , word_in[15]);
  not (_11387_, \oc8051_gm_cxrom_1.cell1.valid );
  or (_11388_, _11387_, \oc8051_gm_cxrom_1.cell1.data [7]);
  and (_11389_, _11388_, _11386_);
  or (_11390_, _11389_, rst);
  or (_11391_, \oc8051_gm_cxrom_1.cell1.data [7], _13707_);
  and (_13756_, _11391_, _11390_);
  or (_11392_, word_in[8], \oc8051_gm_cxrom_1.cell1.valid );
  or (_11393_, \oc8051_gm_cxrom_1.cell1.data [0], _11387_);
  and (_11394_, _11393_, _11392_);
  or (_11395_, _11394_, rst);
  or (_11396_, \oc8051_gm_cxrom_1.cell1.data [0], _13707_);
  and (_13763_, _11396_, _11395_);
  or (_11397_, word_in[9], \oc8051_gm_cxrom_1.cell1.valid );
  or (_11398_, \oc8051_gm_cxrom_1.cell1.data [1], _11387_);
  and (_11399_, _11398_, _11397_);
  or (_11400_, _11399_, rst);
  or (_11401_, \oc8051_gm_cxrom_1.cell1.data [1], _13707_);
  and (_13767_, _11401_, _11400_);
  or (_11402_, word_in[10], \oc8051_gm_cxrom_1.cell1.valid );
  or (_11403_, \oc8051_gm_cxrom_1.cell1.data [2], _11387_);
  and (_11404_, _11403_, _11402_);
  or (_11405_, _11404_, rst);
  or (_11406_, \oc8051_gm_cxrom_1.cell1.data [2], _13707_);
  and (_13771_, _11406_, _11405_);
  or (_11407_, word_in[11], \oc8051_gm_cxrom_1.cell1.valid );
  or (_11408_, \oc8051_gm_cxrom_1.cell1.data [3], _11387_);
  and (_11409_, _11408_, _11407_);
  or (_11410_, _11409_, rst);
  or (_11411_, \oc8051_gm_cxrom_1.cell1.data [3], _13707_);
  and (_13775_, _11411_, _11410_);
  or (_11412_, word_in[12], \oc8051_gm_cxrom_1.cell1.valid );
  or (_11413_, \oc8051_gm_cxrom_1.cell1.data [4], _11387_);
  and (_11414_, _11413_, _11412_);
  or (_11415_, _11414_, rst);
  or (_11416_, \oc8051_gm_cxrom_1.cell1.data [4], _13707_);
  and (_13779_, _11416_, _11415_);
  or (_11417_, word_in[13], \oc8051_gm_cxrom_1.cell1.valid );
  or (_11418_, \oc8051_gm_cxrom_1.cell1.data [5], _11387_);
  and (_11419_, _11418_, _11417_);
  or (_11420_, _11419_, rst);
  or (_11421_, \oc8051_gm_cxrom_1.cell1.data [5], _13707_);
  and (_13782_, _11421_, _11420_);
  or (_11422_, word_in[14], \oc8051_gm_cxrom_1.cell1.valid );
  or (_11423_, \oc8051_gm_cxrom_1.cell1.data [6], _11387_);
  and (_11424_, _11423_, _11422_);
  or (_11425_, _11424_, rst);
  or (_11426_, \oc8051_gm_cxrom_1.cell1.data [6], _13707_);
  and (_13786_, _11426_, _11425_);
  or (_11427_, \oc8051_gm_cxrom_1.cell2.valid , word_in[23]);
  not (_11428_, \oc8051_gm_cxrom_1.cell2.valid );
  or (_11429_, _11428_, \oc8051_gm_cxrom_1.cell2.data [7]);
  and (_11430_, _11429_, _11427_);
  or (_11431_, _11430_, rst);
  or (_11432_, \oc8051_gm_cxrom_1.cell2.data [7], _13707_);
  and (_13808_, _11432_, _11431_);
  or (_11433_, word_in[16], \oc8051_gm_cxrom_1.cell2.valid );
  or (_11434_, \oc8051_gm_cxrom_1.cell2.data [0], _11428_);
  and (_11435_, _11434_, _11433_);
  or (_11436_, _11435_, rst);
  or (_11437_, \oc8051_gm_cxrom_1.cell2.data [0], _13707_);
  and (_13814_, _11437_, _11436_);
  or (_11438_, word_in[17], \oc8051_gm_cxrom_1.cell2.valid );
  or (_11439_, \oc8051_gm_cxrom_1.cell2.data [1], _11428_);
  and (_11440_, _11439_, _11438_);
  or (_11441_, _11440_, rst);
  or (_11442_, \oc8051_gm_cxrom_1.cell2.data [1], _13707_);
  and (_13818_, _11442_, _11441_);
  or (_11443_, word_in[18], \oc8051_gm_cxrom_1.cell2.valid );
  or (_11444_, \oc8051_gm_cxrom_1.cell2.data [2], _11428_);
  and (_11445_, _11444_, _11443_);
  or (_11446_, _11445_, rst);
  or (_11447_, \oc8051_gm_cxrom_1.cell2.data [2], _13707_);
  and (_13822_, _11447_, _11446_);
  or (_11448_, word_in[19], \oc8051_gm_cxrom_1.cell2.valid );
  or (_11449_, \oc8051_gm_cxrom_1.cell2.data [3], _11428_);
  and (_11450_, _11449_, _11448_);
  or (_11451_, _11450_, rst);
  or (_11452_, \oc8051_gm_cxrom_1.cell2.data [3], _13707_);
  and (_00012_, _11452_, _11451_);
  or (_11453_, word_in[20], \oc8051_gm_cxrom_1.cell2.valid );
  or (_11454_, \oc8051_gm_cxrom_1.cell2.data [4], _11428_);
  and (_11455_, _11454_, _11453_);
  or (_11456_, _11455_, rst);
  or (_11457_, \oc8051_gm_cxrom_1.cell2.data [4], _13707_);
  and (_00016_, _11457_, _11456_);
  or (_11458_, word_in[21], \oc8051_gm_cxrom_1.cell2.valid );
  or (_11459_, \oc8051_gm_cxrom_1.cell2.data [5], _11428_);
  and (_11460_, _11459_, _11458_);
  or (_11461_, _11460_, rst);
  or (_11462_, \oc8051_gm_cxrom_1.cell2.data [5], _13707_);
  and (_00020_, _11462_, _11461_);
  or (_11463_, word_in[22], \oc8051_gm_cxrom_1.cell2.valid );
  or (_11464_, \oc8051_gm_cxrom_1.cell2.data [6], _11428_);
  and (_11465_, _11464_, _11463_);
  or (_11466_, _11465_, rst);
  or (_11467_, \oc8051_gm_cxrom_1.cell2.data [6], _13707_);
  and (_00024_, _11467_, _11466_);
  or (_11468_, \oc8051_gm_cxrom_1.cell3.valid , word_in[31]);
  not (_11469_, \oc8051_gm_cxrom_1.cell3.valid );
  or (_11470_, _11469_, \oc8051_gm_cxrom_1.cell3.data [7]);
  and (_11471_, _11470_, _11468_);
  or (_11472_, _11471_, rst);
  or (_11473_, \oc8051_gm_cxrom_1.cell3.data [7], _13707_);
  and (_00045_, _11473_, _11472_);
  or (_11474_, word_in[24], \oc8051_gm_cxrom_1.cell3.valid );
  or (_11475_, \oc8051_gm_cxrom_1.cell3.data [0], _11469_);
  and (_11476_, _11475_, _11474_);
  or (_11477_, _11476_, rst);
  or (_11478_, \oc8051_gm_cxrom_1.cell3.data [0], _13707_);
  and (_00052_, _11478_, _11477_);
  or (_11479_, word_in[25], \oc8051_gm_cxrom_1.cell3.valid );
  or (_11480_, \oc8051_gm_cxrom_1.cell3.data [1], _11469_);
  and (_11481_, _11480_, _11479_);
  or (_11482_, _11481_, rst);
  or (_11483_, \oc8051_gm_cxrom_1.cell3.data [1], _13707_);
  and (_00056_, _11483_, _11482_);
  or (_11484_, word_in[26], \oc8051_gm_cxrom_1.cell3.valid );
  or (_11485_, \oc8051_gm_cxrom_1.cell3.data [2], _11469_);
  and (_11486_, _11485_, _11484_);
  or (_11487_, _11486_, rst);
  or (_11488_, \oc8051_gm_cxrom_1.cell3.data [2], _13707_);
  and (_00059_, _11488_, _11487_);
  or (_11489_, word_in[27], \oc8051_gm_cxrom_1.cell3.valid );
  or (_11490_, \oc8051_gm_cxrom_1.cell3.data [3], _11469_);
  and (_11491_, _11490_, _11489_);
  or (_11492_, _11491_, rst);
  or (_11493_, \oc8051_gm_cxrom_1.cell3.data [3], _13707_);
  and (_00063_, _11493_, _11492_);
  or (_11494_, word_in[28], \oc8051_gm_cxrom_1.cell3.valid );
  or (_11495_, \oc8051_gm_cxrom_1.cell3.data [4], _11469_);
  and (_11496_, _11495_, _11494_);
  or (_11497_, _11496_, rst);
  or (_11498_, \oc8051_gm_cxrom_1.cell3.data [4], _13707_);
  and (_00067_, _11498_, _11497_);
  or (_11499_, word_in[29], \oc8051_gm_cxrom_1.cell3.valid );
  or (_11500_, \oc8051_gm_cxrom_1.cell3.data [5], _11469_);
  and (_11501_, _11500_, _11499_);
  or (_11502_, _11501_, rst);
  or (_11503_, \oc8051_gm_cxrom_1.cell3.data [5], _13707_);
  and (_00071_, _11503_, _11502_);
  or (_11504_, word_in[30], \oc8051_gm_cxrom_1.cell3.valid );
  or (_11505_, \oc8051_gm_cxrom_1.cell3.data [6], _11469_);
  and (_11506_, _11505_, _11504_);
  or (_11507_, _11506_, rst);
  or (_11508_, \oc8051_gm_cxrom_1.cell3.data [6], _13707_);
  and (_00075_, _11508_, _11507_);
  or (_11509_, \oc8051_gm_cxrom_1.cell4.valid , word_in[39]);
  not (_11510_, \oc8051_gm_cxrom_1.cell4.valid );
  or (_11511_, _11510_, \oc8051_gm_cxrom_1.cell4.data [7]);
  and (_11512_, _11511_, _11509_);
  or (_11513_, _11512_, rst);
  or (_11514_, \oc8051_gm_cxrom_1.cell4.data [7], _13707_);
  and (_00096_, _11514_, _11513_);
  or (_11515_, word_in[32], \oc8051_gm_cxrom_1.cell4.valid );
  or (_11516_, \oc8051_gm_cxrom_1.cell4.data [0], _11510_);
  and (_11517_, _11516_, _11515_);
  or (_11518_, _11517_, rst);
  or (_11519_, \oc8051_gm_cxrom_1.cell4.data [0], _13707_);
  and (_00103_, _11519_, _11518_);
  or (_11520_, word_in[33], \oc8051_gm_cxrom_1.cell4.valid );
  or (_11521_, \oc8051_gm_cxrom_1.cell4.data [1], _11510_);
  and (_11522_, _11521_, _11520_);
  or (_11523_, _11522_, rst);
  or (_11524_, \oc8051_gm_cxrom_1.cell4.data [1], _13707_);
  and (_00107_, _11524_, _11523_);
  or (_11525_, word_in[34], \oc8051_gm_cxrom_1.cell4.valid );
  or (_11526_, \oc8051_gm_cxrom_1.cell4.data [2], _11510_);
  and (_11527_, _11526_, _11525_);
  or (_11528_, _11527_, rst);
  or (_11529_, \oc8051_gm_cxrom_1.cell4.data [2], _13707_);
  and (_00111_, _11529_, _11528_);
  or (_11530_, word_in[35], \oc8051_gm_cxrom_1.cell4.valid );
  or (_11531_, \oc8051_gm_cxrom_1.cell4.data [3], _11510_);
  and (_11532_, _11531_, _11530_);
  or (_11533_, _11532_, rst);
  or (_11534_, \oc8051_gm_cxrom_1.cell4.data [3], _13707_);
  and (_00114_, _11534_, _11533_);
  or (_11535_, word_in[36], \oc8051_gm_cxrom_1.cell4.valid );
  or (_11536_, \oc8051_gm_cxrom_1.cell4.data [4], _11510_);
  and (_11537_, _11536_, _11535_);
  or (_11538_, _11537_, rst);
  or (_11539_, \oc8051_gm_cxrom_1.cell4.data [4], _13707_);
  and (_00118_, _11539_, _11538_);
  or (_11540_, word_in[37], \oc8051_gm_cxrom_1.cell4.valid );
  or (_11541_, \oc8051_gm_cxrom_1.cell4.data [5], _11510_);
  and (_11542_, _11541_, _11540_);
  or (_11543_, _11542_, rst);
  or (_11544_, \oc8051_gm_cxrom_1.cell4.data [5], _13707_);
  and (_00122_, _11544_, _11543_);
  or (_11545_, word_in[38], \oc8051_gm_cxrom_1.cell4.valid );
  or (_11546_, \oc8051_gm_cxrom_1.cell4.data [6], _11510_);
  and (_11547_, _11546_, _11545_);
  or (_11548_, _11547_, rst);
  or (_11549_, \oc8051_gm_cxrom_1.cell4.data [6], _13707_);
  and (_00126_, _11549_, _11548_);
  or (_11550_, \oc8051_gm_cxrom_1.cell5.valid , word_in[47]);
  not (_11551_, \oc8051_gm_cxrom_1.cell5.valid );
  or (_11552_, _11551_, \oc8051_gm_cxrom_1.cell5.data [7]);
  and (_11553_, _11552_, _11550_);
  or (_11554_, _11553_, rst);
  or (_11555_, \oc8051_gm_cxrom_1.cell5.data [7], _13707_);
  and (_00146_, _11555_, _11554_);
  or (_11556_, word_in[40], \oc8051_gm_cxrom_1.cell5.valid );
  or (_11557_, \oc8051_gm_cxrom_1.cell5.data [0], _11551_);
  and (_11558_, _11557_, _11556_);
  or (_11559_, _11558_, rst);
  or (_11560_, \oc8051_gm_cxrom_1.cell5.data [0], _13707_);
  and (_00153_, _11560_, _11559_);
  or (_11561_, word_in[41], \oc8051_gm_cxrom_1.cell5.valid );
  or (_11562_, \oc8051_gm_cxrom_1.cell5.data [1], _11551_);
  and (_11563_, _11562_, _11561_);
  or (_11564_, _11563_, rst);
  or (_11565_, \oc8051_gm_cxrom_1.cell5.data [1], _13707_);
  and (_00156_, _11565_, _11564_);
  or (_11566_, word_in[42], \oc8051_gm_cxrom_1.cell5.valid );
  or (_11567_, \oc8051_gm_cxrom_1.cell5.data [2], _11551_);
  and (_11568_, _11567_, _11566_);
  or (_11569_, _11568_, rst);
  or (_11570_, \oc8051_gm_cxrom_1.cell5.data [2], _13707_);
  and (_00160_, _11570_, _11569_);
  or (_11571_, word_in[43], \oc8051_gm_cxrom_1.cell5.valid );
  or (_11572_, \oc8051_gm_cxrom_1.cell5.data [3], _11551_);
  and (_11573_, _11572_, _11571_);
  or (_11574_, _11573_, rst);
  or (_11575_, \oc8051_gm_cxrom_1.cell5.data [3], _13707_);
  and (_00163_, _11575_, _11574_);
  or (_11576_, word_in[44], \oc8051_gm_cxrom_1.cell5.valid );
  or (_11577_, \oc8051_gm_cxrom_1.cell5.data [4], _11551_);
  and (_11578_, _11577_, _11576_);
  or (_11579_, _11578_, rst);
  or (_11580_, \oc8051_gm_cxrom_1.cell5.data [4], _13707_);
  and (_00167_, _11580_, _11579_);
  or (_11581_, word_in[45], \oc8051_gm_cxrom_1.cell5.valid );
  or (_11582_, \oc8051_gm_cxrom_1.cell5.data [5], _11551_);
  and (_11583_, _11582_, _11581_);
  or (_11584_, _11583_, rst);
  or (_11585_, \oc8051_gm_cxrom_1.cell5.data [5], _13707_);
  and (_00171_, _11585_, _11584_);
  or (_11587_, word_in[46], \oc8051_gm_cxrom_1.cell5.valid );
  or (_11588_, \oc8051_gm_cxrom_1.cell5.data [6], _11551_);
  and (_11589_, _11588_, _11587_);
  or (_11590_, _11589_, rst);
  or (_11592_, \oc8051_gm_cxrom_1.cell5.data [6], _13707_);
  and (_00174_, _11592_, _11590_);
  or (_11593_, \oc8051_gm_cxrom_1.cell6.valid , word_in[55]);
  not (_11594_, \oc8051_gm_cxrom_1.cell6.valid );
  or (_11595_, _11594_, \oc8051_gm_cxrom_1.cell6.data [7]);
  and (_11597_, _11595_, _11593_);
  or (_11598_, _11597_, rst);
  or (_11599_, \oc8051_gm_cxrom_1.cell6.data [7], _13707_);
  and (_00194_, _11599_, _11598_);
  or (_11600_, word_in[48], \oc8051_gm_cxrom_1.cell6.valid );
  or (_11602_, \oc8051_gm_cxrom_1.cell6.data [0], _11594_);
  and (_11603_, _11602_, _11600_);
  or (_11604_, _11603_, rst);
  or (_11605_, \oc8051_gm_cxrom_1.cell6.data [0], _13707_);
  and (_00200_, _11605_, _11604_);
  or (_11607_, word_in[49], \oc8051_gm_cxrom_1.cell6.valid );
  or (_11608_, \oc8051_gm_cxrom_1.cell6.data [1], _11594_);
  and (_11609_, _11608_, _11607_);
  or (_11610_, _11609_, rst);
  or (_11611_, \oc8051_gm_cxrom_1.cell6.data [1], _13707_);
  and (_00204_, _11611_, _11610_);
  or (_11613_, word_in[50], \oc8051_gm_cxrom_1.cell6.valid );
  or (_11614_, \oc8051_gm_cxrom_1.cell6.data [2], _11594_);
  and (_11615_, _11614_, _11613_);
  or (_11616_, _11615_, rst);
  or (_11618_, \oc8051_gm_cxrom_1.cell6.data [2], _13707_);
  and (_00207_, _11618_, _11616_);
  or (_11620_, word_in[51], \oc8051_gm_cxrom_1.cell6.valid );
  or (_11621_, \oc8051_gm_cxrom_1.cell6.data [3], _11594_);
  and (_11622_, _11621_, _11620_);
  or (_11623_, _11622_, rst);
  or (_11624_, \oc8051_gm_cxrom_1.cell6.data [3], _13707_);
  and (_00211_, _11624_, _11623_);
  or (_11625_, word_in[52], \oc8051_gm_cxrom_1.cell6.valid );
  or (_11627_, \oc8051_gm_cxrom_1.cell6.data [4], _11594_);
  and (_11628_, _11627_, _11625_);
  or (_11629_, _11628_, rst);
  or (_11631_, \oc8051_gm_cxrom_1.cell6.data [4], _13707_);
  and (_00215_, _11631_, _11629_);
  or (_11632_, word_in[53], \oc8051_gm_cxrom_1.cell6.valid );
  or (_11634_, \oc8051_gm_cxrom_1.cell6.data [5], _11594_);
  and (_11635_, _11634_, _11632_);
  or (_11636_, _11635_, rst);
  or (_11638_, \oc8051_gm_cxrom_1.cell6.data [5], _13707_);
  and (_00218_, _11638_, _11636_);
  or (_11639_, word_in[54], \oc8051_gm_cxrom_1.cell6.valid );
  or (_11641_, \oc8051_gm_cxrom_1.cell6.data [6], _11594_);
  and (_11642_, _11641_, _11639_);
  or (_11643_, _11642_, rst);
  or (_11645_, \oc8051_gm_cxrom_1.cell6.data [6], _13707_);
  and (_00222_, _11645_, _11643_);
  or (_11646_, \oc8051_gm_cxrom_1.cell7.valid , word_in[63]);
  not (_11648_, \oc8051_gm_cxrom_1.cell7.valid );
  or (_11649_, _11648_, \oc8051_gm_cxrom_1.cell7.data [7]);
  and (_11651_, _11649_, _11646_);
  or (_11652_, _11651_, rst);
  or (_11653_, \oc8051_gm_cxrom_1.cell7.data [7], _13707_);
  and (_00241_, _11653_, _11652_);
  or (_11654_, word_in[56], \oc8051_gm_cxrom_1.cell7.valid );
  or (_11655_, \oc8051_gm_cxrom_1.cell7.data [0], _11648_);
  and (_11656_, _11655_, _11654_);
  or (_11658_, _11656_, rst);
  or (_11659_, \oc8051_gm_cxrom_1.cell7.data [0], _13707_);
  and (_00248_, _11659_, _11658_);
  or (_11661_, word_in[57], \oc8051_gm_cxrom_1.cell7.valid );
  or (_11662_, \oc8051_gm_cxrom_1.cell7.data [1], _11648_);
  and (_11663_, _11662_, _11661_);
  or (_11665_, _11663_, rst);
  or (_11666_, \oc8051_gm_cxrom_1.cell7.data [1], _13707_);
  and (_00251_, _11666_, _11665_);
  or (_11668_, word_in[58], \oc8051_gm_cxrom_1.cell7.valid );
  or (_11669_, \oc8051_gm_cxrom_1.cell7.data [2], _11648_);
  and (_11670_, _11669_, _11668_);
  or (_11672_, _11670_, rst);
  or (_11673_, \oc8051_gm_cxrom_1.cell7.data [2], _13707_);
  and (_00255_, _11673_, _11672_);
  or (_11675_, word_in[59], \oc8051_gm_cxrom_1.cell7.valid );
  or (_11676_, \oc8051_gm_cxrom_1.cell7.data [3], _11648_);
  and (_11677_, _11676_, _11675_);
  or (_11679_, _11677_, rst);
  or (_11680_, \oc8051_gm_cxrom_1.cell7.data [3], _13707_);
  and (_00259_, _11680_, _11679_);
  or (_11682_, word_in[60], \oc8051_gm_cxrom_1.cell7.valid );
  or (_11683_, \oc8051_gm_cxrom_1.cell7.data [4], _11648_);
  and (_11684_, _11683_, _11682_);
  or (_11685_, _11684_, rst);
  or (_11687_, \oc8051_gm_cxrom_1.cell7.data [4], _13707_);
  and (_00262_, _11687_, _11685_);
  or (_11688_, word_in[61], \oc8051_gm_cxrom_1.cell7.valid );
  or (_11690_, \oc8051_gm_cxrom_1.cell7.data [5], _11648_);
  and (_11691_, _11690_, _11688_);
  or (_11692_, _11691_, rst);
  or (_11694_, \oc8051_gm_cxrom_1.cell7.data [5], _13707_);
  and (_00266_, _11694_, _11692_);
  or (_11695_, word_in[62], \oc8051_gm_cxrom_1.cell7.valid );
  or (_11697_, \oc8051_gm_cxrom_1.cell7.data [6], _11648_);
  and (_11698_, _11697_, _11695_);
  or (_11699_, _11698_, rst);
  or (_11701_, \oc8051_gm_cxrom_1.cell7.data [6], _13707_);
  and (_00269_, _11701_, _11699_);
  or (_11702_, \oc8051_gm_cxrom_1.cell8.valid , word_in[71]);
  not (_11704_, \oc8051_gm_cxrom_1.cell8.valid );
  or (_11705_, _11704_, \oc8051_gm_cxrom_1.cell8.data [7]);
  and (_11706_, _11705_, _11702_);
  or (_11708_, _11706_, rst);
  or (_11709_, \oc8051_gm_cxrom_1.cell8.data [7], _13707_);
  and (_00282_, _11709_, _11708_);
  or (_11711_, word_in[64], \oc8051_gm_cxrom_1.cell8.valid );
  or (_11712_, \oc8051_gm_cxrom_1.cell8.data [0], _11704_);
  and (_11713_, _11712_, _11711_);
  or (_11714_, _11713_, rst);
  or (_11715_, \oc8051_gm_cxrom_1.cell8.data [0], _13707_);
  and (_00287_, _11715_, _11714_);
  or (_11717_, word_in[65], \oc8051_gm_cxrom_1.cell8.valid );
  or (_11718_, \oc8051_gm_cxrom_1.cell8.data [1], _11704_);
  and (_11719_, _11718_, _11717_);
  or (_11721_, _11719_, rst);
  or (_11722_, \oc8051_gm_cxrom_1.cell8.data [1], _13707_);
  and (_00291_, _11722_, _11721_);
  or (_11724_, word_in[66], \oc8051_gm_cxrom_1.cell8.valid );
  or (_11725_, \oc8051_gm_cxrom_1.cell8.data [2], _11704_);
  and (_11726_, _11725_, _11724_);
  or (_11728_, _11726_, rst);
  or (_11729_, \oc8051_gm_cxrom_1.cell8.data [2], _13707_);
  and (_00294_, _11729_, _11728_);
  or (_11731_, word_in[67], \oc8051_gm_cxrom_1.cell8.valid );
  or (_11732_, \oc8051_gm_cxrom_1.cell8.data [3], _11704_);
  and (_11733_, _11732_, _11731_);
  or (_11735_, _11733_, rst);
  or (_11736_, \oc8051_gm_cxrom_1.cell8.data [3], _13707_);
  and (_00297_, _11736_, _11735_);
  or (_11738_, word_in[68], \oc8051_gm_cxrom_1.cell8.valid );
  or (_11739_, \oc8051_gm_cxrom_1.cell8.data [4], _11704_);
  and (_11741_, _11739_, _11738_);
  or (_11742_, _11741_, rst);
  or (_11743_, \oc8051_gm_cxrom_1.cell8.data [4], _13707_);
  and (_00300_, _11743_, _11742_);
  or (_11745_, word_in[69], \oc8051_gm_cxrom_1.cell8.valid );
  or (_11746_, \oc8051_gm_cxrom_1.cell8.data [5], _11704_);
  and (_11747_, _11746_, _11745_);
  or (_11749_, _11747_, rst);
  or (_11750_, \oc8051_gm_cxrom_1.cell8.data [5], _13707_);
  and (_00304_, _11750_, _11749_);
  or (_11752_, word_in[70], \oc8051_gm_cxrom_1.cell8.valid );
  or (_11753_, \oc8051_gm_cxrom_1.cell8.data [6], _11704_);
  and (_11754_, _11753_, _11752_);
  or (_11756_, _11754_, rst);
  or (_11757_, \oc8051_gm_cxrom_1.cell8.data [6], _13707_);
  and (_00307_, _11757_, _11756_);
  or (_11759_, \oc8051_gm_cxrom_1.cell9.valid , word_in[79]);
  not (_11760_, \oc8051_gm_cxrom_1.cell9.valid );
  or (_11761_, _11760_, \oc8051_gm_cxrom_1.cell9.data [7]);
  and (_11763_, _11761_, _11759_);
  or (_11764_, _11763_, rst);
  or (_11765_, \oc8051_gm_cxrom_1.cell9.data [7], _13707_);
  and (_00322_, _11765_, _11764_);
  or (_11767_, word_in[72], \oc8051_gm_cxrom_1.cell9.valid );
  or (_11769_, \oc8051_gm_cxrom_1.cell9.data [0], _11760_);
  and (_11770_, _11769_, _11767_);
  or (_11771_, _11770_, rst);
  or (_11772_, \oc8051_gm_cxrom_1.cell9.data [0], _13707_);
  and (_00327_, _11772_, _11771_);
  or (_11774_, word_in[73], \oc8051_gm_cxrom_1.cell9.valid );
  or (_11775_, \oc8051_gm_cxrom_1.cell9.data [1], _11760_);
  and (_11777_, _11775_, _11774_);
  or (_11778_, _11777_, rst);
  or (_11779_, \oc8051_gm_cxrom_1.cell9.data [1], _13707_);
  and (_00331_, _11779_, _11778_);
  or (_11781_, word_in[74], \oc8051_gm_cxrom_1.cell9.valid );
  or (_11782_, \oc8051_gm_cxrom_1.cell9.data [2], _11760_);
  and (_11784_, _11782_, _11781_);
  or (_11785_, _11784_, rst);
  or (_11786_, \oc8051_gm_cxrom_1.cell9.data [2], _13707_);
  and (_00334_, _11786_, _11785_);
  or (_11788_, word_in[75], \oc8051_gm_cxrom_1.cell9.valid );
  or (_11789_, \oc8051_gm_cxrom_1.cell9.data [3], _11760_);
  and (_11791_, _11789_, _11788_);
  or (_11792_, _11791_, rst);
  or (_11793_, \oc8051_gm_cxrom_1.cell9.data [3], _13707_);
  and (_00337_, _11793_, _11792_);
  or (_11795_, word_in[76], \oc8051_gm_cxrom_1.cell9.valid );
  or (_11797_, \oc8051_gm_cxrom_1.cell9.data [4], _11760_);
  and (_11798_, _11797_, _11795_);
  or (_11799_, _11798_, rst);
  or (_11800_, \oc8051_gm_cxrom_1.cell9.data [4], _13707_);
  and (_00340_, _11800_, _11799_);
  or (_11802_, word_in[77], \oc8051_gm_cxrom_1.cell9.valid );
  or (_11803_, \oc8051_gm_cxrom_1.cell9.data [5], _11760_);
  and (_11805_, _11803_, _11802_);
  or (_11806_, _11805_, rst);
  or (_11807_, \oc8051_gm_cxrom_1.cell9.data [5], _13707_);
  and (_00344_, _11807_, _11806_);
  or (_11809_, word_in[78], \oc8051_gm_cxrom_1.cell9.valid );
  or (_11810_, \oc8051_gm_cxrom_1.cell9.data [6], _11760_);
  and (_11812_, _11810_, _11809_);
  or (_11813_, _11812_, rst);
  or (_11814_, \oc8051_gm_cxrom_1.cell9.data [6], _13707_);
  and (_00347_, _11814_, _11813_);
  or (_11816_, \oc8051_gm_cxrom_1.cell10.valid , word_in[87]);
  not (_11817_, \oc8051_gm_cxrom_1.cell10.valid );
  or (_11819_, _11817_, \oc8051_gm_cxrom_1.cell10.data [7]);
  and (_11820_, _11819_, _11816_);
  or (_11821_, _11820_, rst);
  or (_11823_, \oc8051_gm_cxrom_1.cell10.data [7], _13707_);
  and (_00364_, _11823_, _11821_);
  or (_11825_, word_in[80], \oc8051_gm_cxrom_1.cell10.valid );
  or (_11826_, \oc8051_gm_cxrom_1.cell10.data [0], _11817_);
  and (_11827_, _11826_, _11825_);
  or (_11828_, _11827_, rst);
  or (_11829_, \oc8051_gm_cxrom_1.cell10.data [0], _13707_);
  and (_00369_, _11829_, _11828_);
  or (_11830_, word_in[81], \oc8051_gm_cxrom_1.cell10.valid );
  or (_11832_, \oc8051_gm_cxrom_1.cell10.data [1], _11817_);
  and (_11833_, _11832_, _11830_);
  or (_11834_, _11833_, rst);
  or (_11836_, \oc8051_gm_cxrom_1.cell10.data [1], _13707_);
  and (_00373_, _11836_, _11834_);
  or (_11837_, word_in[82], \oc8051_gm_cxrom_1.cell10.valid );
  or (_11839_, \oc8051_gm_cxrom_1.cell10.data [2], _11817_);
  and (_11840_, _11839_, _11837_);
  or (_11841_, _11840_, rst);
  or (_11843_, \oc8051_gm_cxrom_1.cell10.data [2], _13707_);
  and (_00376_, _11843_, _11841_);
  or (_11844_, word_in[83], \oc8051_gm_cxrom_1.cell10.valid );
  or (_11846_, \oc8051_gm_cxrom_1.cell10.data [3], _11817_);
  and (_11847_, _11846_, _11844_);
  or (_11848_, _11847_, rst);
  or (_11850_, \oc8051_gm_cxrom_1.cell10.data [3], _13707_);
  and (_00379_, _11850_, _11848_);
  or (_11851_, word_in[84], \oc8051_gm_cxrom_1.cell10.valid );
  or (_11853_, \oc8051_gm_cxrom_1.cell10.data [4], _11817_);
  and (_11854_, _11853_, _11851_);
  or (_11856_, _11854_, rst);
  or (_11857_, \oc8051_gm_cxrom_1.cell10.data [4], _13707_);
  and (_00382_, _11857_, _11856_);
  or (_11858_, word_in[85], \oc8051_gm_cxrom_1.cell10.valid );
  or (_11860_, \oc8051_gm_cxrom_1.cell10.data [5], _11817_);
  and (_11861_, _11860_, _11858_);
  or (_11862_, _11861_, rst);
  or (_11864_, \oc8051_gm_cxrom_1.cell10.data [5], _13707_);
  and (_00386_, _11864_, _11862_);
  or (_11865_, word_in[86], \oc8051_gm_cxrom_1.cell10.valid );
  or (_11867_, \oc8051_gm_cxrom_1.cell10.data [6], _11817_);
  and (_11868_, _11867_, _11865_);
  or (_11869_, _11868_, rst);
  or (_11871_, \oc8051_gm_cxrom_1.cell10.data [6], _13707_);
  and (_00389_, _11871_, _11869_);
  or (_11872_, \oc8051_gm_cxrom_1.cell11.valid , word_in[95]);
  not (_11874_, \oc8051_gm_cxrom_1.cell11.valid );
  or (_11875_, _11874_, \oc8051_gm_cxrom_1.cell11.data [7]);
  and (_11876_, _11875_, _11872_);
  or (_11878_, _11876_, rst);
  or (_11879_, \oc8051_gm_cxrom_1.cell11.data [7], _13707_);
  and (_00406_, _11879_, _11878_);
  or (_11881_, word_in[88], \oc8051_gm_cxrom_1.cell11.valid );
  or (_11882_, \oc8051_gm_cxrom_1.cell11.data [0], _11874_);
  and (_11884_, _11882_, _11881_);
  or (_11885_, _11884_, rst);
  or (_11886_, \oc8051_gm_cxrom_1.cell11.data [0], _13707_);
  and (_00411_, _11886_, _11885_);
  or (_11888_, word_in[89], \oc8051_gm_cxrom_1.cell11.valid );
  or (_11889_, \oc8051_gm_cxrom_1.cell11.data [1], _11874_);
  and (_11890_, _11889_, _11888_);
  or (_11892_, _11890_, rst);
  or (_11893_, \oc8051_gm_cxrom_1.cell11.data [1], _13707_);
  and (_00415_, _11893_, _11892_);
  or (_11895_, word_in[90], \oc8051_gm_cxrom_1.cell11.valid );
  or (_11896_, \oc8051_gm_cxrom_1.cell11.data [2], _11874_);
  and (_11897_, _11896_, _11895_);
  or (_11899_, _11897_, rst);
  or (_11900_, \oc8051_gm_cxrom_1.cell11.data [2], _13707_);
  and (_00418_, _11900_, _11899_);
  or (_11902_, word_in[91], \oc8051_gm_cxrom_1.cell11.valid );
  or (_11903_, \oc8051_gm_cxrom_1.cell11.data [3], _11874_);
  and (_11904_, _11903_, _11902_);
  or (_11906_, _11904_, rst);
  or (_11907_, \oc8051_gm_cxrom_1.cell11.data [3], _13707_);
  and (_00421_, _11907_, _11906_);
  or (_11909_, word_in[92], \oc8051_gm_cxrom_1.cell11.valid );
  or (_11910_, \oc8051_gm_cxrom_1.cell11.data [4], _11874_);
  and (_11912_, _11910_, _11909_);
  or (_11913_, _11912_, rst);
  or (_11914_, \oc8051_gm_cxrom_1.cell11.data [4], _13707_);
  and (_00424_, _11914_, _11913_);
  or (_11916_, word_in[93], \oc8051_gm_cxrom_1.cell11.valid );
  or (_11917_, \oc8051_gm_cxrom_1.cell11.data [5], _11874_);
  and (_11918_, _11917_, _11916_);
  or (_11920_, _11918_, rst);
  or (_11921_, \oc8051_gm_cxrom_1.cell11.data [5], _13707_);
  and (_00428_, _11921_, _11920_);
  or (_11923_, word_in[94], \oc8051_gm_cxrom_1.cell11.valid );
  or (_11924_, \oc8051_gm_cxrom_1.cell11.data [6], _11874_);
  and (_11925_, _11924_, _11923_);
  or (_11927_, _11925_, rst);
  or (_11928_, \oc8051_gm_cxrom_1.cell11.data [6], _13707_);
  and (_00431_, _11928_, _11927_);
  or (_11930_, \oc8051_gm_cxrom_1.cell12.valid , word_in[103]);
  not (_11931_, \oc8051_gm_cxrom_1.cell12.valid );
  or (_11932_, _11931_, \oc8051_gm_cxrom_1.cell12.data [7]);
  and (_11934_, _11932_, _11930_);
  or (_11935_, _11934_, rst);
  or (_11936_, \oc8051_gm_cxrom_1.cell12.data [7], _13707_);
  and (_00450_, _11936_, _11935_);
  or (_11938_, word_in[96], \oc8051_gm_cxrom_1.cell12.valid );
  or (_11940_, \oc8051_gm_cxrom_1.cell12.data [0], _11931_);
  and (_11941_, _11940_, _11938_);
  or (_11942_, _11941_, rst);
  or (_11943_, \oc8051_gm_cxrom_1.cell12.data [0], _13707_);
  and (_00456_, _11943_, _11942_);
  or (_11945_, word_in[97], \oc8051_gm_cxrom_1.cell12.valid );
  or (_11946_, \oc8051_gm_cxrom_1.cell12.data [1], _11931_);
  and (_11947_, _11946_, _11945_);
  or (_11949_, _11947_, rst);
  or (_11950_, \oc8051_gm_cxrom_1.cell12.data [1], _13707_);
  and (_00459_, _11950_, _11949_);
  or (_11952_, word_in[98], \oc8051_gm_cxrom_1.cell12.valid );
  or (_11953_, \oc8051_gm_cxrom_1.cell12.data [2], _11931_);
  and (_11954_, _11953_, _11952_);
  or (_11956_, _11954_, rst);
  or (_11957_, \oc8051_gm_cxrom_1.cell12.data [2], _13707_);
  and (_00463_, _11957_, _11956_);
  or (_11959_, word_in[99], \oc8051_gm_cxrom_1.cell12.valid );
  or (_11960_, \oc8051_gm_cxrom_1.cell12.data [3], _11931_);
  and (_11961_, _11960_, _11959_);
  or (_11963_, _11961_, rst);
  or (_11964_, \oc8051_gm_cxrom_1.cell12.data [3], _13707_);
  and (_00466_, _11964_, _11963_);
  or (_11966_, word_in[100], \oc8051_gm_cxrom_1.cell12.valid );
  or (_11967_, \oc8051_gm_cxrom_1.cell12.data [4], _11931_);
  and (_11969_, _11967_, _11966_);
  or (_11970_, _11969_, rst);
  or (_11971_, \oc8051_gm_cxrom_1.cell12.data [4], _13707_);
  and (_00470_, _11971_, _11970_);
  or (_11973_, word_in[101], \oc8051_gm_cxrom_1.cell12.valid );
  or (_11974_, \oc8051_gm_cxrom_1.cell12.data [5], _11931_);
  and (_11975_, _11974_, _11973_);
  or (_11977_, _11975_, rst);
  or (_11978_, \oc8051_gm_cxrom_1.cell12.data [5], _13707_);
  and (_00473_, _11978_, _11977_);
  or (_11980_, word_in[102], \oc8051_gm_cxrom_1.cell12.valid );
  or (_11981_, \oc8051_gm_cxrom_1.cell12.data [6], _11931_);
  and (_11982_, _11981_, _11980_);
  or (_11984_, _11982_, rst);
  or (_11985_, \oc8051_gm_cxrom_1.cell12.data [6], _13707_);
  and (_00477_, _11985_, _11984_);
  or (_11987_, \oc8051_gm_cxrom_1.cell13.valid , word_in[111]);
  not (_11988_, \oc8051_gm_cxrom_1.cell13.valid );
  or (_11989_, _11988_, \oc8051_gm_cxrom_1.cell13.data [7]);
  and (_11991_, _11989_, _11987_);
  or (_11992_, _11991_, rst);
  or (_11993_, \oc8051_gm_cxrom_1.cell13.data [7], _13707_);
  and (_00496_, _11993_, _11992_);
  or (_11995_, word_in[104], \oc8051_gm_cxrom_1.cell13.valid );
  or (_11997_, \oc8051_gm_cxrom_1.cell13.data [0], _11988_);
  and (_11998_, _11997_, _11995_);
  or (_11999_, _11998_, rst);
  or (_12000_, \oc8051_gm_cxrom_1.cell13.data [0], _13707_);
  and (_00503_, _12000_, _11999_);
  or (_12002_, word_in[105], \oc8051_gm_cxrom_1.cell13.valid );
  or (_12003_, \oc8051_gm_cxrom_1.cell13.data [1], _11988_);
  and (_12005_, _12003_, _12002_);
  or (_12006_, _12005_, rst);
  or (_12007_, \oc8051_gm_cxrom_1.cell13.data [1], _13707_);
  and (_00506_, _12007_, _12006_);
  or (_12009_, word_in[106], \oc8051_gm_cxrom_1.cell13.valid );
  or (_12010_, \oc8051_gm_cxrom_1.cell13.data [2], _11988_);
  and (_12012_, _12010_, _12009_);
  or (_12013_, _12012_, rst);
  or (_12014_, \oc8051_gm_cxrom_1.cell13.data [2], _13707_);
  and (_00510_, _12014_, _12013_);
  or (_12016_, word_in[107], \oc8051_gm_cxrom_1.cell13.valid );
  or (_12017_, \oc8051_gm_cxrom_1.cell13.data [3], _11988_);
  and (_12019_, _12017_, _12016_);
  or (_12020_, _12019_, rst);
  or (_12021_, \oc8051_gm_cxrom_1.cell13.data [3], _13707_);
  and (_00514_, _12021_, _12020_);
  or (_12023_, word_in[108], \oc8051_gm_cxrom_1.cell13.valid );
  or (_12025_, \oc8051_gm_cxrom_1.cell13.data [4], _11988_);
  and (_12026_, _12025_, _12023_);
  or (_12027_, _12026_, rst);
  or (_12028_, \oc8051_gm_cxrom_1.cell13.data [4], _13707_);
  and (_00517_, _12028_, _12027_);
  or (_12030_, word_in[109], \oc8051_gm_cxrom_1.cell13.valid );
  or (_12031_, \oc8051_gm_cxrom_1.cell13.data [5], _11988_);
  and (_12033_, _12031_, _12030_);
  or (_12034_, _12033_, rst);
  or (_12035_, \oc8051_gm_cxrom_1.cell13.data [5], _13707_);
  and (_00521_, _12035_, _12034_);
  or (_12037_, word_in[110], \oc8051_gm_cxrom_1.cell13.valid );
  or (_12038_, \oc8051_gm_cxrom_1.cell13.data [6], _11988_);
  and (_12040_, _12038_, _12037_);
  or (_12041_, _12040_, rst);
  or (_12042_, \oc8051_gm_cxrom_1.cell13.data [6], _13707_);
  and (_00524_, _12042_, _12041_);
  or (_12044_, \oc8051_gm_cxrom_1.cell14.valid , word_in[119]);
  not (_12045_, \oc8051_gm_cxrom_1.cell14.valid );
  or (_12047_, _12045_, \oc8051_gm_cxrom_1.cell14.data [7]);
  and (_12048_, _12047_, _12044_);
  or (_12049_, _12048_, rst);
  or (_12051_, \oc8051_gm_cxrom_1.cell14.data [7], _13707_);
  and (_13825_[7], _12051_, _12049_);
  or (_12052_, word_in[112], \oc8051_gm_cxrom_1.cell14.valid );
  or (_12053_, \oc8051_gm_cxrom_1.cell14.data [0], _12045_);
  and (_12054_, _12053_, _12052_);
  or (_12055_, _12054_, rst);
  or (_12056_, \oc8051_gm_cxrom_1.cell14.data [0], _13707_);
  and (_13825_[0], _12056_, _12055_);
  or (_12057_, word_in[113], \oc8051_gm_cxrom_1.cell14.valid );
  or (_12058_, \oc8051_gm_cxrom_1.cell14.data [1], _12045_);
  and (_12059_, _12058_, _12057_);
  or (_12060_, _12059_, rst);
  or (_12061_, \oc8051_gm_cxrom_1.cell14.data [1], _13707_);
  and (_13825_[1], _12061_, _12060_);
  or (_12062_, word_in[114], \oc8051_gm_cxrom_1.cell14.valid );
  or (_12063_, \oc8051_gm_cxrom_1.cell14.data [2], _12045_);
  and (_12064_, _12063_, _12062_);
  or (_12065_, _12064_, rst);
  or (_12066_, \oc8051_gm_cxrom_1.cell14.data [2], _13707_);
  and (_13825_[2], _12066_, _12065_);
  or (_12067_, word_in[115], \oc8051_gm_cxrom_1.cell14.valid );
  or (_12068_, \oc8051_gm_cxrom_1.cell14.data [3], _12045_);
  and (_12069_, _12068_, _12067_);
  or (_12070_, _12069_, rst);
  or (_12071_, \oc8051_gm_cxrom_1.cell14.data [3], _13707_);
  and (_13825_[3], _12071_, _12070_);
  or (_12072_, word_in[116], \oc8051_gm_cxrom_1.cell14.valid );
  or (_12073_, \oc8051_gm_cxrom_1.cell14.data [4], _12045_);
  and (_12074_, _12073_, _12072_);
  or (_12075_, _12074_, rst);
  or (_12076_, \oc8051_gm_cxrom_1.cell14.data [4], _13707_);
  and (_13825_[4], _12076_, _12075_);
  or (_12077_, word_in[117], \oc8051_gm_cxrom_1.cell14.valid );
  or (_12078_, \oc8051_gm_cxrom_1.cell14.data [5], _12045_);
  and (_12079_, _12078_, _12077_);
  or (_12080_, _12079_, rst);
  or (_12081_, \oc8051_gm_cxrom_1.cell14.data [5], _13707_);
  and (_13825_[5], _12081_, _12080_);
  or (_12082_, word_in[118], \oc8051_gm_cxrom_1.cell14.valid );
  or (_12083_, \oc8051_gm_cxrom_1.cell14.data [6], _12045_);
  and (_12084_, _12083_, _12082_);
  or (_12085_, _12084_, rst);
  or (_12086_, \oc8051_gm_cxrom_1.cell14.data [6], _13707_);
  and (_13825_[6], _12086_, _12085_);
  or (_12087_, \oc8051_gm_cxrom_1.cell15.valid , word_in[127]);
  not (_12088_, \oc8051_gm_cxrom_1.cell15.valid );
  or (_12089_, _12088_, \oc8051_gm_cxrom_1.cell15.data [7]);
  and (_12090_, _12089_, _12087_);
  or (_12091_, _12090_, rst);
  or (_12092_, \oc8051_gm_cxrom_1.cell15.data [7], _13707_);
  and (_13826_[7], _12092_, _12091_);
  or (_12093_, word_in[120], \oc8051_gm_cxrom_1.cell15.valid );
  or (_12094_, \oc8051_gm_cxrom_1.cell15.data [0], _12088_);
  and (_12095_, _12094_, _12093_);
  or (_12096_, _12095_, rst);
  or (_12097_, \oc8051_gm_cxrom_1.cell15.data [0], _13707_);
  and (_13826_[0], _12097_, _12096_);
  or (_12098_, word_in[121], \oc8051_gm_cxrom_1.cell15.valid );
  or (_12099_, \oc8051_gm_cxrom_1.cell15.data [1], _12088_);
  and (_12100_, _12099_, _12098_);
  or (_12101_, _12100_, rst);
  or (_12102_, \oc8051_gm_cxrom_1.cell15.data [1], _13707_);
  and (_13826_[1], _12102_, _12101_);
  or (_12103_, word_in[122], \oc8051_gm_cxrom_1.cell15.valid );
  or (_12104_, \oc8051_gm_cxrom_1.cell15.data [2], _12088_);
  and (_12105_, _12104_, _12103_);
  or (_12106_, _12105_, rst);
  or (_12107_, \oc8051_gm_cxrom_1.cell15.data [2], _13707_);
  and (_13826_[2], _12107_, _12106_);
  or (_12108_, word_in[123], \oc8051_gm_cxrom_1.cell15.valid );
  or (_12109_, \oc8051_gm_cxrom_1.cell15.data [3], _12088_);
  and (_12110_, _12109_, _12108_);
  or (_12111_, _12110_, rst);
  or (_12112_, \oc8051_gm_cxrom_1.cell15.data [3], _13707_);
  and (_13826_[3], _12112_, _12111_);
  or (_12113_, word_in[124], \oc8051_gm_cxrom_1.cell15.valid );
  or (_12114_, \oc8051_gm_cxrom_1.cell15.data [4], _12088_);
  and (_12115_, _12114_, _12113_);
  or (_12116_, _12115_, rst);
  or (_12117_, \oc8051_gm_cxrom_1.cell15.data [4], _13707_);
  and (_13826_[4], _12117_, _12116_);
  or (_12118_, word_in[125], \oc8051_gm_cxrom_1.cell15.valid );
  or (_12119_, \oc8051_gm_cxrom_1.cell15.data [5], _12088_);
  and (_12120_, _12119_, _12118_);
  or (_12121_, _12120_, rst);
  or (_12122_, \oc8051_gm_cxrom_1.cell15.data [5], _13707_);
  and (_13826_[5], _12122_, _12121_);
  or (_12123_, word_in[126], \oc8051_gm_cxrom_1.cell15.valid );
  or (_12124_, \oc8051_gm_cxrom_1.cell15.data [6], _12088_);
  and (_12125_, _12124_, _12123_);
  or (_12126_, _12125_, rst);
  or (_12127_, \oc8051_gm_cxrom_1.cell15.data [6], _13707_);
  and (_13826_[6], _12127_, _12126_);
  nor (_13913_[2], _08909_, rst);
  and (_12128_, _08527_, _13707_);
  nand (_12129_, _12128_, _08754_);
  nor (_12130_, _08804_, _08769_);
  or (_13914_[2], _12130_, _12129_);
  not (_12131_, _08689_);
  and (_12132_, _08714_, _12131_);
  not (_12133_, _08665_);
  and (_12134_, _08590_, _08566_);
  not (_12135_, _08638_);
  nor (_12136_, _12135_, _08614_);
  and (_12137_, _12136_, _12134_);
  and (_12138_, _12137_, _12133_);
  and (_12139_, _12138_, _12132_);
  not (_12140_, _08714_);
  and (_12141_, _12140_, _08689_);
  not (_12142_, _08590_);
  nor (_12143_, _12142_, _08566_);
  and (_12144_, _12143_, _12136_);
  and (_12145_, _12144_, _08665_);
  and (_12146_, _12145_, _12141_);
  or (_12147_, _12146_, _12139_);
  and (_12148_, _08714_, _08689_);
  and (_12149_, _08741_, _12133_);
  nor (_12150_, _08741_, _12133_);
  nor (_12151_, _12150_, _12149_);
  and (_12152_, _12151_, _12148_);
  and (_12153_, _12152_, _12144_);
  not (_12154_, _08741_);
  nor (_12155_, _08714_, _08689_);
  and (_12156_, _12155_, _12154_);
  and (_12157_, _12156_, _12144_);
  or (_12158_, _12157_, _12153_);
  nor (_12159_, _12133_, _08590_);
  and (_12160_, _12155_, _08741_);
  and (_12161_, _12160_, _12159_);
  and (_12162_, _12143_, _08614_);
  nor (_12163_, _08741_, _08665_);
  and (_12164_, _12155_, _12163_);
  and (_12165_, _12164_, _12162_);
  or (_12166_, _12165_, _12161_);
  and (_12167_, _12155_, _12150_);
  and (_12168_, _12167_, _12162_);
  not (_12169_, _08614_);
  and (_12170_, _12134_, _12169_);
  and (_12171_, _12150_, _12132_);
  and (_12172_, _12171_, _12170_);
  or (_12173_, _12172_, _12168_);
  or (_12174_, _12173_, _12166_);
  or (_12175_, _12174_, _12158_);
  or (_12176_, _12175_, _12147_);
  and (_12177_, _12141_, _12149_);
  and (_12178_, _12177_, _12144_);
  and (_12179_, _12148_, _12150_);
  and (_12180_, _12179_, _12144_);
  and (_12181_, _12143_, _12169_);
  not (_12182_, _12181_);
  and (_12183_, _12141_, _12163_);
  nor (_12184_, _12183_, _12135_);
  nor (_12185_, _12184_, _12182_);
  or (_12186_, _12185_, _12180_);
  nor (_12187_, _12186_, _12178_);
  and (_12188_, _12149_, _12132_);
  and (_12189_, _12144_, _12188_);
  and (_12190_, _12132_, _08741_);
  and (_12191_, _12162_, _12135_);
  and (_12192_, _12191_, _12190_);
  and (_12193_, _12162_, _08638_);
  and (_12194_, _12148_, _08741_);
  and (_12195_, _12194_, _12193_);
  or (_12196_, _12195_, _12192_);
  or (_12197_, _12196_, _12189_);
  and (_12198_, _12150_, _12141_);
  and (_12199_, _12191_, _12198_);
  and (_12200_, _12148_, _12154_);
  and (_12201_, _12193_, _12200_);
  or (_12202_, _12201_, _12199_);
  and (_12203_, _12160_, _08665_);
  and (_12204_, _12170_, _12135_);
  and (_12205_, _12204_, _12203_);
  and (_12206_, _12132_, _12154_);
  not (_12207_, _12206_);
  and (_12208_, _08665_, _08614_);
  and (_12209_, _12208_, _12134_);
  nor (_12210_, _12209_, _12159_);
  nor (_12211_, _12210_, _12207_);
  or (_12212_, _12211_, _12205_);
  or (_12213_, _12212_, _12202_);
  nor (_12214_, _12213_, _12197_);
  nand (_12215_, _12214_, _12187_);
  or (_12216_, _12215_, _12176_);
  and (_12217_, _12216_, _08528_);
  not (_12218_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_12219_, _08526_, _06841_);
  and (_12220_, _12219_, _08846_);
  nor (_12221_, _12220_, _12218_);
  or (_12222_, _12221_, rst);
  or (_13915_[1], _12222_, _12217_);
  nand (_12223_, _08689_, _08521_);
  or (_12224_, _08521_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and (_12225_, _12224_, _13707_);
  and (_13916_[7], _12225_, _12223_);
  and (_12226_, \oc8051_top_1.oc8051_sfr1.wait_data , _13707_);
  and (_12227_, _12226_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_12228_, _08902_, _08755_);
  and (_12229_, _08886_, _08821_);
  and (_12230_, _12229_, _08669_);
  or (_12231_, _12230_, _12228_);
  and (_12232_, _08824_, _08804_);
  or (_12233_, _12232_, _08852_);
  or (_12234_, _12233_, _08817_);
  and (_12235_, _08782_, _08769_);
  and (_12236_, _08886_, _08790_);
  or (_12237_, _12236_, _12235_);
  nor (_12238_, _12237_, _12234_);
  nand (_12239_, _12238_, _08839_);
  or (_12240_, _12239_, _12231_);
  and (_12241_, _12240_, _12128_);
  or (_13917_, _12241_, _12227_);
  and (_12242_, _08746_, _08759_);
  nor (_12243_, _08670_, _08595_);
  and (_12244_, _12243_, _12242_);
  and (_12245_, _12244_, _08695_);
  or (_12246_, _12245_, _08872_);
  and (_12247_, _08619_, _08596_);
  and (_12248_, _12247_, _08790_);
  or (_12249_, _12248_, _12246_);
  and (_12250_, _08804_, _08822_);
  or (_12251_, _12250_, _08887_);
  or (_12252_, _12251_, _12249_);
  and (_12253_, _12252_, _08527_);
  and (_12254_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_12255_, \oc8051_top_1.oc8051_decoder1.state [0], _06841_);
  and (_12256_, _12255_, _12218_);
  and (_12257_, _08906_, _12256_);
  or (_12258_, _12257_, _12254_);
  or (_12259_, _12258_, _12253_);
  and (_13918_[1], _12259_, _13707_);
  and (_12260_, _12226_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and (_12261_, _08902_, _08773_);
  or (_12262_, _08782_, _08773_);
  and (_12263_, _12262_, _08646_);
  or (_12264_, _12263_, _12261_);
  and (_12265_, _12247_, _08800_);
  or (_12266_, _12265_, _12264_);
  nor (_12267_, _08669_, _08595_);
  and (_12268_, _12267_, _08772_);
  and (_12269_, _12262_, _08775_);
  or (_12270_, _12269_, _12268_);
  or (_12271_, _12270_, _08880_);
  and (_12272_, _12267_, _08748_);
  and (_12273_, _08902_, _08721_);
  or (_12274_, _12273_, _12272_);
  or (_12275_, _12274_, _12251_);
  or (_12276_, _12275_, _12271_);
  or (_12277_, _12276_, _12266_);
  and (_12278_, _12277_, _12128_);
  or (_13919_[1], _12278_, _12260_);
  and (_12279_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_12280_, _08825_, _08527_);
  or (_12281_, _12280_, _12279_);
  or (_12282_, _12281_, _12257_);
  and (_13920_[2], _12282_, _13707_);
  not (_12283_, _12130_);
  and (_12284_, _12283_, _08755_);
  nor (_12285_, _12284_, _12229_);
  not (_12286_, _12285_);
  and (_12287_, _12286_, _12256_);
  or (_12288_, _12287_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_12289_, _08768_, _08645_);
  and (_12290_, _08772_, _08770_);
  nor (_12291_, _12290_, _12289_);
  nor (_12292_, _12291_, _08669_);
  and (_12293_, _12230_, _08523_);
  or (_12294_, _12293_, _12292_);
  and (_12295_, _12294_, _08846_);
  or (_12296_, _12295_, _12288_);
  or (_12297_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2], _06841_);
  and (_12298_, _12297_, _13707_);
  and (_13921_[2], _12298_, _12296_);
  and (_12299_, _12226_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  or (_12300_, _12268_, _08887_);
  and (_12301_, _08782_, _08775_);
  or (_12302_, _12301_, _08810_);
  or (_12303_, _12302_, _12300_);
  and (_12304_, _08770_, _08748_);
  or (_12305_, _12265_, _12235_);
  or (_12306_, _12305_, _12304_);
  or (_12307_, _08800_, _08790_);
  and (_12308_, _12307_, _08750_);
  or (_12309_, _12245_, _08791_);
  or (_12310_, _12309_, _12308_);
  or (_12311_, _12310_, _12306_);
  or (_12312_, _12311_, _12303_);
  and (_12313_, _12312_, _12128_);
  or (_13922_[1], _12313_, _12299_);
  and (_12314_, _12226_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  or (_12315_, _12248_, _08805_);
  and (_12316_, _08886_, _08763_);
  and (_12317_, _12247_, _08788_);
  or (_12318_, _12317_, _12316_);
  or (_12319_, _12318_, _12315_);
  or (_12320_, _12319_, _12270_);
  and (_12321_, _08782_, _08750_);
  and (_12322_, _12242_, _08751_);
  or (_12323_, _12322_, _08866_);
  or (_12324_, _12323_, _12321_);
  and (_12325_, _08902_, _08797_);
  or (_12326_, _08809_, _08798_);
  or (_12327_, _12326_, _12325_);
  or (_12328_, _12327_, _12324_);
  or (_12329_, _12328_, _12320_);
  nor (_12330_, _08879_, _08828_);
  not (_12331_, _12330_);
  not (_12332_, _08815_);
  and (_12333_, _08788_, _08775_);
  or (_12334_, _12333_, _12244_);
  or (_12335_, _12334_, _12332_);
  or (_12336_, _12335_, _12331_);
  or (_12337_, _12336_, _12266_);
  or (_12338_, _12337_, _12329_);
  and (_12339_, _12338_, _12128_);
  or (_13923_[3], _12339_, _12314_);
  and (_12340_, _08764_, _08750_);
  and (_12341_, _12267_, _08821_);
  and (_12342_, _12247_, _08764_);
  or (_12343_, _12342_, _12341_);
  or (_12344_, _12343_, _12340_);
  and (_12345_, _08764_, _08775_);
  or (_12346_, _12345_, _08876_);
  or (_12347_, _12346_, _12344_);
  and (_12348_, _12247_, _08822_);
  or (_12349_, _12348_, _08906_);
  or (_12350_, _12349_, _12347_);
  and (_12351_, _12350_, _12128_);
  nor (_12352_, _08905_, _08523_);
  and (_12353_, \oc8051_top_1.oc8051_sfr1.wait_data , \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or (_12354_, _12353_, _12352_);
  and (_12355_, _12354_, _13707_);
  or (_13924_[1], _12355_, _12351_);
  or (_12356_, _08791_, _08783_);
  not (_12357_, _08818_);
  or (_12358_, _12263_, _12357_);
  or (_12359_, _12358_, _12356_);
  and (_12360_, _08800_, _08770_);
  nor (_12361_, _08746_, _08719_);
  and (_12362_, _12361_, _08670_);
  and (_12363_, _12362_, _08646_);
  or (_12364_, _12363_, _08801_);
  or (_12365_, _12364_, _08798_);
  or (_12366_, _12365_, _12360_);
  or (_12367_, _12366_, _08830_);
  or (_12368_, _12367_, _12359_);
  or (_12369_, _08870_, _08777_);
  or (_12370_, _12369_, _08832_);
  or (_12371_, _12370_, _12246_);
  and (_12372_, _08875_, _12361_);
  or (_12373_, _12372_, _08879_);
  or (_12374_, _12373_, _08752_);
  and (_12375_, _12289_, _08670_);
  and (_12376_, _12267_, _12361_);
  or (_12377_, _12376_, _12375_);
  and (_12378_, _08824_, _08775_);
  or (_12379_, _12378_, _12377_);
  or (_12380_, _12379_, _12374_);
  or (_12381_, _12380_, _12371_);
  or (_12382_, _12381_, _12270_);
  or (_12383_, _12382_, _12368_);
  and (_12384_, _12383_, _08527_);
  and (_12385_, \oc8051_top_1.oc8051_decoder1.wr , \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_12386_, _08848_, _08849_);
  or (_12387_, _12360_, _12375_);
  and (_12388_, _12387_, _08848_);
  or (_12389_, _12388_, _12257_);
  or (_12390_, _12389_, _12386_);
  or (_12391_, _12390_, _12385_);
  or (_12392_, _12391_, _12384_);
  and (_13925_, _12392_, _13707_);
  and (_13913_[0], _08898_, _13707_);
  nor (_13913_[1], _08858_, rst);
  nand (_13914_[0], _12286_, _12128_);
  nand (_12393_, _12229_, _12128_);
  not (_12394_, _08804_);
  or (_12395_, _12129_, _12394_);
  and (_13914_[1], _12395_, _12393_);
  or (_12396_, _12201_, \oc8051_top_1.oc8051_decoder1.state [1]);
  or (_12397_, _12396_, _12192_);
  or (_12398_, _12397_, _12139_);
  and (_12399_, _12398_, _12220_);
  nor (_12400_, _12219_, _08846_);
  or (_12401_, _12400_, rst);
  or (_13915_[0], _12401_, _12399_);
  nand (_12402_, _08638_, _08521_);
  or (_12403_, _08521_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and (_12404_, _12403_, _13707_);
  and (_13916_[0], _12404_, _12402_);
  not (_12405_, _08521_);
  or (_12406_, _08614_, _12405_);
  or (_12407_, _08521_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and (_12408_, _12407_, _13707_);
  and (_13916_[1], _12408_, _12406_);
  or (_12409_, _08566_, _12405_);
  or (_12410_, _08521_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and (_12411_, _12410_, _13707_);
  and (_13916_[2], _12411_, _12409_);
  nand (_12412_, _08590_, _08521_);
  or (_12413_, _08521_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and (_12414_, _12413_, _13707_);
  and (_13916_[3], _12414_, _12412_);
  or (_12415_, _08665_, _12405_);
  or (_12416_, _08521_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and (_12417_, _12416_, _13707_);
  and (_13916_[4], _12417_, _12415_);
  nand (_12418_, _08741_, _08521_);
  or (_12419_, _08521_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and (_12420_, _12419_, _13707_);
  and (_13916_[5], _12420_, _12418_);
  nand (_12421_, _08714_, _08521_);
  or (_12422_, _08521_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and (_12423_, _12422_, _13707_);
  and (_13916_[6], _12423_, _12421_);
  and (_12424_, _12267_, _08761_);
  or (_12425_, _12424_, _12345_);
  or (_12426_, _12425_, _12344_);
  and (_12427_, _12247_, _08797_);
  or (_12428_, _12427_, _12250_);
  or (_12429_, _08782_, _08772_);
  and (_12430_, _12429_, _08902_);
  or (_12431_, _12430_, _12428_);
  or (_12432_, _12431_, _12426_);
  or (_12433_, _08864_, _08756_);
  or (_12434_, _12333_, _12228_);
  or (_12435_, _12434_, _12433_);
  and (_12436_, _12243_, _08761_);
  and (_12437_, _08750_, _08822_);
  or (_12438_, _12348_, _12437_);
  or (_12439_, _12438_, _12436_);
  or (_12440_, _08887_, _08866_);
  or (_12441_, _12440_, _12439_);
  or (_12442_, _12441_, _12435_);
  and (_12443_, _12247_, _08762_);
  and (_12444_, _08754_, _08670_);
  and (_12445_, _12444_, _08902_);
  and (_12446_, _08762_, _08750_);
  or (_12447_, _12446_, _12445_);
  or (_12448_, _12447_, _12443_);
  and (_12449_, _08902_, _08808_);
  and (_12450_, _08755_, _08775_);
  or (_12451_, _12450_, _12449_);
  or (_12452_, _12451_, _12318_);
  or (_12453_, _12452_, _12448_);
  or (_12454_, _12453_, _12442_);
  or (_12455_, _12454_, _12432_);
  and (_12456_, _12455_, _08527_);
  and (_12457_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_12458_, _12457_, _12287_);
  or (_12459_, _12458_, _12456_);
  and (_13918_[0], _12459_, _13707_);
  and (_12460_, _12226_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  or (_12461_, _08797_, _08788_);
  and (_12462_, _12461_, _08770_);
  or (_12463_, _12428_, _12334_);
  or (_12464_, _12463_, _12462_);
  nor (_12465_, _12272_, _08878_);
  not (_12466_, _12465_);
  or (_12467_, _12466_, _12273_);
  or (_12468_, _12467_, _08792_);
  or (_12469_, _12468_, _12231_);
  or (_12470_, _08788_, _08765_);
  and (_12471_, _12470_, _08902_);
  or (_12472_, _12471_, _12324_);
  or (_12473_, _12472_, _12469_);
  or (_12474_, _12473_, _12464_);
  and (_12475_, _12474_, _12128_);
  or (_13919_[0], _12475_, _12460_);
  or (_12476_, _12375_, _08870_);
  or (_12477_, _12476_, _12378_);
  or (_12478_, _12477_, _08832_);
  or (_12479_, _12478_, _12368_);
  and (_12480_, _12479_, _08527_);
  and (_12481_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_12482_, _12481_, _12390_);
  or (_12483_, _12482_, _12480_);
  and (_13920_[0], _12483_, _13707_);
  and (_12484_, _08827_, _08669_);
  or (_12485_, _12484_, _08872_);
  or (_12486_, _12485_, _12374_);
  or (_12487_, _12486_, _12292_);
  and (_12488_, _12487_, _08527_);
  and (_12489_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_12490_, _12489_, _12389_);
  or (_12491_, _12490_, _12488_);
  and (_13920_[1], _12491_, _13707_);
  or (_12492_, _12461_, _08808_);
  and (_12493_, _12492_, _08902_);
  or (_12494_, _12493_, _12292_);
  or (_12495_, _12341_, _08869_);
  or (_12496_, _12229_, _08904_);
  and (_12497_, _12342_, _08670_);
  or (_12498_, _12497_, _12443_);
  or (_12499_, _12498_, _12496_);
  or (_12500_, _12499_, _12495_);
  or (_12501_, _12500_, _12494_);
  and (_12502_, _08902_, _08790_);
  or (_12503_, _12348_, _12316_);
  or (_12504_, _12503_, _12502_);
  or (_12505_, _12504_, _12425_);
  and (_12506_, _12247_, _08802_);
  or (_12507_, _12506_, _12228_);
  or (_12508_, _12445_, _08903_);
  or (_12509_, _12508_, _12430_);
  or (_12510_, _12509_, _12507_);
  and (_12511_, _12444_, _08646_);
  and (_12512_, _12342_, _08669_);
  or (_12513_, _12512_, _08888_);
  or (_12514_, _12513_, _12511_);
  and (_12515_, _08832_, _08643_);
  or (_12516_, _12376_, _12437_);
  or (_12517_, _12516_, _12372_);
  or (_12518_, _12517_, _12515_);
  or (_12519_, _12518_, _12514_);
  or (_12520_, _12519_, _12510_);
  or (_12521_, _12520_, _12505_);
  or (_12522_, _12521_, _12501_);
  and (_12523_, _12522_, _08527_);
  and (_12524_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_12525_, _12287_, _12352_);
  or (_12526_, _12525_, _12524_);
  or (_12527_, _12526_, _12523_);
  and (_13921_[0], _12527_, _13707_);
  or (_12528_, _08904_, _12437_);
  or (_12529_, _12363_, _12250_);
  or (_12530_, _12529_, _12528_);
  or (_12531_, _08873_, _08775_);
  and (_12532_, _12531_, _12444_);
  or (_12533_, _12532_, _08832_);
  or (_12534_, _12533_, _12530_);
  or (_12535_, _08891_, _08766_);
  or (_12536_, _12535_, _12534_);
  or (_12537_, _08828_, _08798_);
  and (_12538_, _12537_, _08644_);
  or (_12539_, _12538_, _12495_);
  or (_12540_, _12539_, _12536_);
  or (_12541_, _12510_, _12505_);
  or (_12542_, _12541_, _12540_);
  and (_12543_, _12542_, _08527_);
  and (_12544_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_12545_, _12544_, _12525_);
  or (_12546_, _12545_, _12543_);
  and (_13921_[1], _12546_, _13707_);
  and (_12547_, _12226_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  and (_12548_, _12316_, _08747_);
  and (_12549_, _12548_, _08670_);
  or (_12550_, _12549_, _12303_);
  not (_12551_, _10034_);
  or (_12552_, _12348_, _12551_);
  and (_12553_, _08886_, _08772_);
  and (_12554_, _12553_, _08670_);
  and (_12555_, _12235_, _08644_);
  or (_12556_, _12555_, _12554_);
  or (_12557_, _12556_, _12552_);
  or (_12558_, _12557_, _12550_);
  and (_12559_, _08902_, _08782_);
  or (_12560_, _12559_, _12265_);
  or (_12561_, _12356_, _12308_);
  or (_12562_, _12561_, _12560_);
  and (_12563_, _08886_, _08802_);
  or (_12564_, _12563_, _12497_);
  or (_12565_, _12341_, _12245_);
  and (_12566_, _12340_, _08670_);
  or (_12567_, _12566_, _12565_);
  or (_12568_, _12567_, _12564_);
  and (_12569_, _08836_, _08775_);
  or (_12570_, _12569_, _12437_);
  nor (_12571_, _12570_, _08823_);
  nand (_12572_, _12571_, _10035_);
  or (_12573_, _12572_, _12568_);
  or (_12574_, _12573_, _12562_);
  or (_12575_, _12574_, _12558_);
  and (_12576_, _12575_, _12128_);
  or (_13922_[0], _12576_, _12547_);
  or (_12577_, _12322_, _12248_);
  or (_12578_, _12321_, _08813_);
  or (_12579_, _12578_, _12577_);
  or (_12580_, _12244_, _10128_);
  or (_12581_, _12580_, _08887_);
  or (_12582_, _12581_, _12513_);
  or (_12583_, _12582_, _12579_);
  or (_12584_, _12499_, _12327_);
  or (_12585_, _12584_, _12583_);
  or (_12586_, _12549_, _12559_);
  or (_12587_, _08869_, _08833_);
  or (_12588_, _12554_, _12425_);
  or (_12589_, _12588_, _12587_);
  or (_12590_, _12589_, _12586_);
  or (_12591_, _12590_, _12585_);
  or (_12592_, _08904_, _08523_);
  or (_12593_, \oc8051_top_1.oc8051_decoder1.alu_op [0], _06841_);
  and (_12594_, _12593_, _13707_);
  and (_12595_, _12594_, _12592_);
  and (_13923_[0], _12595_, _12591_);
  and (_12596_, _12226_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  nor (_12597_, _12443_, _08832_);
  not (_12598_, _12597_);
  nor (_12599_, _12598_, _08831_);
  or (_12600_, _12248_, _08877_);
  or (_12601_, _12600_, _12565_);
  or (_12602_, _08904_, _08814_);
  or (_12603_, _12348_, _12272_);
  or (_12604_, _12603_, _12602_);
  or (_12605_, _12604_, _12507_);
  nor (_12606_, _12605_, _12601_);
  nand (_12607_, _12606_, _12599_);
  and (_12608_, _08769_, _08802_);
  or (_12609_, _12608_, _12445_);
  or (_12610_, _12446_, _12424_);
  or (_12611_, _12610_, _12548_);
  or (_12612_, _12611_, _12609_);
  or (_12613_, _12612_, _12271_);
  or (_12614_, _12613_, _12266_);
  or (_12615_, _12614_, _12607_);
  nor (_12616_, \oc8051_top_1.oc8051_sfr1.wait_data , rst);
  and (_12617_, _12616_, _12592_);
  and (_12618_, _12617_, _12615_);
  or (_13923_[1], _12618_, _12596_);
  or (_12619_, _12610_, _12598_);
  or (_12620_, _12619_, _12609_);
  or (_12621_, _08879_, _08872_);
  nor (_12622_, _12621_, _12553_);
  nand (_12623_, _12622_, _10034_);
  or (_12624_, _12560_, _12309_);
  or (_12625_, _12624_, _12623_);
  or (_12626_, _12270_, _12264_);
  or (_12627_, _12626_, _12625_);
  or (_12628_, _12627_, _12620_);
  and (_12629_, _12628_, _08527_);
  and (_12630_, \oc8051_top_1.oc8051_decoder1.alu_op [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_12631_, _08903_, _06841_);
  or (_12632_, _12631_, _12630_);
  or (_12633_, _12632_, _12629_);
  and (_13923_[2], _12633_, _13707_);
  and (_12634_, _12226_, \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  or (_12635_, _12552_, _12347_);
  or (_12636_, _12635_, _12556_);
  not (_12637_, _08768_);
  or (_12638_, _08886_, _12637_);
  and (_12639_, _12638_, _08802_);
  nor (_12640_, _12236_, _08784_);
  nand (_12641_, _12640_, _10035_);
  or (_12642_, _12641_, _12639_);
  or (_12643_, _12642_, _12586_);
  or (_12644_, _12643_, _12636_);
  and (_12645_, _12644_, _12128_);
  or (_13924_[0], _12645_, _12634_);
  nor (_13910_[7], _08689_, rst);
  nor (_13911_[7], _10265_, rst);
  and (_12646_, _10128_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [7]);
  and (_12647_, _08533_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  and (_12648_, _08545_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and (_12649_, _08537_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor (_12650_, _12649_, _12648_);
  and (_12651_, _08557_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_12652_, _08552_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_12653_, _12652_, _12651_);
  and (_12654_, _08548_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_12655_, _08541_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor (_12656_, _12655_, _12654_);
  and (_12657_, _12656_, _12653_);
  and (_12658_, _12657_, _12650_);
  nor (_12659_, _12658_, _08533_);
  nor (_12660_, _12659_, _12647_);
  nor (_12661_, _12660_, _10128_);
  nor (_12662_, _12661_, _12646_);
  nor (_13912_[7], _12662_, rst);
  nor (_13910_[0], _08638_, rst);
  and (_13910_[1], _08614_, _13707_);
  and (_13910_[2], _08566_, _13707_);
  nor (_13910_[3], _08590_, rst);
  and (_13910_[4], _08665_, _13707_);
  nor (_13910_[5], _08741_, rst);
  nor (_13910_[6], _08714_, rst);
  nor (_13911_[0], _10319_, rst);
  nor (_13911_[1], _10479_, rst);
  nor (_13911_[2], _10144_, rst);
  nor (_13911_[3], _10367_, rst);
  nor (_13911_[4], _10526_, rst);
  nor (_13911_[5], _10191_, rst);
  nor (_13911_[6], _10423_, rst);
  and (_12663_, _10128_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [0]);
  and (_12664_, _08533_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  and (_12665_, _08545_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and (_12666_, _08537_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_12667_, _12666_, _12665_);
  and (_12668_, _08557_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_12669_, _08552_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_12670_, _12669_, _12668_);
  and (_12671_, _08548_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_12672_, _08541_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor (_12673_, _12672_, _12671_);
  and (_12674_, _12673_, _12670_);
  and (_12675_, _12674_, _12667_);
  nor (_12676_, _12675_, _08533_);
  nor (_12677_, _12676_, _12664_);
  nor (_12678_, _12677_, _10128_);
  nor (_12679_, _12678_, _12663_);
  nor (_13912_[0], _12679_, rst);
  and (_12680_, _10128_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [1]);
  and (_12681_, _08533_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  and (_12682_, _08557_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_12683_, _08537_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_12684_, _12683_, _12682_);
  and (_12685_, _08548_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_12686_, _08541_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nor (_12687_, _12686_, _12685_);
  and (_12688_, _12687_, _12684_);
  and (_12689_, _08545_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and (_12690_, _08552_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_12691_, _12690_, _12689_);
  and (_12692_, _12691_, _12688_);
  nor (_12693_, _12692_, _08533_);
  nor (_12694_, _12693_, _12681_);
  nor (_12695_, _12694_, _10128_);
  nor (_12696_, _12695_, _12680_);
  nor (_13912_[1], _12696_, rst);
  and (_12697_, _10128_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [2]);
  and (_12698_, _08533_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  and (_12699_, _08545_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and (_12700_, _08537_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_12701_, _12700_, _12699_);
  and (_12702_, _08557_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_12703_, _08552_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_12704_, _12703_, _12702_);
  and (_12705_, _08548_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_12706_, _08541_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor (_12707_, _12706_, _12705_);
  and (_12708_, _12707_, _12704_);
  and (_12709_, _12708_, _12701_);
  nor (_12710_, _12709_, _08533_);
  nor (_12711_, _12710_, _12698_);
  nor (_12712_, _12711_, _10128_);
  nor (_12713_, _12712_, _12697_);
  nor (_13912_[2], _12713_, rst);
  and (_12714_, _10128_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [3]);
  and (_12715_, _08533_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  and (_12716_, _08545_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and (_12717_, _08537_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_12718_, _12717_, _12716_);
  and (_12719_, _08557_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_12720_, _08552_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_12721_, _12720_, _12719_);
  and (_12722_, _08548_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_12723_, _08541_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor (_12724_, _12723_, _12722_);
  and (_12725_, _12724_, _12721_);
  and (_12726_, _12725_, _12718_);
  nor (_12727_, _12726_, _08533_);
  nor (_12728_, _12727_, _12715_);
  nor (_12729_, _12728_, _10128_);
  nor (_12730_, _12729_, _12714_);
  nor (_13912_[3], _12730_, rst);
  and (_12731_, _10128_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [4]);
  and (_12732_, _08533_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  and (_12733_, _08548_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_12734_, _08552_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_12735_, _12734_, _12733_);
  and (_12736_, _08545_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and (_12737_, _08541_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor (_12738_, _12737_, _12736_);
  and (_12739_, _08537_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  and (_12740_, _08557_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nor (_12741_, _12740_, _12739_);
  and (_12742_, _12741_, _12738_);
  and (_12743_, _12742_, _12735_);
  nor (_12744_, _12743_, _08533_);
  nor (_12745_, _12744_, _12732_);
  nor (_12746_, _12745_, _10128_);
  nor (_12747_, _12746_, _12731_);
  nor (_13912_[4], _12747_, rst);
  and (_12748_, _10128_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [5]);
  and (_12749_, _08533_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  and (_12750_, _08548_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_12751_, _08552_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_12752_, _12751_, _12750_);
  and (_12753_, _08545_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and (_12754_, _08541_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor (_12755_, _12754_, _12753_);
  and (_12756_, _08537_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  and (_12757_, _08557_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  nor (_12758_, _12757_, _12756_);
  and (_12759_, _12758_, _12755_);
  and (_12760_, _12759_, _12752_);
  nor (_12761_, _12760_, _08533_);
  nor (_12762_, _12761_, _12749_);
  nor (_12763_, _12762_, _10128_);
  nor (_12764_, _12763_, _12748_);
  nor (_13912_[5], _12764_, rst);
  and (_12765_, _10128_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [6]);
  and (_12766_, _08533_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  and (_12767_, _08557_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_12768_, _08537_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor (_12769_, _12768_, _12767_);
  and (_12770_, _08548_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_12771_, _08541_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor (_12772_, _12771_, _12770_);
  and (_12773_, _12772_, _12769_);
  and (_12774_, _08545_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and (_12775_, _08552_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_12776_, _12775_, _12774_);
  and (_12777_, _12776_, _12773_);
  nor (_12778_, _12777_, _08533_);
  nor (_12779_, _12778_, _12766_);
  nor (_12780_, _12779_, _10128_);
  nor (_12781_, _12780_, _12765_);
  nor (_13912_[6], _12781_, rst);
  and (_12782_, _08528_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  or (_12783_, _12782_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nand (_12784_, _12782_, _07092_);
  and (_12785_, _12784_, _13707_);
  and (_13927_[15], _12785_, _12783_);
  not (_12786_, _12782_);
  or (_12787_, _12786_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  and (_00002_, _12782_, _13707_);
  and (_12788_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _13707_);
  or (_12789_, _12788_, _00002_);
  and (_13928_[15], _12789_, _12787_);
  nor (_13929_, _10271_, rst);
  and (_13930_, \oc8051_top_1.oc8051_memory_interface1.dstb_o , _13707_);
  nor (_13931_[4], _10531_, rst);
  and (_13932_[7], _10250_, _13707_);
  and (_12790_, _10271_, _07695_);
  nor (_12791_, _10271_, _07695_);
  or (_12792_, _12791_, _12790_);
  not (_12793_, _10429_);
  nor (_12794_, _12793_, _07666_);
  and (_12795_, _12793_, _07666_);
  or (_12796_, _12795_, _12794_);
  or (_12797_, _12796_, _12792_);
  nor (_12798_, _10537_, _07724_);
  and (_12799_, _10537_, _07724_);
  or (_12800_, _12799_, _12798_);
  and (_12801_, _10199_, _09489_);
  nor (_12802_, _10199_, _09489_);
  or (_12803_, _12802_, _12801_);
  or (_12804_, _12803_, _12800_);
  or (_12805_, _12804_, _12797_);
  and (_12806_, _10372_, _10045_);
  nor (_12807_, _10372_, _10045_);
  or (_12808_, _12807_, _12806_);
  nor (_12809_, _12808_, _12805_);
  or (_12810_, _10324_, _07738_);
  nand (_12811_, _10324_, _07738_);
  and (_12812_, _12811_, _12810_);
  nor (_12813_, _12812_, _09680_);
  and (_12814_, _10485_, _08235_);
  nor (_12815_, _10485_, _08235_);
  or (_12816_, _12815_, _12814_);
  or (_12817_, _10149_, _07761_);
  nand (_12818_, _10149_, _07761_);
  and (_12819_, _12818_, _12817_);
  nor (_12820_, _12819_, _12816_);
  and (_12821_, _12820_, _12813_);
  and (_12822_, _12821_, _12809_);
  nor (_12823_, _07694_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_12824_, _12823_, _12822_);
  not (_12825_, _12824_);
  nor (_12826_, _08839_, _12255_);
  and (_12827_, _08507_, _08008_);
  and (_12828_, _12827_, _12826_);
  and (_12829_, _12828_, _12809_);
  and (_12830_, _08195_, _07822_);
  nand (_12831_, _12830_, _08249_);
  nor (_12832_, _12831_, _08312_);
  and (_12833_, _12832_, _08380_);
  and (_12834_, _12833_, _08459_);
  and (_12835_, _10203_, _10218_);
  nor (_12836_, _12835_, _12255_);
  or (_12837_, _12836_, _08853_);
  nor (_12838_, _12837_, _08074_);
  and (_12839_, _12838_, _12834_);
  and (_12840_, _12839_, _07876_);
  and (_12841_, _12826_, _07854_);
  nor (_12842_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_12843_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_12844_, _12843_, _12842_);
  nor (_12845_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor (_12846_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_12847_, _12846_, _12845_);
  and (_12848_, _12847_, _12844_);
  and (_12849_, _12848_, _08895_);
  or (_12850_, _12826_, _08746_);
  and (_12851_, _12850_, _08853_);
  and (_12852_, _12851_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or (_12853_, _12852_, _12849_);
  or (_12854_, _12853_, _12841_);
  nor (_12855_, _12854_, _12840_);
  or (_12856_, _12506_, _08810_);
  nor (_12857_, _12856_, _12301_);
  or (_12858_, _08808_, _08836_);
  or (_12859_, _12858_, _08762_);
  nand (_12860_, _12859_, _08804_);
  and (_12861_, _12860_, _12465_);
  nand (_12862_, _12861_, _12857_);
  nand (_12863_, _12862_, _12855_);
  nor (_12864_, _08849_, _10217_);
  nand (_12865_, _08852_, _08669_);
  and (_12866_, _12865_, _12864_);
  or (_12867_, _12866_, _12855_);
  nor (_12868_, _08619_, _08571_);
  and (_12869_, _08644_, _08595_);
  and (_12870_, _12869_, _12868_);
  and (_12871_, _12870_, _08808_);
  nor (_12872_, _12871_, _12232_);
  and (_12873_, _12872_, _12867_);
  and (_12874_, _12873_, _12863_);
  or (_12875_, _12874_, _10204_);
  nor (_12876_, _12291_, _08522_);
  not (_12877_, _12876_);
  and (_12878_, _12877_, _08854_);
  and (_12879_, _12878_, _12875_);
  or (_12880_, _09507_, _09501_);
  and (_12881_, _12880_, _08895_);
  not (_12882_, _09378_);
  or (_12883_, _09388_, _12882_);
  or (_12884_, _12883_, _09383_);
  and (_12885_, _12884_, _12851_);
  or (_12886_, _12885_, _12881_);
  nor (_12887_, _12886_, _12879_);
  not (_12888_, _12887_);
  nor (_12889_, _12888_, _12829_);
  and (_12890_, _12889_, _12825_);
  nor (_12891_, _08855_, rst);
  and (_13935_, _12891_, _12890_);
  and (_13936_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _13707_);
  nor (_12892_, \oc8051_top_1.oc8051_memory_interface1.dstb_o , rst);
  and (_12893_, _12892_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [7]);
  and (_12894_, _13930_, xram_data_in_reg[7]);
  or (_13937_[7], _12894_, _12893_);
  nor (_12895_, _08555_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_12896_, _12895_, _10128_);
  nor (_12897_, _12896_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  not (_12898_, _12897_);
  and (_12899_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and (_12900_, _12899_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and (_12901_, _12900_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and (_12902_, _12901_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_12903_, _12902_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and (_12904_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9], \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_12905_, _12904_, _12903_);
  and (_12906_, _12905_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_12907_, _12906_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and (_12908_, _12907_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and (_12909_, _12908_, _12898_);
  and (_12910_, _12909_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and (_12911_, _12910_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or (_12912_, _12911_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nand (_12913_, _12911_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_12914_, _12913_, _12912_);
  or (_12915_, _12914_, _12890_);
  and (_12916_, _12915_, _13707_);
  nor (_12917_, _12856_, _12466_);
  nand (_12918_, _12917_, _12835_);
  nand (_12919_, _12918_, _08848_);
  and (_12920_, _12290_, _08523_);
  and (_12921_, _08834_, _08523_);
  or (_12922_, _12921_, _12920_);
  nor (_12923_, _12922_, _08855_);
  and (_12924_, _12923_, _12919_);
  and (_12925_, _12924_, _10265_);
  not (_12926_, _12662_);
  nor (_12927_, _12924_, _12926_);
  nor (_12928_, _12927_, _12925_);
  not (_12929_, _12928_);
  and (_12930_, _12928_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor (_12931_, _12928_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_12932_, _12924_, _10423_);
  not (_12933_, _12781_);
  nor (_12934_, _12924_, _12933_);
  nor (_12935_, _12934_, _12932_);
  and (_12936_, _12935_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  not (_12937_, _12936_);
  nor (_12938_, _12935_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_12939_, _12938_, _12936_);
  and (_12940_, _12924_, _10191_);
  not (_12941_, _12764_);
  nor (_12942_, _12924_, _12941_);
  nor (_12943_, _12942_, _12940_);
  nor (_12944_, _12943_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_12945_, _12943_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_12946_, _12924_, _10526_);
  not (_12947_, _12747_);
  nor (_12948_, _12924_, _12947_);
  nor (_12949_, _12948_, _12946_);
  nand (_12950_, _12949_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_12951_, _12924_, _10367_);
  not (_12952_, _12730_);
  nor (_12953_, _12924_, _12952_);
  nor (_12954_, _12953_, _12951_);
  nor (_12955_, _12954_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_12956_, _12954_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_12957_, _12924_, _10144_);
  not (_12958_, _12713_);
  nor (_12959_, _12924_, _12958_);
  nor (_12960_, _12959_, _12957_);
  and (_12961_, _12960_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nand (_12962_, _12924_, _10479_);
  not (_12963_, _12696_);
  or (_12964_, _12924_, _12963_);
  nand (_12965_, _12964_, _12962_);
  or (_12966_, _12965_, _07119_);
  and (_12967_, _12924_, _10319_);
  not (_12968_, _12679_);
  nor (_12969_, _12924_, _12968_);
  nor (_12970_, _12969_, _12967_);
  and (_12971_, _12970_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nand (_12972_, _12965_, _07119_);
  and (_12973_, _12972_, _12966_);
  and (_12974_, _12973_, _12971_);
  not (_12975_, _12974_);
  nand (_12976_, _12975_, _12966_);
  nor (_12977_, _12960_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nor (_12978_, _12977_, _12961_);
  and (_12979_, _12978_, _12976_);
  or (_12980_, _12979_, _12961_);
  nor (_12981_, _12980_, _12956_);
  nor (_12982_, _12981_, _12955_);
  or (_12983_, _12949_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_12984_, _12983_, _12950_);
  nand (_12985_, _12984_, _12982_);
  nand (_12986_, _12985_, _12950_);
  nor (_12987_, _12986_, _12945_);
  nor (_12988_, _12987_, _12944_);
  nand (_12989_, _12988_, _12939_);
  and (_12990_, _12989_, _12937_);
  nor (_12991_, _12990_, _12931_);
  or (_12992_, _12991_, _12930_);
  and (_12993_, \oc8051_top_1.oc8051_memory_interface1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_12994_, _12993_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_12995_, _12994_, _12992_);
  and (_12996_, _12995_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_12997_, _12996_, _12929_);
  and (_12998_, _12997_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_12999_, _12992_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_13000_, _12999_, _07121_);
  and (_13001_, _13000_, _07140_);
  and (_13002_, _12928_, _07021_);
  nand (_13003_, _13002_, _13001_);
  nor (_13004_, _13003_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  or (_13005_, _13004_, _12998_);
  nor (_13006_, _12928_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_13007_, _12928_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_13008_, _13007_, _13006_);
  nand (_13009_, _13008_, _13005_);
  nor (_13010_, _12928_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_13011_, _12928_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  or (_13012_, _13011_, _13010_);
  or (_13013_, _13012_, _13009_);
  or (_13014_, _13013_, _07092_);
  nand (_13015_, _13013_, _07092_);
  nor (_13016_, _12466_, _08852_);
  and (_13017_, _13016_, _12872_);
  and (_13018_, _12857_, _12835_);
  and (_13019_, _13018_, _13017_);
  nor (_13020_, _13019_, _10204_);
  nor (_13021_, _13020_, _12921_);
  and (_13022_, _08888_, _08848_);
  nor (_13023_, _13022_, _12876_);
  not (_13024_, _13023_);
  and (_13025_, _13024_, _12924_);
  nor (_13026_, _13025_, _13021_);
  and (_13027_, _13026_, _13015_);
  and (_13028_, _13027_, _13014_);
  and (_13029_, _08855_, _08002_);
  and (_13030_, _13022_, _09129_);
  not (_13031_, _13020_);
  and (_13032_, _13023_, _12924_);
  and (_13033_, _13032_, _13031_);
  and (_13034_, _13033_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_13035_, _12920_, _10266_);
  or (_13036_, _13035_, _13034_);
  and (_13037_, \oc8051_top_1.oc8051_memory_interface1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_13038_, _13037_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_13039_, \oc8051_top_1.oc8051_memory_interface1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_13040_, \oc8051_top_1.oc8051_memory_interface1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_13041_, _13040_, _13039_);
  and (_13042_, _13041_, _13038_);
  and (_13043_, _13042_, _12994_);
  and (_13044_, _13043_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_13045_, _13044_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_13046_, _13045_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nand (_13047_, _13046_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand (_13048_, _13047_, _07092_);
  or (_13049_, _13047_, _07092_);
  and (_13050_, _13049_, _13048_);
  and (_13051_, _13025_, _13031_);
  and (_13052_, _13051_, _13050_);
  or (_13053_, _13052_, _13036_);
  nor (_13054_, _13053_, _13030_);
  nand (_13055_, _13054_, _12890_);
  or (_13056_, _13055_, _13029_);
  or (_13057_, _13056_, _13028_);
  and (_13938_[15], _13057_, _12916_);
  and (_13058_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _13707_);
  and (_13059_, _13058_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  not (_13060_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_13061_, _08527_, _13060_);
  not (_13062_, _13061_);
  not (_13063_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  not (_13064_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  not (_13065_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  not (_13066_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  not (_13067_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  not (_13068_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  not (_13069_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  not (_13070_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  not (_13071_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  not (_13072_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_13073_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4], \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_13074_, _13073_, _13072_);
  and (_13075_, _13074_, _13071_);
  and (_13076_, _13075_, _13070_);
  and (_13077_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_13078_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_13079_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_13080_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  nor (_13081_, _13080_, _13078_);
  and (_13082_, _13081_, _13079_);
  nor (_13083_, _13082_, _13078_);
  nor (_13084_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_13085_, _13084_, _13077_);
  not (_13086_, _13085_);
  nor (_13087_, _13086_, _13083_);
  nor (_13088_, _13087_, _13077_);
  and (_13089_, _13088_, _13076_);
  and (_13090_, _13089_, _13069_);
  and (_13091_, _13090_, _13068_);
  and (_13092_, _13091_, _13067_);
  and (_13093_, _13092_, _13066_);
  and (_13094_, _13093_, _13065_);
  and (_13095_, _13094_, _13064_);
  and (_13096_, _13095_, _13063_);
  nor (_13097_, _13096_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_13098_, _13096_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nor (_13099_, _13098_, _13097_);
  nor (_13100_, _13095_, _13063_);
  nor (_13101_, _13100_, _13096_);
  not (_13102_, _13101_);
  nor (_13103_, _13094_, _13064_);
  or (_13104_, _13103_, _13095_);
  nor (_13105_, _13093_, _13065_);
  nor (_13106_, _13105_, _13094_);
  not (_13107_, _13106_);
  nor (_13108_, _13092_, _13066_);
  nor (_13109_, _13108_, _13093_);
  not (_13110_, _13109_);
  nor (_13111_, _13091_, _13067_);
  nor (_13112_, _13111_, _13092_);
  not (_13113_, _13112_);
  nor (_13114_, _13090_, _13068_);
  or (_13115_, _13114_, _13091_);
  and (_13116_, _13088_, _13075_);
  nor (_13117_, _13116_, _13070_);
  nor (_13118_, _13117_, _13089_);
  not (_13119_, _13118_);
  and (_13120_, _13088_, _13074_);
  nor (_13121_, _13120_, _13071_);
  nor (_13122_, _13121_, _13116_);
  not (_13123_, _13122_);
  and (_13124_, _13088_, _13073_);
  nor (_13125_, _13124_, _13072_);
  nor (_13126_, _13125_, _13120_);
  not (_13127_, _13126_);
  not (_13128_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_13129_, _13088_, _13128_);
  nor (_13130_, _13088_, _13128_);
  nor (_13131_, _13130_, _13129_);
  not (_13132_, _13131_);
  not (_13133_, _12145_);
  and (_13134_, _12210_, _13133_);
  nor (_13135_, _13134_, _12207_);
  not (_13136_, _13135_);
  and (_13137_, _12179_, _12137_);
  not (_13138_, _13137_);
  not (_13139_, _12204_);
  nor (_13140_, _12200_, _12164_);
  nor (_13141_, _13140_, _13139_);
  not (_13142_, _12137_);
  and (_13143_, _08741_, _08665_);
  and (_13144_, _13143_, _12132_);
  nor (_13145_, _13144_, _12198_);
  nor (_13146_, _13145_, _13142_);
  nor (_13147_, _13146_, _13141_);
  and (_13148_, _13147_, _13138_);
  and (_13149_, _13148_, _12187_);
  and (_13150_, _13149_, _13136_);
  and (_13151_, _13143_, _12141_);
  and (_13152_, _13151_, _12170_);
  nor (_13153_, _13152_, _12193_);
  and (_13154_, _12163_, _12132_);
  or (_13155_, _13144_, _13154_);
  nor (_13156_, _13155_, _13151_);
  nor (_13157_, _13156_, _13153_);
  not (_13158_, _12193_);
  and (_13159_, _12155_, _12149_);
  nor (_13160_, _13159_, _12171_);
  nor (_13161_, _12203_, _12198_);
  and (_13162_, _13161_, _13160_);
  nor (_13163_, _13162_, _13158_);
  nor (_13164_, _13163_, _13157_);
  and (_13165_, _12200_, _12138_);
  not (_13166_, _13154_);
  nor (_13167_, _12198_, _12188_);
  and (_13168_, _13167_, _13166_);
  nor (_13169_, _13168_, _08590_);
  nor (_13170_, _13169_, _13165_);
  and (_13171_, _13170_, _13164_);
  nor (_13172_, _13167_, _13139_);
  not (_13173_, _13172_);
  and (_13174_, _12141_, _12154_);
  and (_13175_, _12209_, _13174_);
  not (_13176_, _13175_);
  and (_13177_, _12133_, _08614_);
  and (_13178_, _13177_, _12132_);
  and (_13179_, _13178_, _12134_);
  nor (_13180_, _13179_, _12161_);
  and (_13181_, _13180_, _13176_);
  and (_13182_, _13181_, _13173_);
  and (_13183_, _12191_, _12177_);
  and (_13184_, _12193_, _12188_);
  nor (_13185_, _13184_, _13183_);
  and (_13186_, _13185_, _13182_);
  not (_13187_, _12194_);
  nor (_13188_, _12204_, _12193_);
  nor (_13189_, _13188_, _13187_);
  nor (_13190_, _13189_, _12146_);
  and (_13191_, _13190_, _13186_);
  and (_13192_, _13191_, _13171_);
  nor (_13193_, _12205_, _12153_);
  nand (_13194_, _12172_, _12135_);
  and (_13195_, _12171_, _12137_);
  and (_13196_, _12191_, _13151_);
  nor (_13197_, _13196_, _13195_);
  and (_13198_, _13197_, _13194_);
  and (_13199_, _13198_, _13193_);
  nor (_13200_, _12177_, _12167_);
  nor (_13201_, _13159_, _13144_);
  and (_13202_, _13201_, _13200_);
  nor (_13203_, _13202_, _13139_);
  nor (_13204_, _12162_, _12170_);
  and (_13205_, _12177_, _08638_);
  nor (_13206_, _13205_, _12183_);
  nor (_13207_, _13206_, _13204_);
  nor (_13208_, _13207_, _13203_);
  and (_13209_, _13144_, _12144_);
  not (_13210_, _12144_);
  nor (_13211_, _12160_, _12188_);
  and (_13212_, _13211_, _13166_);
  nor (_13213_, _13212_, _13210_);
  nor (_13214_, _13213_, _13209_);
  and (_13215_, _13214_, _13208_);
  and (_13216_, _13215_, _13199_);
  and (_13217_, _13216_, _13192_);
  and (_13218_, _13217_, _13150_);
  nor (_13219_, _13081_, _13079_);
  nor (_13220_, _13219_, _13082_);
  not (_13221_, _13220_);
  nor (_13222_, _13221_, _13218_);
  not (_13223_, _13222_);
  and (_13224_, _12141_, _12133_);
  and (_13225_, _13224_, _12191_);
  or (_13226_, _13172_, _12195_);
  or (_13227_, _13226_, _13225_);
  or (_13228_, _12211_, _12180_);
  or (_13229_, _13228_, _13209_);
  nor (_13230_, _13229_, _13227_);
  nand (_13231_, _13230_, _13199_);
  nor (_13232_, _13231_, _13218_);
  not (_13233_, _13232_);
  nor (_13234_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_13235_, _13234_, _13079_);
  and (_13236_, _13235_, _13233_);
  and (_13237_, _13221_, _13218_);
  nor (_13238_, _13237_, _13222_);
  nand (_13239_, _13238_, _13236_);
  and (_13240_, _13239_, _13223_);
  not (_13241_, _13240_);
  and (_13242_, _13086_, _13083_);
  nor (_13243_, _13242_, _13087_);
  and (_13244_, _13243_, _13241_);
  and (_13245_, _13244_, _13132_);
  not (_13246_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_13247_, _13129_, _13246_);
  or (_13248_, _13247_, _13124_);
  and (_13249_, _13248_, _13245_);
  and (_13250_, _13249_, _13127_);
  and (_13251_, _13250_, _13123_);
  and (_13252_, _13251_, _13119_);
  nor (_13253_, _13089_, _13069_);
  or (_13254_, _13253_, _13090_);
  and (_13255_, _13254_, _13252_);
  and (_13256_, _13255_, _13115_);
  and (_13257_, _13256_, _13113_);
  and (_13258_, _13257_, _13110_);
  and (_13259_, _13258_, _13107_);
  and (_13260_, _13259_, _13104_);
  and (_13261_, _13260_, _13102_);
  or (_13262_, _13261_, _13099_);
  nand (_13263_, _13261_, _13099_);
  and (_13264_, _13263_, _13262_);
  or (_13265_, _13264_, _13062_);
  or (_13266_, _13061_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor (_13267_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , rst);
  and (_13268_, _13267_, _13266_);
  and (_13269_, _13268_, _13265_);
  or (_13939_[15], _13269_, _13059_);
  nor (_13270_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , rst);
  and (_13940_, _13270_, \oc8051_top_1.oc8051_memory_interface1.int_ack_buff );
  and (_13941_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , _13707_);
  and (_13271_, \oc8051_top_1.oc8051_rom1.ea_int , _08524_);
  nand (_13272_, _13271_, _08527_);
  and (_13942_, _13272_, _13941_);
  and (_13943_[7], \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _13707_);
  nor (_13273_, _12897_, _10128_);
  nor (_13274_, _13218_, _08535_);
  not (_13275_, _13274_);
  nor (_13276_, _13232_, _08539_);
  and (_13277_, _13218_, _08535_);
  nor (_13278_, _13277_, _13274_);
  nand (_13279_, _13278_, _13276_);
  and (_13280_, _13279_, _13275_);
  nor (_13281_, _13280_, _10128_);
  and (_13282_, _13281_, _08534_);
  nor (_13283_, _13281_, _08534_);
  nor (_13284_, _13283_, _13282_);
  nor (_13285_, _13284_, _13273_);
  and (_13286_, _08536_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_13287_, _13286_, _13273_);
  and (_13288_, _13287_, _13231_);
  or (_13289_, _13288_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_13290_, _13289_, _13285_);
  and (_13944_[2], _13290_, _13707_);
  and (_13291_, _08708_, _08608_);
  not (_13292_, _08659_);
  and (_13293_, _08683_, _13292_);
  and (_13294_, _13293_, _13291_);
  not (_13295_, _08634_);
  and (_13296_, _08737_, _13295_);
  and (_13297_, _08528_, _13707_);
  nand (_13298_, _13297_, _08561_);
  nor (_13299_, _13298_, _08586_);
  and (_13300_, _13299_, _13296_);
  and (_13947_, _13300_, _13294_);
  not (_13301_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  and (_13302_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [7]);
  or (_13303_, _13302_, _13301_);
  or (_13304_, \oc8051_top_1.oc8051_memory_interface1.cdata [7], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  and (_13305_, _13304_, _13707_);
  and (_13948_[7], _13305_, _13303_);
  and (_13949_, \oc8051_top_1.oc8051_memory_interface1.istb_t , _13707_);
  not (_13306_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and (_13307_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_13308_, _13307_, _13306_);
  and (_13309_, _13307_, _13306_);
  nor (_13310_, _13309_, _13308_);
  not (_13311_, _13310_);
  and (_13312_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and (_13313_, _13312_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_13314_, _13312_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_13315_, _13314_, _13313_);
  or (_13316_, _13315_, _13307_);
  and (_13317_, _13316_, _13311_);
  nor (_13318_, _13308_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and (_13319_, _13308_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  or (_13320_, _13319_, _13318_);
  or (_13321_, _13313_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  and (_13951_[3], _13321_, _13707_);
  and (_13322_, _13951_[3], _13320_);
  and (_13950_, _13322_, _13317_);
  not (_13323_, \oc8051_top_1.oc8051_rom1.ea_int );
  nor (_13324_, _12897_, _13323_);
  and (_13325_, _13324_, \oc8051_top_1.oc8051_rom1.data_o [31]);
  not (_13326_, _13324_);
  and (_13327_, _13326_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  or (_13328_, _13327_, _13325_);
  and (_13952_[31], _13328_, _13707_);
  and (_13329_, _13324_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and (_13330_, _13326_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  or (_13331_, _13330_, _13329_);
  and (_13953_[31], _13331_, _13707_);
  not (_13332_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  nor (_13333_, \oc8051_top_1.oc8051_decoder1.mem_act [2], \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  nor (_13334_, _13333_, _13332_);
  and (_13335_, \oc8051_top_1.oc8051_decoder1.mem_act [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_13336_, _13335_, _13333_);
  or (_13337_, _13336_, _13334_);
  and (_13954_[7], _13337_, _13707_);
  and (_13338_, \oc8051_top_1.oc8051_decoder1.mem_act [2], \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  not (_13339_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_13340_, \oc8051_top_1.oc8051_decoder1.mem_act [0], _13339_);
  or (_13341_, _13340_, _13338_);
  and (_13955_, _13341_, _12892_);
  and (_13956_, _13333_, _13707_);
  not (_13342_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  nor (_13343_, _13333_, _13342_);
  not (_13344_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  and (_13345_, _13344_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  and (_13346_, _13345_, _13333_);
  or (_13347_, _13346_, _13343_);
  and (_13957_[15], _13347_, _13707_);
  or (_13348_, _13339_, \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and (_13958_, _13348_, _12892_);
  nor (_13349_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  and (_13350_, _13349_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_13351_, \oc8051_top_1.oc8051_memory_interface1.istb_t , \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or (_13352_, _13351_, _13350_);
  and (_13959_, _13352_, _13707_);
  and (_13353_, _13323_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or (_13354_, _13353_, _13350_);
  and (_13960_, _13354_, _13707_);
  not (_13355_, _13350_);
  or (_13356_, _13355_, _09129_);
  or (_13357_, _13350_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [15]);
  and (_13358_, _13357_, _13707_);
  and (_13961_[15], _13358_, _13356_);
  or (_13359_, _12782_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nand (_13360_, _12782_, _07171_);
  and (_13361_, _13360_, _13707_);
  and (_13927_[0], _13361_, _13359_);
  or (_13362_, _12782_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nand (_13363_, _12782_, _07119_);
  and (_13364_, _13363_, _13707_);
  and (_13927_[1], _13364_, _13362_);
  or (_13365_, _12782_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nand (_13366_, _12782_, _07138_);
  and (_13367_, _13366_, _13707_);
  and (_13927_[2], _13367_, _13365_);
  or (_13368_, _12782_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nand (_13369_, _12782_, _07019_);
  and (_13370_, _13369_, _13707_);
  and (_13927_[3], _13370_, _13368_);
  or (_13371_, _12782_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  nand (_13372_, _12782_, _06859_);
  and (_13373_, _13372_, _13707_);
  and (_13927_[4], _13373_, _13371_);
  or (_13374_, _12782_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nand (_13375_, _12782_, _07038_);
  and (_13376_, _13375_, _13707_);
  and (_13927_[5], _13376_, _13374_);
  or (_13377_, _12782_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  nand (_13378_, _12782_, _07060_);
  and (_13379_, _13378_, _13707_);
  and (_13927_[6], _13379_, _13377_);
  or (_13380_, _12782_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  nand (_13381_, _12782_, _07094_);
  and (_13382_, _13381_, _13707_);
  and (_13927_[7], _13382_, _13380_);
  or (_13383_, _12782_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nand (_13384_, _12782_, _07173_);
  and (_13385_, _13384_, _13707_);
  and (_13927_[8], _13385_, _13383_);
  or (_13386_, _12782_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nand (_13387_, _12782_, _07121_);
  and (_13388_, _13387_, _13707_);
  and (_13927_[9], _13388_, _13386_);
  or (_13389_, _12782_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nand (_13390_, _12782_, _07140_);
  and (_13391_, _13390_, _13707_);
  and (_13927_[10], _13391_, _13389_);
  or (_13392_, _12782_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nand (_13393_, _12782_, _07021_);
  and (_13394_, _13393_, _13707_);
  and (_13927_[11], _13394_, _13392_);
  or (_13395_, _12782_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nand (_13396_, _12782_, _06865_);
  and (_13397_, _13396_, _13707_);
  and (_13927_[12], _13397_, _13395_);
  or (_13398_, _12782_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nand (_13399_, _12782_, _07040_);
  and (_13400_, _13399_, _13707_);
  and (_13927_[13], _13400_, _13398_);
  or (_13401_, _12782_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nand (_13402_, _12782_, _07062_);
  and (_13403_, _13402_, _13707_);
  and (_13927_[14], _13403_, _13401_);
  or (_13404_, _12786_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_13405_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _13707_);
  or (_13406_, _13405_, _00002_);
  and (_13928_[0], _13406_, _13404_);
  or (_13407_, _12786_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_13408_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _13707_);
  or (_13409_, _13408_, _00002_);
  and (_13928_[1], _13409_, _13407_);
  or (_13410_, _12786_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_13411_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _13707_);
  or (_13412_, _13411_, _00002_);
  and (_13928_[2], _13412_, _13410_);
  or (_13413_, _12786_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_13414_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _13707_);
  or (_13415_, _13414_, _00002_);
  and (_13928_[3], _13415_, _13413_);
  or (_13416_, _12786_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  and (_13417_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _13707_);
  or (_13418_, _13417_, _00002_);
  and (_13928_[4], _13418_, _13416_);
  or (_13419_, _12786_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  and (_13420_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _13707_);
  or (_13421_, _13420_, _00002_);
  and (_13928_[5], _13421_, _13419_);
  or (_13422_, _12786_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  and (_13423_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _13707_);
  or (_13424_, _13423_, _00002_);
  and (_13928_[6], _13424_, _13422_);
  or (_13425_, _12786_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  and (_13426_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _13707_);
  or (_13427_, _13426_, _00002_);
  and (_13928_[7], _13427_, _13425_);
  or (_13428_, _12786_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  and (_13429_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _13707_);
  or (_13430_, _13429_, _00002_);
  and (_13928_[8], _13430_, _13428_);
  or (_13431_, _12786_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and (_13432_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _13707_);
  or (_13433_, _13432_, _00002_);
  and (_13928_[9], _13433_, _13431_);
  or (_13434_, _12786_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  and (_13435_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _13707_);
  or (_13436_, _13435_, _00002_);
  and (_13928_[10], _13436_, _13434_);
  or (_13437_, _12786_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and (_13438_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _13707_);
  or (_13439_, _13438_, _00002_);
  and (_13928_[11], _13439_, _13437_);
  or (_13440_, _12786_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  and (_13441_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _13707_);
  or (_13442_, _13441_, _00002_);
  and (_13928_[12], _13442_, _13440_);
  or (_13443_, _12786_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and (_13444_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _13707_);
  or (_13445_, _13444_, _00002_);
  and (_13928_[13], _13445_, _13443_);
  or (_13446_, _12786_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  and (_13447_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _13707_);
  or (_13448_, _13447_, _00002_);
  and (_13928_[14], _13448_, _13446_);
  and (_13449_, _13326_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_13450_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [0]);
  and (_13451_, _13450_, _13324_);
  or (_13452_, _13451_, _13449_);
  and (_13952_[0], _13452_, _13707_);
  and (_13453_, _13326_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_13454_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [1]);
  and (_13455_, _13454_, _13324_);
  or (_13456_, _13455_, _13453_);
  and (_13952_[1], _13456_, _13707_);
  and (_13457_, _13326_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_13458_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [2]);
  and (_13459_, _13458_, _13324_);
  or (_13460_, _13459_, _13457_);
  and (_13952_[2], _13460_, _13707_);
  and (_13461_, _13326_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_13462_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [3]);
  and (_13463_, _13462_, _13324_);
  or (_13464_, _13463_, _13461_);
  and (_13952_[3], _13464_, _13707_);
  and (_13465_, _13326_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_13466_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [4]);
  and (_13467_, _13466_, _13324_);
  or (_13468_, _13467_, _13465_);
  and (_13952_[4], _13468_, _13707_);
  and (_13469_, _13326_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_13470_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [5]);
  and (_13471_, _13470_, _13324_);
  or (_13472_, _13471_, _13469_);
  and (_13952_[5], _13472_, _13707_);
  and (_13473_, _13324_, \oc8051_top_1.oc8051_rom1.data_o [6]);
  and (_13474_, _13326_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  or (_13475_, _13474_, _13473_);
  and (_13952_[6], _13475_, _13707_);
  and (_13476_, _13326_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_13477_, _13324_, _13302_);
  or (_13478_, _13477_, _13476_);
  and (_13952_[7], _13478_, _13707_);
  and (_13479_, _13324_, \oc8051_top_1.oc8051_rom1.data_o [8]);
  and (_13480_, _13326_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  or (_13481_, _13480_, _13479_);
  and (_13952_[8], _13481_, _13707_);
  and (_13482_, _13324_, \oc8051_top_1.oc8051_rom1.data_o [9]);
  and (_13483_, _13326_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  or (_13484_, _13483_, _13482_);
  and (_13952_[9], _13484_, _13707_);
  and (_13485_, _13324_, \oc8051_top_1.oc8051_rom1.data_o [10]);
  and (_13486_, _13326_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  or (_13487_, _13486_, _13485_);
  and (_13952_[10], _13487_, _13707_);
  and (_13488_, _13324_, \oc8051_top_1.oc8051_rom1.data_o [11]);
  and (_13489_, _13326_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  or (_13490_, _13489_, _13488_);
  and (_13952_[11], _13490_, _13707_);
  and (_13491_, _13324_, \oc8051_top_1.oc8051_rom1.data_o [12]);
  and (_13492_, _13326_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  or (_13493_, _13492_, _13491_);
  and (_13952_[12], _13493_, _13707_);
  and (_13494_, _13324_, \oc8051_top_1.oc8051_rom1.data_o [13]);
  and (_13495_, _13326_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  or (_13496_, _13495_, _13494_);
  and (_13952_[13], _13496_, _13707_);
  and (_13497_, _13324_, \oc8051_top_1.oc8051_rom1.data_o [14]);
  and (_13498_, _13326_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  or (_13499_, _13498_, _13497_);
  and (_13952_[14], _13499_, _13707_);
  and (_13500_, _13324_, \oc8051_top_1.oc8051_rom1.data_o [15]);
  and (_13501_, _13326_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  or (_13502_, _13501_, _13500_);
  and (_13952_[15], _13502_, _13707_);
  and (_13503_, _13324_, \oc8051_top_1.oc8051_rom1.data_o [16]);
  and (_13504_, _13326_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  or (_13505_, _13504_, _13503_);
  and (_13952_[16], _13505_, _13707_);
  and (_13506_, _13324_, \oc8051_top_1.oc8051_rom1.data_o [17]);
  and (_13507_, _13326_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  or (_13508_, _13507_, _13506_);
  and (_13952_[17], _13508_, _13707_);
  and (_13509_, _13324_, \oc8051_top_1.oc8051_rom1.data_o [18]);
  and (_13510_, _13326_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  or (_13511_, _13510_, _13509_);
  and (_13952_[18], _13511_, _13707_);
  and (_13512_, _13324_, \oc8051_top_1.oc8051_rom1.data_o [19]);
  and (_13513_, _13326_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  or (_13514_, _13513_, _13512_);
  and (_13952_[19], _13514_, _13707_);
  and (_13515_, _13324_, \oc8051_top_1.oc8051_rom1.data_o [20]);
  and (_13516_, _13326_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  or (_13517_, _13516_, _13515_);
  and (_13952_[20], _13517_, _13707_);
  and (_13518_, _13324_, \oc8051_top_1.oc8051_rom1.data_o [21]);
  and (_13519_, _13326_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  or (_13520_, _13519_, _13518_);
  and (_13952_[21], _13520_, _13707_);
  and (_13521_, _13324_, \oc8051_top_1.oc8051_rom1.data_o [22]);
  and (_13522_, _13326_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  or (_13523_, _13522_, _13521_);
  and (_13952_[22], _13523_, _13707_);
  and (_13524_, _13324_, \oc8051_top_1.oc8051_rom1.data_o [23]);
  and (_13525_, _13326_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  or (_13526_, _13525_, _13524_);
  and (_13952_[23], _13526_, _13707_);
  and (_13527_, _13324_, \oc8051_top_1.oc8051_rom1.data_o [24]);
  and (_13528_, _13326_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  or (_13529_, _13528_, _13527_);
  and (_13952_[24], _13529_, _13707_);
  and (_13530_, _13324_, \oc8051_top_1.oc8051_rom1.data_o [25]);
  and (_13531_, _13326_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  or (_13532_, _13531_, _13530_);
  and (_13952_[25], _13532_, _13707_);
  and (_13533_, _13324_, \oc8051_top_1.oc8051_rom1.data_o [26]);
  and (_13534_, _13326_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  or (_13535_, _13534_, _13533_);
  and (_13952_[26], _13535_, _13707_);
  and (_13536_, _13324_, \oc8051_top_1.oc8051_rom1.data_o [27]);
  and (_13537_, _13326_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  or (_13538_, _13537_, _13536_);
  and (_13952_[27], _13538_, _13707_);
  and (_13539_, _13324_, \oc8051_top_1.oc8051_rom1.data_o [28]);
  and (_13540_, _13326_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  or (_13541_, _13540_, _13539_);
  and (_13952_[28], _13541_, _13707_);
  and (_13542_, _13324_, \oc8051_top_1.oc8051_rom1.data_o [29]);
  and (_13543_, _13326_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  or (_13544_, _13543_, _13542_);
  and (_13952_[29], _13544_, _13707_);
  and (_13545_, _13324_, \oc8051_top_1.oc8051_rom1.data_o [30]);
  and (_13546_, _13326_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  or (_13547_, _13546_, _13545_);
  and (_13952_[30], _13547_, _13707_);
  nor (_13931_[0], _08643_, rst);
  nor (_13931_[1], _08619_, rst);
  and (_13931_[2], _08571_, _13707_);
  nor (_13931_[3], _10047_, rst);
  and (_13932_[0], _10299_, _13707_);
  and (_13932_[1], _10457_, _13707_);
  and (_13932_[2], _10114_, _13707_);
  and (_13932_[3], _10346_, _13707_);
  and (_13932_[4], _10509_, _13707_);
  and (_13932_[5], _10173_, _13707_);
  and (_13932_[6], _10406_, _13707_);
  and (_13548_, _12892_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [0]);
  and (_13549_, _13930_, xram_data_in_reg[0]);
  or (_13937_[0], _13549_, _13548_);
  and (_13550_, _12892_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [1]);
  and (_13551_, _13930_, xram_data_in_reg[1]);
  or (_13937_[1], _13551_, _13550_);
  and (_13552_, _12892_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [2]);
  and (_13553_, _13930_, xram_data_in_reg[2]);
  or (_13937_[2], _13553_, _13552_);
  and (_13554_, _12892_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [3]);
  and (_13555_, _13930_, xram_data_in_reg[3]);
  or (_13937_[3], _13555_, _13554_);
  and (_13556_, _12892_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [4]);
  and (_13557_, _13930_, xram_data_in_reg[4]);
  or (_13937_[4], _13557_, _13556_);
  and (_13558_, _12892_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [5]);
  and (_13559_, _13930_, xram_data_in_reg[5]);
  or (_13937_[5], _13559_, _13558_);
  and (_13560_, _12892_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [6]);
  and (_13561_, _13930_, xram_data_in_reg[6]);
  or (_13937_[6], _13561_, _13560_);
  or (_13562_, _12890_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and (_13563_, _13562_, _13707_);
  or (_13564_, _13033_, _13022_);
  and (_13565_, _13564_, _08106_);
  or (_13566_, _12970_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  not (_13567_, _12971_);
  and (_13568_, _13026_, _13567_);
  and (_13569_, _13568_, _13566_);
  and (_13570_, _12920_, _12968_);
  and (_13571_, _08855_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and (_13572_, _13051_, _10320_);
  or (_13573_, _13572_, _13571_);
  or (_13574_, _13573_, _13570_);
  nor (_13575_, _13574_, _13569_);
  nand (_13576_, _13575_, _12890_);
  or (_13577_, _13576_, _13565_);
  and (_13938_[0], _13577_, _13563_);
  or (_13578_, _12890_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  and (_13579_, _13578_, _13707_);
  and (_13580_, _13564_, _08166_);
  or (_13581_, _12973_, _12971_);
  and (_13582_, _13026_, _12975_);
  and (_13583_, _13582_, _13581_);
  and (_13584_, _12920_, _12963_);
  and (_13585_, _08855_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  and (_13586_, _13051_, _10480_);
  or (_13587_, _13586_, _13585_);
  or (_13588_, _13587_, _13584_);
  nor (_13589_, _13588_, _13583_);
  nand (_13590_, _13589_, _12890_);
  or (_13591_, _13590_, _13580_);
  and (_13938_[1], _13591_, _13579_);
  not (_13592_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_13593_, _12897_, _13592_);
  and (_13594_, _12897_, _13592_);
  nor (_13595_, _13594_, _13593_);
  or (_13596_, _13595_, _12890_);
  and (_13597_, _13596_, _13707_);
  and (_13598_, _13564_, _08224_);
  or (_13599_, _12978_, _12976_);
  not (_13600_, _12979_);
  and (_13601_, _13026_, _13600_);
  and (_13602_, _13601_, _13599_);
  and (_13603_, _12920_, _12958_);
  and (_13604_, _08855_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and (_13605_, _13051_, _10145_);
  or (_13606_, _13605_, _13604_);
  or (_13607_, _13606_, _13603_);
  nor (_13608_, _13607_, _13602_);
  nand (_13609_, _13608_, _12890_);
  or (_13610_, _13609_, _13598_);
  and (_13938_[2], _13610_, _13597_);
  and (_13611_, _13593_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_13612_, _13593_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_13613_, _13612_, _13611_);
  or (_13614_, _13613_, _12890_);
  and (_13615_, _13614_, _13707_);
  and (_13616_, _13564_, _08288_);
  not (_13617_, _12980_);
  or (_13618_, _12955_, _12956_);
  nand (_13619_, _13618_, _13617_);
  or (_13620_, _13618_, _13617_);
  and (_13621_, _13620_, _13026_);
  and (_13622_, _13621_, _13619_);
  and (_13623_, _12920_, _12952_);
  and (_13624_, _08855_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_13625_, _13051_, _10368_);
  or (_13626_, _13625_, _13624_);
  or (_13627_, _13626_, _13623_);
  nor (_13628_, _13627_, _13622_);
  nand (_13629_, _13628_, _12890_);
  or (_13630_, _13629_, _13616_);
  and (_13938_[3], _13630_, _13615_);
  and (_13631_, _12900_, _12898_);
  nor (_13632_, _13611_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_13633_, _13632_, _13631_);
  or (_13634_, _13633_, _12890_);
  and (_13635_, _13634_, _13707_);
  and (_13636_, _13564_, _08354_);
  or (_13637_, _12984_, _12982_);
  and (_13638_, _13026_, _12985_);
  and (_13639_, _13638_, _13637_);
  and (_13640_, _13051_, _10527_);
  and (_13641_, _12920_, _12947_);
  and (_13642_, _08855_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or (_13643_, _13642_, _13641_);
  or (_13644_, _13643_, _13640_);
  nor (_13645_, _13644_, _13639_);
  nand (_13646_, _13645_, _12890_);
  or (_13647_, _13646_, _13636_);
  and (_13938_[4], _13647_, _13635_);
  and (_13648_, _12901_, _12898_);
  not (_13649_, _13648_);
  or (_13650_, _13631_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and (_13651_, _13650_, _13649_);
  or (_13652_, _13651_, _12890_);
  and (_13653_, _13652_, _13707_);
  and (_13654_, _13564_, _08428_);
  or (_13655_, _12944_, _12945_);
  not (_13656_, _13655_);
  nand (_13657_, _13656_, _12986_);
  or (_13658_, _13656_, _12986_);
  and (_13659_, _13658_, _13026_);
  and (_13660_, _13659_, _13657_);
  and (_13661_, _12920_, _12941_);
  and (_13662_, _08855_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and (_13663_, _13051_, _10192_);
  or (_13664_, _13663_, _13662_);
  or (_13665_, _13664_, _13661_);
  nor (_13666_, _13665_, _13660_);
  nand (_13667_, _13666_, _12890_);
  or (_13668_, _13667_, _13654_);
  and (_13938_[5], _13668_, _13653_);
  nor (_13669_, _13648_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_13670_, _13648_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor (_13671_, _13670_, _13669_);
  or (_13672_, _13671_, _12890_);
  and (_13673_, _13672_, _13707_);
  and (_13674_, _13564_, _08500_);
  or (_13675_, _12988_, _12939_);
  and (_13676_, _13026_, _12989_);
  nand (_13677_, _13676_, _13675_);
  and (_13678_, _12920_, _12933_);
  and (_13679_, _08855_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_13680_, _13051_, _10424_);
  or (_13681_, _13680_, _13679_);
  nor (_13682_, _13681_, _13678_);
  and (_13683_, _13682_, _13677_);
  nand (_13684_, _13683_, _12890_);
  or (_13686_, _13684_, _13674_);
  and (_13938_[6], _13686_, _13673_);
  nor (_13689_, _13670_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and (_13691_, _13670_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  or (_13693_, _13691_, _13689_);
  nor (_13695_, _13693_, _12890_);
  and (_13697_, _13564_, _08002_);
  or (_13698_, _12930_, _12931_);
  nand (_13699_, _13698_, _12990_);
  or (_13700_, _13698_, _12990_);
  and (_13701_, _13700_, _13026_);
  and (_13702_, _13701_, _13699_);
  and (_13703_, _13051_, _10266_);
  and (_13705_, _12920_, _12926_);
  and (_13706_, _08855_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  or (_13708_, _13706_, _13705_);
  or (_13709_, _13708_, _13703_);
  or (_13710_, _13709_, _13702_);
  or (_13712_, _13710_, _13697_);
  and (_13713_, _13712_, _12890_);
  or (_13714_, _13713_, _13695_);
  and (_13938_[7], _13714_, _13707_);
  nand (_13716_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7], \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or (_13717_, _13716_, _13069_);
  nor (_13719_, _13717_, _13649_);
  nor (_13720_, _13691_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor (_13721_, _13720_, _13719_);
  or (_13723_, _13721_, _12890_);
  and (_13724_, _13723_, _13707_);
  and (_13725_, _12836_, _08507_);
  and (_13727_, _13725_, _08008_);
  and (_13728_, _13727_, _12809_);
  and (_13729_, _12822_, _07695_);
  and (_13731_, _13729_, _08004_);
  and (_13732_, _08853_, _08746_);
  and (_13733_, _12884_, _13732_);
  and (_13735_, _08804_, _08787_);
  and (_13736_, _13735_, _08848_);
  and (_13737_, _12880_, _13736_);
  or (_13738_, _13737_, _12879_);
  or (_13739_, _13738_, _13733_);
  or (_13740_, _13739_, _13731_);
  or (_13741_, _13740_, _13728_);
  and (_13742_, _08804_, _08523_);
  and (_13743_, _13742_, _08764_);
  nor (_13744_, _13020_, _13743_);
  not (_13745_, _13743_);
  and (_13746_, _08847_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and (_13747_, _13746_, _08771_);
  nor (_13748_, _12920_, _13747_);
  and (_13749_, _13748_, _12919_);
  and (_13750_, _13749_, _13745_);
  and (_13751_, _12871_, _08848_);
  nor (_13752_, _13751_, _12876_);
  not (_13753_, _13752_);
  and (_13754_, _13753_, _13750_);
  nor (_13755_, _13754_, _13744_);
  and (_13757_, _12992_, _07173_);
  nor (_13758_, _12992_, _07173_);
  nor (_13760_, _13758_, _13757_);
  or (_13761_, _13760_, _12929_);
  nand (_13762_, _13760_, _12929_);
  and (_13764_, _13762_, _13761_);
  and (_13765_, _13764_, _13755_);
  and (_13766_, _13747_, _08106_);
  and (_13768_, _13033_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_13769_, _12920_, _10320_);
  and (_13770_, _13051_, _12154_);
  or (_13772_, _13770_, _13769_);
  or (_13773_, _13772_, _13768_);
  and (_13774_, _13751_, _09165_);
  or (_13776_, _13774_, _13773_);
  or (_13777_, _13776_, _13766_);
  or (_13778_, _13777_, _13765_);
  or (_13780_, _13778_, _13741_);
  and (_13938_[8], _13780_, _13724_);
  or (_13781_, _13719_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  nand (_13783_, _13719_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and (_13784_, _13783_, _13781_);
  or (_13785_, _13784_, _12890_);
  and (_13787_, _13785_, _13707_);
  and (_13788_, _12992_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_13789_, _13788_, _12929_);
  and (_13790_, _12999_, _12928_);
  nor (_13791_, _13790_, _13789_);
  nand (_13792_, _13791_, _07121_);
  or (_13793_, _13791_, _07121_);
  and (_13794_, _13793_, _13026_);
  and (_13795_, _13794_, _13792_);
  and (_13796_, _08855_, _08166_);
  not (_13797_, _13022_);
  nor (_13798_, _13797_, _09198_);
  and (_13799_, _13033_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and (_13800_, _12920_, _10480_);
  and (_13801_, _13051_, _12140_);
  or (_13802_, _13801_, _13800_);
  or (_13803_, _13802_, _13799_);
  nor (_13804_, _13803_, _13798_);
  nand (_13805_, _13804_, _12890_);
  or (_13806_, _13805_, _13796_);
  or (_13807_, _13806_, _13795_);
  and (_13938_[9], _13807_, _13787_);
  and (_13809_, _12905_, _12898_);
  nor (_13811_, _13809_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_13812_, _13809_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor (_13813_, _13812_, _13811_);
  or (_13815_, _13813_, _12890_);
  and (_13816_, _13815_, _13707_);
  and (_13817_, _13000_, _12928_);
  and (_13819_, _13789_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor (_13820_, _13819_, _13817_);
  nand (_13821_, _13820_, _07140_);
  or (_13823_, _13820_, _07140_);
  and (_13824_, _13823_, _13026_);
  and (_00011_, _13824_, _13821_);
  and (_00013_, _08855_, _08224_);
  not (_00014_, _12890_);
  nor (_00015_, _13797_, _09228_);
  and (_00017_, _13033_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_00018_, _12920_, _10145_);
  and (_00019_, _13051_, _12131_);
  or (_00021_, _00019_, _00018_);
  or (_00022_, _00021_, _00017_);
  or (_00023_, _00022_, _00015_);
  or (_00025_, _00023_, _00014_);
  or (_00026_, _00025_, _00013_);
  or (_00027_, _00026_, _00011_);
  and (_13938_[10], _00027_, _13816_);
  nor (_00028_, _13812_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and (_00029_, _13812_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor (_00030_, _00029_, _00028_);
  or (_00031_, _00030_, _12890_);
  and (_00032_, _00031_, _13707_);
  and (_00033_, _12995_, _12929_);
  and (_00034_, _13001_, _12928_);
  nor (_00035_, _00034_, _00033_);
  nand (_00036_, _00035_, _07021_);
  or (_00037_, _00035_, _07021_);
  and (_00038_, _00037_, _13026_);
  and (_00039_, _00038_, _00036_);
  and (_00040_, _08855_, _08288_);
  nor (_00041_, _13797_, _09258_);
  and (_00042_, _12920_, _10368_);
  and (_00043_, _13033_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor (_00044_, _13043_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_00046_, _00044_, _13044_);
  and (_00047_, _00046_, _13051_);
  or (_00049_, _00047_, _00043_);
  or (_00050_, _00049_, _00042_);
  or (_00051_, _00050_, _00041_);
  or (_00053_, _00051_, _00014_);
  or (_00054_, _00053_, _00040_);
  or (_00055_, _00054_, _00039_);
  and (_13938_[11], _00055_, _00032_);
  or (_00057_, _00029_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nand (_00058_, _00029_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and (_00060_, _00058_, _00057_);
  or (_00061_, _00060_, _12890_);
  and (_00062_, _00061_, _13707_);
  not (_00064_, _12997_);
  and (_00065_, _13003_, _00064_);
  or (_00066_, _00065_, _06865_);
  nand (_00068_, _00065_, _06865_);
  and (_00069_, _00068_, _13026_);
  and (_00070_, _00069_, _00066_);
  and (_00072_, _08855_, _08354_);
  nor (_00073_, _13797_, _09290_);
  and (_00074_, _12920_, _10527_);
  and (_00076_, _13033_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor (_00077_, _13044_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_00078_, _00077_, _13045_);
  and (_00079_, _00078_, _13051_);
  or (_00080_, _00079_, _00076_);
  or (_00081_, _00080_, _00074_);
  nor (_00082_, _00081_, _00073_);
  nand (_00083_, _00082_, _12890_);
  or (_00084_, _00083_, _00072_);
  or (_00085_, _00084_, _00070_);
  and (_13938_[12], _00085_, _00062_);
  and (_00086_, _13005_, _07040_);
  nor (_00087_, _13005_, _07040_);
  or (_00088_, _00087_, _00086_);
  and (_00089_, _00088_, _13026_);
  and (_00090_, _08855_, _08428_);
  nor (_00091_, _13797_, _09324_);
  and (_00092_, _13033_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and (_00093_, _12920_, _10192_);
  or (_00094_, _00093_, _00092_);
  nor (_00095_, _13045_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_00097_, _00095_, _13046_);
  and (_00098_, _00097_, _13051_);
  or (_00100_, _00098_, _00094_);
  or (_00101_, _00100_, _00091_);
  or (_00102_, _00101_, _00090_);
  or (_00104_, _00102_, _00089_);
  or (_00105_, _00104_, _13741_);
  nor (_00106_, _12909_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or (_00108_, _00106_, _12910_);
  nand (_00109_, _00108_, _13741_);
  and (_00110_, _00109_, _13707_);
  and (_13938_[13], _00110_, _00105_);
  and (_00112_, _08855_, _08500_);
  nor (_00113_, _13797_, _09353_);
  and (_00115_, _12920_, _10424_);
  and (_00116_, _13033_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or (_00117_, _13046_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_00119_, _00117_, _13047_);
  and (_00120_, _00119_, _13051_);
  or (_00121_, _00120_, _00116_);
  or (_00123_, _00121_, _00115_);
  or (_00124_, _00123_, _00113_);
  or (_00125_, _00124_, _00112_);
  and (_00127_, _13009_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor (_00128_, _13009_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  or (_00129_, _00128_, _00127_);
  and (_00130_, _00129_, _13026_);
  or (_00131_, _00130_, _00125_);
  or (_00132_, _00131_, _13741_);
  nor (_00133_, _12910_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or (_00134_, _00133_, _12911_);
  nand (_00135_, _00134_, _13741_);
  and (_00136_, _00135_, _13707_);
  and (_13938_[14], _00136_, _00132_);
  and (_00137_, _13058_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nor (_00138_, _13235_, _13233_);
  nor (_00139_, _00138_, _13236_);
  or (_00140_, _00139_, _13062_);
  or (_00141_, _13061_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_00142_, _00141_, _13267_);
  and (_00143_, _00142_, _00140_);
  or (_13939_[0], _00143_, _00137_);
  and (_00144_, _13058_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or (_00145_, _13238_, _13236_);
  and (_00147_, _00145_, _13239_);
  or (_00148_, _00147_, _13062_);
  or (_00150_, _13061_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_00151_, _00150_, _13267_);
  and (_00152_, _00151_, _00148_);
  or (_13939_[1], _00152_, _00144_);
  and (_00154_, _13058_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_00155_, _13243_, _13241_);
  nor (_00157_, _00155_, _13244_);
  or (_00158_, _00157_, _13062_);
  or (_00159_, _13061_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_00161_, _00159_, _13267_);
  and (_00162_, _00161_, _00158_);
  or (_13939_[2], _00162_, _00154_);
  and (_00164_, _13058_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_00165_, _13244_, _13132_);
  nor (_00166_, _00165_, _13245_);
  or (_00168_, _00166_, _13062_);
  or (_00169_, _13061_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_00170_, _00169_, _13267_);
  and (_00172_, _00170_, _00168_);
  or (_13939_[3], _00172_, _00164_);
  nor (_00173_, _13248_, _13245_);
  nor (_00175_, _00173_, _13249_);
  or (_00176_, _00175_, _13062_);
  or (_00177_, _13061_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_00178_, _00177_, _13267_);
  and (_00179_, _00178_, _00176_);
  and (_00180_, _13058_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or (_13939_[4], _00180_, _00179_);
  or (_00181_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5], _08524_);
  and (_00182_, _00181_, _13707_);
  or (_00183_, _13249_, _13127_);
  nor (_00184_, _13250_, _13062_);
  and (_00185_, _00184_, _00183_);
  nor (_00186_, _13061_, _07038_);
  or (_00187_, _00186_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_00188_, _00187_, _00185_);
  and (_13939_[5], _00188_, _00182_);
  nor (_00189_, _13250_, _13123_);
  nor (_00190_, _00189_, _13251_);
  or (_00191_, _00190_, _13062_);
  or (_00192_, _13061_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_00193_, _00192_, _13267_);
  and (_00195_, _00193_, _00191_);
  and (_00196_, _13058_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or (_13939_[6], _00196_, _00195_);
  and (_00198_, _13058_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor (_00199_, _13251_, _13119_);
  nor (_00201_, _00199_, _13252_);
  or (_00202_, _00201_, _13062_);
  or (_00203_, _13061_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_00205_, _00203_, _13267_);
  and (_00206_, _00205_, _00202_);
  or (_13939_[7], _00206_, _00198_);
  and (_00208_, _13058_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor (_00209_, _13254_, _13252_);
  nor (_00210_, _00209_, _13255_);
  or (_00212_, _00210_, _13062_);
  or (_00213_, _13061_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_00214_, _00213_, _13267_);
  and (_00216_, _00214_, _00212_);
  or (_13939_[8], _00216_, _00208_);
  nor (_00217_, _13255_, _13115_);
  nor (_00219_, _00217_, _13256_);
  or (_00220_, _00219_, _13062_);
  or (_00221_, _13061_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_00223_, _00221_, _13267_);
  and (_00224_, _00223_, _00220_);
  and (_00225_, _13058_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  or (_13939_[9], _00225_, _00224_);
  nor (_00226_, _13256_, _13113_);
  nor (_00227_, _00226_, _13257_);
  or (_00228_, _00227_, _13062_);
  or (_00229_, _13061_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_00230_, _00229_, _13267_);
  and (_00231_, _00230_, _00228_);
  and (_00232_, _13058_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  or (_13939_[10], _00232_, _00231_);
  nor (_00233_, _13257_, _13110_);
  nor (_00234_, _00233_, _13258_);
  or (_00235_, _00234_, _13062_);
  or (_00236_, _13061_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_00237_, _00236_, _13267_);
  and (_00238_, _00237_, _00235_);
  and (_00239_, _13058_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  or (_13939_[11], _00239_, _00238_);
  nor (_00240_, _13258_, _13107_);
  nor (_00242_, _00240_, _13259_);
  or (_00243_, _00242_, _13062_);
  or (_00245_, _13061_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_00246_, _00245_, _13267_);
  and (_00247_, _00246_, _00243_);
  and (_00249_, _13058_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  or (_13939_[12], _00249_, _00247_);
  nor (_00250_, _13259_, _13104_);
  nor (_00252_, _00250_, _13260_);
  or (_00253_, _00252_, _13062_);
  or (_00254_, _13061_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_00256_, _00254_, _13267_);
  and (_00257_, _00256_, _00253_);
  and (_00258_, _13058_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or (_13939_[13], _00258_, _00257_);
  nor (_00260_, _13260_, _13102_);
  nor (_00261_, _00260_, _13261_);
  or (_00263_, _00261_, _13062_);
  or (_00264_, _13061_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_00265_, _00264_, _13267_);
  and (_00267_, _00265_, _00263_);
  and (_00268_, _13058_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or (_13939_[14], _00268_, _00267_);
  and (_13943_[0], \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], _13707_);
  and (_13943_[1], \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], _13707_);
  and (_13943_[2], \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _13707_);
  and (_13943_[3], \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], _13707_);
  and (_13943_[4], \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _13707_);
  and (_13943_[5], \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], _13707_);
  and (_13943_[6], \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _13707_);
  nor (_00270_, _13232_, _10128_);
  nand (_00271_, _00270_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  or (_00272_, _00270_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_00273_, _00272_, _13267_);
  and (_13944_[0], _00273_, _00271_);
  or (_00274_, _13278_, _13276_);
  and (_00275_, _00274_, _13279_);
  or (_00276_, _00275_, _10128_);
  or (_00277_, _08527_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_00278_, _00277_, _13267_);
  and (_13944_[1], _00278_, _00276_);
  or (_00279_, _13450_, _13301_);
  or (_00280_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  and (_00281_, _00280_, _13707_);
  and (_13948_[0], _00281_, _00279_);
  or (_00283_, _13454_, _13301_);
  or (_00285_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  and (_00286_, _00285_, _13707_);
  and (_13948_[1], _00286_, _00283_);
  or (_00288_, _13458_, _13301_);
  or (_00289_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  and (_00290_, _00289_, _13707_);
  and (_13948_[2], _00290_, _00288_);
  or (_00292_, _13462_, _13301_);
  or (_00293_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  and (_00295_, _00293_, _13707_);
  and (_13948_[3], _00295_, _00292_);
  or (_00296_, _13466_, _13301_);
  or (_00298_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  and (_00299_, _00298_, _13707_);
  and (_13948_[4], _00299_, _00296_);
  or (_00301_, _13470_, _13301_);
  or (_00302_, \oc8051_top_1.oc8051_memory_interface1.cdata [5], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  and (_00303_, _00302_, _13707_);
  and (_13948_[5], _00303_, _00301_);
  and (_00305_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [6]);
  or (_00306_, _00305_, _13301_);
  or (_00308_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  and (_00309_, _00308_, _13707_);
  and (_13948_[6], _00309_, _00306_);
  and (_13951_[0], _13310_, _13707_);
  nor (_13951_[1], _13320_, rst);
  and (_13951_[2], _13316_, _13707_);
  and (_00310_, _13324_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_00311_, _13326_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  or (_00312_, _00311_, _00310_);
  and (_13953_[0], _00312_, _13707_);
  and (_00313_, _13324_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_00314_, _13326_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  or (_00315_, _00314_, _00313_);
  and (_13953_[1], _00315_, _13707_);
  and (_00316_, _13324_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_00317_, _13326_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  or (_00318_, _00317_, _00316_);
  and (_13953_[2], _00318_, _13707_);
  and (_00319_, _13324_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_00320_, _13326_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  or (_00321_, _00320_, _00319_);
  and (_13953_[3], _00321_, _13707_);
  and (_00323_, _13324_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_00325_, _13326_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  or (_00326_, _00325_, _00323_);
  and (_13953_[4], _00326_, _13707_);
  and (_00328_, _13324_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_00329_, _13326_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  or (_00330_, _00329_, _00328_);
  and (_13953_[5], _00330_, _13707_);
  and (_00332_, _13324_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_00333_, _13326_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  or (_00335_, _00333_, _00332_);
  and (_13953_[6], _00335_, _13707_);
  and (_00336_, _13324_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_00338_, _13326_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  or (_00339_, _00338_, _00336_);
  and (_13953_[7], _00339_, _13707_);
  and (_00341_, _13324_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_00342_, _13326_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  or (_00343_, _00342_, _00341_);
  and (_13953_[8], _00343_, _13707_);
  and (_00345_, _13324_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_00346_, _13326_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  or (_00348_, _00346_, _00345_);
  and (_13953_[9], _00348_, _13707_);
  and (_00349_, _13324_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_00350_, _13326_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  or (_00351_, _00350_, _00349_);
  and (_13953_[10], _00351_, _13707_);
  and (_00352_, _13324_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_00353_, _13326_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  or (_00354_, _00353_, _00352_);
  and (_13953_[11], _00354_, _13707_);
  and (_00355_, _13324_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_00356_, _13326_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  or (_00357_, _00356_, _00355_);
  and (_13953_[12], _00357_, _13707_);
  and (_00358_, _13324_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_00359_, _13326_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  or (_00360_, _00359_, _00358_);
  and (_13953_[13], _00360_, _13707_);
  and (_00361_, _13324_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_00362_, _13326_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  or (_00363_, _00362_, _00361_);
  and (_13953_[14], _00363_, _13707_);
  and (_00365_, _13324_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_00367_, _13326_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  or (_00368_, _00367_, _00365_);
  and (_13953_[15], _00368_, _13707_);
  and (_00370_, _13324_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_00371_, _13326_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  or (_00372_, _00371_, _00370_);
  and (_13953_[16], _00372_, _13707_);
  and (_00374_, _13324_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_00375_, _13326_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  or (_00377_, _00375_, _00374_);
  and (_13953_[17], _00377_, _13707_);
  and (_00378_, _13324_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_00380_, _13326_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  or (_00381_, _00380_, _00378_);
  and (_13953_[18], _00381_, _13707_);
  and (_00383_, _13324_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_00384_, _13326_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  or (_00385_, _00384_, _00383_);
  and (_13953_[19], _00385_, _13707_);
  and (_00387_, _13324_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_00388_, _13326_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  or (_00390_, _00388_, _00387_);
  and (_13953_[20], _00390_, _13707_);
  and (_00391_, _13324_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_00392_, _13326_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  or (_00393_, _00392_, _00391_);
  and (_13953_[21], _00393_, _13707_);
  and (_00394_, _13324_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_00395_, _13326_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  or (_00396_, _00395_, _00394_);
  and (_13953_[22], _00396_, _13707_);
  and (_00397_, _13324_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_00398_, _13326_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  or (_00399_, _00398_, _00397_);
  and (_13953_[23], _00399_, _13707_);
  and (_00400_, _13324_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and (_00401_, _13326_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  or (_00402_, _00401_, _00400_);
  and (_13953_[24], _00402_, _13707_);
  and (_00403_, _13324_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and (_00404_, _13326_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  or (_00405_, _00404_, _00403_);
  and (_13953_[25], _00405_, _13707_);
  and (_00407_, _13324_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and (_00409_, _13326_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  or (_00410_, _00409_, _00407_);
  and (_13953_[26], _00410_, _13707_);
  and (_00412_, _13324_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and (_00413_, _13326_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  or (_00414_, _00413_, _00412_);
  and (_13953_[27], _00414_, _13707_);
  and (_00416_, _13324_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and (_00417_, _13326_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  or (_00419_, _00417_, _00416_);
  and (_13953_[28], _00419_, _13707_);
  and (_00420_, _13324_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and (_00422_, _13326_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  or (_00423_, _00422_, _00420_);
  and (_13953_[29], _00423_, _13707_);
  and (_00425_, _13324_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and (_00426_, _13326_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  or (_00427_, _00426_, _00425_);
  and (_13953_[30], _00427_, _13707_);
  not (_00429_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  nor (_00430_, _13333_, _00429_);
  and (_00432_, \oc8051_top_1.oc8051_decoder1.mem_act [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and (_00433_, _00432_, _13333_);
  or (_00434_, _00433_, _00430_);
  and (_13954_[0], _00434_, _13707_);
  not (_00435_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  nor (_00436_, _13333_, _00435_);
  and (_00437_, \oc8051_top_1.oc8051_decoder1.mem_act [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_00438_, _00437_, _13333_);
  or (_00439_, _00438_, _00436_);
  and (_13954_[1], _00439_, _13707_);
  not (_00440_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  nor (_00441_, _13333_, _00440_);
  and (_00442_, \oc8051_top_1.oc8051_decoder1.mem_act [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_00443_, _00442_, _13333_);
  or (_00444_, _00443_, _00441_);
  and (_13954_[2], _00444_, _13707_);
  not (_00445_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  nor (_00446_, _13333_, _00445_);
  and (_00447_, \oc8051_top_1.oc8051_decoder1.mem_act [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_00448_, _00447_, _13333_);
  or (_00449_, _00448_, _00446_);
  and (_13954_[3], _00449_, _13707_);
  not (_00451_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  nor (_00453_, _13333_, _00451_);
  and (_00454_, \oc8051_top_1.oc8051_decoder1.mem_act [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_00455_, _00454_, _13333_);
  or (_00457_, _00455_, _00453_);
  and (_13954_[4], _00457_, _13707_);
  not (_00458_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  nor (_00460_, _13333_, _00458_);
  and (_00461_, \oc8051_top_1.oc8051_decoder1.mem_act [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_00462_, _00461_, _13333_);
  or (_00464_, _00462_, _00460_);
  and (_13954_[5], _00464_, _13707_);
  not (_00465_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  nor (_00467_, _13333_, _00465_);
  and (_00468_, \oc8051_top_1.oc8051_decoder1.mem_act [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_00469_, _00468_, _13333_);
  or (_00471_, _00469_, _00467_);
  and (_13954_[6], _00471_, _13707_);
  not (_00472_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  nor (_00474_, _13333_, _00472_);
  or (_00475_, _10299_, _13344_);
  or (_00476_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_00478_, _00476_, _13333_);
  and (_00479_, _00478_, _00475_);
  or (_00480_, _00479_, _00474_);
  and (_13957_[0], _00480_, _13707_);
  not (_00481_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  nor (_00482_, _13333_, _00481_);
  or (_00483_, _10457_, _13344_);
  or (_00484_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_00485_, _00484_, _13333_);
  and (_00486_, _00485_, _00483_);
  or (_00487_, _00486_, _00482_);
  and (_13957_[1], _00487_, _13707_);
  not (_00488_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  nor (_00489_, _13333_, _00488_);
  or (_00490_, _10114_, _13344_);
  or (_00491_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_00492_, _00491_, _13333_);
  and (_00493_, _00492_, _00490_);
  or (_00494_, _00493_, _00489_);
  and (_13957_[2], _00494_, _13707_);
  not (_00495_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  nor (_00497_, _13333_, _00495_);
  or (_00498_, _10346_, _13344_);
  or (_00500_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_00501_, _00500_, _13333_);
  and (_00502_, _00501_, _00498_);
  or (_00504_, _00502_, _00497_);
  and (_13957_[3], _00504_, _13707_);
  not (_00505_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  nor (_00507_, _13333_, _00505_);
  or (_00508_, _10509_, _13344_);
  or (_00509_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_00511_, _00509_, _13333_);
  and (_00512_, _00511_, _00508_);
  or (_00513_, _00512_, _00507_);
  and (_13957_[4], _00513_, _13707_);
  not (_00515_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  nor (_00516_, _13333_, _00515_);
  or (_00518_, _10173_, _13344_);
  or (_00519_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_00520_, _00519_, _13333_);
  and (_00522_, _00520_, _00518_);
  or (_00523_, _00522_, _00516_);
  and (_13957_[5], _00523_, _13707_);
  not (_00525_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  nor (_00526_, _13333_, _00525_);
  or (_00527_, _10406_, _13344_);
  or (_00528_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_00529_, _00528_, _13333_);
  and (_00530_, _00529_, _00527_);
  or (_00531_, _00530_, _00526_);
  and (_13957_[6], _00531_, _13707_);
  not (_00532_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  nor (_00533_, _13333_, _00532_);
  or (_00534_, _10250_, _13344_);
  or (_00535_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_00536_, _00535_, _13333_);
  and (_00537_, _00536_, _00534_);
  or (_00538_, _00537_, _00533_);
  and (_13957_[7], _00538_, _13707_);
  not (_00539_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  nor (_00540_, _13333_, _00539_);
  and (_00541_, _13344_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and (_00542_, _00541_, _13333_);
  or (_00543_, _00542_, _00540_);
  and (_13957_[8], _00543_, _13707_);
  not (_00544_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  nor (_00546_, _13333_, _00544_);
  and (_00547_, _13344_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  and (_00548_, _00547_, _13333_);
  or (_00549_, _00548_, _00546_);
  and (_13957_[9], _00549_, _13707_);
  not (_00550_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  nor (_00551_, _13333_, _00550_);
  and (_00552_, _13344_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  and (_00553_, _00552_, _13333_);
  or (_00554_, _00553_, _00551_);
  and (_13957_[10], _00554_, _13707_);
  not (_00555_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  nor (_00556_, _13333_, _00555_);
  and (_00557_, _13344_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  and (_00558_, _00557_, _13333_);
  or (_00559_, _00558_, _00556_);
  and (_13957_[11], _00559_, _13707_);
  not (_00560_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  nor (_00561_, _13333_, _00560_);
  and (_00562_, _13344_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  and (_00563_, _00562_, _13333_);
  or (_00564_, _00563_, _00561_);
  and (_13957_[12], _00564_, _13707_);
  not (_00565_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  nor (_00566_, _13333_, _00565_);
  and (_00567_, _13344_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  and (_00568_, _00567_, _13333_);
  or (_00569_, _00568_, _00566_);
  and (_13957_[13], _00569_, _13707_);
  not (_00570_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  nor (_00571_, _13333_, _00570_);
  and (_00572_, _13344_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  and (_00573_, _00572_, _13333_);
  or (_00574_, _00573_, _00571_);
  and (_13957_[14], _00574_, _13707_);
  nand (_00575_, _13350_, _08105_);
  or (_00576_, _13350_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  and (_00577_, _00576_, _13707_);
  and (_13961_[0], _00577_, _00575_);
  or (_00578_, _13355_, _08166_);
  or (_00579_, _13350_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1]);
  and (_00580_, _00579_, _13707_);
  and (_13961_[1], _00580_, _00578_);
  nand (_00581_, _13350_, _08223_);
  or (_00582_, _13350_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2]);
  and (_00583_, _00582_, _13707_);
  and (_13961_[2], _00583_, _00581_);
  or (_00584_, _13355_, _08288_);
  or (_00585_, _13350_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3]);
  and (_00586_, _00585_, _13707_);
  and (_13961_[3], _00586_, _00584_);
  or (_00587_, _13355_, _08354_);
  or (_00588_, _13350_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [4]);
  and (_00589_, _00588_, _13707_);
  and (_13961_[4], _00589_, _00587_);
  or (_00590_, _13355_, _08428_);
  or (_00591_, _13350_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [5]);
  and (_00592_, _00591_, _13707_);
  and (_13961_[5], _00592_, _00590_);
  nand (_00593_, _13350_, _08499_);
  or (_00594_, _13350_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [6]);
  and (_00595_, _00594_, _13707_);
  and (_13961_[6], _00595_, _00593_);
  nand (_00596_, _13350_, _08001_);
  or (_00597_, _13350_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [7]);
  and (_00598_, _00597_, _13707_);
  and (_13961_[7], _00598_, _00596_);
  or (_00599_, _13355_, _09165_);
  or (_00600_, _13350_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [8]);
  and (_00601_, _00600_, _13707_);
  and (_13961_[8], _00601_, _00599_);
  nand (_00602_, _13350_, _09198_);
  or (_00603_, _13350_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [9]);
  and (_00604_, _00603_, _13707_);
  and (_13961_[9], _00604_, _00602_);
  nand (_00605_, _13350_, _09228_);
  or (_00606_, _13350_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [10]);
  and (_00607_, _00606_, _13707_);
  and (_13961_[10], _00607_, _00605_);
  nand (_00608_, _13350_, _09258_);
  or (_00609_, _13350_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [11]);
  and (_00610_, _00609_, _13707_);
  and (_13961_[11], _00610_, _00608_);
  nand (_00611_, _13350_, _09290_);
  or (_00612_, _13350_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [12]);
  and (_00613_, _00612_, _13707_);
  and (_13961_[12], _00613_, _00611_);
  nand (_00614_, _13350_, _09324_);
  or (_00615_, _13350_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [13]);
  and (_00616_, _00615_, _13707_);
  and (_13961_[13], _00616_, _00614_);
  nand (_00617_, _13350_, _09353_);
  or (_00618_, _13350_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [14]);
  and (_00619_, _00618_, _13707_);
  and (_13961_[14], _00619_, _00617_);
  nor (_13926_, _10041_, rst);
  nor (_00620_, _10429_, _10271_);
  nor (_00621_, _10537_, _10200_);
  and (_00622_, _00621_, _10372_);
  and (_00623_, _00622_, _00620_);
  not (_00624_, _00623_);
  nor (_00625_, _12793_, _10271_);
  and (_00626_, _00625_, _10372_);
  nor (_00627_, _10373_, _10271_);
  nor (_00628_, _10429_, _10199_);
  and (_00629_, _00628_, _00627_);
  nor (_00630_, _00629_, _00626_);
  nand (_00631_, _00630_, _00624_);
  not (_00632_, _09387_);
  and (_00633_, _08761_, _08775_);
  not (_00634_, _00633_);
  nor (_00635_, _12268_, _08774_);
  and (_00636_, _00635_, _00634_);
  nor (_00637_, _08789_, _08783_);
  and (_00638_, _00637_, _00636_);
  nor (_00639_, _12331_, _12269_);
  and (_00640_, _00639_, _00638_);
  and (_00641_, _08760_, _08751_);
  not (_00642_, _00641_);
  nor (_00643_, _12446_, _12333_);
  and (_00644_, _00643_, _00642_);
  and (_00645_, _00644_, _12599_);
  and (_00646_, _00645_, _00640_);
  and (_00647_, _00646_, _08820_);
  nor (_00648_, _00647_, _08522_);
  not (_00649_, _00648_);
  and (_00650_, _00649_, _00626_);
  nor (_00651_, _00650_, _00632_);
  and (_00652_, _00651_, _12809_);
  and (_00653_, _00652_, _00631_);
  and (_00654_, _00627_, _10537_);
  and (_00655_, _00654_, _00628_);
  and (_00656_, _00655_, _09487_);
  and (_00657_, _00631_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_00658_, _00657_, _12822_);
  nand (_00659_, _00658_, _08059_);
  not (_00660_, _10149_);
  nand (_00661_, _09555_, _09553_);
  nand (_00662_, _09569_, _00661_);
  or (_00663_, _09569_, _00661_);
  nand (_00664_, _00663_, _00662_);
  nand (_00665_, _09524_, _09523_);
  nand (_00666_, _09544_, _00665_);
  or (_00667_, _09544_, _00665_);
  and (_00668_, _00667_, _00666_);
  nand (_00669_, _00668_, _00664_);
  or (_00670_, _00668_, _00664_);
  nand (_00671_, _00670_, _00669_);
  nand (_00672_, _09593_, _09581_);
  or (_00673_, _09593_, _09581_);
  nand (_00674_, _00673_, _00672_);
  nand (_00675_, _09604_, _09602_);
  nand (_00676_, _00675_, _09514_);
  or (_00677_, _00675_, _09514_);
  and (_00678_, _00677_, _00676_);
  nand (_00679_, _00678_, _00674_);
  or (_00680_, _00678_, _00674_);
  nand (_00681_, _00680_, _00679_);
  nand (_00682_, _00681_, _00671_);
  or (_00683_, _00681_, _00671_);
  nand (_00684_, _00683_, _00682_);
  or (_00685_, _00684_, _00660_);
  and (_00686_, _10324_, _10485_);
  or (_00687_, _10149_, _09459_);
  and (_00688_, _00687_, _00686_);
  and (_00689_, _00688_, _00685_);
  nor (_00690_, _10324_, _10485_);
  and (_00691_, _00690_, _10149_);
  and (_00692_, _00691_, _09448_);
  or (_00693_, _10149_, _09468_);
  not (_00694_, _10485_);
  nor (_00695_, _10324_, _00694_);
  or (_00696_, _00660_, _09405_);
  and (_00697_, _00696_, _00695_);
  and (_00698_, _00697_, _00693_);
  and (_00699_, _00690_, _00660_);
  and (_00700_, _00699_, _09398_);
  or (_00701_, _00700_, _00698_);
  or (_00702_, _00701_, _00692_);
  or (_00703_, _00660_, _09441_);
  and (_00704_, _10324_, _00694_);
  or (_00705_, _10149_, _09484_);
  and (_00706_, _00705_, _00704_);
  and (_00707_, _00706_, _00703_);
  or (_00708_, _00707_, _00702_);
  or (_00709_, _00708_, _00689_);
  and (_00710_, _00709_, _00623_);
  or (_00711_, _10149_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nand (_00712_, _10149_, _08108_);
  and (_00713_, _00712_, _00686_);
  and (_00714_, _00713_, _00711_);
  and (_00715_, _00691_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  or (_00716_, _00715_, _00714_);
  nor (_00717_, _10149_, _08430_);
  and (_00718_, _10149_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  or (_00719_, _00718_, _00717_);
  and (_00720_, _00719_, _00695_);
  nor (_00721_, _10149_, _08502_);
  and (_00722_, _10149_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or (_00723_, _00722_, _00721_);
  and (_00724_, _00723_, _00704_);
  and (_00725_, _00699_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  or (_00726_, _00725_, _00724_);
  or (_00727_, _00726_, _00720_);
  or (_00728_, _00727_, _00716_);
  and (_00729_, _00728_, _00629_);
  or (_00730_, _12782_, p1in_reg[0]);
  or (_00731_, _12786_, p1_in[0]);
  and (_00732_, _00731_, _00730_);
  or (_00733_, _00732_, _00648_);
  or (_00734_, _00649_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and (_00735_, _00734_, _00733_);
  or (_00736_, _00735_, _00660_);
  or (_00737_, _12782_, p1in_reg[4]);
  or (_00738_, _12786_, p1_in[4]);
  and (_00739_, _00738_, _00737_);
  or (_00740_, _00739_, _00648_);
  or (_00741_, _00649_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_00742_, _00741_, _00740_);
  or (_00743_, _00742_, _10149_);
  and (_00744_, _00743_, _00686_);
  and (_00745_, _00744_, _00736_);
  or (_00746_, _12782_, p1in_reg[3]);
  or (_00747_, _12786_, p1_in[3]);
  and (_00748_, _00747_, _00746_);
  or (_00749_, _00748_, _00648_);
  or (_00750_, _00649_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_00751_, _00750_, _00749_);
  and (_00752_, _00751_, _00691_);
  or (_00753_, _00752_, _00745_);
  or (_00754_, _12782_, p1in_reg[5]);
  or (_00755_, _12786_, p1_in[5]);
  and (_00756_, _00755_, _00754_);
  or (_00757_, _00756_, _00648_);
  or (_00758_, _00649_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_00759_, _00758_, _00757_);
  and (_00760_, _00759_, _00660_);
  or (_00761_, _12782_, p1in_reg[1]);
  or (_00762_, _12786_, p1_in[1]);
  and (_00763_, _00762_, _00761_);
  or (_00764_, _00763_, _00648_);
  or (_00765_, _00649_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_00766_, _00765_, _00764_);
  and (_00767_, _00766_, _10149_);
  or (_00768_, _00767_, _00760_);
  and (_00769_, _00768_, _00695_);
  or (_00770_, _12782_, p1in_reg[6]);
  or (_00771_, _12786_, p1_in[6]);
  and (_00772_, _00771_, _00770_);
  or (_00773_, _00772_, _00648_);
  or (_00774_, _00649_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_00775_, _00774_, _00773_);
  and (_00776_, _00775_, _00660_);
  or (_00777_, _12782_, p1in_reg[2]);
  or (_00778_, _12786_, p1_in[2]);
  and (_00779_, _00778_, _00777_);
  or (_00780_, _00779_, _00648_);
  nand (_00781_, _00648_, _09792_);
  and (_00782_, _00781_, _00780_);
  and (_00783_, _00782_, _10149_);
  or (_00784_, _00783_, _00776_);
  and (_00785_, _00784_, _00704_);
  or (_00786_, _12782_, p1in_reg[7]);
  or (_00787_, _12786_, p1_in[7]);
  and (_00788_, _00787_, _00786_);
  or (_00789_, _00788_, _00648_);
  nand (_00790_, _00648_, _09627_);
  and (_00791_, _00790_, _00789_);
  and (_00792_, _00791_, _00699_);
  or (_00793_, _00792_, _00785_);
  or (_00794_, _00793_, _00769_);
  or (_00795_, _00794_, _00753_);
  and (_00796_, _00626_, _10199_);
  and (_00797_, _00796_, _00795_);
  or (_00798_, _00797_, _00729_);
  and (_00799_, _00798_, _10538_);
  nor (_00800_, _10149_, _06893_);
  and (_00801_, _10149_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_00802_, _00801_, _00800_);
  and (_00803_, _00802_, _00686_);
  and (_00804_, _00699_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_00805_, _00804_, _00803_);
  nor (_00806_, _10149_, _06929_);
  and (_00807_, _10149_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_00808_, _00807_, _00806_);
  and (_00809_, _00808_, _00695_);
  nor (_00810_, _10149_, _07013_);
  and (_00811_, _10149_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_00812_, _00811_, _00810_);
  and (_00813_, _00812_, _00704_);
  and (_00814_, _00691_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_00815_, _00814_, _00813_);
  or (_00816_, _00815_, _00809_);
  or (_00817_, _00816_, _00805_);
  and (_00818_, _00817_, _00655_);
  or (_00819_, _00818_, _00658_);
  or (_00820_, _12782_, p3in_reg[7]);
  or (_00821_, _12786_, p3_in[7]);
  and (_00822_, _00821_, _00820_);
  or (_00823_, _00822_, _00648_);
  nand (_00824_, _00648_, _09655_);
  and (_00825_, _00824_, _00823_);
  and (_00826_, _00825_, _00699_);
  or (_00827_, _12782_, p3in_reg[0]);
  or (_00828_, _12786_, p3_in[0]);
  and (_00829_, _00828_, _00827_);
  or (_00830_, _00829_, _00648_);
  or (_00831_, _00649_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and (_00832_, _00831_, _00830_);
  or (_00833_, _00832_, _00660_);
  or (_00834_, _12782_, p3in_reg[4]);
  or (_00835_, _12786_, p3_in[4]);
  and (_00836_, _00835_, _00834_);
  or (_00837_, _00836_, _00648_);
  or (_00838_, _00649_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_00839_, _00838_, _00837_);
  or (_00840_, _00839_, _10149_);
  and (_00841_, _00840_, _00686_);
  and (_00842_, _00841_, _00833_);
  or (_00843_, _12782_, p3in_reg[3]);
  or (_00844_, _12786_, p3_in[3]);
  and (_00845_, _00844_, _00843_);
  or (_00846_, _00845_, _00648_);
  or (_00847_, _00649_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_00848_, _00847_, _00846_);
  and (_00849_, _00848_, _00691_);
  or (_00850_, _00849_, _00842_);
  or (_00851_, _00850_, _00826_);
  or (_00852_, _12782_, p3in_reg[6]);
  or (_00853_, _12786_, p3_in[6]);
  and (_00854_, _00853_, _00852_);
  or (_00855_, _00854_, _00648_);
  or (_00856_, _00649_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and (_00857_, _00856_, _00855_);
  and (_00858_, _00857_, _00660_);
  or (_00859_, _12782_, p3in_reg[2]);
  or (_00860_, _12786_, p3_in[2]);
  and (_00861_, _00860_, _00859_);
  or (_00862_, _00861_, _00648_);
  nand (_00863_, _00648_, _09960_);
  and (_00864_, _00863_, _00862_);
  and (_00865_, _00864_, _10149_);
  or (_00866_, _00865_, _00858_);
  and (_00867_, _00866_, _00704_);
  or (_00868_, _12782_, p3in_reg[5]);
  or (_00869_, _12786_, p3_in[5]);
  and (_00870_, _00869_, _00868_);
  or (_00871_, _00870_, _00648_);
  or (_00872_, _00649_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_00873_, _00872_, _00871_);
  and (_00874_, _00873_, _00660_);
  or (_00875_, _12782_, p3in_reg[1]);
  or (_00876_, _12786_, p3_in[1]);
  and (_00877_, _00876_, _00875_);
  or (_00878_, _00877_, _00648_);
  or (_00879_, _00649_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_00880_, _00879_, _00878_);
  and (_00881_, _00880_, _10149_);
  or (_00882_, _00881_, _00874_);
  and (_00883_, _00882_, _00695_);
  or (_00884_, _00883_, _00867_);
  or (_00885_, _00884_, _00851_);
  and (_00886_, _10429_, _10200_);
  and (_00887_, _00886_, _10538_);
  and (_00888_, _00887_, _00627_);
  and (_00889_, _00888_, _00885_);
  or (_00890_, _12782_, p2in_reg[7]);
  or (_00891_, _12786_, p2_in[7]);
  and (_00892_, _00891_, _00890_);
  or (_00893_, _00892_, _00648_);
  nand (_00894_, _00648_, _09647_);
  and (_00895_, _00894_, _00893_);
  and (_00896_, _00895_, _00699_);
  or (_00897_, _12782_, p2in_reg[0]);
  or (_00898_, _12786_, p2_in[0]);
  and (_00899_, _00898_, _00897_);
  or (_00900_, _00899_, _00648_);
  or (_00901_, _00649_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and (_00902_, _00901_, _00900_);
  or (_00903_, _00902_, _00660_);
  or (_00904_, _12782_, p2in_reg[4]);
  or (_00905_, _12786_, p2_in[4]);
  and (_00906_, _00905_, _00904_);
  or (_00907_, _00906_, _00648_);
  or (_00908_, _00649_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_00909_, _00908_, _00907_);
  or (_00910_, _00909_, _10149_);
  and (_00911_, _00910_, _00686_);
  and (_00912_, _00911_, _00903_);
  or (_00913_, _12782_, p2in_reg[3]);
  or (_00914_, _12786_, p2_in[3]);
  and (_00915_, _00914_, _00913_);
  or (_00916_, _00915_, _00648_);
  or (_00917_, _00649_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_00918_, _00917_, _00916_);
  and (_00919_, _00918_, _00691_);
  or (_00920_, _00919_, _00912_);
  or (_00921_, _00920_, _00896_);
  or (_00922_, _12782_, p2in_reg[6]);
  or (_00923_, _12786_, p2_in[6]);
  and (_00924_, _00923_, _00922_);
  or (_00925_, _00924_, _00648_);
  or (_00926_, _00649_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_00927_, _00926_, _00925_);
  and (_00928_, _00927_, _00660_);
  or (_00929_, _12782_, p2in_reg[2]);
  or (_00930_, _12786_, p2_in[2]);
  and (_00931_, _00930_, _00929_);
  or (_00932_, _00931_, _00648_);
  nand (_00933_, _00648_, _09877_);
  and (_00934_, _00933_, _00932_);
  and (_00935_, _00934_, _10149_);
  or (_00936_, _00935_, _00928_);
  and (_00937_, _00936_, _00704_);
  or (_00938_, _12782_, p2in_reg[5]);
  or (_00939_, _12786_, p2_in[5]);
  and (_00940_, _00939_, _00938_);
  or (_00941_, _00940_, _00648_);
  or (_00942_, _00649_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_00943_, _00942_, _00941_);
  and (_00944_, _00943_, _00660_);
  or (_00945_, _12782_, p2in_reg[1]);
  or (_00946_, _12786_, p2_in[1]);
  and (_00947_, _00946_, _00945_);
  or (_00948_, _00947_, _00648_);
  or (_00949_, _00649_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_00950_, _00949_, _00948_);
  and (_00951_, _00950_, _10149_);
  or (_00952_, _00951_, _00944_);
  and (_00953_, _00952_, _00695_);
  or (_00954_, _00953_, _00937_);
  or (_00955_, _00954_, _00921_);
  and (_00956_, _00886_, _00654_);
  and (_00957_, _00956_, _00955_);
  or (_00958_, _00957_, _00889_);
  and (_00959_, _10537_, _10199_);
  and (_00960_, _00959_, _00626_);
  or (_00961_, _12782_, p0in_reg[7]);
  or (_00962_, _12786_, p0_in[7]);
  and (_00963_, _00962_, _00961_);
  or (_00964_, _00963_, _00648_);
  nand (_00965_, _00648_, _09617_);
  and (_00966_, _00965_, _00964_);
  and (_00967_, _00966_, _00699_);
  or (_00968_, _12782_, p0in_reg[3]);
  or (_00969_, _12786_, p0_in[3]);
  and (_00970_, _00969_, _00968_);
  or (_00971_, _00970_, _00648_);
  or (_00972_, _00649_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_00973_, _00972_, _00971_);
  and (_00974_, _00973_, _00691_);
  or (_00975_, _00974_, _00967_);
  or (_00976_, _12782_, p0in_reg[0]);
  or (_00977_, _12786_, p0_in[0]);
  and (_00978_, _00977_, _00976_);
  or (_00979_, _00978_, _00648_);
  or (_00980_, _00649_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  and (_00981_, _00980_, _00979_);
  or (_00982_, _00981_, _00660_);
  or (_00983_, _12782_, p0in_reg[4]);
  or (_00984_, _12786_, p0_in[4]);
  and (_00985_, _00984_, _00983_);
  or (_00986_, _00985_, _00648_);
  or (_00987_, _00649_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_00988_, _00987_, _00986_);
  or (_00989_, _00988_, _10149_);
  and (_00990_, _00989_, _00686_);
  and (_00991_, _00990_, _00982_);
  or (_00992_, _12782_, p0in_reg[6]);
  or (_00993_, _12786_, p0_in[6]);
  and (_00994_, _00993_, _00992_);
  or (_00995_, _00994_, _00648_);
  nand (_00996_, _00648_, _09751_);
  and (_00997_, _00996_, _00995_);
  and (_00998_, _00997_, _00660_);
  or (_00999_, _12782_, p0in_reg[2]);
  or (_01000_, _12786_, p0_in[2]);
  and (_01001_, _01000_, _00999_);
  or (_01002_, _01001_, _00648_);
  nand (_01003_, _00648_, _09707_);
  and (_01004_, _01003_, _01002_);
  and (_01005_, _01004_, _10149_);
  or (_01006_, _01005_, _00998_);
  and (_01007_, _01006_, _00704_);
  or (_01008_, _12782_, p0in_reg[5]);
  or (_01009_, _12786_, p0_in[5]);
  and (_01010_, _01009_, _01008_);
  or (_01011_, _01010_, _00648_);
  or (_01012_, _00649_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_01013_, _01012_, _01011_);
  and (_01014_, _01013_, _00660_);
  or (_01015_, _12782_, p0in_reg[1]);
  or (_01016_, _12786_, p0_in[1]);
  and (_01018_, _01016_, _01015_);
  or (_01019_, _01018_, _00648_);
  or (_01020_, _00649_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_01021_, _01020_, _01019_);
  and (_01022_, _01021_, _10149_);
  or (_01023_, _01022_, _01014_);
  and (_01024_, _01023_, _00695_);
  or (_01025_, _01024_, _01007_);
  or (_01026_, _01025_, _00991_);
  or (_01027_, _01026_, _00975_);
  and (_01028_, _01027_, _00960_);
  or (_01029_, _01028_, _00958_);
  or (_01030_, _01029_, _00819_);
  or (_01031_, _01030_, _00799_);
  or (_01032_, _01031_, _00710_);
  and (_01033_, _01032_, _00659_);
  or (_01034_, _01033_, _00656_);
  and (_01035_, _10149_, _09525_);
  and (_01036_, _00660_, _09581_);
  or (_01037_, _01036_, _01035_);
  and (_01038_, _01037_, _00686_);
  and (_01039_, _10149_, _09556_);
  and (_01040_, _00660_, _09605_);
  or (_01041_, _01040_, _01039_);
  and (_01042_, _01041_, _00704_);
  and (_01043_, _10149_, _09544_);
  and (_01044_, _00660_, _09593_);
  or (_01045_, _01044_, _01043_);
  and (_01046_, _01045_, _00695_);
  and (_01047_, _00699_, _09514_);
  and (_01049_, _00691_, _09569_);
  or (_01050_, _01049_, _01047_);
  or (_01051_, _01050_, _01046_);
  or (_01052_, _01051_, _01042_);
  nor (_01053_, _01052_, _01038_);
  nand (_01054_, _01053_, _00656_);
  and (_01055_, _01054_, _01034_);
  or (_01056_, _01055_, _00653_);
  or (_01057_, _10149_, _10383_);
  nand (_01058_, _10149_, _08960_);
  and (_01059_, _01058_, _00704_);
  and (_01060_, _01059_, _01057_);
  or (_01061_, _10149_, _10487_);
  nand (_01062_, _10149_, _08975_);
  and (_01063_, _01062_, _00686_);
  and (_01064_, _01063_, _01061_);
  or (_01065_, _01064_, _01060_);
  and (_01066_, _00691_, _10326_);
  not (_01067_, _08997_);
  and (_01068_, _00699_, _01067_);
  and (_01070_, _10149_, _10436_);
  nor (_01071_, _10149_, _08937_);
  or (_01072_, _01071_, _01070_);
  and (_01073_, _01072_, _00695_);
  or (_01074_, _01073_, _01068_);
  or (_01075_, _01074_, _01066_);
  nor (_01076_, _01075_, _01065_);
  nand (_01077_, _01076_, _00653_);
  and (_01078_, _01077_, _13707_);
  and (_13967_, _01078_, _01056_);
  and (_01079_, _00959_, _00625_);
  and (_01080_, _10372_, _10149_);
  and (_01081_, _01080_, _00690_);
  and (_01082_, _01081_, _01079_);
  and (_01083_, _01082_, _09048_);
  and (_01084_, _01080_, _00686_);
  and (_01085_, _01084_, _00620_);
  and (_01086_, _01085_, _00621_);
  and (_01087_, _01086_, _12882_);
  nor (_01088_, _01087_, _01083_);
  nor (_01089_, _01088_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_01090_, _01089_);
  or (_01091_, _09498_, _09487_);
  and (_01092_, _10537_, _10200_);
  and (_01093_, _01092_, _01085_);
  and (_01094_, _01093_, _01091_);
  not (_01095_, _09500_);
  nor (_01096_, _00699_, _01095_);
  and (_01097_, _01096_, _12809_);
  nor (_01098_, _01097_, _01094_);
  and (_01099_, _01098_, _12825_);
  and (_01100_, _01099_, _01090_);
  and (_01101_, _01080_, _00704_);
  and (_01102_, _01101_, _01079_);
  and (_01103_, _01102_, _09048_);
  or (_01104_, _01103_, rst);
  nor (_13968_, _01104_, _01100_);
  nand (_01105_, _01103_, _08001_);
  or (_01106_, _01100_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  nor (_01107_, _10537_, _10199_);
  and (_01108_, _01107_, _01085_);
  and (_01109_, _01108_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_01110_, _01093_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_01111_, _01110_, _01109_);
  and (_01112_, _01086_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  and (_01113_, _01084_, _00625_);
  and (_01114_, _01113_, _00621_);
  and (_01115_, _01114_, _00791_);
  or (_01116_, _01115_, _01112_);
  or (_01117_, _01116_, _01111_);
  and (_01118_, _01113_, _01092_);
  and (_01119_, _01118_, _00895_);
  and (_01120_, _01113_, _01107_);
  and (_01121_, _01120_, _00825_);
  or (_01122_, _01121_, _01119_);
  and (_01123_, _01102_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_01124_, _01082_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_01125_, _01124_, _01123_);
  and (_01126_, _01080_, _00695_);
  and (_01127_, _01126_, _01079_);
  and (_01128_, _01127_, _08999_);
  and (_01129_, _01084_, _01079_);
  and (_01130_, _01129_, _00966_);
  or (_01131_, _01130_, _01128_);
  or (_01132_, _01131_, _01125_);
  or (_01133_, _01132_, _01122_);
  nor (_01134_, _01133_, _01117_);
  nand (_01135_, _01134_, _01100_);
  and (_01136_, _01135_, _01106_);
  or (_01137_, _01136_, _01103_);
  and (_01138_, _01137_, _13707_);
  and (_13969_[7], _01138_, _01105_);
  and (_01139_, _01086_, _00684_);
  and (_01140_, _01118_, _00902_);
  and (_01141_, _01093_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and (_01142_, _01120_, _00832_);
  or (_01143_, _01142_, _01141_);
  or (_01144_, _01143_, _01140_);
  and (_01145_, _01082_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and (_01146_, _01127_, _10302_);
  or (_01147_, _01146_, _01145_);
  and (_01148_, _01102_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_01149_, _01129_, _00981_);
  or (_01150_, _01149_, _01148_);
  or (_01151_, _01150_, _01147_);
  and (_01152_, _01108_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  and (_01153_, _01114_, _00735_);
  or (_01154_, _01153_, _01152_);
  or (_01155_, _01154_, _01151_);
  nor (_01156_, _01155_, _01144_);
  nand (_01157_, _01156_, _01100_);
  or (_01158_, _01157_, _01139_);
  or (_01159_, _01100_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  and (_01160_, _01159_, _01158_);
  or (_01161_, _01160_, _01103_);
  nand (_01162_, _01103_, _08105_);
  and (_01163_, _01162_, _13707_);
  and (_13969_[0], _01163_, _01161_);
  nand (_01164_, _01103_, _09168_);
  or (_01165_, _01100_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  and (_01166_, _01093_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_01167_, _01086_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  or (_01168_, _01167_, _01166_);
  and (_01169_, _01108_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_01170_, _01114_, _00766_);
  or (_01171_, _01170_, _01169_);
  or (_01172_, _01171_, _01168_);
  and (_01173_, _01118_, _00950_);
  and (_01174_, _01120_, _00880_);
  or (_01175_, _01174_, _01173_);
  and (_01176_, _01082_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  and (_01177_, _01129_, _01021_);
  or (_01178_, _01177_, _01176_);
  and (_01179_, _01102_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_01180_, _01127_, _10460_);
  or (_01181_, _01180_, _01179_);
  or (_01182_, _01181_, _01178_);
  or (_01183_, _01182_, _01175_);
  nor (_01184_, _01183_, _01172_);
  nand (_01185_, _01184_, _01100_);
  and (_01186_, _01185_, _01165_);
  or (_01187_, _01186_, _01103_);
  and (_01188_, _01187_, _13707_);
  and (_13969_[1], _01188_, _01164_);
  nand (_01189_, _01103_, _08223_);
  or (_01190_, _01100_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  and (_01191_, _01086_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  and (_01192_, _01118_, _00934_);
  or (_01193_, _01192_, _01191_);
  and (_01194_, _01108_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_01195_, _01114_, _00782_);
  or (_01196_, _01195_, _01194_);
  or (_01197_, _01196_, _01193_);
  and (_01198_, _01082_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  and (_01199_, _01127_, _10119_);
  or (_01200_, _01199_, _01198_);
  and (_01201_, _01102_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_01202_, _01129_, _01004_);
  or (_01203_, _01202_, _01201_);
  or (_01204_, _01203_, _01200_);
  and (_01205_, _01093_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_01206_, _01120_, _00864_);
  or (_01207_, _01206_, _01205_);
  or (_01208_, _01207_, _01204_);
  nor (_01209_, _01208_, _01197_);
  nand (_01210_, _01209_, _01100_);
  and (_01211_, _01210_, _01190_);
  or (_01212_, _01211_, _01103_);
  and (_01213_, _01212_, _13707_);
  and (_13969_[2], _01213_, _01189_);
  nand (_01214_, _01103_, _09231_);
  or (_01215_, _01100_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  and (_01216_, _01108_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_01217_, _01086_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  or (_01218_, _01217_, _01216_);
  and (_01219_, _01093_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_01220_, _01114_, _00751_);
  or (_01221_, _01220_, _01219_);
  or (_01222_, _01221_, _01218_);
  and (_01223_, _01118_, _00918_);
  and (_01224_, _01120_, _00848_);
  or (_01225_, _01224_, _01223_);
  and (_01226_, _01127_, _10349_);
  and (_01227_, _01129_, _00973_);
  or (_01228_, _01227_, _01226_);
  and (_01229_, _01102_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_01230_, _01082_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_01231_, _01230_, _01229_);
  or (_01232_, _01231_, _01228_);
  or (_01233_, _01232_, _01225_);
  nor (_01234_, _01233_, _01222_);
  nand (_01235_, _01234_, _01100_);
  and (_01236_, _01235_, _01215_);
  or (_01237_, _01236_, _01103_);
  and (_01238_, _01237_, _13707_);
  and (_13969_[3], _01238_, _01214_);
  nand (_01239_, _01103_, _09261_);
  or (_01240_, _01100_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  and (_01241_, _01108_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_01242_, _01093_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or (_01243_, _01242_, _01241_);
  and (_01244_, _01086_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_01245_, _01114_, _00742_);
  or (_01246_, _01245_, _01244_);
  or (_01247_, _01246_, _01243_);
  and (_01248_, _01118_, _00909_);
  and (_01249_, _01120_, _00839_);
  or (_01250_, _01249_, _01248_);
  and (_01251_, _01127_, _10511_);
  and (_01252_, _01129_, _00988_);
  or (_01253_, _01252_, _01251_);
  and (_01254_, _01102_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_01255_, _01082_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or (_01256_, _01255_, _01254_);
  or (_01257_, _01256_, _01253_);
  or (_01258_, _01257_, _01250_);
  nor (_01259_, _01258_, _01247_);
  nand (_01260_, _01259_, _01100_);
  and (_01261_, _01260_, _01240_);
  or (_01262_, _01261_, _01103_);
  and (_01263_, _01262_, _13707_);
  and (_13969_[4], _01263_, _01239_);
  nand (_01264_, _01103_, _09293_);
  or (_01265_, _01100_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  and (_01266_, _01108_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_01267_, _01086_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  or (_01268_, _01267_, _01266_);
  and (_01269_, _01093_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_01270_, _01114_, _00759_);
  or (_01271_, _01270_, _01269_);
  or (_01272_, _01271_, _01268_);
  and (_01273_, _01118_, _00943_);
  and (_01274_, _01120_, _00873_);
  or (_01275_, _01274_, _01273_);
  and (_01276_, _01102_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_01277_, _01129_, _01013_);
  or (_01278_, _01277_, _01276_);
  and (_01279_, _01082_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  and (_01280_, _01127_, _10175_);
  or (_01281_, _01280_, _01279_);
  or (_01282_, _01281_, _01278_);
  or (_01283_, _01282_, _01275_);
  nor (_01284_, _01283_, _01272_);
  nand (_01285_, _01284_, _01100_);
  and (_01286_, _01285_, _01265_);
  or (_01287_, _01286_, _01103_);
  and (_01288_, _01287_, _13707_);
  and (_13969_[5], _01288_, _01264_);
  nand (_01289_, _01103_, _08499_);
  or (_01290_, _01100_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  and (_01291_, _01093_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_01292_, _01086_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  or (_01293_, _01292_, _01291_);
  and (_01294_, _01108_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_01295_, _01114_, _00775_);
  or (_01296_, _01295_, _01294_);
  or (_01297_, _01296_, _01293_);
  and (_01298_, _01118_, _00927_);
  and (_01299_, _01120_, _00857_);
  or (_01300_, _01299_, _01298_);
  and (_01301_, _01127_, _10408_);
  and (_01302_, _01129_, _00997_);
  or (_01303_, _01302_, _01301_);
  and (_01304_, _01102_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_01305_, _01082_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_01306_, _01305_, _01304_);
  or (_01307_, _01306_, _01303_);
  or (_01308_, _01307_, _01300_);
  nor (_01309_, _01308_, _01297_);
  nand (_01310_, _01309_, _01100_);
  and (_01311_, _01310_, _01290_);
  or (_01312_, _01311_, _01103_);
  and (_01313_, _01312_, _13707_);
  and (_13969_[6], _01313_, _01289_);
  and (_13963_, _10550_, _13707_);
  and (_13964_[7], _10237_, _13707_);
  nor (_13966_[2], _10149_, rst);
  and (_13964_[0], _10287_, _13707_);
  and (_13964_[1], _10445_, _13707_);
  and (_13964_[2], _10098_, _13707_);
  and (_13964_[3], _10334_, _13707_);
  nor (_13964_[4], _10505_, rst);
  nor (_13964_[5], _10160_, rst);
  nor (_13964_[6], _10393_, rst);
  nor (_13966_[0], _10324_, rst);
  nor (_13966_[1], _10485_, rst);
  nor (_01314_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_01315_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _13301_);
  nor (_01316_, _01315_, _01314_);
  nor (_01317_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_01318_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _13301_);
  nor (_01319_, _01318_, _01317_);
  nor (_01320_, _01319_, _01316_);
  not (_01321_, _01320_);
  nor (_01322_, _13595_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_01323_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _13301_);
  nor (_01324_, _01323_, _01322_);
  and (_01325_, _01324_, _01321_);
  nor (_01326_, _01324_, _01321_);
  nor (_01327_, _01326_, _01325_);
  nor (_01328_, _13613_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_01329_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _13301_);
  nor (_01330_, _01329_, _01328_);
  not (_01331_, _01330_);
  and (_01332_, _01331_, _01325_);
  nor (_01333_, _01331_, _01325_);
  nor (_01334_, _01333_, _01332_);
  nor (_01335_, _01334_, _01327_);
  and (_01336_, _01319_, _01316_);
  and (_01337_, _01336_, _01335_);
  and (_01338_, _01337_, _11820_);
  not (_01339_, _01316_);
  and (_01340_, _01319_, _01339_);
  and (_01341_, _01340_, _01335_);
  and (_01342_, _01341_, _11763_);
  or (_01343_, _01342_, _01338_);
  nor (_01344_, _01319_, _01339_);
  and (_01345_, _01344_, _01335_);
  and (_01346_, _01345_, _11706_);
  and (_01347_, _01324_, _01320_);
  and (_01348_, _01331_, _01347_);
  and (_01349_, _01348_, _11651_);
  or (_01350_, _01349_, _01346_);
  or (_01351_, _01350_, _01343_);
  and (_01352_, _01331_, _01326_);
  and (_01353_, _01352_, _11471_);
  and (_01354_, _01331_, _01327_);
  and (_01355_, _01354_, _01340_);
  and (_01356_, _01355_, _11553_);
  and (_01357_, _01354_, _01336_);
  and (_01358_, _01357_, _11597_);
  or (_01359_, _01358_, _01356_);
  or (_01360_, _01359_, _01353_);
  and (_01361_, _01354_, _01344_);
  and (_01362_, _01361_, _11512_);
  not (_01363_, _01327_);
  and (_01364_, _01334_, _01363_);
  and (_01365_, _01340_, _01364_);
  and (_01366_, _01365_, _11389_);
  or (_01367_, _01366_, _01362_);
  or (_01368_, _01367_, _01360_);
  or (_01369_, _01368_, _01351_);
  and (_01370_, _01336_, _01333_);
  and (_01371_, _01370_, _12048_);
  and (_01372_, _01340_, _01333_);
  and (_01373_, _01372_, _11991_);
  or (_01374_, _01373_, _01371_);
  and (_01375_, _01330_, _01326_);
  and (_01376_, _01375_, _11876_);
  and (_01377_, _01344_, _01333_);
  and (_01378_, _01377_, _11934_);
  or (_01379_, _01378_, _01376_);
  or (_01380_, _01379_, _01374_);
  and (_01381_, _01330_, _01347_);
  and (_01382_, _01381_, _12090_);
  and (_01383_, _01364_, _01336_);
  and (_01384_, _01383_, _11430_);
  and (_01385_, _01364_, _01344_);
  and (_01386_, _01385_, _11348_);
  or (_01387_, _01386_, _01384_);
  or (_01388_, _01387_, _01382_);
  or (_01389_, _01388_, _01380_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [31], _01389_, _01369_);
  and (_01390_, _01372_, _11876_);
  and (_01391_, _01370_, _11934_);
  or (_01392_, _01391_, _01390_);
  and (_01393_, _01385_, _12048_);
  or (_01394_, _01393_, _01392_);
  and (_01395_, _01337_, _11706_);
  and (_01396_, _01365_, _12090_);
  or (_01397_, _01396_, _01395_);
  or (_01398_, _01397_, _01394_);
  and (_01399_, _01348_, _11553_);
  and (_01400_, _01355_, _11471_);
  and (_01401_, _01357_, _11512_);
  or (_01402_, _01401_, _01400_);
  or (_01403_, _01402_, _01399_);
  and (_01404_, _01352_, _11389_);
  and (_01405_, _01345_, _11597_);
  or (_01406_, _01405_, _01404_);
  or (_01407_, _01406_, _01403_);
  or (_01408_, _01407_, _01398_);
  and (_01409_, _01381_, _11991_);
  and (_01410_, _01383_, _11348_);
  and (_01411_, _01361_, _11430_);
  or (_01412_, _01411_, _01410_);
  and (_01413_, _01341_, _11651_);
  and (_01414_, _01375_, _11763_);
  and (_01415_, _01377_, _11820_);
  or (_01416_, _01415_, _01414_);
  or (_01417_, _01416_, _01413_);
  or (_01418_, _01417_, _01412_);
  or (_01419_, _01418_, _01409_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [15], _01419_, _01408_);
  and (_01420_, _01337_, _11763_);
  and (_01421_, _01385_, _12090_);
  and (_01422_, _01365_, _11348_);
  or (_01423_, _01422_, _01421_);
  or (_01424_, _01423_, _01420_);
  and (_01425_, _01355_, _11512_);
  and (_01426_, _01348_, _11597_);
  and (_01427_, _01352_, _11430_);
  or (_01428_, _01427_, _01426_);
  and (_01429_, _01381_, _12048_);
  and (_01430_, _01375_, _11820_);
  or (_01431_, _01430_, _01429_);
  or (_01432_, _01431_, _01428_);
  or (_01433_, _01432_, _01425_);
  and (_01434_, _01357_, _11553_);
  and (_01435_, _01361_, _11471_);
  or (_01436_, _01435_, _01434_);
  or (_01437_, _01436_, _01433_);
  and (_01438_, _01341_, _11706_);
  and (_01439_, _01370_, _11991_);
  and (_01440_, _01372_, _11934_);
  and (_01441_, _01377_, _11876_);
  or (_01442_, _01441_, _01440_);
  or (_01443_, _01442_, _01439_);
  or (_01444_, _01443_, _01438_);
  and (_01445_, _01383_, _11389_);
  and (_01446_, _01345_, _11651_);
  or (_01447_, _01446_, _01445_);
  or (_01448_, _01447_, _01444_);
  or (_01449_, _01448_, _01437_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [23], _01449_, _01424_);
  and (_01450_, _01341_, _11597_);
  and (_01451_, _01365_, _12048_);
  and (_01452_, _01345_, _11553_);
  or (_01453_, _01452_, _01451_);
  or (_01454_, _01453_, _01450_);
  and (_01455_, _01361_, _11389_);
  and (_01456_, _01375_, _11706_);
  and (_01457_, _01348_, _11512_);
  or (_01458_, _01457_, _01456_);
  and (_01459_, _01381_, _11934_);
  and (_01460_, _01352_, _11348_);
  or (_01461_, _01460_, _01459_);
  or (_01462_, _01461_, _01458_);
  or (_01463_, _01462_, _01455_);
  and (_01464_, _01355_, _11430_);
  and (_01465_, _01357_, _11471_);
  or (_01466_, _01465_, _01464_);
  or (_01467_, _01466_, _01463_);
  and (_01468_, _01337_, _11651_);
  and (_01469_, _01370_, _11876_);
  and (_01470_, _01377_, _11763_);
  and (_01471_, _01372_, _11820_);
  or (_01472_, _01471_, _01470_);
  or (_01473_, _01472_, _01469_);
  or (_01474_, _01473_, _01468_);
  and (_01475_, _01383_, _12090_);
  and (_01476_, _01385_, _11991_);
  or (_01477_, _01476_, _01475_);
  or (_01478_, _01477_, _01474_);
  or (_01479_, _01478_, _01467_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [7], _01479_, _01454_);
  and (_01480_, _01365_, _11394_);
  and (_01481_, _01337_, _11827_);
  and (_01482_, _01341_, _11770_);
  or (_01483_, _01482_, _01481_);
  or (_01484_, _01483_, _01480_);
  and (_01485_, _01355_, _11558_);
  and (_01486_, _01357_, _11603_);
  or (_01487_, _01486_, _01485_);
  and (_01488_, _01361_, _11517_);
  and (_01489_, _01375_, _11884_);
  and (_01490_, _01348_, _11656_);
  or (_01491_, _01490_, _01489_);
  and (_01492_, _01381_, _12095_);
  and (_01493_, _01352_, _11476_);
  or (_01494_, _01493_, _01492_);
  or (_01495_, _01494_, _01491_);
  or (_01496_, _01495_, _01488_);
  or (_01497_, _01496_, _01487_);
  and (_01498_, _01385_, _11353_);
  and (_01499_, _01383_, _11435_);
  or (_01500_, _01499_, _01498_);
  and (_01501_, _01345_, _11713_);
  and (_01502_, _01377_, _11941_);
  and (_01503_, _01370_, _12054_);
  and (_01504_, _01372_, _11998_);
  or (_01505_, _01504_, _01503_);
  or (_01506_, _01505_, _01502_);
  or (_01507_, _01506_, _01501_);
  or (_01508_, _01507_, _01500_);
  or (_01509_, _01508_, _01497_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [24], _01509_, _01484_);
  and (_01510_, _01337_, _11833_);
  and (_01511_, _01383_, _11440_);
  and (_01512_, _01341_, _11777_);
  or (_01513_, _01512_, _01511_);
  or (_01514_, _01513_, _01510_);
  and (_01515_, _01357_, _11609_);
  and (_01516_, _01381_, _12100_);
  and (_01517_, _01348_, _11663_);
  or (_01518_, _01517_, _01516_);
  and (_01519_, _01352_, _11481_);
  and (_01520_, _01375_, _11890_);
  or (_01521_, _01520_, _01519_);
  or (_01522_, _01521_, _01518_);
  or (_01523_, _01522_, _01515_);
  and (_01524_, _01355_, _11563_);
  and (_01525_, _01361_, _11522_);
  or (_01526_, _01525_, _01524_);
  or (_01527_, _01526_, _01523_);
  and (_01528_, _01345_, _11719_);
  and (_01529_, _01370_, _12059_);
  and (_01530_, _01372_, _12005_);
  or (_01531_, _01530_, _01529_);
  and (_01532_, _01377_, _11947_);
  or (_01533_, _01532_, _01531_);
  or (_01534_, _01533_, _01528_);
  and (_01535_, _01385_, _11358_);
  and (_01536_, _01365_, _11399_);
  or (_01537_, _01536_, _01535_);
  or (_01538_, _01537_, _01534_);
  or (_01539_, _01538_, _01527_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [25], _01539_, _01514_);
  and (_01540_, _01345_, _11726_);
  and (_01541_, _01337_, _11840_);
  and (_01542_, _01341_, _11784_);
  or (_01543_, _01542_, _01541_);
  or (_01544_, _01543_, _01540_);
  and (_01545_, _01355_, _11568_);
  and (_01546_, _01357_, _11615_);
  or (_01547_, _01546_, _01545_);
  and (_01548_, _01361_, _11527_);
  and (_01549_, _01348_, _11670_);
  and (_01550_, _01352_, _11486_);
  or (_01551_, _01550_, _01549_);
  and (_01552_, _01381_, _12105_);
  and (_01553_, _01375_, _11897_);
  or (_01554_, _01553_, _01552_);
  or (_01555_, _01554_, _01551_);
  or (_01556_, _01555_, _01548_);
  or (_01557_, _01556_, _01547_);
  and (_01558_, _01383_, _11445_);
  and (_01559_, _01377_, _11954_);
  and (_01560_, _01372_, _12012_);
  and (_01561_, _01370_, _12064_);
  or (_01562_, _01561_, _01560_);
  or (_01563_, _01562_, _01559_);
  or (_01564_, _01563_, _01558_);
  and (_01565_, _01385_, _11363_);
  and (_01566_, _01365_, _11404_);
  or (_01567_, _01566_, _01565_);
  or (_01568_, _01567_, _01564_);
  or (_01569_, _01568_, _01557_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [26], _01569_, _01544_);
  and (_01570_, _01345_, _11733_);
  and (_01571_, _01337_, _11847_);
  and (_01572_, _01341_, _11791_);
  or (_01573_, _01572_, _01571_);
  or (_01574_, _01573_, _01570_);
  and (_01575_, _01357_, _11622_);
  and (_01576_, _01355_, _11573_);
  or (_01577_, _01576_, _01575_);
  and (_01578_, _01361_, _11532_);
  and (_01579_, _01348_, _11677_);
  and (_01580_, _01352_, _11491_);
  or (_01581_, _01580_, _01579_);
  and (_01582_, _01381_, _12110_);
  and (_01583_, _01375_, _11904_);
  or (_01584_, _01583_, _01582_);
  or (_01585_, _01584_, _01581_);
  or (_01586_, _01585_, _01578_);
  or (_01587_, _01586_, _01577_);
  and (_01588_, _01383_, _11450_);
  and (_01589_, _01377_, _11961_);
  and (_01590_, _01372_, _12019_);
  and (_01591_, _01370_, _12069_);
  or (_01592_, _01591_, _01590_);
  or (_01593_, _01592_, _01589_);
  or (_01594_, _01593_, _01588_);
  and (_01595_, _01385_, _11368_);
  and (_01596_, _01365_, _11409_);
  or (_01597_, _01596_, _01595_);
  or (_01598_, _01597_, _01594_);
  or (_01599_, _01598_, _01587_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [27], _01599_, _01574_);
  and (_01600_, _01345_, _11741_);
  and (_01601_, _01341_, _11798_);
  and (_01602_, _01337_, _11854_);
  or (_01603_, _01602_, _01601_);
  or (_01604_, _01603_, _01600_);
  and (_01605_, _01375_, _11912_);
  and (_01606_, _01370_, _12074_);
  and (_01607_, _01372_, _12026_);
  or (_01608_, _01607_, _01606_);
  or (_01609_, _01608_, _01605_);
  and (_01610_, _01348_, _11684_);
  and (_01611_, _01377_, _11969_);
  or (_01612_, _01611_, _01610_);
  or (_01613_, _01612_, _01609_);
  or (_01614_, _01613_, _01604_);
  and (_01615_, _01365_, _11414_);
  and (_01616_, _01357_, _11628_);
  and (_01617_, _01355_, _11578_);
  or (_01618_, _01617_, _01616_);
  and (_01619_, _01352_, _11496_);
  and (_01620_, _01361_, _11537_);
  or (_01621_, _01620_, _01619_);
  or (_01622_, _01621_, _01618_);
  or (_01623_, _01622_, _01615_);
  and (_01624_, _01381_, _12115_);
  and (_01625_, _01383_, _11455_);
  and (_01626_, _01385_, _11373_);
  or (_01627_, _01626_, _01625_);
  or (_01628_, _01627_, _01624_);
  or (_01629_, _01628_, _01623_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [28], _01629_, _01614_);
  and (_01630_, _01345_, _11747_);
  and (_01631_, _01337_, _11861_);
  and (_01632_, _01341_, _11805_);
  or (_01633_, _01632_, _01631_);
  or (_01634_, _01633_, _01630_);
  and (_01635_, _01357_, _11635_);
  and (_01636_, _01348_, _11691_);
  and (_01637_, _01352_, _11501_);
  or (_01638_, _01637_, _01636_);
  and (_01639_, _01381_, _12120_);
  and (_01640_, _01375_, _11918_);
  or (_01641_, _01640_, _01639_);
  or (_01642_, _01641_, _01638_);
  or (_01643_, _01642_, _01635_);
  and (_01644_, _01355_, _11583_);
  and (_01645_, _01361_, _11542_);
  or (_01646_, _01645_, _01644_);
  or (_01647_, _01646_, _01643_);
  and (_01648_, _01383_, _11460_);
  and (_01649_, _01370_, _12079_);
  and (_01650_, _01372_, _12033_);
  or (_01651_, _01650_, _01649_);
  and (_01652_, _01377_, _11975_);
  or (_01653_, _01652_, _01651_);
  or (_01654_, _01653_, _01648_);
  and (_01655_, _01385_, _11378_);
  and (_01656_, _01365_, _11419_);
  or (_01657_, _01656_, _01655_);
  or (_01658_, _01657_, _01654_);
  or (_01659_, _01658_, _01647_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [29], _01659_, _01634_);
  and (_01660_, _01345_, _11754_);
  and (_01661_, _01337_, _11868_);
  and (_01662_, _01341_, _11812_);
  or (_01663_, _01662_, _01661_);
  or (_01664_, _01663_, _01660_);
  and (_01665_, _01355_, _11589_);
  and (_01666_, _01357_, _11642_);
  or (_01667_, _01666_, _01665_);
  and (_01668_, _01361_, _11547_);
  and (_01669_, _01348_, _11698_);
  and (_01670_, _01352_, _11506_);
  or (_01671_, _01670_, _01669_);
  and (_01672_, _01381_, _12125_);
  and (_01673_, _01375_, _11925_);
  or (_01674_, _01673_, _01672_);
  or (_01675_, _01674_, _01671_);
  or (_01676_, _01675_, _01668_);
  or (_01677_, _01676_, _01667_);
  and (_01678_, _01383_, _11465_);
  and (_01679_, _01370_, _12084_);
  and (_01680_, _01372_, _12040_);
  or (_01681_, _01680_, _01679_);
  and (_01682_, _01377_, _11982_);
  or (_01683_, _01682_, _01681_);
  or (_01684_, _01683_, _01678_);
  and (_01685_, _01385_, _11383_);
  and (_01686_, _01365_, _11424_);
  or (_01687_, _01686_, _01685_);
  or (_01688_, _01687_, _01684_);
  or (_01689_, _01688_, _01677_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [30], _01689_, _01664_);
  and (_01690_, _01385_, _12054_);
  and (_01691_, _01370_, _11941_);
  and (_01692_, _01372_, _11884_);
  or (_01693_, _01692_, _01691_);
  or (_01694_, _01693_, _01690_);
  and (_01695_, _01365_, _12095_);
  and (_01696_, _01341_, _11656_);
  or (_01697_, _01696_, _01695_);
  or (_01698_, _01697_, _01694_);
  and (_01699_, _01357_, _11517_);
  and (_01700_, _01355_, _11476_);
  or (_01701_, _01700_, _01699_);
  and (_01702_, _01348_, _11558_);
  or (_01703_, _01702_, _01701_);
  and (_01704_, _01352_, _11394_);
  and (_01705_, _01345_, _11603_);
  or (_01706_, _01705_, _01704_);
  or (_01707_, _01706_, _01703_);
  or (_01708_, _01707_, _01698_);
  and (_01709_, _01381_, _11998_);
  and (_01710_, _01361_, _11435_);
  and (_01711_, _01383_, _11353_);
  or (_01712_, _01711_, _01710_);
  and (_01713_, _01337_, _11713_);
  and (_01714_, _01375_, _11770_);
  and (_01715_, _01377_, _11827_);
  or (_01716_, _01715_, _01714_);
  or (_01717_, _01716_, _01713_);
  or (_01718_, _01717_, _01712_);
  or (_01719_, _01718_, _01709_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [8], _01719_, _01708_);
  and (_01720_, _01365_, _12100_);
  and (_01721_, _01385_, _12059_);
  and (_01722_, _01341_, _11663_);
  or (_01723_, _01722_, _01721_);
  or (_01724_, _01723_, _01720_);
  and (_01725_, _01355_, _11481_);
  and (_01726_, _01375_, _11777_);
  and (_01727_, _01348_, _11563_);
  or (_01728_, _01727_, _01726_);
  and (_01729_, _01381_, _12005_);
  and (_01730_, _01352_, _11399_);
  or (_01731_, _01730_, _01729_);
  or (_01732_, _01731_, _01728_);
  or (_01733_, _01732_, _01725_);
  and (_01734_, _01361_, _11440_);
  and (_01735_, _01357_, _11522_);
  or (_01736_, _01735_, _01734_);
  or (_01737_, _01736_, _01733_);
  and (_01738_, _01337_, _11719_);
  and (_01739_, _01372_, _11890_);
  and (_01740_, _01370_, _11947_);
  and (_01741_, _01377_, _11833_);
  or (_01742_, _01741_, _01740_);
  or (_01743_, _01742_, _01739_);
  or (_01744_, _01743_, _01738_);
  and (_01745_, _01383_, _11358_);
  and (_01746_, _01345_, _11609_);
  or (_01747_, _01746_, _01745_);
  or (_01748_, _01747_, _01744_);
  or (_01749_, _01748_, _01737_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [9], _01749_, _01724_);
  and (_01750_, _01372_, _11897_);
  and (_01751_, _01370_, _11954_);
  or (_01752_, _01751_, _01750_);
  and (_01753_, _01385_, _12064_);
  or (_01754_, _01753_, _01752_);
  and (_01755_, _01341_, _11670_);
  and (_01756_, _01365_, _12105_);
  or (_01757_, _01756_, _01755_);
  or (_01758_, _01757_, _01754_);
  and (_01759_, _01348_, _11568_);
  and (_01760_, _01355_, _11486_);
  and (_01761_, _01357_, _11527_);
  or (_01762_, _01761_, _01760_);
  or (_01763_, _01762_, _01759_);
  and (_01764_, _01352_, _11404_);
  and (_01765_, _01345_, _11615_);
  or (_01766_, _01765_, _01764_);
  or (_01767_, _01766_, _01763_);
  or (_01768_, _01767_, _01758_);
  and (_01769_, _01381_, _12012_);
  and (_01770_, _01383_, _11363_);
  and (_01771_, _01361_, _11445_);
  or (_01772_, _01771_, _01770_);
  and (_01773_, _01337_, _11726_);
  and (_01774_, _01375_, _11784_);
  and (_01775_, _01377_, _11840_);
  or (_01776_, _01775_, _01774_);
  or (_01777_, _01776_, _01773_);
  or (_01778_, _01777_, _01772_);
  or (_01779_, _01778_, _01769_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [10], _01779_, _01768_);
  and (_01780_, _01372_, _11904_);
  and (_01781_, _01370_, _11961_);
  or (_01782_, _01781_, _01780_);
  and (_01783_, _01385_, _12069_);
  or (_01784_, _01783_, _01782_);
  and (_01785_, _01337_, _11733_);
  and (_01786_, _01365_, _12110_);
  or (_01787_, _01786_, _01785_);
  or (_01788_, _01787_, _01784_);
  and (_01789_, _01348_, _11573_);
  and (_01790_, _01355_, _11491_);
  and (_01791_, _01357_, _11532_);
  or (_01792_, _01791_, _01790_);
  or (_01793_, _01792_, _01789_);
  and (_01794_, _01352_, _11409_);
  and (_01795_, _01345_, _11622_);
  or (_01796_, _01795_, _01794_);
  or (_01797_, _01796_, _01793_);
  or (_01798_, _01797_, _01788_);
  and (_01799_, _01381_, _12019_);
  and (_01800_, _01383_, _11368_);
  and (_01801_, _01361_, _11450_);
  or (_01802_, _01801_, _01800_);
  and (_01803_, _01341_, _11677_);
  and (_01804_, _01375_, _11791_);
  and (_01805_, _01377_, _11847_);
  or (_01806_, _01805_, _01804_);
  or (_01807_, _01806_, _01803_);
  or (_01808_, _01807_, _01802_);
  or (_01809_, _01808_, _01799_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [11], _01809_, _01798_);
  and (_01810_, _01341_, _11684_);
  and (_01811_, _01365_, _12115_);
  and (_01812_, _01383_, _11373_);
  or (_01813_, _01812_, _01811_);
  or (_01814_, _01813_, _01810_);
  and (_01815_, _01357_, _11537_);
  and (_01816_, _01375_, _11798_);
  and (_01817_, _01381_, _12026_);
  or (_01818_, _01817_, _01816_);
  and (_01819_, _01348_, _11578_);
  and (_01820_, _01352_, _11414_);
  or (_01821_, _01820_, _01819_);
  or (_01822_, _01821_, _01818_);
  or (_01823_, _01822_, _01815_);
  and (_01824_, _01355_, _11496_);
  and (_01825_, _01361_, _11455_);
  or (_01826_, _01825_, _01824_);
  or (_01827_, _01826_, _01823_);
  and (_01828_, _01337_, _11741_);
  and (_01829_, _01377_, _11854_);
  and (_01830_, _01370_, _11969_);
  and (_01831_, _01372_, _11912_);
  or (_01832_, _01831_, _01830_);
  or (_01833_, _01832_, _01829_);
  or (_01834_, _01833_, _01828_);
  and (_01835_, _01385_, _12074_);
  and (_01836_, _01345_, _11628_);
  or (_01837_, _01836_, _01835_);
  or (_01838_, _01837_, _01834_);
  or (_01839_, _01838_, _01827_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [12], _01839_, _01814_);
  and (_01840_, _01385_, _12079_);
  and (_01841_, _01370_, _11975_);
  and (_01842_, _01372_, _11918_);
  or (_01843_, _01842_, _01841_);
  or (_01844_, _01843_, _01840_);
  and (_01845_, _01365_, _12120_);
  and (_01846_, _01337_, _11747_);
  or (_01847_, _01846_, _01845_);
  or (_01848_, _01847_, _01844_);
  and (_01849_, _01357_, _11542_);
  and (_01850_, _01355_, _11501_);
  or (_01851_, _01850_, _01849_);
  and (_01852_, _01348_, _11583_);
  or (_01853_, _01852_, _01851_);
  and (_01854_, _01352_, _11419_);
  and (_01855_, _01345_, _11635_);
  or (_01856_, _01855_, _01854_);
  or (_01857_, _01856_, _01853_);
  or (_01858_, _01857_, _01848_);
  and (_01859_, _01381_, _12033_);
  and (_01860_, _01361_, _11460_);
  and (_01861_, _01383_, _11378_);
  or (_01862_, _01861_, _01860_);
  and (_01863_, _01341_, _11691_);
  and (_01864_, _01375_, _11805_);
  and (_01865_, _01377_, _11861_);
  or (_01866_, _01865_, _01864_);
  or (_01867_, _01866_, _01863_);
  or (_01868_, _01867_, _01862_);
  or (_01869_, _01868_, _01859_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [13], _01869_, _01858_);
  and (_01870_, _01337_, _11754_);
  and (_01871_, _01341_, _11698_);
  and (_01872_, _01385_, _12084_);
  or (_01873_, _01872_, _01871_);
  or (_01874_, _01873_, _01870_);
  and (_01875_, _01355_, _11506_);
  and (_01876_, _01375_, _11812_);
  and (_01877_, _01348_, _11589_);
  or (_01878_, _01877_, _01876_);
  and (_01879_, _01381_, _12040_);
  and (_01880_, _01352_, _11424_);
  or (_01881_, _01880_, _01879_);
  or (_01882_, _01881_, _01878_);
  or (_01883_, _01882_, _01875_);
  and (_01884_, _01361_, _11465_);
  and (_01885_, _01357_, _11547_);
  or (_01886_, _01885_, _01884_);
  or (_01887_, _01886_, _01883_);
  and (_01888_, _01365_, _12125_);
  and (_01889_, _01377_, _11868_);
  and (_01890_, _01370_, _11982_);
  and (_01891_, _01372_, _11925_);
  or (_01892_, _01891_, _01890_);
  or (_01893_, _01892_, _01889_);
  or (_01894_, _01893_, _01888_);
  and (_01895_, _01383_, _11383_);
  and (_01896_, _01345_, _11642_);
  or (_01897_, _01896_, _01895_);
  or (_01898_, _01897_, _01894_);
  or (_01899_, _01898_, _01887_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [14], _01899_, _01874_);
  and (_01900_, _01341_, _11713_);
  and (_01901_, _01365_, _11353_);
  and (_01902_, _01345_, _11656_);
  or (_01903_, _01902_, _01901_);
  or (_01904_, _01903_, _01900_);
  and (_01905_, _01355_, _11517_);
  and (_01906_, _01348_, _11603_);
  and (_01907_, _01381_, _12054_);
  or (_01908_, _01907_, _01906_);
  and (_01909_, _01352_, _11435_);
  and (_01910_, _01375_, _11827_);
  or (_01911_, _01910_, _01909_);
  or (_01912_, _01911_, _01908_);
  or (_01913_, _01912_, _01905_);
  and (_01914_, _01357_, _11558_);
  and (_01915_, _01361_, _11476_);
  or (_01916_, _01915_, _01914_);
  or (_01917_, _01916_, _01913_);
  and (_01918_, _01337_, _11770_);
  and (_01919_, _01370_, _11998_);
  and (_01920_, _01372_, _11941_);
  and (_01921_, _01377_, _11884_);
  or (_01922_, _01921_, _01920_);
  or (_01923_, _01922_, _01919_);
  or (_01924_, _01923_, _01918_);
  and (_01925_, _01385_, _12095_);
  and (_01926_, _01383_, _11394_);
  or (_01927_, _01926_, _01925_);
  or (_01928_, _01927_, _01924_);
  or (_01929_, _01928_, _01917_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [16], _01929_, _01904_);
  and (_01930_, _01385_, _12100_);
  and (_01931_, _01365_, _11358_);
  and (_01932_, _01341_, _11719_);
  or (_01933_, _01932_, _01931_);
  or (_01934_, _01933_, _01930_);
  and (_01935_, _01355_, _11522_);
  and (_01936_, _01348_, _11609_);
  and (_01937_, _01381_, _12059_);
  or (_01938_, _01937_, _01936_);
  and (_01939_, _01352_, _11440_);
  and (_01940_, _01375_, _11833_);
  or (_01941_, _01940_, _01939_);
  or (_01942_, _01941_, _01938_);
  or (_01943_, _01942_, _01935_);
  and (_01944_, _01357_, _11563_);
  and (_01945_, _01361_, _11481_);
  or (_01946_, _01945_, _01944_);
  or (_01947_, _01946_, _01943_);
  and (_01948_, _01337_, _11777_);
  and (_01949_, _01370_, _12005_);
  and (_01950_, _01372_, _11947_);
  and (_01951_, _01377_, _11890_);
  or (_01952_, _01951_, _01950_);
  or (_01953_, _01952_, _01949_);
  or (_01954_, _01953_, _01948_);
  and (_01955_, _01383_, _11399_);
  and (_01956_, _01345_, _11663_);
  or (_01957_, _01956_, _01955_);
  or (_01958_, _01957_, _01954_);
  or (_01959_, _01958_, _01947_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [17], _01959_, _01934_);
  and (_01960_, _01385_, _12105_);
  and (_01961_, _01337_, _11784_);
  and (_01962_, _01345_, _11670_);
  or (_01963_, _01962_, _01961_);
  or (_01964_, _01963_, _01960_);
  and (_01965_, _01355_, _11527_);
  and (_01966_, _01375_, _11840_);
  and (_01967_, _01348_, _11615_);
  or (_01968_, _01967_, _01966_);
  and (_01969_, _01381_, _12064_);
  and (_01970_, _01352_, _11445_);
  or (_01971_, _01970_, _01969_);
  or (_01972_, _01971_, _01968_);
  or (_01973_, _01972_, _01965_);
  and (_01974_, _01357_, _11568_);
  and (_01975_, _01361_, _11486_);
  or (_01976_, _01975_, _01974_);
  or (_01977_, _01976_, _01973_);
  and (_01978_, _01365_, _11363_);
  and (_01979_, _01370_, _12012_);
  and (_01980_, _01377_, _11897_);
  and (_01981_, _01372_, _11954_);
  or (_01982_, _01981_, _01980_);
  or (_01983_, _01982_, _01979_);
  or (_01984_, _01983_, _01978_);
  and (_01985_, _01341_, _11726_);
  and (_01986_, _01383_, _11404_);
  or (_01987_, _01986_, _01985_);
  or (_01988_, _01987_, _01984_);
  or (_01989_, _01988_, _01977_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [18], _01989_, _01964_);
  and (_01990_, _01370_, _12019_);
  and (_01991_, _01377_, _11904_);
  and (_01992_, _01372_, _11961_);
  or (_01993_, _01992_, _01991_);
  or (_01994_, _01993_, _01990_);
  and (_01995_, _01385_, _12110_);
  and (_01996_, _01341_, _11733_);
  or (_01997_, _01996_, _01995_);
  or (_01998_, _01997_, _01994_);
  and (_01999_, _01361_, _11491_);
  and (_02000_, _01348_, _11622_);
  and (_02001_, _01357_, _11573_);
  or (_02002_, _02001_, _02000_);
  or (_02003_, _02002_, _01999_);
  and (_02004_, _01383_, _11409_);
  and (_02005_, _01355_, _11532_);
  or (_02006_, _02005_, _02004_);
  or (_02007_, _02006_, _02003_);
  or (_02008_, _02007_, _01998_);
  and (_02009_, _01345_, _11677_);
  and (_02010_, _01337_, _11791_);
  and (_02011_, _01375_, _11847_);
  or (_02012_, _02011_, _02010_);
  or (_02013_, _02012_, _02009_);
  and (_02014_, _01381_, _12069_);
  and (_02015_, _01352_, _11450_);
  and (_02016_, _01365_, _11368_);
  or (_02017_, _02016_, _02015_);
  or (_02018_, _02017_, _02014_);
  or (_02019_, _02018_, _02013_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [19], _02019_, _02008_);
  and (_02020_, _01383_, _11414_);
  and (_02021_, _01365_, _11373_);
  and (_02022_, _01337_, _11798_);
  or (_02023_, _02022_, _02021_);
  or (_02024_, _02023_, _02020_);
  and (_02025_, _01355_, _11537_);
  and (_02026_, _01348_, _11628_);
  and (_02027_, _01381_, _12074_);
  or (_02028_, _02027_, _02026_);
  and (_02029_, _01352_, _11455_);
  and (_02030_, _01375_, _11854_);
  or (_02031_, _02030_, _02029_);
  or (_02032_, _02031_, _02028_);
  or (_02033_, _02032_, _02025_);
  and (_02034_, _01357_, _11578_);
  and (_02035_, _01361_, _11496_);
  or (_02036_, _02035_, _02034_);
  or (_02037_, _02036_, _02033_);
  and (_02038_, _01341_, _11741_);
  and (_02039_, _01370_, _12026_);
  and (_02040_, _01372_, _11969_);
  and (_02041_, _01377_, _11912_);
  or (_02042_, _02041_, _02040_);
  or (_02043_, _02042_, _02039_);
  or (_02044_, _02043_, _02038_);
  and (_02045_, _01385_, _12115_);
  and (_02046_, _01345_, _11684_);
  or (_02047_, _02046_, _02045_);
  or (_02048_, _02047_, _02044_);
  or (_02049_, _02048_, _02037_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [20], _02049_, _02024_);
  and (_02050_, _01337_, _11805_);
  and (_02051_, _01385_, _12120_);
  and (_02052_, _01365_, _11378_);
  or (_02053_, _02052_, _02051_);
  or (_02054_, _02053_, _02050_);
  and (_02055_, _01355_, _11542_);
  and (_02056_, _01348_, _11635_);
  and (_02057_, _01352_, _11460_);
  or (_02058_, _02057_, _02056_);
  and (_02059_, _01381_, _12079_);
  and (_02060_, _01375_, _11861_);
  or (_02061_, _02060_, _02059_);
  or (_02062_, _02061_, _02058_);
  or (_02063_, _02062_, _02055_);
  and (_02064_, _01357_, _11583_);
  and (_02065_, _01361_, _11501_);
  or (_02066_, _02065_, _02064_);
  or (_02067_, _02066_, _02063_);
  and (_02068_, _01345_, _11691_);
  and (_02069_, _01370_, _12033_);
  and (_02070_, _01372_, _11975_);
  and (_02071_, _01377_, _11918_);
  or (_02072_, _02071_, _02070_);
  or (_02073_, _02072_, _02069_);
  or (_02074_, _02073_, _02068_);
  and (_02075_, _01383_, _11419_);
  and (_02076_, _01341_, _11747_);
  or (_02077_, _02076_, _02075_);
  or (_02078_, _02077_, _02074_);
  or (_02079_, _02078_, _02067_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [21], _02079_, _02054_);
  and (_02080_, _01337_, _11812_);
  and (_02081_, _01365_, _11383_);
  and (_02082_, _01341_, _11754_);
  or (_02083_, _02082_, _02081_);
  or (_02084_, _02083_, _02080_);
  and (_02085_, _01355_, _11547_);
  and (_02086_, _01348_, _11642_);
  and (_02087_, _01352_, _11465_);
  or (_02088_, _02087_, _02086_);
  and (_02089_, _01375_, _11868_);
  and (_02090_, _01381_, _12084_);
  or (_02091_, _02090_, _02089_);
  or (_02092_, _02091_, _02088_);
  or (_02093_, _02092_, _02085_);
  and (_02094_, _01357_, _11589_);
  and (_02095_, _01361_, _11506_);
  or (_02096_, _02095_, _02094_);
  or (_02097_, _02096_, _02093_);
  and (_02098_, _01345_, _11698_);
  and (_02099_, _01370_, _12040_);
  and (_02100_, _01372_, _11982_);
  and (_02101_, _01377_, _11925_);
  or (_02102_, _02101_, _02100_);
  or (_02103_, _02102_, _02099_);
  or (_02104_, _02103_, _02098_);
  and (_02105_, _01385_, _12125_);
  and (_02106_, _01383_, _11424_);
  or (_02107_, _02106_, _02105_);
  or (_02108_, _02107_, _02104_);
  or (_02109_, _02108_, _02097_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [22], _02109_, _02084_);
  and (_02110_, _01345_, _11558_);
  and (_02111_, _01337_, _11656_);
  and (_02112_, _01385_, _11998_);
  or (_02113_, _02112_, _02111_);
  or (_02114_, _02113_, _02110_);
  and (_02115_, _01355_, _11435_);
  and (_02116_, _01361_, _11394_);
  or (_02117_, _02116_, _02115_);
  and (_02118_, _01357_, _11476_);
  and (_02119_, _01352_, _11353_);
  and (_02120_, _01348_, _11517_);
  or (_02121_, _02120_, _02119_);
  and (_02122_, _01375_, _11713_);
  and (_02123_, _01381_, _11941_);
  or (_02124_, _02123_, _02122_);
  or (_02125_, _02124_, _02121_);
  or (_02126_, _02125_, _02118_);
  or (_02127_, _02126_, _02117_);
  and (_02128_, _01383_, _12095_);
  and (_02129_, _01377_, _11770_);
  and (_02130_, _01372_, _11827_);
  and (_02131_, _01370_, _11884_);
  or (_02132_, _02131_, _02130_);
  or (_02133_, _02132_, _02129_);
  or (_02134_, _02133_, _02128_);
  and (_02135_, _01341_, _11603_);
  and (_02136_, _01365_, _12054_);
  or (_02137_, _02136_, _02135_);
  or (_02138_, _02137_, _02134_);
  or (_02139_, _02138_, _02127_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [0], _02139_, _02114_);
  and (_02140_, _01385_, _12005_);
  and (_02141_, _01383_, _12100_);
  and (_02142_, _01345_, _11563_);
  or (_02143_, _02142_, _02141_);
  or (_02144_, _02143_, _02140_);
  and (_02145_, _01361_, _11399_);
  and (_02146_, _01348_, _11522_);
  and (_02147_, _01381_, _11947_);
  or (_02148_, _02147_, _02146_);
  and (_02149_, _01352_, _11358_);
  and (_02150_, _01375_, _11719_);
  or (_02151_, _02150_, _02149_);
  or (_02152_, _02151_, _02148_);
  or (_02153_, _02152_, _02145_);
  and (_02154_, _01355_, _11440_);
  and (_02155_, _01357_, _11481_);
  or (_02156_, _02155_, _02154_);
  or (_02157_, _02156_, _02153_);
  and (_02158_, _01337_, _11663_);
  and (_02159_, _01377_, _11777_);
  and (_02160_, _01372_, _11833_);
  and (_02161_, _01370_, _11890_);
  or (_02162_, _02161_, _02160_);
  or (_02163_, _02162_, _02159_);
  or (_02164_, _02163_, _02158_);
  and (_02165_, _01341_, _11609_);
  and (_02166_, _01365_, _12059_);
  or (_02167_, _02166_, _02165_);
  or (_02168_, _02167_, _02164_);
  or (_02169_, _02168_, _02157_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [1], _02169_, _02144_);
  and (_02170_, _01337_, _11670_);
  and (_02171_, _01345_, _11568_);
  and (_02172_, _01385_, _12012_);
  or (_02173_, _02172_, _02171_);
  or (_02174_, _02173_, _02170_);
  and (_02175_, _01361_, _11404_);
  and (_02176_, _01355_, _11445_);
  or (_02177_, _02176_, _02175_);
  and (_02178_, _01357_, _11486_);
  and (_02179_, _01352_, _11363_);
  and (_02180_, _01348_, _11527_);
  or (_02181_, _02180_, _02179_);
  and (_02182_, _01375_, _11726_);
  and (_02183_, _01381_, _11954_);
  or (_02184_, _02183_, _02182_);
  or (_02185_, _02184_, _02181_);
  or (_02186_, _02185_, _02178_);
  or (_02187_, _02186_, _02177_);
  and (_02188_, _01383_, _12105_);
  and (_02189_, _01372_, _11840_);
  and (_02190_, _01377_, _11784_);
  or (_02191_, _02190_, _02189_);
  and (_02192_, _01370_, _11897_);
  or (_02193_, _02192_, _02191_);
  or (_02194_, _02193_, _02188_);
  and (_02195_, _01341_, _11615_);
  and (_02196_, _01365_, _12064_);
  or (_02197_, _02196_, _02195_);
  or (_02198_, _02197_, _02194_);
  or (_02199_, _02198_, _02187_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [2], _02199_, _02174_);
  and (_02200_, _01383_, _12110_);
  and (_02201_, _01337_, _11677_);
  and (_02202_, _01345_, _11573_);
  or (_02203_, _02202_, _02201_);
  or (_02204_, _02203_, _02200_);
  and (_02205_, _01355_, _11450_);
  and (_02206_, _01352_, _11368_);
  and (_02207_, _01348_, _11532_);
  or (_02208_, _02207_, _02206_);
  and (_02209_, _01381_, _11961_);
  and (_02210_, _01375_, _11733_);
  or (_02211_, _02210_, _02209_);
  or (_02212_, _02211_, _02208_);
  or (_02213_, _02212_, _02205_);
  and (_02214_, _01361_, _11409_);
  and (_02215_, _01357_, _11491_);
  or (_02216_, _02215_, _02214_);
  or (_02217_, _02216_, _02213_);
  and (_02218_, _01365_, _12069_);
  and (_02219_, _01372_, _11847_);
  and (_02220_, _01370_, _11904_);
  and (_02221_, _01377_, _11791_);
  or (_02222_, _02221_, _02220_);
  or (_02223_, _02222_, _02219_);
  or (_02224_, _02223_, _02218_);
  and (_02225_, _01385_, _12019_);
  and (_02226_, _01341_, _11622_);
  or (_02227_, _02226_, _02225_);
  or (_02228_, _02227_, _02224_);
  or (_02229_, _02228_, _02217_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [3], _02229_, _02204_);
  and (_02230_, _01385_, _12026_);
  and (_02231_, _01383_, _12115_);
  and (_02232_, _01345_, _11578_);
  or (_02233_, _02232_, _02231_);
  or (_02234_, _02233_, _02230_);
  and (_02235_, _01361_, _11414_);
  and (_02236_, _01348_, _11537_);
  and (_02237_, _01381_, _11969_);
  or (_02238_, _02237_, _02236_);
  and (_02239_, _01352_, _11373_);
  and (_02240_, _01375_, _11741_);
  or (_02241_, _02240_, _02239_);
  or (_02242_, _02241_, _02238_);
  or (_02243_, _02242_, _02235_);
  and (_02244_, _01355_, _11455_);
  and (_02245_, _01357_, _11496_);
  or (_02246_, _02245_, _02244_);
  or (_02247_, _02246_, _02243_);
  and (_02248_, _01337_, _11684_);
  and (_02249_, _01377_, _11798_);
  and (_02250_, _01372_, _11854_);
  and (_02251_, _01370_, _11912_);
  or (_02252_, _02251_, _02250_);
  or (_02253_, _02252_, _02249_);
  or (_02254_, _02253_, _02248_);
  and (_02255_, _01341_, _11628_);
  and (_02256_, _01365_, _12074_);
  or (_02257_, _02256_, _02255_);
  or (_02258_, _02257_, _02254_);
  or (_02259_, _02258_, _02247_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [4], _02259_, _02234_);
  and (_02260_, _01337_, _11691_);
  and (_02261_, _01383_, _12120_);
  and (_02262_, _01345_, _11583_);
  or (_02263_, _02262_, _02261_);
  or (_02264_, _02263_, _02260_);
  and (_02265_, _01355_, _11460_);
  and (_02266_, _01375_, _11747_);
  and (_02267_, _01348_, _11542_);
  or (_02268_, _02267_, _02266_);
  and (_02269_, _01381_, _11975_);
  and (_02270_, _01352_, _11378_);
  or (_02271_, _02270_, _02269_);
  or (_02272_, _02271_, _02268_);
  or (_02273_, _02272_, _02265_);
  and (_02274_, _01361_, _11419_);
  and (_02275_, _01357_, _11501_);
  or (_02276_, _02275_, _02274_);
  or (_02277_, _02276_, _02273_);
  and (_02278_, _01365_, _12079_);
  and (_02279_, _01372_, _11861_);
  and (_02280_, _01370_, _11918_);
  and (_02281_, _01377_, _11805_);
  or (_02282_, _02281_, _02280_);
  or (_02283_, _02282_, _02279_);
  or (_02284_, _02283_, _02278_);
  and (_02285_, _01385_, _12033_);
  and (_02286_, _01341_, _11635_);
  or (_02287_, _02286_, _02285_);
  or (_02288_, _02287_, _02284_);
  or (_02289_, _02288_, _02277_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [5], _02289_, _02264_);
  and (_02290_, _01385_, _12040_);
  and (_02291_, _01383_, _12125_);
  and (_02292_, _01345_, _11589_);
  or (_02293_, _02292_, _02291_);
  or (_02294_, _02293_, _02290_);
  and (_02295_, _01355_, _11465_);
  and (_02296_, _01352_, _11383_);
  and (_02297_, _01375_, _11754_);
  or (_02298_, _02297_, _02296_);
  and (_02299_, _01348_, _11547_);
  and (_02300_, _01381_, _11982_);
  or (_02301_, _02300_, _02299_);
  or (_02302_, _02301_, _02298_);
  or (_02303_, _02302_, _02295_);
  and (_02304_, _01361_, _11424_);
  and (_02305_, _01357_, _11506_);
  or (_02306_, _02305_, _02304_);
  or (_02307_, _02306_, _02303_);
  and (_02308_, _01365_, _12084_);
  and (_02309_, _01372_, _11868_);
  and (_02310_, _01377_, _11812_);
  and (_02311_, _01370_, _11925_);
  or (_02312_, _02311_, _02310_);
  or (_02313_, _02312_, _02309_);
  or (_02314_, _02313_, _02308_);
  and (_02315_, _01341_, _11642_);
  and (_02316_, _01337_, _11698_);
  or (_02317_, _02316_, _02315_);
  or (_02318_, _02317_, _02314_);
  or (_02319_, _02318_, _02307_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [6], _02319_, _02294_);
  not (_02320_, _11363_);
  or (_02321_, \oc8051_golden_model_1.PC [1], \oc8051_golden_model_1.PC [0]);
  or (_02322_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [3]);
  or (_02323_, _02322_, _02321_);
  or (_02324_, _02323_, _02320_);
  not (_02325_, _11445_);
  not (_02326_, \oc8051_golden_model_1.PC [0]);
  nand (_02327_, \oc8051_golden_model_1.PC [1], _02326_);
  or (_02328_, _02327_, _02322_);
  or (_02329_, _02328_, _02325_);
  and (_02330_, _02329_, _02324_);
  not (_02331_, _12064_);
  and (_02332_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [3]);
  not (_02333_, _02332_);
  or (_02334_, _02333_, _02327_);
  or (_02335_, _02334_, _02331_);
  not (_02336_, _11954_);
  or (_02337_, _02333_, _02321_);
  or (_02338_, _02337_, _02336_);
  and (_02339_, _02338_, _02335_);
  and (_02340_, _02339_, _02330_);
  not (_02341_, _11568_);
  not (_02342_, \oc8051_golden_model_1.PC [3]);
  and (_02343_, \oc8051_golden_model_1.PC [2], _02342_);
  not (_02344_, _02343_);
  or (_02345_, \oc8051_golden_model_1.PC [1], _02326_);
  or (_02346_, _02345_, _02344_);
  or (_02347_, _02346_, _02341_);
  not (_02348_, _11615_);
  or (_02349_, _02344_, _02327_);
  or (_02350_, _02349_, _02348_);
  and (_02351_, _02350_, _02347_);
  not (_02352_, _11897_);
  and (_02353_, \oc8051_golden_model_1.PC [1], \oc8051_golden_model_1.PC [0]);
  not (_02354_, _02353_);
  or (_02355_, \oc8051_golden_model_1.PC [2], _02342_);
  or (_02356_, _02355_, _02354_);
  or (_02357_, _02356_, _02352_);
  not (_02358_, _11726_);
  or (_02359_, _02355_, _02321_);
  or (_02360_, _02359_, _02358_);
  and (_02361_, _02360_, _02357_);
  and (_02362_, _02361_, _02351_);
  and (_02363_, _02362_, _02340_);
  not (_02364_, _11486_);
  or (_02365_, _02354_, _02322_);
  or (_02366_, _02365_, _02364_);
  not (_02367_, _11404_);
  or (_02368_, _02345_, _02322_);
  or (_02369_, _02368_, _02367_);
  and (_02370_, _02369_, _02366_);
  not (_02371_, _11840_);
  or (_02372_, _02355_, _02327_);
  or (_02373_, _02372_, _02371_);
  and (_02374_, _02353_, _02343_);
  nand (_02375_, _02374_, _11670_);
  and (_02376_, _02375_, _02373_);
  and (_02377_, _02376_, _02370_);
  and (_02378_, _02353_, _02332_);
  nand (_02379_, _02378_, _12105_);
  not (_02380_, _12012_);
  or (_02381_, _02345_, _02333_);
  or (_02382_, _02381_, _02380_);
  and (_02383_, _02382_, _02379_);
  not (_02384_, _11784_);
  or (_02385_, _02355_, _02345_);
  or (_02386_, _02385_, _02384_);
  not (_02387_, _11527_);
  or (_02388_, _02344_, _02321_);
  or (_02389_, _02388_, _02387_);
  and (_02390_, _02389_, _02386_);
  and (_02391_, _02390_, _02383_);
  and (_02392_, _02391_, _02377_);
  nand (_02393_, _02392_, _02363_);
  not (_02394_, _11961_);
  or (_02395_, _02337_, _02394_);
  not (_02396_, _11733_);
  or (_02397_, _02359_, _02396_);
  and (_02398_, _02397_, _02395_);
  not (_02399_, _11904_);
  or (_02400_, _02356_, _02399_);
  not (_02401_, _11532_);
  or (_02402_, _02388_, _02401_);
  and (_02403_, _02402_, _02400_);
  and (_02404_, _02403_, _02398_);
  not (_02405_, _11847_);
  or (_02406_, _02372_, _02405_);
  not (_02407_, _11409_);
  or (_02408_, _02368_, _02407_);
  and (_02409_, _02408_, _02406_);
  not (_02410_, _12019_);
  or (_02411_, _02381_, _02410_);
  not (_02412_, _11791_);
  or (_02413_, _02385_, _02412_);
  and (_02414_, _02413_, _02411_);
  and (_02415_, _02414_, _02409_);
  and (_02416_, _02415_, _02404_);
  not (_02417_, _12069_);
  or (_02418_, _02334_, _02417_);
  not (_02419_, _11491_);
  or (_02420_, _02365_, _02419_);
  and (_02421_, _02420_, _02418_);
  nand (_02422_, _02378_, _12110_);
  nand (_02423_, _02374_, _11677_);
  and (_02424_, _02423_, _02422_);
  and (_02425_, _02424_, _02421_);
  not (_02426_, _11573_);
  or (_02427_, _02346_, _02426_);
  not (_02428_, _11450_);
  or (_02429_, _02328_, _02428_);
  and (_02430_, _02429_, _02427_);
  not (_02431_, _11622_);
  or (_02432_, _02349_, _02431_);
  not (_02433_, _11368_);
  or (_02434_, _02323_, _02433_);
  and (_02435_, _02434_, _02432_);
  and (_02436_, _02435_, _02430_);
  and (_02437_, _02436_, _02425_);
  and (_02438_, _02437_, _02416_);
  and (_02439_, _02438_, _02393_);
  not (_02440_, _11941_);
  or (_02441_, _02337_, _02440_);
  not (_02442_, _11713_);
  or (_02443_, _02359_, _02442_);
  and (_02444_, _02443_, _02441_);
  not (_02445_, _11884_);
  or (_02446_, _02356_, _02445_);
  not (_02447_, _11394_);
  or (_02448_, _02368_, _02447_);
  and (_02449_, _02448_, _02446_);
  and (_02450_, _02449_, _02444_);
  not (_02451_, _11827_);
  or (_02452_, _02372_, _02451_);
  not (_02453_, _11353_);
  or (_02454_, _02323_, _02453_);
  and (_02455_, _02454_, _02452_);
  not (_02456_, _11998_);
  or (_02457_, _02381_, _02456_);
  not (_02458_, _11770_);
  or (_02459_, _02385_, _02458_);
  and (_02460_, _02459_, _02457_);
  and (_02461_, _02460_, _02455_);
  and (_02462_, _02461_, _02450_);
  not (_02463_, _12054_);
  or (_02464_, _02334_, _02463_);
  not (_02465_, _11558_);
  or (_02466_, _02346_, _02465_);
  and (_02467_, _02466_, _02464_);
  nand (_02468_, _02378_, _12095_);
  not (_02469_, _11603_);
  or (_02470_, _02349_, _02469_);
  and (_02471_, _02470_, _02468_);
  and (_02472_, _02471_, _02467_);
  not (_02473_, _11517_);
  or (_02474_, _02388_, _02473_);
  not (_02475_, _11435_);
  or (_02476_, _02328_, _02475_);
  and (_02477_, _02476_, _02474_);
  nand (_02478_, _02374_, _11656_);
  not (_02479_, _11476_);
  or (_02480_, _02365_, _02479_);
  and (_02481_, _02480_, _02478_);
  and (_02482_, _02481_, _02477_);
  and (_02483_, _02482_, _02472_);
  nand (_02484_, _02483_, _02462_);
  not (_02485_, _11522_);
  or (_02486_, _02388_, _02485_);
  not (_02487_, _11358_);
  or (_02488_, _02323_, _02487_);
  and (_02489_, _02488_, _02486_);
  not (_02490_, _11719_);
  or (_02491_, _02359_, _02490_);
  not (_02492_, _11481_);
  or (_02493_, _02365_, _02492_);
  and (_02494_, _02493_, _02491_);
  and (_02495_, _02494_, _02489_);
  not (_02496_, _11609_);
  or (_02497_, _02349_, _02496_);
  not (_02498_, _11440_);
  or (_02499_, _02328_, _02498_);
  and (_02500_, _02499_, _02497_);
  not (_02501_, _11563_);
  or (_02502_, _02346_, _02501_);
  not (_02503_, _11399_);
  or (_02504_, _02368_, _02503_);
  and (_02505_, _02504_, _02502_);
  and (_02506_, _02505_, _02500_);
  and (_02507_, _02506_, _02495_);
  not (_02508_, _12005_);
  or (_02509_, _02381_, _02508_);
  not (_02510_, _12059_);
  or (_02511_, _02334_, _02510_);
  and (_02512_, _02511_, _02509_);
  not (_02513_, _11947_);
  or (_02514_, _02337_, _02513_);
  nand (_02515_, _02374_, _11663_);
  and (_02516_, _02515_, _02514_);
  and (_02517_, _02516_, _02512_);
  not (_02518_, _11890_);
  or (_02519_, _02356_, _02518_);
  not (_02520_, _11777_);
  or (_02521_, _02385_, _02520_);
  and (_02522_, _02521_, _02519_);
  nand (_02523_, _02378_, _12100_);
  not (_02524_, _11833_);
  or (_02525_, _02372_, _02524_);
  and (_02526_, _02525_, _02523_);
  and (_02527_, _02526_, _02522_);
  and (_02528_, _02527_, _02517_);
  and (_02529_, _02528_, _02507_);
  and (_02530_, _02529_, _02484_);
  and (_02531_, _02530_, _02439_);
  not (_02532_, _11496_);
  or (_02533_, _02365_, _02532_);
  not (_02534_, _11373_);
  or (_02535_, _02323_, _02534_);
  and (_02536_, _02535_, _02533_);
  not (_02537_, _12074_);
  or (_02538_, _02334_, _02537_);
  not (_02539_, _11969_);
  or (_02540_, _02337_, _02539_);
  and (_02541_, _02540_, _02538_);
  and (_02542_, _02541_, _02536_);
  not (_02543_, _11578_);
  or (_02544_, _02346_, _02543_);
  not (_02545_, _11628_);
  or (_02546_, _02349_, _02545_);
  and (_02547_, _02546_, _02544_);
  not (_02548_, _11912_);
  or (_02549_, _02356_, _02548_);
  not (_02550_, _11741_);
  or (_02551_, _02359_, _02550_);
  and (_02552_, _02551_, _02549_);
  and (_02553_, _02552_, _02547_);
  and (_02554_, _02553_, _02542_);
  not (_02555_, _11414_);
  or (_02556_, _02368_, _02555_);
  not (_02557_, _11455_);
  or (_02558_, _02328_, _02557_);
  and (_02559_, _02558_, _02556_);
  not (_02560_, _11854_);
  or (_02561_, _02372_, _02560_);
  nand (_02562_, _02374_, _11684_);
  and (_02563_, _02562_, _02561_);
  and (_02564_, _02563_, _02559_);
  nand (_02565_, _02378_, _12115_);
  not (_02566_, _12026_);
  or (_02567_, _02381_, _02566_);
  and (_02568_, _02567_, _02565_);
  not (_02569_, _11798_);
  or (_02570_, _02385_, _02569_);
  not (_02571_, _11537_);
  or (_02572_, _02388_, _02571_);
  and (_02573_, _02572_, _02570_);
  and (_02574_, _02573_, _02568_);
  and (_02575_, _02574_, _02564_);
  and (_02576_, _02575_, _02554_);
  not (_02577_, _11583_);
  or (_02578_, _02346_, _02577_);
  not (_02579_, _11501_);
  or (_02580_, _02365_, _02579_);
  and (_02581_, _02580_, _02578_);
  not (_02582_, _12079_);
  or (_02583_, _02334_, _02582_);
  not (_02584_, _11747_);
  or (_02585_, _02359_, _02584_);
  and (_02586_, _02585_, _02583_);
  and (_02587_, _02586_, _02581_);
  not (_02588_, _12033_);
  or (_02589_, _02381_, _02588_);
  not (_02590_, _11975_);
  or (_02591_, _02337_, _02590_);
  and (_02592_, _02591_, _02589_);
  not (_02593_, _11861_);
  or (_02594_, _02372_, _02593_);
  not (_02595_, _11419_);
  or (_02596_, _02368_, _02595_);
  and (_02597_, _02596_, _02594_);
  and (_02598_, _02597_, _02592_);
  and (_02599_, _02598_, _02587_);
  not (_02600_, _11635_);
  or (_02601_, _02349_, _02600_);
  not (_02602_, _11542_);
  or (_02603_, _02388_, _02602_);
  and (_02604_, _02603_, _02601_);
  nand (_02605_, _02374_, _11691_);
  not (_02606_, _11378_);
  or (_02607_, _02323_, _02606_);
  and (_02608_, _02607_, _02605_);
  and (_02609_, _02608_, _02604_);
  nand (_02610_, _02378_, _12120_);
  not (_02611_, _11918_);
  or (_02612_, _02356_, _02611_);
  and (_02613_, _02612_, _02610_);
  not (_02614_, _11805_);
  or (_02615_, _02385_, _02614_);
  not (_02616_, _11460_);
  or (_02617_, _02328_, _02616_);
  and (_02618_, _02617_, _02615_);
  and (_02619_, _02618_, _02613_);
  and (_02620_, _02619_, _02609_);
  and (_02621_, _02620_, _02599_);
  and (_02622_, _02621_, _02576_);
  not (_02623_, _11547_);
  or (_02624_, _02388_, _02623_);
  not (_02625_, _11383_);
  or (_02626_, _02323_, _02625_);
  and (_02627_, _02626_, _02624_);
  not (_02628_, _11754_);
  or (_02629_, _02359_, _02628_);
  not (_02630_, _11506_);
  or (_02631_, _02365_, _02630_);
  and (_02632_, _02631_, _02629_);
  and (_02633_, _02632_, _02627_);
  not (_02634_, _11642_);
  or (_02635_, _02349_, _02634_);
  not (_02636_, _11465_);
  or (_02637_, _02328_, _02636_);
  and (_02638_, _02637_, _02635_);
  not (_02639_, _11589_);
  or (_02640_, _02346_, _02639_);
  not (_02641_, _11424_);
  or (_02642_, _02368_, _02641_);
  and (_02643_, _02642_, _02640_);
  and (_02644_, _02643_, _02638_);
  and (_02645_, _02644_, _02633_);
  nand (_02646_, _02378_, _12125_);
  not (_02647_, _11925_);
  or (_02648_, _02356_, _02647_);
  and (_02649_, _02648_, _02646_);
  not (_02650_, _12084_);
  or (_02651_, _02334_, _02650_);
  nand (_02652_, _02374_, _11698_);
  and (_02653_, _02652_, _02651_);
  and (_02654_, _02653_, _02649_);
  not (_02655_, _11982_);
  or (_02656_, _02337_, _02655_);
  not (_02657_, _11868_);
  or (_02658_, _02372_, _02657_);
  and (_02659_, _02658_, _02656_);
  not (_02660_, _12040_);
  or (_02661_, _02381_, _02660_);
  not (_02662_, _11812_);
  or (_02663_, _02385_, _02662_);
  and (_02664_, _02663_, _02661_);
  and (_02665_, _02664_, _02659_);
  and (_02666_, _02665_, _02654_);
  and (_02667_, _02666_, _02645_);
  not (_02668_, _11706_);
  or (_02669_, _02359_, _02668_);
  not (_02670_, _11430_);
  or (_02671_, _02328_, _02670_);
  and (_02672_, _02671_, _02669_);
  not (_02673_, _11991_);
  or (_02674_, _02381_, _02673_);
  not (_02675_, _11876_);
  or (_02676_, _02356_, _02675_);
  and (_02677_, _02676_, _02674_);
  and (_02678_, _02677_, _02672_);
  not (_02679_, _11820_);
  or (_02680_, _02372_, _02679_);
  not (_02681_, _11348_);
  or (_02682_, _02323_, _02681_);
  and (_02683_, _02682_, _02680_);
  not (_02684_, _11763_);
  or (_02685_, _02385_, _02684_);
  not (_02686_, _11471_);
  or (_02687_, _02365_, _02686_);
  and (_02688_, _02687_, _02685_);
  and (_02689_, _02688_, _02683_);
  and (_02690_, _02689_, _02678_);
  nand (_02691_, _02378_, _12090_);
  not (_02692_, _11553_);
  or (_02693_, _02346_, _02692_);
  and (_02694_, _02693_, _02691_);
  not (_02695_, _12048_);
  or (_02696_, _02334_, _02695_);
  nand (_02697_, _02374_, _11651_);
  and (_02698_, _02697_, _02696_);
  and (_02699_, _02698_, _02694_);
  not (_02700_, _11934_);
  or (_02701_, _02337_, _02700_);
  not (_02702_, _11512_);
  or (_02703_, _02388_, _02702_);
  and (_02704_, _02703_, _02701_);
  not (_02705_, _11597_);
  or (_02706_, _02349_, _02705_);
  not (_02707_, _11389_);
  or (_02708_, _02368_, _02707_);
  and (_02709_, _02708_, _02706_);
  and (_02710_, _02709_, _02704_);
  and (_02711_, _02710_, _02699_);
  and (_02712_, _02711_, _02690_);
  and (_02713_, _02712_, _02667_);
  and (_02714_, _02713_, _02622_);
  nand (_02715_, _02714_, _02531_);
  and (_02716_, _02715_, XRAM_DATA_OUT_abstr[7]);
  or (_02717_, _02716_, _12786_);
  or (_02718_, _12782_, \oc8051_golden_model_1.XRAM_DATA_OUT [7]);
  and (_02719_, _02718_, _13707_);
  and (_13851_[7], _02719_, _02717_);
  and (_02720_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [1]);
  and (_02721_, _02720_, \oc8051_golden_model_1.PC [3]);
  and (_02722_, _02721_, \oc8051_golden_model_1.PC [4]);
  and (_02723_, _02722_, \oc8051_golden_model_1.PC [5]);
  and (_02724_, _02723_, \oc8051_golden_model_1.PC [6]);
  and (_02725_, _02724_, \oc8051_golden_model_1.PC [7]);
  and (_02726_, _02725_, \oc8051_golden_model_1.PC [8]);
  and (_02727_, _02726_, \oc8051_golden_model_1.PC [9]);
  and (_02728_, _02727_, \oc8051_golden_model_1.PC [10]);
  and (_02729_, _02728_, \oc8051_golden_model_1.PC [11]);
  and (_02730_, _02729_, \oc8051_golden_model_1.PC [12]);
  and (_02731_, _02730_, \oc8051_golden_model_1.PC [13]);
  and (_02732_, _02731_, \oc8051_golden_model_1.PC [14]);
  nor (_02733_, _02732_, \oc8051_golden_model_1.PC [15]);
  and (_02734_, _02732_, \oc8051_golden_model_1.PC [15]);
  or (_02735_, _02734_, _02733_);
  nor (_02736_, _02735_, _02715_);
  and (_02737_, _02715_, PC_abstr[15]);
  nor (_02738_, _02737_, _02736_);
  nand (_02739_, _02738_, _12782_);
  or (_02740_, _12782_, \oc8051_golden_model_1.PC [15]);
  and (_02741_, _02740_, _13707_);
  and (_13839_[15], _02741_, _02739_);
  and (_02742_, _02715_, XRAM_ADDR_abstr[15]);
  or (_02743_, _02742_, _12786_);
  or (_02744_, _12782_, \oc8051_golden_model_1.XRAM_ADDR [15]);
  and (_02745_, _02744_, _13707_);
  and (_13850_[15], _02745_, _02743_);
  and (_13849_[7], \oc8051_golden_model_1.TMOD [7], _13707_);
  and (_13848_[7], \oc8051_golden_model_1.TL1 [7], _13707_);
  and (_13847_[7], \oc8051_golden_model_1.TL0 [7], _13707_);
  and (_13846_[7], \oc8051_golden_model_1.TH1 [7], _13707_);
  and (_13845_[7], \oc8051_golden_model_1.TH0 [7], _13707_);
  and (_13844_[7], \oc8051_golden_model_1.TCON [7], _13707_);
  or (_02747_, _12782_, \oc8051_golden_model_1.SP [7]);
  and (_02748_, _02747_, _13707_);
  and (_02749_, _02715_, SP_abstr[7]);
  or (_02750_, _02749_, _12786_);
  and (_02751_, _02353_, \oc8051_golden_model_1.PC [2]);
  nor (_02752_, _02751_, _02342_);
  nor (_02753_, _02752_, _02374_);
  or (_02754_, _02715_, _02753_);
  nand (_02755_, _02715_, RD_ROM_1_ABSTR_ADDR[3]);
  and (_02756_, _02755_, _02754_);
  nand (_02757_, _02715_, RD_ROM_1_ABSTR_ADDR[2]);
  and (_02758_, _02714_, _02531_);
  nor (_02759_, _02353_, \oc8051_golden_model_1.PC [2]);
  nor (_02760_, _02759_, _02751_);
  nand (_02761_, _02760_, _02758_);
  nand (_02762_, _02761_, _02757_);
  or (_02763_, _02762_, _02756_);
  or (_02764_, _02715_, _02326_);
  or (_02765_, _02758_, RD_ROM_1_ABSTR_ADDR[0]);
  nand (_02766_, _02765_, _02764_);
  and (_02767_, _02354_, _02321_);
  nand (_02768_, _02767_, _02758_);
  nand (_02769_, _02715_, RD_ROM_1_ABSTR_ADDR[1]);
  and (_02770_, _02769_, _02768_);
  or (_02771_, _02770_, _02766_);
  or (_02772_, _02771_, _02763_);
  or (_02773_, _02772_, _02352_);
  and (_02774_, _02765_, _02764_);
  nand (_02775_, _02769_, _02768_);
  or (_02776_, _02775_, _02774_);
  nand (_02777_, _02755_, _02754_);
  or (_02778_, _02762_, _02777_);
  or (_02779_, _02778_, _02776_);
  or (_02780_, _02779_, _02320_);
  and (_02781_, _02780_, _02773_);
  and (_02782_, _02761_, _02757_);
  or (_02783_, _02782_, _02756_);
  nor (_02784_, _02783_, _02771_);
  nand (_02785_, _02784_, _12105_);
  or (_02786_, _02775_, _02766_);
  or (_02787_, _02782_, _02777_);
  or (_02788_, _02787_, _02786_);
  or (_02789_, _02788_, _02341_);
  and (_02790_, _02789_, _02785_);
  and (_02791_, _02790_, _02781_);
  or (_02792_, _02770_, _02774_);
  or (_02793_, _02792_, _02763_);
  or (_02794_, _02793_, _02371_);
  or (_02795_, _02786_, _02763_);
  or (_02796_, _02795_, _02384_);
  and (_02797_, _02796_, _02794_);
  or (_02798_, _02792_, _02783_);
  or (_02799_, _02798_, _02331_);
  or (_02800_, _02778_, _02771_);
  or (_02801_, _02800_, _02364_);
  and (_02802_, _02801_, _02799_);
  and (_02803_, _02802_, _02797_);
  and (_02804_, _02803_, _02791_);
  not (_02805_, _11670_);
  or (_02806_, _02787_, _02771_);
  or (_02807_, _02806_, _02805_);
  or (_02808_, _02787_, _02792_);
  or (_02809_, _02808_, _02348_);
  and (_02810_, _02809_, _02807_);
  or (_02811_, _02787_, _02776_);
  or (_02812_, _02811_, _02387_);
  or (_02813_, _02786_, _02778_);
  or (_02814_, _02813_, _02367_);
  and (_02815_, _02814_, _02812_);
  and (_02816_, _02815_, _02810_);
  or (_02817_, _02776_, _02763_);
  or (_02818_, _02817_, _02358_);
  or (_02819_, _02792_, _02778_);
  or (_02820_, _02819_, _02325_);
  and (_02821_, _02820_, _02818_);
  or (_02822_, _02786_, _02783_);
  or (_02823_, _02822_, _02380_);
  or (_02824_, _02783_, _02776_);
  or (_02825_, _02824_, _02336_);
  and (_02826_, _02825_, _02823_);
  and (_02827_, _02826_, _02821_);
  and (_02828_, _02827_, _02816_);
  and (_02829_, _02828_, _02804_);
  or (_02830_, _02811_, _02401_);
  or (_02831_, _02800_, _02419_);
  and (_02832_, _02831_, _02830_);
  or (_02833_, _02798_, _02417_);
  or (_02834_, _02817_, _02396_);
  and (_02835_, _02834_, _02833_);
  and (_02836_, _02835_, _02832_);
  or (_02837_, _02808_, _02431_);
  or (_02838_, _02788_, _02426_);
  and (_02839_, _02838_, _02837_);
  or (_02840_, _02819_, _02428_);
  or (_02841_, _02813_, _02407_);
  and (_02842_, _02841_, _02840_);
  and (_02843_, _02842_, _02839_);
  and (_02844_, _02843_, _02836_);
  or (_02845_, _02824_, _02394_);
  or (_02846_, _02772_, _02399_);
  and (_02847_, _02846_, _02845_);
  nand (_02848_, _02784_, _12110_);
  or (_02849_, _02822_, _02410_);
  and (_02850_, _02849_, _02848_);
  and (_02851_, _02850_, _02847_);
  or (_02852_, _02793_, _02405_);
  or (_02853_, _02795_, _02412_);
  and (_02854_, _02853_, _02852_);
  not (_02855_, _11677_);
  or (_02856_, _02806_, _02855_);
  or (_02857_, _02779_, _02433_);
  and (_02858_, _02857_, _02856_);
  and (_02859_, _02858_, _02854_);
  and (_02860_, _02859_, _02851_);
  and (_02861_, _02860_, _02844_);
  and (_02862_, _02861_, _02829_);
  or (_02863_, _02772_, _02548_);
  or (_02864_, _02793_, _02560_);
  and (_02865_, _02864_, _02863_);
  or (_02866_, _02824_, _02539_);
  or (_02867_, _02795_, _02569_);
  and (_02868_, _02867_, _02866_);
  and (_02869_, _02868_, _02865_);
  not (_02870_, _11684_);
  or (_02871_, _02806_, _02870_);
  or (_02872_, _02808_, _02545_);
  and (_02873_, _02872_, _02871_);
  or (_02874_, _02811_, _02571_);
  or (_02875_, _02819_, _02557_);
  and (_02876_, _02875_, _02874_);
  and (_02877_, _02876_, _02873_);
  and (_02878_, _02877_, _02869_);
  or (_02879_, _02822_, _02566_);
  or (_02880_, _02779_, _02534_);
  and (_02881_, _02880_, _02879_);
  or (_02882_, _02817_, _02550_);
  or (_02883_, _02800_, _02532_);
  and (_02884_, _02883_, _02882_);
  and (_02885_, _02884_, _02881_);
  nand (_02886_, _02784_, _12115_);
  or (_02887_, _02813_, _02555_);
  and (_02888_, _02887_, _02886_);
  or (_02889_, _02798_, _02537_);
  or (_02890_, _02788_, _02543_);
  and (_02891_, _02890_, _02889_);
  and (_02892_, _02891_, _02888_);
  and (_02893_, _02892_, _02885_);
  and (_02894_, _02893_, _02878_);
  or (_02895_, _02824_, _02655_);
  or (_02896_, _02772_, _02647_);
  and (_02897_, _02896_, _02895_);
  or (_02898_, _02808_, _02634_);
  or (_02899_, _02788_, _02639_);
  and (_02900_, _02899_, _02898_);
  and (_02901_, _02900_, _02897_);
  or (_02902_, _02798_, _02650_);
  or (_02903_, _02822_, _02660_);
  and (_02904_, _02903_, _02902_);
  or (_02905_, _02793_, _02657_);
  or (_02906_, _02795_, _02662_);
  and (_02907_, _02906_, _02905_);
  and (_02908_, _02907_, _02904_);
  and (_02909_, _02908_, _02901_);
  or (_02910_, _02779_, _02625_);
  or (_02911_, _02819_, _02636_);
  and (_02912_, _02911_, _02910_);
  not (_02913_, _11698_);
  or (_02914_, _02806_, _02913_);
  or (_02915_, _02811_, _02623_);
  and (_02916_, _02915_, _02914_);
  and (_02917_, _02916_, _02912_);
  nand (_02918_, _02784_, _12125_);
  or (_02919_, _02817_, _02628_);
  and (_02920_, _02919_, _02918_);
  or (_02921_, _02800_, _02630_);
  or (_02922_, _02813_, _02641_);
  and (_02923_, _02922_, _02921_);
  and (_02924_, _02923_, _02920_);
  and (_02925_, _02924_, _02917_);
  and (_02926_, _02925_, _02909_);
  or (_02927_, _02772_, _02675_);
  or (_02928_, _02779_, _02681_);
  and (_02929_, _02928_, _02927_);
  nand (_02930_, _02784_, _12090_);
  or (_02931_, _02788_, _02692_);
  and (_02932_, _02931_, _02930_);
  and (_02933_, _02932_, _02929_);
  or (_02934_, _02793_, _02679_);
  or (_02935_, _02795_, _02684_);
  and (_02936_, _02935_, _02934_);
  or (_02937_, _02798_, _02695_);
  or (_02938_, _02819_, _02670_);
  and (_02939_, _02938_, _02937_);
  and (_02940_, _02939_, _02936_);
  and (_02941_, _02940_, _02933_);
  not (_02942_, _11651_);
  or (_02943_, _02806_, _02942_);
  or (_02944_, _02808_, _02705_);
  and (_02945_, _02944_, _02943_);
  or (_02946_, _02811_, _02702_);
  or (_02948_, _02813_, _02707_);
  and (_02949_, _02948_, _02946_);
  and (_02950_, _02949_, _02945_);
  or (_02951_, _02817_, _02668_);
  or (_02952_, _02800_, _02686_);
  and (_02953_, _02952_, _02951_);
  or (_02954_, _02822_, _02673_);
  or (_02955_, _02824_, _02700_);
  and (_02956_, _02955_, _02954_);
  and (_02957_, _02956_, _02953_);
  and (_02958_, _02957_, _02950_);
  nand (_02959_, _02958_, _02941_);
  and (_02960_, _02959_, _02926_);
  not (_02961_, _11691_);
  or (_02962_, _02806_, _02961_);
  or (_02963_, _02800_, _02579_);
  and (_02964_, _02963_, _02962_);
  or (_02965_, _02793_, _02593_);
  or (_02966_, _02817_, _02584_);
  and (_02967_, _02966_, _02965_);
  and (_02968_, _02967_, _02964_);
  or (_02969_, _02819_, _02616_);
  or (_02970_, _02813_, _02595_);
  and (_02971_, _02970_, _02969_);
  or (_02972_, _02788_, _02577_);
  or (_02973_, _02811_, _02602_);
  and (_02974_, _02973_, _02972_);
  and (_02975_, _02974_, _02971_);
  and (_02976_, _02975_, _02968_);
  or (_02977_, _02798_, _02582_);
  or (_02978_, _02795_, _02614_);
  and (_02979_, _02978_, _02977_);
  or (_02980_, _02822_, _02588_);
  or (_02981_, _02772_, _02611_);
  and (_02982_, _02981_, _02980_);
  and (_02983_, _02982_, _02979_);
  or (_02984_, _02808_, _02600_);
  or (_02985_, _02779_, _02606_);
  and (_02986_, _02985_, _02984_);
  nand (_02987_, _02784_, _12120_);
  or (_02988_, _02824_, _02590_);
  and (_02989_, _02988_, _02987_);
  and (_02990_, _02989_, _02986_);
  and (_02991_, _02990_, _02983_);
  nand (_02992_, _02991_, _02976_);
  not (_02993_, _02992_);
  and (_02994_, _02993_, _02960_);
  and (_02995_, _02994_, _02894_);
  nand (_02996_, _02784_, _12095_);
  or (_02997_, _02800_, _02479_);
  and (_02998_, _02997_, _02996_);
  or (_02999_, _02822_, _02456_);
  or (_03000_, _02817_, _02442_);
  and (_03001_, _03000_, _02999_);
  and (_03002_, _03001_, _02998_);
  or (_03003_, _02772_, _02445_);
  not (_03004_, _11656_);
  or (_03005_, _02806_, _03004_);
  and (_03006_, _03005_, _03003_);
  or (_03007_, _02808_, _02469_);
  or (_03009_, _02813_, _02447_);
  and (_03010_, _03009_, _03007_);
  and (_03011_, _03010_, _03006_);
  and (_03012_, _03011_, _03002_);
  or (_03013_, _02798_, _02463_);
  or (_03014_, _02824_, _02440_);
  and (_03015_, _03014_, _03013_);
  or (_03016_, _02795_, _02458_);
  or (_03017_, _02819_, _02475_);
  and (_03018_, _03017_, _03016_);
  and (_03020_, _03018_, _03015_);
  or (_03021_, _02793_, _02451_);
  or (_03022_, _02811_, _02473_);
  and (_03023_, _03022_, _03021_);
  or (_03024_, _02788_, _02465_);
  or (_03025_, _02779_, _02453_);
  and (_03026_, _03025_, _03024_);
  and (_03027_, _03026_, _03023_);
  and (_03028_, _03027_, _03020_);
  and (_03029_, _03028_, _03012_);
  not (_03030_, _03029_);
  nand (_03031_, _02784_, _12100_);
  or (_03032_, _02772_, _02518_);
  and (_03033_, _03032_, _03031_);
  or (_03034_, _02808_, _02496_);
  or (_03035_, _02779_, _02487_);
  and (_03036_, _03035_, _03034_);
  and (_03037_, _03036_, _03033_);
  or (_03038_, _02793_, _02524_);
  or (_03039_, _02795_, _02520_);
  and (_03041_, _03039_, _03038_);
  or (_03042_, _02798_, _02510_);
  or (_03043_, _02824_, _02513_);
  and (_03044_, _03043_, _03042_);
  and (_03045_, _03044_, _03041_);
  and (_03046_, _03045_, _03037_);
  or (_03047_, _02811_, _02485_);
  or (_03048_, _02800_, _02492_);
  and (_03049_, _03048_, _03047_);
  not (_03050_, _11663_);
  or (_03051_, _02806_, _03050_);
  or (_03052_, _02788_, _02501_);
  and (_03053_, _03052_, _03051_);
  and (_03054_, _03053_, _03049_);
  or (_03055_, _02819_, _02498_);
  or (_03056_, _02813_, _02503_);
  and (_03057_, _03056_, _03055_);
  or (_03058_, _02822_, _02508_);
  or (_03059_, _02817_, _02490_);
  and (_03060_, _03059_, _03058_);
  and (_03062_, _03060_, _03057_);
  and (_03063_, _03062_, _03054_);
  and (_03064_, _03063_, _03046_);
  and (_03065_, _03064_, _03030_);
  and (_03066_, _03065_, _02995_);
  and (_03067_, _03066_, _02862_);
  not (_03068_, _03067_);
  nand (_03069_, _02860_, _02844_);
  and (_03070_, _03069_, _02758_);
  and (_03071_, _02715_, RD_IRAM_0_ABSTR_ADDR[3]);
  nor (_03072_, _03071_, _03070_);
  not (_03073_, _03072_);
  and (_03074_, _02715_, RD_IRAM_0_ABSTR_ADDR[2]);
  nor (_03075_, _02829_, _02715_);
  nor (_03076_, _03075_, _03074_);
  not (_03077_, _03076_);
  and (_03078_, _02715_, RD_IRAM_0_ABSTR_ADDR[1]);
  not (_03079_, _03078_);
  or (_03080_, _03064_, _02715_);
  and (_03081_, _03080_, _03079_);
  not (_03083_, _03081_);
  and (_03084_, _02715_, RD_IRAM_0_ABSTR_ADDR[0]);
  not (_03085_, _03084_);
  or (_03086_, _03029_, _02715_);
  and (_03087_, _03086_, _03085_);
  and (_03088_, _03087_, \oc8051_golden_model_1.IRAM[0] [7]);
  nand (_03089_, _03086_, _03085_);
  and (_03090_, _03089_, \oc8051_golden_model_1.IRAM[1] [7]);
  nor (_03091_, _03090_, _03088_);
  nor (_03092_, _03091_, _03083_);
  and (_03094_, _03087_, \oc8051_golden_model_1.IRAM[2] [7]);
  and (_03095_, _03089_, \oc8051_golden_model_1.IRAM[3] [7]);
  or (_03096_, _03095_, _03094_);
  and (_03097_, _03096_, _03083_);
  nor (_03098_, _03097_, _03092_);
  nor (_03099_, _03098_, _03077_);
  and (_03100_, _03087_, \oc8051_golden_model_1.IRAM[4] [7]);
  and (_03101_, _03089_, \oc8051_golden_model_1.IRAM[5] [7]);
  or (_03102_, _03101_, _03100_);
  and (_03103_, _03102_, _03081_);
  and (_03105_, _03087_, \oc8051_golden_model_1.IRAM[6] [7]);
  and (_03106_, _03089_, \oc8051_golden_model_1.IRAM[7] [7]);
  or (_03107_, _03106_, _03105_);
  and (_03108_, _03107_, _03083_);
  nor (_03109_, _03108_, _03103_);
  nor (_03110_, _03109_, _03076_);
  nor (_03111_, _03110_, _03099_);
  nor (_03112_, _03111_, _03073_);
  and (_03113_, _03087_, \oc8051_golden_model_1.IRAM[8] [7]);
  and (_03114_, _03089_, \oc8051_golden_model_1.IRAM[9] [7]);
  or (_03116_, _03114_, _03113_);
  and (_03117_, _03116_, _03081_);
  and (_03118_, _03087_, \oc8051_golden_model_1.IRAM[10] [7]);
  and (_03119_, _03089_, \oc8051_golden_model_1.IRAM[11] [7]);
  or (_03120_, _03119_, _03118_);
  and (_03121_, _03120_, _03083_);
  nor (_03122_, _03121_, _03117_);
  nor (_03123_, _03122_, _03077_);
  and (_03124_, _03087_, \oc8051_golden_model_1.IRAM[12] [7]);
  and (_03125_, _03089_, \oc8051_golden_model_1.IRAM[13] [7]);
  or (_03127_, _03125_, _03124_);
  and (_03128_, _03127_, _03081_);
  and (_03129_, _03087_, \oc8051_golden_model_1.IRAM[14] [7]);
  and (_03130_, _03089_, \oc8051_golden_model_1.IRAM[15] [7]);
  or (_03131_, _03130_, _03129_);
  and (_03132_, _03131_, _03083_);
  nor (_03133_, _03132_, _03128_);
  nor (_03134_, _03133_, _03076_);
  nor (_03135_, _03134_, _03123_);
  nor (_03136_, _03135_, _03072_);
  nor (_03138_, _03136_, _03112_);
  nor (_03139_, _03138_, _02959_);
  not (_03140_, _03139_);
  and (_03141_, _03069_, _02829_);
  not (_03142_, _03064_);
  and (_03143_, _03142_, _03029_);
  and (_03144_, _03143_, _02995_);
  and (_03145_, _03144_, _03141_);
  and (_03146_, _03145_, \oc8051_golden_model_1.TL0 [7]);
  not (_03147_, _03146_);
  and (_03149_, _03064_, _03029_);
  and (_03150_, _03149_, _02862_);
  not (_03151_, _02959_);
  nor (_03152_, _03151_, _02926_);
  and (_03153_, _03152_, _03150_);
  nor (_03154_, _02992_, _02894_);
  and (_03155_, _03154_, _03153_);
  and (_03156_, _03155_, \oc8051_golden_model_1.PSW [7]);
  not (_03157_, _03156_);
  not (_03158_, \oc8051_golden_model_1.ACC [7]);
  nand (_03161_, _03152_, _03150_);
  and (_03162_, _02992_, _02894_);
  not (_03163_, _03162_);
  or (_03164_, _03163_, _03161_);
  nor (_03165_, _03164_, _03158_);
  and (_03166_, _03154_, _02960_);
  and (_03167_, _03141_, _03065_);
  and (_03168_, _03167_, _03166_);
  and (_03169_, _03168_, \oc8051_golden_model_1.SBUF [7]);
  nor (_03170_, _03169_, _03165_);
  and (_03172_, _03170_, _03157_);
  and (_03173_, _03172_, _03147_);
  nor (_03174_, _03064_, _03029_);
  and (_03175_, _03174_, _02995_);
  and (_03176_, _03175_, _03141_);
  and (_03177_, _03176_, \oc8051_golden_model_1.TL1 [7]);
  and (_03178_, _03144_, _02862_);
  and (_03179_, _03178_, \oc8051_golden_model_1.DPL [7]);
  nor (_03180_, _03179_, _03177_);
  and (_03181_, _03180_, _03173_);
  and (_03182_, _03067_, \oc8051_golden_model_1.SP [7]);
  not (_03183_, _03182_);
  and (_03184_, _03167_, _02995_);
  and (_03185_, _03184_, \oc8051_golden_model_1.TMOD [7]);
  nor (_03186_, _02861_, _02829_);
  and (_03187_, _03186_, _03066_);
  and (_03188_, _03187_, \oc8051_golden_model_1.TH1 [7]);
  nor (_03189_, _03188_, _03185_);
  and (_03190_, _03189_, _03183_);
  nor (_03191_, _02993_, _02894_);
  and (_03192_, _03191_, _03153_);
  and (_03193_, _03192_, \oc8051_golden_model_1.B [7]);
  and (_03194_, _03149_, _03141_);
  and (_03195_, _03194_, _03166_);
  and (_03196_, _03195_, \oc8051_golden_model_1.SCON [7]);
  nor (_03197_, _03196_, _03193_);
  and (_03198_, _03166_, _03150_);
  and (_03199_, _03198_, \oc8051_golden_model_1.P1 [7]);
  and (_03200_, _03194_, _02995_);
  and (_03201_, _03200_, \oc8051_golden_model_1.TCON [7]);
  nor (_03202_, _03201_, _03199_);
  and (_03203_, _03202_, _03197_);
  and (_03204_, _03191_, _02960_);
  and (_03205_, _03204_, _03194_);
  and (_03206_, _03205_, \oc8051_golden_model_1.IP [7]);
  and (_03207_, _03162_, _02960_);
  and (_03208_, _03207_, _03150_);
  and (_03209_, _03208_, \oc8051_golden_model_1.P2 [7]);
  nor (_03210_, _03209_, _03206_);
  and (_03211_, _03207_, _03194_);
  and (_03212_, _03211_, \oc8051_golden_model_1.IE [7]);
  and (_03213_, _03204_, _03150_);
  and (_03214_, _03213_, \oc8051_golden_model_1.P3 [7]);
  nor (_03215_, _03214_, _03212_);
  and (_03216_, _03215_, _03210_);
  and (_03217_, _03150_, _02995_);
  and (_03218_, _03217_, \oc8051_golden_model_1.P0 [7]);
  and (_03219_, _03186_, _03149_);
  and (_03220_, _03219_, _02995_);
  and (_03221_, _03220_, \oc8051_golden_model_1.TH0 [7]);
  nor (_03222_, _03221_, _03218_);
  and (_03223_, _03222_, _03216_);
  and (_03224_, _03223_, _03203_);
  and (_03225_, _03224_, _03190_);
  nor (_03226_, _03069_, _02829_);
  and (_03227_, _03226_, _03175_);
  and (_03228_, _03227_, \oc8051_golden_model_1.PCON [7]);
  and (_03229_, _03175_, _02862_);
  and (_03230_, _03229_, \oc8051_golden_model_1.DPH [7]);
  nor (_03231_, _03230_, _03228_);
  and (_03232_, _03231_, _03225_);
  and (_03233_, _03232_, _03181_);
  and (_03234_, _03233_, _03140_);
  and (_03235_, _03087_, \oc8051_golden_model_1.IRAM[0] [6]);
  and (_03236_, _03089_, \oc8051_golden_model_1.IRAM[1] [6]);
  or (_03237_, _03236_, _03235_);
  and (_03238_, _03237_, _03081_);
  and (_03239_, _03087_, \oc8051_golden_model_1.IRAM[2] [6]);
  and (_03240_, _03089_, \oc8051_golden_model_1.IRAM[3] [6]);
  or (_03241_, _03240_, _03239_);
  and (_03242_, _03241_, _03083_);
  nor (_03243_, _03242_, _03238_);
  nor (_03244_, _03243_, _03077_);
  and (_03245_, _03087_, \oc8051_golden_model_1.IRAM[4] [6]);
  and (_03246_, _03089_, \oc8051_golden_model_1.IRAM[5] [6]);
  or (_03247_, _03246_, _03245_);
  and (_03248_, _03247_, _03081_);
  and (_03249_, _03087_, \oc8051_golden_model_1.IRAM[6] [6]);
  and (_03250_, _03089_, \oc8051_golden_model_1.IRAM[7] [6]);
  or (_03251_, _03250_, _03249_);
  and (_03252_, _03251_, _03083_);
  nor (_03253_, _03252_, _03248_);
  nor (_03254_, _03253_, _03076_);
  nor (_03255_, _03254_, _03244_);
  nor (_03256_, _03255_, _03073_);
  and (_03257_, _03087_, \oc8051_golden_model_1.IRAM[8] [6]);
  and (_03258_, _03089_, \oc8051_golden_model_1.IRAM[9] [6]);
  or (_03259_, _03258_, _03257_);
  and (_03260_, _03259_, _03081_);
  and (_03261_, _03087_, \oc8051_golden_model_1.IRAM[10] [6]);
  and (_03262_, _03089_, \oc8051_golden_model_1.IRAM[11] [6]);
  or (_03263_, _03262_, _03261_);
  and (_03264_, _03263_, _03083_);
  nor (_03265_, _03264_, _03260_);
  nor (_03266_, _03265_, _03077_);
  and (_03267_, _03087_, \oc8051_golden_model_1.IRAM[12] [6]);
  and (_03268_, _03089_, \oc8051_golden_model_1.IRAM[13] [6]);
  or (_03269_, _03268_, _03267_);
  and (_03270_, _03269_, _03081_);
  and (_03271_, _03087_, \oc8051_golden_model_1.IRAM[14] [6]);
  and (_03272_, _03089_, \oc8051_golden_model_1.IRAM[15] [6]);
  or (_03273_, _03272_, _03271_);
  and (_03274_, _03273_, _03083_);
  nor (_03275_, _03274_, _03270_);
  nor (_03276_, _03275_, _03076_);
  nor (_03277_, _03276_, _03266_);
  nor (_03278_, _03277_, _03072_);
  nor (_03279_, _03278_, _03256_);
  nor (_03280_, _03279_, _02959_);
  not (_03281_, _03280_);
  and (_03282_, _03145_, \oc8051_golden_model_1.TL0 [6]);
  not (_03283_, _03282_);
  and (_03284_, _03220_, \oc8051_golden_model_1.TH0 [6]);
  not (_03285_, _03284_);
  and (_03286_, _03195_, \oc8051_golden_model_1.SCON [6]);
  and (_03287_, _03168_, \oc8051_golden_model_1.SBUF [6]);
  nor (_03288_, _03287_, _03286_);
  and (_03289_, _03288_, _03285_);
  and (_03290_, _03289_, _03283_);
  and (_03291_, _03176_, \oc8051_golden_model_1.TL1 [6]);
  and (_03292_, _03178_, \oc8051_golden_model_1.DPL [6]);
  nor (_03293_, _03292_, _03291_);
  and (_03294_, _03293_, _03290_);
  and (_03295_, _03067_, \oc8051_golden_model_1.SP [6]);
  not (_03296_, _03295_);
  and (_03297_, _03184_, \oc8051_golden_model_1.TMOD [6]);
  and (_03298_, _03187_, \oc8051_golden_model_1.TH1 [6]);
  nor (_03299_, _03298_, _03297_);
  and (_03300_, _03299_, _03296_);
  and (_03301_, _03192_, \oc8051_golden_model_1.B [6]);
  and (_03302_, _03198_, \oc8051_golden_model_1.P1 [6]);
  nor (_03303_, _03302_, _03301_);
  and (_03304_, _03200_, \oc8051_golden_model_1.TCON [6]);
  and (_03305_, _03217_, \oc8051_golden_model_1.P0 [6]);
  nor (_03306_, _03305_, _03304_);
  and (_03307_, _03306_, _03303_);
  and (_03308_, _03205_, \oc8051_golden_model_1.IP [6]);
  and (_03309_, _03208_, \oc8051_golden_model_1.P2 [6]);
  nor (_03310_, _03309_, _03308_);
  and (_03311_, _03211_, \oc8051_golden_model_1.IE [6]);
  and (_03312_, _03213_, \oc8051_golden_model_1.P3 [6]);
  nor (_03313_, _03312_, _03311_);
  and (_03314_, _03313_, _03310_);
  not (_03315_, \oc8051_golden_model_1.ACC [6]);
  nor (_03316_, _03164_, _03315_);
  and (_03317_, _03155_, \oc8051_golden_model_1.PSW [6]);
  nor (_03318_, _03317_, _03316_);
  and (_03319_, _03318_, _03314_);
  and (_03320_, _03319_, _03307_);
  and (_03321_, _03320_, _03300_);
  and (_03322_, _03227_, \oc8051_golden_model_1.PCON [6]);
  and (_03323_, _03229_, \oc8051_golden_model_1.DPH [6]);
  nor (_03324_, _03323_, _03322_);
  and (_03325_, _03324_, _03321_);
  and (_03326_, _03325_, _03294_);
  and (_03327_, _03326_, _03281_);
  not (_03328_, _03327_);
  and (_03329_, _03087_, \oc8051_golden_model_1.IRAM[0] [5]);
  and (_03330_, _03089_, \oc8051_golden_model_1.IRAM[1] [5]);
  or (_03331_, _03330_, _03329_);
  and (_03332_, _03331_, _03081_);
  and (_03333_, _03087_, \oc8051_golden_model_1.IRAM[2] [5]);
  and (_03334_, _03089_, \oc8051_golden_model_1.IRAM[3] [5]);
  or (_03335_, _03334_, _03333_);
  and (_03336_, _03335_, _03083_);
  nor (_03337_, _03336_, _03332_);
  nor (_03338_, _03337_, _03077_);
  and (_03339_, _03087_, \oc8051_golden_model_1.IRAM[4] [5]);
  and (_03340_, _03089_, \oc8051_golden_model_1.IRAM[5] [5]);
  or (_03341_, _03340_, _03339_);
  and (_03342_, _03341_, _03081_);
  and (_03343_, _03087_, \oc8051_golden_model_1.IRAM[6] [5]);
  and (_03344_, _03089_, \oc8051_golden_model_1.IRAM[7] [5]);
  or (_03345_, _03344_, _03343_);
  and (_03346_, _03345_, _03083_);
  nor (_03347_, _03346_, _03342_);
  nor (_03348_, _03347_, _03076_);
  nor (_03349_, _03348_, _03338_);
  nor (_03350_, _03349_, _03073_);
  and (_03351_, _03087_, \oc8051_golden_model_1.IRAM[8] [5]);
  and (_03352_, _03089_, \oc8051_golden_model_1.IRAM[9] [5]);
  or (_03353_, _03352_, _03351_);
  and (_03354_, _03353_, _03081_);
  and (_03355_, _03087_, \oc8051_golden_model_1.IRAM[10] [5]);
  and (_03356_, _03089_, \oc8051_golden_model_1.IRAM[11] [5]);
  or (_03357_, _03356_, _03355_);
  and (_03358_, _03357_, _03083_);
  nor (_03359_, _03358_, _03354_);
  nor (_03360_, _03359_, _03077_);
  and (_03361_, _03087_, \oc8051_golden_model_1.IRAM[12] [5]);
  and (_03363_, _03089_, \oc8051_golden_model_1.IRAM[13] [5]);
  or (_03364_, _03363_, _03361_);
  and (_03365_, _03364_, _03081_);
  and (_03366_, _03087_, \oc8051_golden_model_1.IRAM[14] [5]);
  and (_03367_, _03089_, \oc8051_golden_model_1.IRAM[15] [5]);
  or (_03368_, _03367_, _03366_);
  and (_03369_, _03368_, _03083_);
  nor (_03370_, _03369_, _03365_);
  nor (_03371_, _03370_, _03076_);
  nor (_03372_, _03371_, _03360_);
  nor (_03373_, _03372_, _03072_);
  nor (_03374_, _03373_, _03350_);
  nor (_03375_, _03374_, _02959_);
  not (_03376_, _03375_);
  and (_03377_, _03178_, \oc8051_golden_model_1.DPL [5]);
  not (_03378_, _03377_);
  and (_03379_, _03195_, \oc8051_golden_model_1.SCON [5]);
  not (_03380_, _03379_);
  and (_03381_, _03200_, \oc8051_golden_model_1.TCON [5]);
  and (_03382_, _03220_, \oc8051_golden_model_1.TH0 [5]);
  nor (_03383_, _03382_, _03381_);
  and (_03384_, _03383_, _03380_);
  and (_03385_, _03384_, _03378_);
  and (_03386_, _03176_, \oc8051_golden_model_1.TL1 [5]);
  and (_03387_, _03145_, \oc8051_golden_model_1.TL0 [5]);
  nor (_03388_, _03387_, _03386_);
  and (_03389_, _03388_, _03385_);
  and (_03390_, _03067_, \oc8051_golden_model_1.SP [5]);
  not (_03391_, _03390_);
  and (_03392_, _03184_, \oc8051_golden_model_1.TMOD [5]);
  and (_03393_, _03187_, \oc8051_golden_model_1.TH1 [5]);
  nor (_03394_, _03393_, _03392_);
  and (_03395_, _03394_, _03391_);
  and (_03396_, _03198_, \oc8051_golden_model_1.P1 [5]);
  and (_03397_, _03217_, \oc8051_golden_model_1.P0 [5]);
  nor (_03398_, _03397_, _03396_);
  and (_03399_, _03192_, \oc8051_golden_model_1.B [5]);
  and (_03400_, _03168_, \oc8051_golden_model_1.SBUF [5]);
  nor (_03401_, _03400_, _03399_);
  and (_03402_, _03401_, _03398_);
  and (_03403_, _03213_, \oc8051_golden_model_1.P3 [5]);
  and (_03404_, _03208_, \oc8051_golden_model_1.P2 [5]);
  nor (_03405_, _03404_, _03403_);
  and (_03406_, _03211_, \oc8051_golden_model_1.IE [5]);
  and (_03407_, _03205_, \oc8051_golden_model_1.IP [5]);
  nor (_03408_, _03407_, _03406_);
  and (_03409_, _03408_, _03405_);
  not (_03410_, \oc8051_golden_model_1.ACC [5]);
  nor (_03411_, _03164_, _03410_);
  and (_03412_, _03155_, \oc8051_golden_model_1.PSW [5]);
  nor (_03413_, _03412_, _03411_);
  and (_03414_, _03413_, _03409_);
  and (_03415_, _03414_, _03402_);
  and (_03416_, _03415_, _03395_);
  and (_03417_, _03227_, \oc8051_golden_model_1.PCON [5]);
  and (_03418_, _03229_, \oc8051_golden_model_1.DPH [5]);
  nor (_03419_, _03418_, _03417_);
  and (_03420_, _03419_, _03416_);
  and (_03421_, _03420_, _03389_);
  and (_03422_, _03421_, _03376_);
  nor (_03423_, _03089_, \oc8051_golden_model_1.IRAM[8] [3]);
  or (_03424_, _03087_, \oc8051_golden_model_1.IRAM[9] [3]);
  nand (_03425_, _03424_, _03081_);
  or (_03426_, _03425_, _03423_);
  not (_03427_, \oc8051_golden_model_1.IRAM[10] [3]);
  and (_03428_, _03087_, _03427_);
  or (_03429_, _03087_, \oc8051_golden_model_1.IRAM[11] [3]);
  nand (_03430_, _03429_, _03083_);
  or (_03431_, _03430_, _03428_);
  nand (_03432_, _03431_, _03426_);
  nand (_03433_, _03432_, _03076_);
  nor (_03434_, _03087_, \oc8051_golden_model_1.IRAM[13] [3]);
  or (_03435_, _03089_, \oc8051_golden_model_1.IRAM[12] [3]);
  nand (_03436_, _03435_, _03081_);
  or (_03437_, _03436_, _03434_);
  not (_03438_, \oc8051_golden_model_1.IRAM[15] [3]);
  and (_03439_, _03089_, _03438_);
  or (_03440_, _03089_, \oc8051_golden_model_1.IRAM[14] [3]);
  nand (_03441_, _03440_, _03083_);
  or (_03442_, _03441_, _03439_);
  nand (_03443_, _03442_, _03437_);
  nand (_03444_, _03443_, _03077_);
  nand (_03445_, _03444_, _03433_);
  nand (_03446_, _03445_, _03073_);
  nor (_03447_, _03087_, \oc8051_golden_model_1.IRAM[1] [3]);
  or (_03448_, _03089_, \oc8051_golden_model_1.IRAM[0] [3]);
  nand (_03449_, _03448_, _03081_);
  or (_03450_, _03449_, _03447_);
  not (_03451_, \oc8051_golden_model_1.IRAM[2] [3]);
  and (_03452_, _03087_, _03451_);
  or (_03453_, _03087_, \oc8051_golden_model_1.IRAM[3] [3]);
  nand (_03454_, _03453_, _03083_);
  or (_03455_, _03454_, _03452_);
  nand (_03456_, _03455_, _03450_);
  nand (_03457_, _03456_, _03076_);
  not (_03458_, \oc8051_golden_model_1.IRAM[5] [3]);
  and (_03459_, _03089_, _03458_);
  or (_03460_, _03089_, \oc8051_golden_model_1.IRAM[4] [3]);
  nand (_03461_, _03460_, _03081_);
  or (_03462_, _03461_, _03459_);
  nor (_03463_, _03089_, \oc8051_golden_model_1.IRAM[6] [3]);
  or (_03464_, _03087_, \oc8051_golden_model_1.IRAM[7] [3]);
  nand (_03465_, _03464_, _03083_);
  or (_03466_, _03465_, _03463_);
  nand (_03467_, _03466_, _03462_);
  nand (_03468_, _03467_, _03077_);
  nand (_03469_, _03468_, _03457_);
  nand (_03470_, _03469_, _03072_);
  nand (_03471_, _03470_, _03446_);
  nand (_03472_, _03471_, _03151_);
  and (_03473_, _03176_, \oc8051_golden_model_1.TL1 [3]);
  not (_03474_, _03473_);
  and (_03475_, _03220_, \oc8051_golden_model_1.TH0 [3]);
  not (_03476_, _03475_);
  and (_03477_, _03192_, \oc8051_golden_model_1.B [3]);
  and (_03478_, _03200_, \oc8051_golden_model_1.TCON [3]);
  nor (_03479_, _03478_, _03477_);
  and (_03480_, _03479_, _03476_);
  and (_03481_, _03480_, _03474_);
  and (_03482_, _03145_, \oc8051_golden_model_1.TL0 [3]);
  and (_03483_, _03178_, \oc8051_golden_model_1.DPL [3]);
  nor (_03484_, _03483_, _03482_);
  and (_03485_, _03484_, _03481_);
  and (_03486_, _03184_, \oc8051_golden_model_1.TMOD [3]);
  nand (_03487_, _03187_, \oc8051_golden_model_1.TH1 [3]);
  nand (_03488_, _03067_, \oc8051_golden_model_1.SP [3]);
  nand (_03489_, _03488_, _03487_);
  nor (_03490_, _03489_, _03486_);
  not (_03491_, \oc8051_golden_model_1.ACC [3]);
  nor (_03492_, _03164_, _03491_);
  and (_03493_, _03198_, \oc8051_golden_model_1.P1 [3]);
  nor (_03494_, _03493_, _03492_);
  and (_03495_, _03155_, \oc8051_golden_model_1.PSW [3]);
  and (_03496_, _03195_, \oc8051_golden_model_1.SCON [3]);
  nor (_03497_, _03496_, _03495_);
  and (_03498_, _03497_, _03494_);
  nand (_03499_, _03213_, \oc8051_golden_model_1.P3 [3]);
  nand (_03500_, _03208_, \oc8051_golden_model_1.P2 [3]);
  and (_03501_, _03500_, _03499_);
  nand (_03502_, _03211_, \oc8051_golden_model_1.IE [3]);
  nand (_03503_, _03205_, \oc8051_golden_model_1.IP [3]);
  and (_03504_, _03503_, _03502_);
  and (_03505_, _03504_, _03501_);
  and (_03506_, _03168_, \oc8051_golden_model_1.SBUF [3]);
  and (_03507_, _03217_, \oc8051_golden_model_1.P0 [3]);
  nor (_03508_, _03507_, _03506_);
  and (_03509_, _03508_, _03505_);
  and (_03510_, _03509_, _03498_);
  and (_03511_, _03510_, _03490_);
  and (_03512_, _03227_, \oc8051_golden_model_1.PCON [3]);
  and (_03513_, _03229_, \oc8051_golden_model_1.DPH [3]);
  nor (_03514_, _03513_, _03512_);
  and (_03515_, _03514_, _03511_);
  and (_03516_, _03515_, _03485_);
  and (_03517_, _03516_, _03472_);
  or (_03518_, _03089_, \oc8051_golden_model_1.IRAM[0] [1]);
  or (_03519_, _03087_, \oc8051_golden_model_1.IRAM[1] [1]);
  and (_03520_, _03519_, _03081_);
  nand (_03521_, _03520_, _03518_);
  or (_03522_, _03089_, \oc8051_golden_model_1.IRAM[2] [1]);
  or (_03523_, _03087_, \oc8051_golden_model_1.IRAM[3] [1]);
  and (_03524_, _03523_, _03083_);
  nand (_03525_, _03524_, _03522_);
  nand (_03526_, _03525_, _03521_);
  nand (_03527_, _03526_, _03076_);
  or (_03528_, _03087_, \oc8051_golden_model_1.IRAM[5] [1]);
  or (_03529_, _03089_, \oc8051_golden_model_1.IRAM[4] [1]);
  and (_03530_, _03529_, _03081_);
  nand (_03531_, _03530_, _03528_);
  or (_03532_, _03089_, \oc8051_golden_model_1.IRAM[6] [1]);
  or (_03533_, _03087_, \oc8051_golden_model_1.IRAM[7] [1]);
  and (_03534_, _03533_, _03083_);
  nand (_03535_, _03534_, _03532_);
  nand (_03536_, _03535_, _03531_);
  nand (_03537_, _03536_, _03077_);
  nand (_03538_, _03537_, _03527_);
  nand (_03539_, _03538_, _03072_);
  or (_03540_, _03087_, \oc8051_golden_model_1.IRAM[9] [1]);
  or (_03541_, _03089_, \oc8051_golden_model_1.IRAM[8] [1]);
  and (_03542_, _03541_, _03081_);
  nand (_03543_, _03542_, _03540_);
  or (_03544_, _03087_, \oc8051_golden_model_1.IRAM[11] [1]);
  or (_03545_, _03089_, \oc8051_golden_model_1.IRAM[10] [1]);
  and (_03546_, _03545_, _03083_);
  nand (_03547_, _03546_, _03544_);
  nand (_03548_, _03547_, _03543_);
  nand (_03549_, _03548_, _03076_);
  or (_03550_, _03089_, \oc8051_golden_model_1.IRAM[12] [1]);
  or (_03551_, _03087_, \oc8051_golden_model_1.IRAM[13] [1]);
  and (_03552_, _03551_, _03081_);
  nand (_03553_, _03552_, _03550_);
  or (_03554_, _03089_, \oc8051_golden_model_1.IRAM[14] [1]);
  or (_03555_, _03087_, \oc8051_golden_model_1.IRAM[15] [1]);
  and (_03556_, _03555_, _03083_);
  nand (_03557_, _03556_, _03554_);
  nand (_03558_, _03557_, _03553_);
  nand (_03559_, _03558_, _03077_);
  nand (_03560_, _03559_, _03549_);
  nand (_03561_, _03560_, _03073_);
  nand (_03562_, _03561_, _03539_);
  nand (_03564_, _03562_, _03151_);
  nand (_03565_, _03145_, \oc8051_golden_model_1.TL0 [1]);
  and (_03566_, _03168_, \oc8051_golden_model_1.SBUF [1]);
  nand (_03567_, _03198_, \oc8051_golden_model_1.P1 [1]);
  nand (_03568_, _03217_, \oc8051_golden_model_1.P0 [1]);
  nand (_03569_, _03568_, _03567_);
  nor (_03570_, _03569_, _03566_);
  and (_03571_, _03570_, _03565_);
  nand (_03572_, _03176_, \oc8051_golden_model_1.TL1 [1]);
  nand (_03573_, _03178_, \oc8051_golden_model_1.DPL [1]);
  and (_03574_, _03573_, _03572_);
  and (_03575_, _03574_, _03571_);
  nand (_03576_, _03184_, \oc8051_golden_model_1.TMOD [1]);
  nand (_03577_, _03187_, \oc8051_golden_model_1.TH1 [1]);
  nand (_03578_, _03067_, \oc8051_golden_model_1.SP [1]);
  and (_03579_, _03578_, _03577_);
  and (_03580_, _03579_, _03576_);
  nand (_03581_, _03195_, \oc8051_golden_model_1.SCON [1]);
  nand (_03582_, _03220_, \oc8051_golden_model_1.TH0 [1]);
  and (_03583_, _03582_, _03581_);
  nand (_03584_, _03192_, \oc8051_golden_model_1.B [1]);
  nand (_03585_, _03200_, \oc8051_golden_model_1.TCON [1]);
  and (_03586_, _03585_, _03584_);
  and (_03587_, _03586_, _03583_);
  nand (_03588_, _03211_, \oc8051_golden_model_1.IE [1]);
  nand (_03589_, _03205_, \oc8051_golden_model_1.IP [1]);
  and (_03590_, _03589_, _03588_);
  nand (_03591_, _03213_, \oc8051_golden_model_1.P3 [1]);
  nand (_03592_, _03208_, \oc8051_golden_model_1.P2 [1]);
  and (_03593_, _03592_, _03591_);
  and (_03594_, _03593_, _03590_);
  not (_03595_, \oc8051_golden_model_1.ACC [1]);
  or (_03596_, _03164_, _03595_);
  not (_03597_, \oc8051_golden_model_1.PSW [1]);
  not (_03598_, _03154_);
  or (_03599_, _03598_, _03161_);
  or (_03600_, _03599_, _03597_);
  and (_03601_, _03600_, _03596_);
  and (_03602_, _03601_, _03594_);
  and (_03603_, _03602_, _03587_);
  and (_03604_, _03603_, _03580_);
  nand (_03605_, _03227_, \oc8051_golden_model_1.PCON [1]);
  nand (_03606_, _03229_, \oc8051_golden_model_1.DPH [1]);
  and (_03607_, _03606_, _03605_);
  and (_03608_, _03607_, _03604_);
  and (_03609_, _03608_, _03575_);
  nand (_03610_, _03609_, _03564_);
  not (_03611_, \oc8051_golden_model_1.IRAM[4] [0]);
  or (_03612_, _03089_, _03611_);
  nand (_03613_, _03089_, \oc8051_golden_model_1.IRAM[5] [0]);
  nand (_03614_, _03613_, _03612_);
  nand (_03615_, _03614_, _03081_);
  nand (_03616_, _03087_, \oc8051_golden_model_1.IRAM[6] [0]);
  not (_03617_, \oc8051_golden_model_1.IRAM[7] [0]);
  or (_03618_, _03087_, _03617_);
  nand (_03619_, _03618_, _03616_);
  nand (_03620_, _03619_, _03083_);
  nand (_03621_, _03620_, _03615_);
  nand (_03622_, _03621_, _03077_);
  not (_03623_, \oc8051_golden_model_1.IRAM[0] [0]);
  or (_03624_, _03089_, _03623_);
  nand (_03625_, _03089_, \oc8051_golden_model_1.IRAM[1] [0]);
  nand (_03626_, _03625_, _03624_);
  nand (_03627_, _03626_, _03081_);
  not (_03628_, \oc8051_golden_model_1.IRAM[3] [0]);
  or (_03629_, _03087_, _03628_);
  nand (_03630_, _03087_, \oc8051_golden_model_1.IRAM[2] [0]);
  nand (_03631_, _03630_, _03629_);
  nand (_03632_, _03631_, _03083_);
  nand (_03633_, _03632_, _03627_);
  nand (_03634_, _03633_, _03076_);
  nand (_03635_, _03634_, _03622_);
  nand (_03636_, _03635_, _03072_);
  or (_03637_, _03089_, \oc8051_golden_model_1.IRAM[8] [0]);
  or (_03638_, _03087_, \oc8051_golden_model_1.IRAM[9] [0]);
  and (_03639_, _03638_, _03081_);
  nand (_03640_, _03639_, _03637_);
  or (_03641_, _03089_, \oc8051_golden_model_1.IRAM[10] [0]);
  or (_03642_, _03087_, \oc8051_golden_model_1.IRAM[11] [0]);
  and (_03643_, _03642_, _03083_);
  nand (_03644_, _03643_, _03641_);
  nand (_03645_, _03644_, _03640_);
  nand (_03646_, _03645_, _03076_);
  or (_03647_, _03087_, \oc8051_golden_model_1.IRAM[13] [0]);
  or (_03648_, _03089_, \oc8051_golden_model_1.IRAM[12] [0]);
  and (_03649_, _03648_, _03081_);
  nand (_03650_, _03649_, _03647_);
  or (_03651_, _03089_, \oc8051_golden_model_1.IRAM[14] [0]);
  or (_03652_, _03087_, \oc8051_golden_model_1.IRAM[15] [0]);
  and (_03653_, _03652_, _03083_);
  nand (_03654_, _03653_, _03651_);
  nand (_03655_, _03654_, _03650_);
  nand (_03656_, _03655_, _03077_);
  nand (_03657_, _03656_, _03646_);
  nand (_03658_, _03657_, _03073_);
  nand (_03659_, _03658_, _03636_);
  nand (_03660_, _03659_, _03151_);
  nand (_03661_, _03145_, \oc8051_golden_model_1.TL0 [0]);
  and (_03662_, _03168_, \oc8051_golden_model_1.SBUF [0]);
  nand (_03663_, _03195_, \oc8051_golden_model_1.SCON [0]);
  nand (_03664_, _03217_, \oc8051_golden_model_1.P0 [0]);
  nand (_03665_, _03664_, _03663_);
  nor (_03666_, _03665_, _03662_);
  and (_03667_, _03666_, _03661_);
  nand (_03668_, _03176_, \oc8051_golden_model_1.TL1 [0]);
  nand (_03669_, _03178_, \oc8051_golden_model_1.DPL [0]);
  and (_03670_, _03669_, _03668_);
  and (_03671_, _03670_, _03667_);
  nand (_03672_, _03067_, \oc8051_golden_model_1.SP [0]);
  nand (_03673_, _03184_, \oc8051_golden_model_1.TMOD [0]);
  nand (_03674_, _03187_, \oc8051_golden_model_1.TH1 [0]);
  and (_03675_, _03674_, _03673_);
  and (_03676_, _03675_, _03672_);
  nand (_03677_, _03155_, \oc8051_golden_model_1.PSW [0]);
  nand (_03678_, _03198_, \oc8051_golden_model_1.P1 [0]);
  and (_03679_, _03678_, _03677_);
  nand (_03680_, _03192_, \oc8051_golden_model_1.B [0]);
  nand (_03681_, _03220_, \oc8051_golden_model_1.TH0 [0]);
  and (_03682_, _03681_, _03680_);
  and (_03683_, _03682_, _03679_);
  nand (_03684_, _03205_, \oc8051_golden_model_1.IP [0]);
  nand (_03685_, _03208_, \oc8051_golden_model_1.P2 [0]);
  and (_03686_, _03685_, _03684_);
  nand (_03687_, _03211_, \oc8051_golden_model_1.IE [0]);
  nand (_03688_, _03213_, \oc8051_golden_model_1.P3 [0]);
  and (_03689_, _03688_, _03687_);
  and (_03690_, _03689_, _03686_);
  not (_03691_, \oc8051_golden_model_1.ACC [0]);
  or (_03692_, _03164_, _03691_);
  nand (_03693_, _03200_, \oc8051_golden_model_1.TCON [0]);
  and (_03694_, _03693_, _03692_);
  and (_03695_, _03694_, _03690_);
  and (_03696_, _03695_, _03683_);
  and (_03697_, _03696_, _03676_);
  nand (_03698_, _03227_, \oc8051_golden_model_1.PCON [0]);
  nand (_03699_, _03229_, \oc8051_golden_model_1.DPH [0]);
  and (_03700_, _03699_, _03698_);
  and (_03701_, _03700_, _03697_);
  and (_03702_, _03701_, _03671_);
  nand (_03703_, _03702_, _03660_);
  and (_03704_, _03703_, _03610_);
  nand (_03705_, _03087_, \oc8051_golden_model_1.IRAM[4] [2]);
  nand (_03706_, _03089_, \oc8051_golden_model_1.IRAM[5] [2]);
  nand (_03707_, _03706_, _03705_);
  nand (_03708_, _03707_, _03081_);
  not (_03709_, \oc8051_golden_model_1.IRAM[6] [2]);
  or (_03710_, _03089_, _03709_);
  not (_03711_, \oc8051_golden_model_1.IRAM[7] [2]);
  or (_03712_, _03087_, _03711_);
  nand (_03713_, _03712_, _03710_);
  nand (_03714_, _03713_, _03083_);
  nand (_03715_, _03714_, _03708_);
  nand (_03716_, _03715_, _03077_);
  nand (_03717_, _03089_, \oc8051_golden_model_1.IRAM[1] [2]);
  nand (_03718_, _03087_, \oc8051_golden_model_1.IRAM[0] [2]);
  nand (_03719_, _03718_, _03717_);
  nand (_03720_, _03719_, _03081_);
  not (_03721_, \oc8051_golden_model_1.IRAM[2] [2]);
  or (_03722_, _03089_, _03721_);
  not (_03723_, \oc8051_golden_model_1.IRAM[3] [2]);
  or (_03724_, _03087_, _03723_);
  nand (_03725_, _03724_, _03722_);
  nand (_03726_, _03725_, _03083_);
  nand (_03727_, _03726_, _03720_);
  nand (_03728_, _03727_, _03076_);
  nand (_03729_, _03728_, _03716_);
  nand (_03730_, _03729_, _03072_);
  or (_03731_, _03089_, \oc8051_golden_model_1.IRAM[8] [2]);
  or (_03732_, _03087_, \oc8051_golden_model_1.IRAM[9] [2]);
  and (_03733_, _03732_, _03081_);
  nand (_03734_, _03733_, _03731_);
  or (_03735_, _03089_, \oc8051_golden_model_1.IRAM[10] [2]);
  or (_03736_, _03087_, \oc8051_golden_model_1.IRAM[11] [2]);
  and (_03737_, _03736_, _03083_);
  nand (_03738_, _03737_, _03735_);
  nand (_03739_, _03738_, _03734_);
  nand (_03740_, _03739_, _03076_);
  or (_03741_, _03087_, \oc8051_golden_model_1.IRAM[13] [2]);
  or (_03742_, _03089_, \oc8051_golden_model_1.IRAM[12] [2]);
  and (_03743_, _03742_, _03081_);
  nand (_03744_, _03743_, _03741_);
  or (_03745_, _03089_, \oc8051_golden_model_1.IRAM[14] [2]);
  or (_03746_, _03087_, \oc8051_golden_model_1.IRAM[15] [2]);
  and (_03747_, _03746_, _03083_);
  nand (_03748_, _03747_, _03745_);
  nand (_03749_, _03748_, _03744_);
  nand (_03750_, _03749_, _03077_);
  nand (_03751_, _03750_, _03740_);
  nand (_03752_, _03751_, _03073_);
  nand (_03753_, _03752_, _03730_);
  nand (_03754_, _03753_, _03151_);
  and (_03755_, _03145_, \oc8051_golden_model_1.TL0 [2]);
  not (_03756_, _03755_);
  and (_03757_, _03168_, \oc8051_golden_model_1.SBUF [2]);
  not (_03758_, \oc8051_golden_model_1.ACC [2]);
  or (_03759_, _03164_, _03758_);
  not (_03760_, \oc8051_golden_model_1.PSW [2]);
  or (_03761_, _03599_, _03760_);
  nand (_03762_, _03761_, _03759_);
  nor (_03763_, _03762_, _03757_);
  and (_03765_, _03763_, _03756_);
  and (_03766_, _03176_, \oc8051_golden_model_1.TL1 [2]);
  and (_03767_, _03178_, \oc8051_golden_model_1.DPL [2]);
  nor (_03768_, _03767_, _03766_);
  and (_03769_, _03768_, _03765_);
  nand (_03770_, _03067_, \oc8051_golden_model_1.SP [2]);
  nand (_03771_, _03184_, \oc8051_golden_model_1.TMOD [2]);
  nand (_03772_, _03187_, \oc8051_golden_model_1.TH1 [2]);
  and (_03773_, _03772_, _03771_);
  and (_03774_, _03773_, _03770_);
  nand (_03775_, _03192_, \oc8051_golden_model_1.B [2]);
  nand (_03776_, _03217_, \oc8051_golden_model_1.P0 [2]);
  and (_03777_, _03776_, _03775_);
  nand (_03778_, _03195_, \oc8051_golden_model_1.SCON [2]);
  nand (_03779_, _03220_, \oc8051_golden_model_1.TH0 [2]);
  and (_03780_, _03779_, _03778_);
  and (_03781_, _03780_, _03777_);
  nand (_03782_, _03211_, \oc8051_golden_model_1.IE [2]);
  nand (_03783_, _03205_, \oc8051_golden_model_1.IP [2]);
  and (_03784_, _03783_, _03782_);
  not (_03785_, \oc8051_golden_model_1.P3 [2]);
  nand (_03786_, _03204_, _03150_);
  or (_03787_, _03786_, _03785_);
  nand (_03788_, _03208_, \oc8051_golden_model_1.P2 [2]);
  and (_03789_, _03788_, _03787_);
  and (_03790_, _03789_, _03784_);
  nand (_03791_, _03200_, \oc8051_golden_model_1.TCON [2]);
  nand (_03792_, _03198_, \oc8051_golden_model_1.P1 [2]);
  and (_03793_, _03792_, _03791_);
  and (_03794_, _03793_, _03790_);
  and (_03795_, _03794_, _03781_);
  and (_03796_, _03795_, _03774_);
  and (_03797_, _03227_, \oc8051_golden_model_1.PCON [2]);
  and (_03798_, _03229_, \oc8051_golden_model_1.DPH [2]);
  nor (_03799_, _03798_, _03797_);
  and (_03800_, _03799_, _03796_);
  and (_03801_, _03800_, _03769_);
  nand (_03802_, _03801_, _03754_);
  nand (_03803_, _03802_, _03704_);
  or (_03804_, _03803_, _03517_);
  and (_03805_, _03087_, \oc8051_golden_model_1.IRAM[4] [4]);
  and (_03806_, _03089_, \oc8051_golden_model_1.IRAM[5] [4]);
  nor (_03807_, _03806_, _03805_);
  nor (_03808_, _03807_, _03083_);
  and (_03809_, _03087_, \oc8051_golden_model_1.IRAM[6] [4]);
  and (_03810_, _03089_, \oc8051_golden_model_1.IRAM[7] [4]);
  nor (_03811_, _03810_, _03809_);
  nor (_03812_, _03811_, _03081_);
  nor (_03813_, _03812_, _03808_);
  nor (_03814_, _03813_, _03076_);
  and (_03815_, _03087_, \oc8051_golden_model_1.IRAM[0] [4]);
  and (_03816_, _03089_, \oc8051_golden_model_1.IRAM[1] [4]);
  nor (_03817_, _03816_, _03815_);
  nor (_03818_, _03817_, _03083_);
  and (_03819_, _03087_, \oc8051_golden_model_1.IRAM[2] [4]);
  and (_03820_, _03089_, \oc8051_golden_model_1.IRAM[3] [4]);
  nor (_03821_, _03820_, _03819_);
  nor (_03822_, _03821_, _03081_);
  nor (_03823_, _03822_, _03818_);
  nor (_03824_, _03823_, _03077_);
  nor (_03825_, _03824_, _03814_);
  nor (_03826_, _03825_, _03073_);
  and (_03827_, _03087_, \oc8051_golden_model_1.IRAM[8] [4]);
  and (_03828_, _03089_, \oc8051_golden_model_1.IRAM[9] [4]);
  or (_03829_, _03828_, _03827_);
  and (_03830_, _03829_, _03081_);
  and (_03831_, _03087_, \oc8051_golden_model_1.IRAM[10] [4]);
  and (_03832_, _03089_, \oc8051_golden_model_1.IRAM[11] [4]);
  or (_03833_, _03832_, _03831_);
  and (_03834_, _03833_, _03083_);
  nor (_03835_, _03834_, _03830_);
  nor (_03836_, _03835_, _03077_);
  and (_03837_, _03087_, \oc8051_golden_model_1.IRAM[12] [4]);
  and (_03838_, _03089_, \oc8051_golden_model_1.IRAM[13] [4]);
  or (_03839_, _03838_, _03837_);
  and (_03840_, _03839_, _03081_);
  and (_03841_, _03087_, \oc8051_golden_model_1.IRAM[14] [4]);
  and (_03842_, _03089_, \oc8051_golden_model_1.IRAM[15] [4]);
  or (_03843_, _03842_, _03841_);
  and (_03844_, _03843_, _03083_);
  nor (_03845_, _03844_, _03840_);
  nor (_03846_, _03845_, _03076_);
  nor (_03847_, _03846_, _03836_);
  nor (_03848_, _03847_, _03072_);
  nor (_03849_, _03848_, _03826_);
  nor (_03850_, _03849_, _02959_);
  not (_03851_, _03850_);
  and (_03852_, _03145_, \oc8051_golden_model_1.TL0 [4]);
  not (_03853_, _03852_);
  and (_03854_, _03198_, \oc8051_golden_model_1.P1 [4]);
  not (_03855_, _03854_);
  and (_03856_, _03195_, \oc8051_golden_model_1.SCON [4]);
  and (_03857_, _03220_, \oc8051_golden_model_1.TH0 [4]);
  nor (_03858_, _03857_, _03856_);
  and (_03859_, _03858_, _03855_);
  and (_03860_, _03859_, _03853_);
  and (_03861_, _03176_, \oc8051_golden_model_1.TL1 [4]);
  and (_03862_, _03178_, \oc8051_golden_model_1.DPL [4]);
  nor (_03863_, _03862_, _03861_);
  and (_03864_, _03863_, _03860_);
  and (_03865_, _03067_, \oc8051_golden_model_1.SP [4]);
  not (_03866_, _03865_);
  and (_03867_, _03184_, \oc8051_golden_model_1.TMOD [4]);
  and (_03868_, _03187_, \oc8051_golden_model_1.TH1 [4]);
  nor (_03869_, _03868_, _03867_);
  and (_03870_, _03869_, _03866_);
  not (_03871_, \oc8051_golden_model_1.ACC [4]);
  nor (_03872_, _03164_, _03871_);
  and (_03873_, _03217_, \oc8051_golden_model_1.P0 [4]);
  nor (_03874_, _03873_, _03872_);
  and (_03875_, _03155_, \oc8051_golden_model_1.PSW [4]);
  and (_03876_, _03200_, \oc8051_golden_model_1.TCON [4]);
  nor (_03877_, _03876_, _03875_);
  and (_03878_, _03877_, _03874_);
  and (_03879_, _03213_, \oc8051_golden_model_1.P3 [4]);
  and (_03880_, _03205_, \oc8051_golden_model_1.IP [4]);
  nor (_03881_, _03880_, _03879_);
  and (_03882_, _03211_, \oc8051_golden_model_1.IE [4]);
  and (_03883_, _03208_, \oc8051_golden_model_1.P2 [4]);
  nor (_03884_, _03883_, _03882_);
  and (_03885_, _03884_, _03881_);
  and (_03886_, _03192_, \oc8051_golden_model_1.B [4]);
  and (_03887_, _03168_, \oc8051_golden_model_1.SBUF [4]);
  nor (_03888_, _03887_, _03886_);
  and (_03889_, _03888_, _03885_);
  and (_03890_, _03889_, _03878_);
  and (_03891_, _03890_, _03870_);
  and (_03892_, _03227_, \oc8051_golden_model_1.PCON [4]);
  and (_03893_, _03229_, \oc8051_golden_model_1.DPH [4]);
  nor (_03894_, _03893_, _03892_);
  and (_03895_, _03894_, _03891_);
  and (_03896_, _03895_, _03864_);
  and (_03897_, _03896_, _03851_);
  or (_03898_, _03897_, _03804_);
  nor (_03899_, _03898_, _03422_);
  nand (_03900_, _03899_, _03328_);
  nand (_03901_, _03900_, _03234_);
  or (_03902_, _03900_, _03234_);
  and (_03903_, _03902_, _03901_);
  or (_03904_, _03903_, _03068_);
  or (_03905_, _03067_, \oc8051_golden_model_1.SP [7]);
  and (_03906_, _03905_, _02758_);
  and (_03907_, _03906_, _03904_);
  or (_03908_, _03907_, _02750_);
  and (_13843_[7], _03908_, _02748_);
  and (_13842_[7], \oc8051_golden_model_1.SCON [7], _13707_);
  and (_13841_[7], \oc8051_golden_model_1.SBUF [7], _13707_);
  and (_13838_[7], \oc8051_golden_model_1.PCON [7], _13707_);
  and (_03909_, _02715_, PSW_abstr[7]);
  or (_03910_, _03903_, _03599_);
  not (_03911_, \oc8051_golden_model_1.PSW [7]);
  and (_03912_, _03599_, _03911_);
  nor (_03913_, _03912_, _02715_);
  and (_03914_, _03913_, _03910_);
  or (_03915_, _03914_, _03909_);
  or (_03916_, _03915_, _12786_);
  or (_03917_, _12782_, \oc8051_golden_model_1.PSW [7]);
  and (_03918_, _03917_, _13707_);
  and (_13840_[7], _03918_, _03916_);
  and (_03919_, _02715_, P3_abstr[7]);
  or (_03920_, _03903_, _03786_);
  or (_03921_, _03213_, \oc8051_golden_model_1.P3 [7]);
  and (_03922_, _03921_, _02758_);
  and (_03923_, _03922_, _03920_);
  or (_03924_, _03923_, _03919_);
  and (_03925_, _03924_, _12782_);
  not (_03926_, \oc8051_golden_model_1.P3 [7]);
  nor (_03927_, _12782_, _03926_);
  or (_03928_, _03927_, rst);
  or (_13837_[7], _03928_, _03925_);
  and (_03929_, _02715_, P2_abstr[7]);
  not (_03930_, _03208_);
  or (_03931_, _03903_, _03930_);
  or (_03932_, _03208_, \oc8051_golden_model_1.P2 [7]);
  and (_03933_, _03932_, _02758_);
  and (_03934_, _03933_, _03931_);
  or (_03935_, _03934_, _03929_);
  and (_03936_, _03935_, _12782_);
  not (_03937_, \oc8051_golden_model_1.P2 [7]);
  nor (_03938_, _12782_, _03937_);
  or (_03939_, _03938_, rst);
  or (_13836_[7], _03939_, _03936_);
  and (_03940_, _02715_, P1_abstr[7]);
  not (_03941_, _03198_);
  or (_03942_, _03903_, _03941_);
  or (_03943_, _03198_, \oc8051_golden_model_1.P1 [7]);
  and (_03944_, _03943_, _02758_);
  and (_03945_, _03944_, _03942_);
  or (_03946_, _03945_, _03940_);
  and (_03947_, _03946_, _12782_);
  not (_03948_, \oc8051_golden_model_1.P1 [7]);
  nor (_03949_, _12782_, _03948_);
  or (_03950_, _03949_, rst);
  or (_13835_[7], _03950_, _03947_);
  and (_03951_, _02715_, P0_abstr[7]);
  not (_03952_, _03217_);
  or (_03953_, _03903_, _03952_);
  or (_03954_, _03217_, \oc8051_golden_model_1.P0 [7]);
  and (_03955_, _03954_, _02758_);
  and (_03956_, _03955_, _03953_);
  or (_03958_, _03956_, _03951_);
  and (_03959_, _03958_, _12782_);
  not (_03960_, \oc8051_golden_model_1.P0 [7]);
  nor (_03961_, _12782_, _03960_);
  or (_03962_, _03961_, rst);
  or (_13834_[7], _03962_, _03959_);
  and (_13833_[7], \oc8051_golden_model_1.IP [7], _13707_);
  and (_13832_[7], \oc8051_golden_model_1.IE [7], _13707_);
  or (_03963_, _12782_, \oc8051_golden_model_1.DPH [7]);
  and (_03964_, _03963_, _13707_);
  and (_03965_, _02715_, DPH_abstr[7]);
  or (_03966_, _03965_, _12786_);
  not (_03967_, _03229_);
  or (_03968_, _03903_, _03967_);
  or (_03969_, _03229_, \oc8051_golden_model_1.DPH [7]);
  and (_03970_, _03969_, _02758_);
  and (_03971_, _03970_, _03968_);
  or (_03972_, _03971_, _03966_);
  and (_13830_[7], _03972_, _03964_);
  or (_03973_, _12782_, \oc8051_golden_model_1.DPL [7]);
  and (_03974_, _03973_, _13707_);
  not (_03975_, _03178_);
  or (_03976_, _03903_, _03975_);
  or (_03977_, _03178_, \oc8051_golden_model_1.DPL [7]);
  and (_03978_, _03977_, _02758_);
  and (_03979_, _03978_, _03976_);
  and (_03980_, _02715_, DPL_abstr[7]);
  or (_03981_, _03980_, _12786_);
  or (_03982_, _03981_, _03979_);
  and (_13831_[7], _03982_, _03974_);
  nor (_03983_, _12782_, _03158_);
  and (_03984_, _03164_, \oc8051_golden_model_1.ACC [7]);
  not (_03985_, _03984_);
  not (_03986_, _03164_);
  nand (_03987_, _03903_, _03986_);
  nand (_03988_, _03987_, _03985_);
  or (_03989_, _03988_, _02715_);
  or (_03990_, _02758_, ACC_abstr[7]);
  and (_03991_, _03990_, _12782_);
  and (_03992_, _03991_, _03989_);
  or (_03993_, _03992_, _03983_);
  and (_13828_[7], _03993_, _13707_);
  or (_03994_, _12782_, \oc8051_golden_model_1.B [7]);
  and (_03995_, _03994_, _13707_);
  not (_03996_, _03192_);
  or (_03997_, _03903_, _03996_);
  or (_03998_, _03192_, \oc8051_golden_model_1.B [7]);
  and (_03999_, _03998_, _02758_);
  and (_04000_, _03999_, _03997_);
  and (_04001_, _02715_, B_abstr[7]);
  or (_04002_, _04001_, _12786_);
  or (_04003_, _04002_, _04000_);
  and (_13829_[7], _04003_, _03995_);
  nor (_04004_, _02959_, _02715_);
  and (_04005_, _04004_, _03029_);
  nor (_04006_, _04004_, WR_ADDR_ABSTR_IRAM_0[0]);
  nor (_04007_, _04006_, _04005_);
  and (_04008_, _04004_, _03064_);
  nor (_04009_, _04004_, WR_ADDR_ABSTR_IRAM_0[1]);
  nor (_04010_, _04009_, _04008_);
  not (_04011_, _00002_);
  and (_04012_, _02715_, WR_COND_ABSTR_IRAM_0);
  nor (_04013_, _04012_, _04004_);
  nor (_04014_, _04013_, _04011_);
  and (_04015_, _04014_, _04010_);
  and (_04016_, _04015_, _04007_);
  and (_04017_, _04004_, _02829_);
  nor (_04018_, _04004_, WR_ADDR_ABSTR_IRAM_0[2]);
  nor (_04019_, _04018_, _04017_);
  and (_04020_, _04004_, _02861_);
  nor (_04021_, _04004_, WR_ADDR_ABSTR_IRAM_0[3]);
  nor (_04022_, _04021_, _04020_);
  and (_04023_, _04022_, _04014_);
  and (_04024_, _04023_, _04019_);
  and (_04025_, _04024_, _04016_);
  or (_04026_, _04025_, \oc8051_golden_model_1.IRAM[15] [7]);
  and (_04027_, _00002_, WR_COND_ABSTR_IRAM_1);
  and (_04028_, _04027_, _02715_);
  and (_04029_, _04028_, WR_ADDR_ABSTR_IRAM_1[2]);
  and (_04030_, _04029_, WR_ADDR_ABSTR_IRAM_1[3]);
  and (_04031_, _04028_, WR_ADDR_ABSTR_IRAM_1[1]);
  and (_04032_, _04031_, WR_ADDR_ABSTR_IRAM_1[0]);
  and (_04033_, _04032_, _04030_);
  not (_04034_, _04033_);
  and (_04035_, _04034_, _04026_);
  not (_04036_, _04025_);
  not (_04037_, _04004_);
  or (_04038_, _04037_, _03903_);
  or (_04039_, _04004_, WR_DATA_ABSTR_IRAM_0[7]);
  and (_04040_, _04039_, _04014_);
  and (_04041_, _04040_, _04038_);
  or (_04042_, _04041_, _04036_);
  and (_04043_, _04042_, _04035_);
  and (_04044_, _04028_, WR_DATA_ABSTR_IRAM_1[7]);
  and (_04045_, _04044_, _04033_);
  or (_13905_[7], _04045_, _04043_);
  and (_04046_, _04014_, _04007_);
  nor (_04047_, _04046_, _04015_);
  and (_04048_, _04019_, _04014_);
  nor (_04049_, _04048_, _04023_);
  and (_04050_, _04049_, _04014_);
  and (_04051_, _04050_, _04047_);
  not (_04052_, _04051_);
  and (_04053_, _03702_, _03660_);
  or (_04054_, _04037_, _04053_);
  or (_04055_, _04004_, WR_DATA_ABSTR_IRAM_0[0]);
  and (_04056_, _04055_, _04014_);
  and (_04057_, _04056_, _04054_);
  or (_04058_, _04057_, _04052_);
  and (_04059_, _04028_, WR_ADDR_ABSTR_IRAM_1[0]);
  nor (_04060_, _04059_, _04031_);
  and (_04061_, _04028_, WR_ADDR_ABSTR_IRAM_1[3]);
  nor (_04062_, _04061_, _04029_);
  and (_04063_, _04062_, _04060_);
  and (_04064_, _04063_, _04028_);
  not (_04065_, _04064_);
  or (_04066_, _04051_, \oc8051_golden_model_1.IRAM[0] [0]);
  and (_04067_, _04066_, _04065_);
  and (_04068_, _04067_, _04058_);
  and (_04069_, _04064_, WR_DATA_ABSTR_IRAM_1[0]);
  or (_13852_, _04069_, _04068_);
  nand (_04070_, _03703_, _03610_);
  or (_04071_, _03703_, _03610_);
  nand (_04072_, _04071_, _04070_);
  nand (_04073_, _04072_, _04004_);
  or (_04074_, _04004_, WR_DATA_ABSTR_IRAM_0[1]);
  and (_04075_, _04074_, _04014_);
  and (_04076_, _04075_, _04073_);
  or (_04077_, _04076_, _04052_);
  or (_04078_, _04051_, \oc8051_golden_model_1.IRAM[0] [1]);
  and (_04079_, _04078_, _04065_);
  and (_04080_, _04079_, _04077_);
  and (_04081_, _04064_, WR_DATA_ABSTR_IRAM_1[1]);
  or (_13853_, _04081_, _04080_);
  or (_04082_, _03802_, _03704_);
  and (_04083_, _04082_, _03803_);
  or (_04084_, _04083_, _04037_);
  or (_04085_, _04004_, WR_DATA_ABSTR_IRAM_0[2]);
  and (_04086_, _04085_, _04014_);
  and (_04087_, _04086_, _04084_);
  or (_04088_, _04087_, _04052_);
  or (_04089_, _04051_, \oc8051_golden_model_1.IRAM[0] [2]);
  and (_04090_, _04089_, _04065_);
  and (_04091_, _04090_, _04088_);
  and (_04092_, _04064_, WR_DATA_ABSTR_IRAM_1[2]);
  or (_13854_, _04092_, _04091_);
  not (_04093_, _03517_);
  and (_04094_, _03802_, _03704_);
  or (_04095_, _04094_, _04093_);
  nand (_04096_, _04095_, _03804_);
  nand (_04097_, _04096_, _04004_);
  or (_04098_, _04004_, WR_DATA_ABSTR_IRAM_0[3]);
  and (_04099_, _04098_, _04014_);
  and (_04100_, _04099_, _04097_);
  or (_04101_, _04100_, _04052_);
  or (_04102_, _04051_, \oc8051_golden_model_1.IRAM[0] [3]);
  and (_04103_, _04102_, _04065_);
  and (_04104_, _04103_, _04101_);
  and (_04105_, _04064_, WR_DATA_ABSTR_IRAM_1[3]);
  or (_13855_, _04105_, _04104_);
  nand (_04106_, _03897_, _03804_);
  nand (_04107_, _04106_, _03898_);
  nand (_04108_, _04107_, _04004_);
  or (_04109_, _04004_, WR_DATA_ABSTR_IRAM_0[4]);
  and (_04110_, _04109_, _04014_);
  and (_04111_, _04110_, _04108_);
  or (_04112_, _04111_, _04052_);
  or (_04113_, _04051_, \oc8051_golden_model_1.IRAM[0] [4]);
  and (_04114_, _04113_, _04065_);
  and (_04115_, _04114_, _04112_);
  and (_04116_, _04064_, WR_DATA_ABSTR_IRAM_1[4]);
  or (_13856_, _04116_, _04115_);
  and (_04117_, _03898_, _03422_);
  nor (_04118_, _04117_, _03899_);
  or (_04119_, _04118_, _04037_);
  or (_04120_, _04004_, WR_DATA_ABSTR_IRAM_0[5]);
  and (_04121_, _04120_, _04014_);
  and (_04122_, _04121_, _04119_);
  or (_04123_, _04122_, _04052_);
  or (_04124_, _04051_, \oc8051_golden_model_1.IRAM[0] [5]);
  and (_04125_, _04124_, _04065_);
  and (_04126_, _04125_, _04123_);
  and (_04127_, _04064_, WR_DATA_ABSTR_IRAM_1[5]);
  or (_13857_, _04127_, _04126_);
  or (_04128_, _03899_, _03328_);
  and (_04129_, _04128_, _03900_);
  or (_04130_, _04129_, _04037_);
  or (_04131_, _04004_, WR_DATA_ABSTR_IRAM_0[6]);
  and (_04132_, _04131_, _04014_);
  and (_04133_, _04132_, _04130_);
  or (_04134_, _04133_, _04052_);
  or (_04135_, _04051_, \oc8051_golden_model_1.IRAM[0] [6]);
  and (_04136_, _04135_, _04065_);
  and (_04137_, _04136_, _04134_);
  and (_04138_, _04064_, WR_DATA_ABSTR_IRAM_1[6]);
  or (_13858_, _04138_, _04137_);
  or (_04139_, _04052_, _04041_);
  or (_04140_, _04051_, \oc8051_golden_model_1.IRAM[0] [7]);
  and (_04141_, _04140_, _04065_);
  and (_04142_, _04141_, _04139_);
  and (_04144_, _04064_, WR_DATA_ABSTR_IRAM_1[7]);
  or (_13859_, _04144_, _04142_);
  not (_04145_, _04010_);
  and (_04146_, _04046_, _04145_);
  and (_04147_, _04146_, _04049_);
  not (_04148_, _04147_);
  or (_04149_, _04148_, _04057_);
  not (_04150_, WR_ADDR_ABSTR_IRAM_1[1]);
  and (_04151_, _04059_, _04150_);
  and (_04152_, _04151_, _04062_);
  not (_04153_, _04152_);
  or (_04154_, _04147_, \oc8051_golden_model_1.IRAM[1] [0]);
  and (_04155_, _04154_, _04153_);
  and (_04156_, _04155_, _04149_);
  and (_04157_, _04028_, WR_DATA_ABSTR_IRAM_1[0]);
  and (_04158_, _04152_, _04157_);
  or (_13860_, _04158_, _04156_);
  or (_04159_, _04148_, _04076_);
  or (_04160_, _04147_, \oc8051_golden_model_1.IRAM[1] [1]);
  and (_04161_, _04160_, _04153_);
  and (_04162_, _04161_, _04159_);
  and (_04163_, _04028_, WR_DATA_ABSTR_IRAM_1[1]);
  and (_04164_, _04163_, _04152_);
  or (_13861_, _04164_, _04162_);
  or (_04165_, _04148_, _04087_);
  or (_04166_, _04147_, \oc8051_golden_model_1.IRAM[1] [2]);
  and (_04167_, _04166_, _04153_);
  and (_04168_, _04167_, _04165_);
  and (_04169_, _04028_, WR_DATA_ABSTR_IRAM_1[2]);
  and (_04170_, _04152_, _04169_);
  or (_13862_, _04170_, _04168_);
  or (_04171_, _04148_, _04100_);
  or (_04172_, _04147_, \oc8051_golden_model_1.IRAM[1] [3]);
  and (_04173_, _04172_, _04153_);
  and (_04174_, _04173_, _04171_);
  and (_04175_, _04028_, WR_DATA_ABSTR_IRAM_1[3]);
  and (_04176_, _04152_, _04175_);
  or (_13863_, _04176_, _04174_);
  or (_04177_, _04148_, _04111_);
  or (_04178_, _04147_, \oc8051_golden_model_1.IRAM[1] [4]);
  and (_04179_, _04178_, _04153_);
  and (_04180_, _04179_, _04177_);
  and (_04181_, _04028_, WR_DATA_ABSTR_IRAM_1[4]);
  and (_04182_, _04181_, _04152_);
  or (_13864_, _04182_, _04180_);
  or (_04183_, _04148_, _04122_);
  or (_04184_, _04147_, \oc8051_golden_model_1.IRAM[1] [5]);
  and (_04185_, _04184_, _04153_);
  and (_04186_, _04185_, _04183_);
  and (_04187_, _04028_, WR_DATA_ABSTR_IRAM_1[5]);
  and (_04188_, _04187_, _04152_);
  or (_13865_, _04188_, _04186_);
  or (_04189_, _04148_, _04133_);
  or (_04190_, _04147_, \oc8051_golden_model_1.IRAM[1] [6]);
  and (_04191_, _04190_, _04153_);
  and (_04192_, _04191_, _04189_);
  and (_04193_, _04028_, WR_DATA_ABSTR_IRAM_1[6]);
  and (_04194_, _04152_, _04193_);
  or (_13866_, _04194_, _04192_);
  or (_04195_, _04148_, _04041_);
  or (_04196_, _04147_, \oc8051_golden_model_1.IRAM[1] [7]);
  and (_04197_, _04196_, _04153_);
  and (_04198_, _04197_, _04195_);
  and (_04199_, _04152_, _04044_);
  or (_13867_, _04199_, _04198_);
  not (_04200_, WR_ADDR_ABSTR_IRAM_1[0]);
  and (_04201_, _04031_, _04200_);
  and (_04202_, _04201_, _04062_);
  and (_04203_, _04202_, _04157_);
  not (_04204_, _04007_);
  and (_04205_, _04015_, _04204_);
  and (_04206_, _04205_, _04049_);
  not (_04207_, _04206_);
  or (_04208_, _04207_, _04057_);
  not (_04209_, _04202_);
  or (_04210_, _04206_, \oc8051_golden_model_1.IRAM[2] [0]);
  and (_04211_, _04210_, _04209_);
  and (_04212_, _04211_, _04208_);
  or (_13868_, _04212_, _04203_);
  or (_04213_, _04207_, _04076_);
  or (_04214_, _04206_, \oc8051_golden_model_1.IRAM[2] [1]);
  and (_04215_, _04214_, _04209_);
  and (_04216_, _04215_, _04213_);
  and (_04217_, _04202_, _04163_);
  or (_13869_, _04217_, _04216_);
  and (_04218_, _04202_, _04169_);
  or (_04219_, _04207_, _04087_);
  or (_04220_, _04206_, \oc8051_golden_model_1.IRAM[2] [2]);
  and (_04221_, _04220_, _04209_);
  and (_04222_, _04221_, _04219_);
  or (_13870_, _04222_, _04218_);
  and (_04223_, _04202_, _04175_);
  or (_04224_, _04207_, _04100_);
  or (_04225_, _04206_, \oc8051_golden_model_1.IRAM[2] [3]);
  and (_04226_, _04225_, _04209_);
  and (_04227_, _04226_, _04224_);
  or (_13871_, _04227_, _04223_);
  or (_04228_, _04207_, _04111_);
  or (_04229_, _04206_, \oc8051_golden_model_1.IRAM[2] [4]);
  and (_04230_, _04229_, _04209_);
  and (_04231_, _04230_, _04228_);
  and (_04232_, _04202_, _04181_);
  or (_13872_, _04232_, _04231_);
  or (_04233_, _04207_, _04122_);
  or (_04234_, _04206_, \oc8051_golden_model_1.IRAM[2] [5]);
  and (_04235_, _04234_, _04209_);
  and (_04236_, _04235_, _04233_);
  and (_04237_, _04202_, _04187_);
  or (_13873_, _04237_, _04236_);
  and (_04238_, _04202_, _04193_);
  or (_04239_, _04207_, _04133_);
  or (_04240_, _04206_, \oc8051_golden_model_1.IRAM[2] [6]);
  and (_04241_, _04240_, _04209_);
  and (_04242_, _04241_, _04239_);
  or (_13874_, _04242_, _04238_);
  or (_04243_, _04207_, _04041_);
  or (_04244_, _04206_, \oc8051_golden_model_1.IRAM[2] [7]);
  and (_04245_, _04244_, _04209_);
  and (_04246_, _04245_, _04243_);
  and (_04247_, _04202_, _04044_);
  or (_13875_, _04247_, _04246_);
  and (_04248_, _04049_, _04016_);
  or (_04249_, _04248_, \oc8051_golden_model_1.IRAM[3] [0]);
  and (_04250_, _04062_, _04032_);
  not (_04251_, _04250_);
  and (_04252_, _04251_, _04249_);
  not (_04253_, _04248_);
  or (_04254_, _04253_, _04057_);
  and (_04255_, _04254_, _04252_);
  and (_04256_, _04250_, _04157_);
  or (_13876_, _04256_, _04255_);
  or (_04257_, _04248_, \oc8051_golden_model_1.IRAM[3] [1]);
  and (_04258_, _04257_, _04251_);
  or (_04259_, _04253_, _04076_);
  and (_04260_, _04259_, _04258_);
  and (_04261_, _04250_, _04163_);
  or (_13877_, _04261_, _04260_);
  or (_04262_, _04248_, \oc8051_golden_model_1.IRAM[3] [2]);
  and (_04263_, _04262_, _04251_);
  or (_04264_, _04253_, _04087_);
  and (_04265_, _04264_, _04263_);
  and (_04266_, _04250_, _04169_);
  or (_13878_, _04266_, _04265_);
  or (_04267_, _04248_, \oc8051_golden_model_1.IRAM[3] [3]);
  and (_04268_, _04267_, _04251_);
  or (_04269_, _04253_, _04100_);
  and (_04270_, _04269_, _04268_);
  and (_04271_, _04250_, _04175_);
  or (_13879_, _04271_, _04270_);
  or (_04272_, _04248_, \oc8051_golden_model_1.IRAM[3] [4]);
  and (_04273_, _04272_, _04251_);
  or (_04274_, _04253_, _04111_);
  and (_04275_, _04274_, _04273_);
  and (_04276_, _04250_, _04181_);
  or (_13880_, _04276_, _04275_);
  or (_04277_, _04248_, \oc8051_golden_model_1.IRAM[3] [5]);
  and (_04278_, _04277_, _04251_);
  or (_04279_, _04253_, _04122_);
  and (_04280_, _04279_, _04278_);
  and (_04281_, _04250_, _04187_);
  or (_13881_, _04281_, _04280_);
  or (_04282_, _04248_, \oc8051_golden_model_1.IRAM[3] [6]);
  and (_04283_, _04282_, _04251_);
  or (_04284_, _04253_, _04133_);
  and (_04285_, _04284_, _04283_);
  and (_04286_, _04250_, _04193_);
  or (_13882_, _04286_, _04285_);
  or (_04287_, _04248_, \oc8051_golden_model_1.IRAM[3] [7]);
  and (_04288_, _04287_, _04251_);
  or (_04289_, _04253_, _04041_);
  and (_04290_, _04289_, _04288_);
  and (_04291_, _04250_, _04044_);
  or (_13883_, _04291_, _04290_);
  not (_04292_, _04022_);
  and (_04293_, _04048_, _04292_);
  and (_04294_, _04293_, _04047_);
  not (_04295_, _04294_);
  or (_04296_, _04295_, _04057_);
  not (_04297_, WR_ADDR_ABSTR_IRAM_1[3]);
  and (_04298_, _04029_, _04297_);
  and (_04299_, _04298_, _04060_);
  not (_04300_, _04299_);
  or (_04301_, _04294_, \oc8051_golden_model_1.IRAM[4] [0]);
  and (_04302_, _04301_, _04300_);
  and (_04303_, _04302_, _04296_);
  and (_04304_, _04299_, _04157_);
  or (_13906_[0], _04304_, _04303_);
  or (_04305_, _04295_, _04076_);
  or (_04306_, _04294_, \oc8051_golden_model_1.IRAM[4] [1]);
  and (_04307_, _04306_, _04300_);
  and (_04308_, _04307_, _04305_);
  and (_04309_, _04299_, _04163_);
  or (_13906_[1], _04309_, _04308_);
  or (_04310_, _04295_, _04087_);
  or (_04311_, _04294_, \oc8051_golden_model_1.IRAM[4] [2]);
  and (_04312_, _04311_, _04300_);
  and (_04313_, _04312_, _04310_);
  and (_04314_, _04299_, _04169_);
  or (_13906_[2], _04314_, _04313_);
  or (_04315_, _04295_, _04100_);
  or (_04317_, _04294_, \oc8051_golden_model_1.IRAM[4] [3]);
  and (_04318_, _04317_, _04300_);
  and (_04319_, _04318_, _04315_);
  and (_04320_, _04299_, _04175_);
  or (_13906_[3], _04320_, _04319_);
  or (_04321_, _04295_, _04111_);
  or (_04322_, _04294_, \oc8051_golden_model_1.IRAM[4] [4]);
  and (_04323_, _04322_, _04300_);
  and (_04324_, _04323_, _04321_);
  and (_04325_, _04299_, _04181_);
  or (_13906_[4], _04325_, _04324_);
  or (_04326_, _04295_, _04122_);
  or (_04327_, _04294_, \oc8051_golden_model_1.IRAM[4] [5]);
  and (_04328_, _04327_, _04300_);
  and (_04329_, _04328_, _04326_);
  and (_04330_, _04299_, _04187_);
  or (_13906_[5], _04330_, _04329_);
  or (_04331_, _04295_, _04133_);
  or (_04332_, _04294_, \oc8051_golden_model_1.IRAM[4] [6]);
  and (_04333_, _04332_, _04300_);
  and (_04334_, _04333_, _04331_);
  and (_04335_, _04299_, _04193_);
  or (_13906_[6], _04335_, _04334_);
  or (_04336_, _04295_, _04041_);
  or (_04337_, _04294_, \oc8051_golden_model_1.IRAM[4] [7]);
  and (_04338_, _04337_, _04300_);
  and (_04339_, _04338_, _04336_);
  and (_04340_, _04299_, _04044_);
  or (_13906_[7], _04340_, _04339_);
  and (_04341_, _04293_, _04146_);
  not (_04342_, _04341_);
  or (_04343_, _04342_, _04057_);
  and (_04344_, _04298_, _04151_);
  not (_04345_, _04344_);
  or (_04346_, _04341_, \oc8051_golden_model_1.IRAM[5] [0]);
  and (_04347_, _04346_, _04345_);
  and (_04348_, _04347_, _04343_);
  and (_04349_, _04344_, _04157_);
  or (_13907_[0], _04349_, _04348_);
  or (_04350_, _04342_, _04076_);
  or (_04351_, _04341_, \oc8051_golden_model_1.IRAM[5] [1]);
  and (_04352_, _04351_, _04345_);
  and (_04353_, _04352_, _04350_);
  and (_04354_, _04344_, _04163_);
  or (_13907_[1], _04354_, _04353_);
  or (_04355_, _04342_, _04087_);
  or (_04356_, _04341_, \oc8051_golden_model_1.IRAM[5] [2]);
  and (_04357_, _04356_, _04345_);
  and (_04358_, _04357_, _04355_);
  and (_04359_, _04344_, _04169_);
  or (_13907_[2], _04359_, _04358_);
  or (_04360_, _04342_, _04100_);
  or (_04361_, _04341_, \oc8051_golden_model_1.IRAM[5] [3]);
  and (_04362_, _04361_, _04345_);
  and (_04363_, _04362_, _04360_);
  and (_04364_, _04344_, _04175_);
  or (_13907_[3], _04364_, _04363_);
  or (_04365_, _04342_, _04111_);
  or (_04366_, _04341_, \oc8051_golden_model_1.IRAM[5] [4]);
  and (_04367_, _04366_, _04345_);
  and (_04368_, _04367_, _04365_);
  and (_04369_, _04344_, _04181_);
  or (_13907_[4], _04369_, _04368_);
  or (_04370_, _04342_, _04122_);
  or (_04371_, _04341_, \oc8051_golden_model_1.IRAM[5] [5]);
  and (_04372_, _04371_, _04345_);
  and (_04373_, _04372_, _04370_);
  and (_04374_, _04344_, _04187_);
  or (_13907_[5], _04374_, _04373_);
  or (_04375_, _04342_, _04133_);
  or (_04376_, _04341_, \oc8051_golden_model_1.IRAM[5] [6]);
  and (_04377_, _04376_, _04345_);
  and (_04378_, _04377_, _04375_);
  and (_04379_, _04344_, _04193_);
  or (_13907_[6], _04379_, _04378_);
  or (_04380_, _04342_, _04041_);
  or (_04381_, _04341_, \oc8051_golden_model_1.IRAM[5] [7]);
  and (_04382_, _04381_, _04345_);
  and (_04383_, _04382_, _04380_);
  and (_04384_, _04344_, _04044_);
  or (_13907_[7], _04384_, _04383_);
  and (_04385_, _04293_, _04205_);
  not (_04386_, _04385_);
  or (_04387_, _04386_, _04057_);
  and (_04388_, _04298_, _04201_);
  not (_04389_, _04388_);
  or (_04390_, _04385_, \oc8051_golden_model_1.IRAM[6] [0]);
  and (_04391_, _04390_, _04389_);
  and (_04392_, _04391_, _04387_);
  and (_04393_, _04388_, _04157_);
  or (_13908_[0], _04393_, _04392_);
  or (_04394_, _04386_, _04076_);
  or (_04395_, _04385_, \oc8051_golden_model_1.IRAM[6] [1]);
  and (_04396_, _04395_, _04389_);
  and (_04397_, _04396_, _04394_);
  and (_04398_, _04388_, _04163_);
  or (_13908_[1], _04398_, _04397_);
  or (_04399_, _04386_, _04087_);
  or (_04400_, _04385_, \oc8051_golden_model_1.IRAM[6] [2]);
  and (_04401_, _04400_, _04389_);
  and (_04403_, _04401_, _04399_);
  and (_04404_, _04388_, _04169_);
  or (_13908_[2], _04404_, _04403_);
  or (_04405_, _04386_, _04100_);
  or (_04406_, _04385_, \oc8051_golden_model_1.IRAM[6] [3]);
  and (_04407_, _04406_, _04389_);
  and (_04408_, _04407_, _04405_);
  and (_04409_, _04388_, _04175_);
  or (_13908_[3], _04409_, _04408_);
  or (_04410_, _04386_, _04111_);
  or (_04411_, _04385_, \oc8051_golden_model_1.IRAM[6] [4]);
  and (_04412_, _04411_, _04389_);
  and (_04413_, _04412_, _04410_);
  and (_04414_, _04388_, _04181_);
  or (_13908_[4], _04414_, _04413_);
  or (_04415_, _04386_, _04122_);
  or (_04416_, _04385_, \oc8051_golden_model_1.IRAM[6] [5]);
  and (_04417_, _04416_, _04389_);
  and (_04418_, _04417_, _04415_);
  and (_04419_, _04388_, _04187_);
  or (_13908_[5], _04419_, _04418_);
  or (_04420_, _04386_, _04133_);
  or (_04421_, _04385_, \oc8051_golden_model_1.IRAM[6] [6]);
  and (_04422_, _04421_, _04389_);
  and (_04423_, _04422_, _04420_);
  and (_04424_, _04388_, _04193_);
  or (_13908_[6], _04424_, _04423_);
  or (_04425_, _04386_, _04041_);
  or (_04426_, _04385_, \oc8051_golden_model_1.IRAM[6] [7]);
  and (_04427_, _04426_, _04389_);
  and (_04428_, _04427_, _04425_);
  and (_04429_, _04388_, _04044_);
  or (_13908_[7], _04429_, _04428_);
  and (_04430_, _04293_, _04016_);
  or (_04431_, _04430_, \oc8051_golden_model_1.IRAM[7] [0]);
  and (_04432_, _04298_, _04032_);
  not (_04433_, _04432_);
  and (_04434_, _04433_, _04431_);
  not (_04435_, _04430_);
  or (_04436_, _04435_, _04057_);
  and (_04437_, _04436_, _04434_);
  and (_04438_, _04432_, _04157_);
  or (_13884_, _04438_, _04437_);
  or (_04439_, _04430_, \oc8051_golden_model_1.IRAM[7] [1]);
  and (_04440_, _04439_, _04433_);
  or (_04441_, _04435_, _04076_);
  and (_04442_, _04441_, _04440_);
  and (_04443_, _04432_, _04163_);
  or (_13885_, _04443_, _04442_);
  or (_04444_, _04430_, \oc8051_golden_model_1.IRAM[7] [2]);
  and (_04445_, _04444_, _04433_);
  or (_04446_, _04435_, _04087_);
  and (_04447_, _04446_, _04445_);
  and (_04448_, _04432_, _04169_);
  or (_13886_, _04448_, _04447_);
  or (_04449_, _04430_, \oc8051_golden_model_1.IRAM[7] [3]);
  and (_04450_, _04449_, _04433_);
  or (_04451_, _04435_, _04100_);
  and (_04452_, _04451_, _04450_);
  and (_04453_, _04432_, _04175_);
  or (_13887_, _04453_, _04452_);
  or (_04454_, _04430_, \oc8051_golden_model_1.IRAM[7] [4]);
  and (_04455_, _04454_, _04433_);
  or (_04456_, _04435_, _04111_);
  and (_04457_, _04456_, _04455_);
  and (_04458_, _04432_, _04181_);
  or (_13888_, _04458_, _04457_);
  or (_04459_, _04430_, \oc8051_golden_model_1.IRAM[7] [5]);
  and (_04460_, _04459_, _04433_);
  or (_04461_, _04435_, _04122_);
  and (_04462_, _04461_, _04460_);
  and (_04463_, _04432_, _04187_);
  or (_13889_, _04463_, _04462_);
  or (_04464_, _04430_, \oc8051_golden_model_1.IRAM[7] [6]);
  and (_04465_, _04464_, _04433_);
  or (_04466_, _04435_, _04133_);
  and (_04467_, _04466_, _04465_);
  and (_04468_, _04432_, _04193_);
  or (_13890_, _04468_, _04467_);
  or (_04469_, _04430_, \oc8051_golden_model_1.IRAM[7] [7]);
  and (_04470_, _04469_, _04433_);
  or (_04471_, _04435_, _04041_);
  and (_04472_, _04471_, _04470_);
  and (_04473_, _04432_, _04044_);
  or (_13891_, _04473_, _04472_);
  not (_04474_, _04019_);
  and (_04475_, _04023_, _04474_);
  and (_04476_, _04475_, _04047_);
  not (_04477_, _04476_);
  or (_04478_, _04477_, _04057_);
  not (_04479_, WR_ADDR_ABSTR_IRAM_1[2]);
  and (_04480_, _04061_, _04479_);
  and (_04481_, _04480_, _04060_);
  not (_04482_, _04481_);
  or (_04483_, _04476_, \oc8051_golden_model_1.IRAM[8] [0]);
  and (_04484_, _04483_, _04482_);
  and (_04485_, _04484_, _04478_);
  and (_04486_, _04481_, _04157_);
  or (_13909_[0], _04486_, _04485_);
  or (_04487_, _04477_, _04076_);
  or (_04489_, _04476_, \oc8051_golden_model_1.IRAM[8] [1]);
  and (_04490_, _04489_, _04482_);
  and (_04491_, _04490_, _04487_);
  and (_04492_, _04481_, _04163_);
  or (_13909_[1], _04492_, _04491_);
  or (_04493_, _04477_, _04087_);
  or (_04494_, _04476_, \oc8051_golden_model_1.IRAM[8] [2]);
  and (_04495_, _04494_, _04482_);
  and (_04496_, _04495_, _04493_);
  and (_04497_, _04481_, _04169_);
  or (_13909_[2], _04497_, _04496_);
  or (_04498_, _04477_, _04100_);
  or (_04499_, _04476_, \oc8051_golden_model_1.IRAM[8] [3]);
  and (_04500_, _04499_, _04482_);
  and (_04501_, _04500_, _04498_);
  and (_04502_, _04481_, _04175_);
  or (_13909_[3], _04502_, _04501_);
  or (_04503_, _04477_, _04111_);
  or (_04504_, _04476_, \oc8051_golden_model_1.IRAM[8] [4]);
  and (_04505_, _04504_, _04482_);
  and (_04506_, _04505_, _04503_);
  and (_04507_, _04481_, _04181_);
  or (_13909_[4], _04507_, _04506_);
  or (_04508_, _04477_, _04122_);
  or (_04509_, _04476_, \oc8051_golden_model_1.IRAM[8] [5]);
  and (_04510_, _04509_, _04482_);
  and (_04511_, _04510_, _04508_);
  and (_04512_, _04481_, _04187_);
  or (_13909_[5], _04512_, _04511_);
  or (_04513_, _04477_, _04133_);
  or (_04514_, _04476_, \oc8051_golden_model_1.IRAM[8] [6]);
  and (_04515_, _04514_, _04482_);
  and (_04516_, _04515_, _04513_);
  and (_04517_, _04481_, _04193_);
  or (_13909_[6], _04517_, _04516_);
  or (_04518_, _04477_, _04041_);
  or (_04519_, _04476_, \oc8051_golden_model_1.IRAM[8] [7]);
  and (_04520_, _04519_, _04482_);
  and (_04521_, _04520_, _04518_);
  and (_04522_, _04481_, _04044_);
  or (_13909_[7], _04522_, _04521_);
  and (_04523_, _04475_, _04146_);
  not (_04524_, _04523_);
  or (_04525_, _04524_, _04057_);
  and (_04526_, _04480_, _04151_);
  not (_04527_, _04526_);
  or (_04528_, _04523_, \oc8051_golden_model_1.IRAM[9] [0]);
  and (_04529_, _04528_, _04527_);
  and (_04530_, _04529_, _04525_);
  and (_04531_, _04526_, _04157_);
  or (_13892_, _04531_, _04530_);
  or (_04532_, _04524_, _04076_);
  or (_04533_, _04523_, \oc8051_golden_model_1.IRAM[9] [1]);
  and (_04534_, _04533_, _04527_);
  and (_04535_, _04534_, _04532_);
  and (_04536_, _04526_, _04163_);
  or (_13893_, _04536_, _04535_);
  or (_04537_, _04524_, _04087_);
  or (_04538_, _04523_, \oc8051_golden_model_1.IRAM[9] [2]);
  and (_04539_, _04538_, _04527_);
  and (_04540_, _04539_, _04537_);
  and (_04541_, _04526_, _04169_);
  or (_13894_, _04541_, _04540_);
  or (_04542_, _04524_, _04100_);
  or (_04543_, _04523_, \oc8051_golden_model_1.IRAM[9] [3]);
  and (_04544_, _04543_, _04527_);
  and (_04545_, _04544_, _04542_);
  and (_04546_, _04526_, _04175_);
  or (_13895_, _04546_, _04545_);
  or (_04547_, _04524_, _04111_);
  or (_04548_, _04523_, \oc8051_golden_model_1.IRAM[9] [4]);
  and (_04549_, _04548_, _04527_);
  and (_04550_, _04549_, _04547_);
  and (_04551_, _04526_, _04181_);
  or (_13896_, _04551_, _04550_);
  or (_04552_, _04524_, _04122_);
  or (_04553_, _04523_, \oc8051_golden_model_1.IRAM[9] [5]);
  and (_04554_, _04553_, _04527_);
  and (_04555_, _04554_, _04552_);
  and (_04556_, _04526_, _04187_);
  or (_13897_, _04556_, _04555_);
  or (_04557_, _04524_, _04133_);
  or (_04558_, _04523_, \oc8051_golden_model_1.IRAM[9] [6]);
  and (_04559_, _04558_, _04527_);
  and (_04560_, _04559_, _04557_);
  and (_04561_, _04526_, _04193_);
  or (_13898_, _04561_, _04560_);
  or (_04562_, _04524_, _04041_);
  or (_04563_, _04523_, \oc8051_golden_model_1.IRAM[9] [7]);
  and (_04564_, _04563_, _04527_);
  and (_04565_, _04564_, _04562_);
  and (_04566_, _04526_, _04044_);
  or (_13899_, _04566_, _04565_);
  and (_04567_, _04475_, _04205_);
  not (_04568_, _04567_);
  or (_04569_, _04568_, _04057_);
  and (_04570_, _04480_, _04201_);
  not (_04571_, _04570_);
  or (_04572_, _04567_, \oc8051_golden_model_1.IRAM[10] [0]);
  and (_04573_, _04572_, _04571_);
  and (_04575_, _04573_, _04569_);
  and (_04576_, _04570_, _04157_);
  or (_13900_[0], _04576_, _04575_);
  or (_04577_, _04568_, _04076_);
  or (_04578_, _04567_, \oc8051_golden_model_1.IRAM[10] [1]);
  and (_04579_, _04578_, _04571_);
  and (_04580_, _04579_, _04577_);
  and (_04581_, _04570_, _04163_);
  or (_13900_[1], _04581_, _04580_);
  or (_04582_, _04568_, _04087_);
  or (_04583_, _04567_, \oc8051_golden_model_1.IRAM[10] [2]);
  and (_04584_, _04583_, _04571_);
  and (_04585_, _04584_, _04582_);
  and (_04586_, _04570_, _04169_);
  or (_13900_[2], _04586_, _04585_);
  or (_04587_, _04568_, _04100_);
  or (_04588_, _04567_, \oc8051_golden_model_1.IRAM[10] [3]);
  and (_04589_, _04588_, _04571_);
  and (_04590_, _04589_, _04587_);
  and (_04591_, _04570_, _04175_);
  or (_13900_[3], _04591_, _04590_);
  or (_04592_, _04568_, _04111_);
  or (_04593_, _04567_, \oc8051_golden_model_1.IRAM[10] [4]);
  and (_04594_, _04593_, _04571_);
  and (_04595_, _04594_, _04592_);
  and (_04596_, _04570_, _04181_);
  or (_13900_[4], _04596_, _04595_);
  or (_04597_, _04568_, _04122_);
  or (_04598_, _04567_, \oc8051_golden_model_1.IRAM[10] [5]);
  and (_04599_, _04598_, _04571_);
  and (_04600_, _04599_, _04597_);
  and (_04601_, _04570_, _04187_);
  or (_13900_[5], _04601_, _04600_);
  or (_04602_, _04568_, _04133_);
  or (_04603_, _04567_, \oc8051_golden_model_1.IRAM[10] [6]);
  and (_04604_, _04603_, _04571_);
  and (_04605_, _04604_, _04602_);
  and (_04606_, _04570_, _04193_);
  or (_13900_[6], _04606_, _04605_);
  or (_04607_, _04568_, _04041_);
  or (_04608_, _04567_, \oc8051_golden_model_1.IRAM[10] [7]);
  and (_04609_, _04608_, _04571_);
  and (_04610_, _04609_, _04607_);
  and (_04611_, _04570_, _04044_);
  or (_13900_[7], _04611_, _04610_);
  and (_04612_, _04475_, _04016_);
  or (_04613_, _04612_, \oc8051_golden_model_1.IRAM[11] [0]);
  and (_04614_, _04480_, _04032_);
  not (_04615_, _04614_);
  and (_04616_, _04615_, _04613_);
  not (_04617_, _04612_);
  or (_04618_, _04617_, _04057_);
  and (_04619_, _04618_, _04616_);
  and (_04620_, _04614_, _04157_);
  or (_13901_[0], _04620_, _04619_);
  or (_04621_, _04612_, \oc8051_golden_model_1.IRAM[11] [1]);
  and (_04622_, _04621_, _04615_);
  or (_04623_, _04617_, _04076_);
  and (_04624_, _04623_, _04622_);
  and (_04625_, _04614_, _04163_);
  or (_13901_[1], _04625_, _04624_);
  or (_04626_, _04612_, \oc8051_golden_model_1.IRAM[11] [2]);
  and (_04627_, _04626_, _04615_);
  or (_04628_, _04617_, _04087_);
  and (_04629_, _04628_, _04627_);
  and (_04630_, _04614_, _04169_);
  or (_13901_[2], _04630_, _04629_);
  or (_04631_, _04612_, \oc8051_golden_model_1.IRAM[11] [3]);
  and (_04632_, _04631_, _04615_);
  or (_04633_, _04617_, _04100_);
  and (_04634_, _04633_, _04632_);
  and (_04635_, _04614_, _04175_);
  or (_13901_[3], _04635_, _04634_);
  or (_04636_, _04612_, \oc8051_golden_model_1.IRAM[11] [4]);
  and (_04637_, _04636_, _04615_);
  or (_04638_, _04617_, _04111_);
  and (_04639_, _04638_, _04637_);
  and (_04640_, _04614_, _04181_);
  or (_13901_[4], _04640_, _04639_);
  or (_04641_, _04612_, \oc8051_golden_model_1.IRAM[11] [5]);
  and (_04642_, _04641_, _04615_);
  or (_04643_, _04617_, _04122_);
  and (_04644_, _04643_, _04642_);
  and (_04645_, _04614_, _04187_);
  or (_13901_[5], _04645_, _04644_);
  or (_04646_, _04612_, \oc8051_golden_model_1.IRAM[11] [6]);
  and (_04647_, _04646_, _04615_);
  or (_04648_, _04617_, _04133_);
  and (_04649_, _04648_, _04647_);
  and (_04650_, _04614_, _04193_);
  or (_13901_[6], _04650_, _04649_);
  or (_04651_, _04612_, \oc8051_golden_model_1.IRAM[11] [7]);
  and (_04652_, _04651_, _04615_);
  or (_04653_, _04617_, _04041_);
  and (_04654_, _04653_, _04652_);
  and (_04655_, _04614_, _04044_);
  or (_13901_[7], _04655_, _04654_);
  and (_04656_, _04060_, _04030_);
  not (_04657_, _04656_);
  and (_04658_, _04047_, _04024_);
  or (_04660_, _04658_, \oc8051_golden_model_1.IRAM[12] [0]);
  and (_04661_, _04660_, _04657_);
  not (_04662_, _04658_);
  or (_04663_, _04662_, _04057_);
  and (_04664_, _04663_, _04661_);
  and (_04665_, _04656_, _04157_);
  or (_13902_[0], _04665_, _04664_);
  or (_04666_, _04658_, \oc8051_golden_model_1.IRAM[12] [1]);
  and (_04667_, _04666_, _04657_);
  or (_04668_, _04662_, _04076_);
  and (_04669_, _04668_, _04667_);
  and (_04670_, _04656_, _04163_);
  or (_13902_[1], _04670_, _04669_);
  or (_04671_, _04658_, \oc8051_golden_model_1.IRAM[12] [2]);
  and (_04672_, _04671_, _04657_);
  or (_04673_, _04662_, _04087_);
  and (_04674_, _04673_, _04672_);
  and (_04675_, _04656_, _04169_);
  or (_13902_[2], _04675_, _04674_);
  or (_04676_, _04658_, \oc8051_golden_model_1.IRAM[12] [3]);
  and (_04677_, _04676_, _04657_);
  or (_04678_, _04662_, _04100_);
  and (_04679_, _04678_, _04677_);
  and (_04680_, _04656_, _04175_);
  or (_13902_[3], _04680_, _04679_);
  or (_04681_, _04658_, \oc8051_golden_model_1.IRAM[12] [4]);
  and (_04682_, _04681_, _04657_);
  or (_04683_, _04662_, _04111_);
  and (_04684_, _04683_, _04682_);
  and (_04685_, _04656_, _04181_);
  or (_13902_[4], _04685_, _04684_);
  or (_04686_, _04658_, \oc8051_golden_model_1.IRAM[12] [5]);
  and (_04687_, _04686_, _04657_);
  or (_04688_, _04662_, _04122_);
  and (_04689_, _04688_, _04687_);
  and (_04690_, _04656_, _04187_);
  or (_13902_[5], _04690_, _04689_);
  or (_04691_, _04658_, \oc8051_golden_model_1.IRAM[12] [6]);
  and (_04692_, _04691_, _04657_);
  or (_04693_, _04662_, _04133_);
  and (_04694_, _04693_, _04692_);
  and (_04695_, _04656_, _04193_);
  or (_13902_[6], _04695_, _04694_);
  or (_04696_, _04658_, \oc8051_golden_model_1.IRAM[12] [7]);
  and (_04697_, _04696_, _04657_);
  or (_04698_, _04662_, _04041_);
  and (_04699_, _04698_, _04697_);
  and (_04700_, _04656_, _04044_);
  or (_13902_[7], _04700_, _04699_);
  and (_04701_, _04151_, _04030_);
  not (_04702_, _04701_);
  and (_04703_, _04146_, _04024_);
  or (_04704_, _04703_, \oc8051_golden_model_1.IRAM[13] [0]);
  and (_04705_, _04704_, _04702_);
  not (_04706_, _04703_);
  or (_04707_, _04706_, _04057_);
  and (_04708_, _04707_, _04705_);
  and (_04709_, _04701_, _04157_);
  or (_13903_[0], _04709_, _04708_);
  or (_04710_, _04703_, \oc8051_golden_model_1.IRAM[13] [1]);
  and (_04711_, _04710_, _04702_);
  or (_04712_, _04706_, _04076_);
  and (_04713_, _04712_, _04711_);
  and (_04714_, _04701_, _04163_);
  or (_13903_[1], _04714_, _04713_);
  or (_04715_, _04703_, \oc8051_golden_model_1.IRAM[13] [2]);
  and (_04716_, _04715_, _04702_);
  or (_04717_, _04706_, _04087_);
  and (_04718_, _04717_, _04716_);
  and (_04719_, _04701_, _04169_);
  or (_13903_[2], _04719_, _04718_);
  or (_04720_, _04703_, \oc8051_golden_model_1.IRAM[13] [3]);
  and (_04721_, _04720_, _04702_);
  or (_04722_, _04706_, _04100_);
  and (_04723_, _04722_, _04721_);
  and (_04724_, _04701_, _04175_);
  or (_13903_[3], _04724_, _04723_);
  or (_04725_, _04703_, \oc8051_golden_model_1.IRAM[13] [4]);
  and (_04726_, _04725_, _04702_);
  or (_04727_, _04706_, _04111_);
  and (_04728_, _04727_, _04726_);
  and (_04729_, _04701_, _04181_);
  or (_13903_[4], _04729_, _04728_);
  or (_04730_, _04703_, \oc8051_golden_model_1.IRAM[13] [5]);
  and (_04731_, _04730_, _04702_);
  or (_04732_, _04706_, _04122_);
  and (_04733_, _04732_, _04731_);
  and (_04734_, _04701_, _04187_);
  or (_13903_[5], _04734_, _04733_);
  or (_04735_, _04703_, \oc8051_golden_model_1.IRAM[13] [6]);
  and (_04736_, _04735_, _04702_);
  or (_04737_, _04706_, _04133_);
  and (_04738_, _04737_, _04736_);
  and (_04739_, _04701_, _04193_);
  or (_13903_[6], _04739_, _04738_);
  or (_04740_, _04703_, \oc8051_golden_model_1.IRAM[13] [7]);
  and (_04741_, _04740_, _04702_);
  or (_04742_, _04706_, _04041_);
  and (_04743_, _04742_, _04741_);
  and (_04744_, _04701_, _04044_);
  or (_13903_[7], _04744_, _04743_);
  and (_04746_, _04201_, _04030_);
  and (_04747_, _04746_, _04157_);
  not (_04748_, _04746_);
  and (_04749_, _04205_, _04024_);
  or (_04750_, _04749_, \oc8051_golden_model_1.IRAM[14] [0]);
  and (_04751_, _04750_, _04748_);
  not (_04752_, _04749_);
  or (_04753_, _04752_, _04057_);
  and (_04754_, _04753_, _04751_);
  or (_13904_[0], _04754_, _04747_);
  or (_04755_, _04749_, \oc8051_golden_model_1.IRAM[14] [1]);
  and (_04756_, _04755_, _04748_);
  or (_04757_, _04752_, _04076_);
  and (_04758_, _04757_, _04756_);
  and (_04759_, _04746_, _04163_);
  or (_13904_[1], _04759_, _04758_);
  and (_04760_, _04746_, _04169_);
  or (_04761_, _04749_, \oc8051_golden_model_1.IRAM[14] [2]);
  and (_04762_, _04761_, _04748_);
  or (_04763_, _04752_, _04087_);
  and (_04764_, _04763_, _04762_);
  or (_13904_[2], _04764_, _04760_);
  and (_04765_, _04746_, _04175_);
  or (_04766_, _04749_, \oc8051_golden_model_1.IRAM[14] [3]);
  and (_04767_, _04766_, _04748_);
  or (_04768_, _04752_, _04100_);
  and (_04769_, _04768_, _04767_);
  or (_13904_[3], _04769_, _04765_);
  and (_04770_, _04746_, _04181_);
  or (_04771_, _04749_, \oc8051_golden_model_1.IRAM[14] [4]);
  and (_04772_, _04771_, _04748_);
  or (_04773_, _04752_, _04111_);
  and (_04774_, _04773_, _04772_);
  or (_13904_[4], _04774_, _04770_);
  or (_04775_, _04749_, \oc8051_golden_model_1.IRAM[14] [5]);
  and (_04776_, _04775_, _04748_);
  or (_04777_, _04752_, _04122_);
  and (_04778_, _04777_, _04776_);
  and (_04779_, _04746_, _04187_);
  or (_13904_[5], _04779_, _04778_);
  and (_04780_, _04746_, _04193_);
  or (_04781_, _04749_, \oc8051_golden_model_1.IRAM[14] [6]);
  and (_04782_, _04781_, _04748_);
  or (_04783_, _04752_, _04133_);
  and (_04784_, _04783_, _04782_);
  or (_13904_[6], _04784_, _04780_);
  and (_04785_, _04746_, _04044_);
  or (_04786_, _04749_, \oc8051_golden_model_1.IRAM[14] [7]);
  and (_04787_, _04786_, _04748_);
  or (_04788_, _04752_, _04041_);
  and (_04789_, _04788_, _04787_);
  or (_13904_[7], _04789_, _04785_);
  or (_04790_, _04025_, \oc8051_golden_model_1.IRAM[15] [0]);
  and (_04791_, _04790_, _04034_);
  or (_04792_, _04057_, _04036_);
  and (_04793_, _04792_, _04791_);
  and (_04794_, _04157_, _04033_);
  or (_13905_[0], _04794_, _04793_);
  or (_04795_, _04025_, \oc8051_golden_model_1.IRAM[15] [1]);
  and (_04796_, _04795_, _04034_);
  or (_04797_, _04076_, _04036_);
  and (_04798_, _04797_, _04796_);
  and (_04799_, _04163_, _04033_);
  or (_13905_[1], _04799_, _04798_);
  or (_04800_, _04025_, \oc8051_golden_model_1.IRAM[15] [2]);
  and (_04801_, _04800_, _04034_);
  or (_04802_, _04087_, _04036_);
  and (_04803_, _04802_, _04801_);
  and (_04804_, _04169_, _04033_);
  or (_13905_[2], _04804_, _04803_);
  or (_04805_, _04025_, \oc8051_golden_model_1.IRAM[15] [3]);
  and (_04806_, _04805_, _04034_);
  or (_04807_, _04100_, _04036_);
  and (_04808_, _04807_, _04806_);
  and (_04809_, _04175_, _04033_);
  or (_13905_[3], _04809_, _04808_);
  or (_04810_, _04025_, \oc8051_golden_model_1.IRAM[15] [4]);
  and (_04811_, _04810_, _04034_);
  or (_04812_, _04111_, _04036_);
  and (_04813_, _04812_, _04811_);
  and (_04814_, _04181_, _04033_);
  or (_13905_[4], _04814_, _04813_);
  or (_04815_, _04025_, \oc8051_golden_model_1.IRAM[15] [5]);
  and (_04816_, _04815_, _04034_);
  or (_04817_, _04122_, _04036_);
  and (_04818_, _04817_, _04816_);
  and (_04819_, _04187_, _04033_);
  or (_13905_[5], _04819_, _04818_);
  or (_04820_, _04025_, \oc8051_golden_model_1.IRAM[15] [6]);
  and (_04821_, _04820_, _04034_);
  or (_04822_, _04133_, _04036_);
  and (_04823_, _04822_, _04821_);
  and (_04824_, _04193_, _04033_);
  or (_13905_[6], _04824_, _04823_);
  or (_04825_, _12782_, \oc8051_golden_model_1.B [0]);
  and (_04826_, _04825_, _13707_);
  and (_04827_, _02715_, B_abstr[0]);
  or (_04828_, _04827_, _12786_);
  or (_04829_, _03192_, \oc8051_golden_model_1.B [0]);
  and (_04831_, _03680_, _02758_);
  and (_04832_, _04831_, _04829_);
  or (_04833_, _04832_, _04828_);
  and (_13829_[0], _04833_, _04826_);
  nand (_04834_, _04072_, _03192_);
  or (_04835_, _03192_, \oc8051_golden_model_1.B [1]);
  and (_04836_, _04835_, _02758_);
  and (_04837_, _04836_, _04834_);
  and (_04838_, _02715_, B_abstr[1]);
  or (_04839_, _04838_, _12786_);
  or (_04840_, _04839_, _04837_);
  or (_04841_, _12782_, \oc8051_golden_model_1.B [1]);
  and (_04842_, _04841_, _13707_);
  and (_13829_[1], _04842_, _04840_);
  or (_04843_, _12782_, \oc8051_golden_model_1.B [2]);
  and (_04844_, _04843_, _13707_);
  and (_04845_, _02715_, B_abstr[2]);
  or (_04846_, _04845_, _12786_);
  or (_04847_, _04083_, _03996_);
  or (_04848_, _03192_, \oc8051_golden_model_1.B [2]);
  and (_04849_, _04848_, _02758_);
  and (_04850_, _04849_, _04847_);
  or (_04851_, _04850_, _04846_);
  and (_13829_[2], _04851_, _04844_);
  nand (_04852_, _04096_, _03192_);
  or (_04853_, _03192_, \oc8051_golden_model_1.B [3]);
  and (_04854_, _04853_, _02758_);
  and (_04855_, _04854_, _04852_);
  and (_04856_, _02715_, B_abstr[3]);
  or (_04857_, _04856_, _12786_);
  or (_04858_, _04857_, _04855_);
  or (_04859_, _12782_, \oc8051_golden_model_1.B [3]);
  and (_04860_, _04859_, _13707_);
  and (_13829_[3], _04860_, _04858_);
  or (_04861_, _12782_, \oc8051_golden_model_1.B [4]);
  and (_04862_, _04861_, _13707_);
  nand (_04863_, _04107_, _03192_);
  or (_04864_, _03192_, \oc8051_golden_model_1.B [4]);
  and (_04865_, _04864_, _02758_);
  and (_04866_, _04865_, _04863_);
  and (_04867_, _02715_, B_abstr[4]);
  or (_04868_, _04867_, _12786_);
  or (_04869_, _04868_, _04866_);
  and (_13829_[4], _04869_, _04862_);
  or (_04870_, _04118_, _03996_);
  or (_04871_, _03192_, \oc8051_golden_model_1.B [5]);
  and (_04872_, _04871_, _02758_);
  and (_04873_, _04872_, _04870_);
  and (_04874_, _02715_, B_abstr[5]);
  or (_04875_, _04874_, _12786_);
  or (_04876_, _04875_, _04873_);
  or (_04877_, _12782_, \oc8051_golden_model_1.B [5]);
  and (_04878_, _04877_, _13707_);
  and (_13829_[5], _04878_, _04876_);
  or (_04879_, _12782_, \oc8051_golden_model_1.B [6]);
  and (_04880_, _04879_, _13707_);
  and (_04881_, _02715_, B_abstr[6]);
  or (_04882_, _04881_, _12786_);
  or (_04883_, _04129_, _03996_);
  or (_04884_, _03192_, \oc8051_golden_model_1.B [6]);
  and (_04885_, _04884_, _02758_);
  and (_04886_, _04885_, _04883_);
  or (_04887_, _04886_, _04882_);
  and (_13829_[6], _04887_, _04880_);
  nor (_04888_, _12782_, _03691_);
  and (_04889_, _03164_, _03691_);
  not (_04890_, _04889_);
  and (_04891_, _04890_, _03692_);
  or (_04892_, _04891_, _02715_);
  or (_04893_, _02758_, ACC_abstr[0]);
  and (_04894_, _04893_, _12782_);
  and (_04895_, _04894_, _04892_);
  or (_04896_, _04895_, _04888_);
  and (_13828_[0], _04896_, _13707_);
  nor (_04897_, _12782_, _03595_);
  and (_04898_, _03164_, \oc8051_golden_model_1.ACC [1]);
  not (_04899_, _04898_);
  or (_04900_, _04072_, _03164_);
  nand (_04901_, _04900_, _04899_);
  or (_04902_, _04901_, _02715_);
  or (_04903_, _02758_, ACC_abstr[1]);
  and (_04904_, _04903_, _12782_);
  and (_04905_, _04904_, _04902_);
  or (_04906_, _04905_, _04897_);
  and (_13828_[1], _04906_, _13707_);
  nor (_04907_, _12782_, _03758_);
  and (_04908_, _03164_, \oc8051_golden_model_1.ACC [2]);
  not (_04909_, _04908_);
  nand (_04910_, _04083_, _03986_);
  and (_04911_, _04910_, _04909_);
  nand (_04912_, _04911_, _02758_);
  or (_04913_, _02758_, ACC_abstr[2]);
  and (_04914_, _04913_, _12782_);
  and (_04915_, _04914_, _04912_);
  or (_04916_, _04915_, _04907_);
  and (_13828_[2], _04916_, _13707_);
  nor (_04917_, _12782_, _03491_);
  and (_04918_, _03164_, \oc8051_golden_model_1.ACC [3]);
  not (_04919_, _04918_);
  or (_04920_, _04096_, _03164_);
  nand (_04922_, _04920_, _04919_);
  or (_04923_, _04922_, _02715_);
  or (_04924_, _02758_, ACC_abstr[3]);
  and (_04925_, _04924_, _12782_);
  and (_04926_, _04925_, _04923_);
  or (_04927_, _04926_, _04917_);
  and (_13828_[3], _04927_, _13707_);
  nor (_04928_, _12782_, _03871_);
  and (_04929_, _03164_, \oc8051_golden_model_1.ACC [4]);
  not (_04930_, _04929_);
  or (_04931_, _04107_, _03164_);
  nand (_04932_, _04931_, _04930_);
  or (_04933_, _04932_, _02715_);
  or (_04934_, _02758_, ACC_abstr[4]);
  and (_04935_, _04934_, _12782_);
  and (_04936_, _04935_, _04933_);
  or (_04937_, _04936_, _04928_);
  and (_13828_[4], _04937_, _13707_);
  nor (_04938_, _12782_, _03410_);
  and (_04939_, _03164_, \oc8051_golden_model_1.ACC [5]);
  and (_04940_, _04118_, _03986_);
  nor (_04941_, _04940_, _04939_);
  nand (_04942_, _04941_, _02758_);
  or (_04943_, _02758_, ACC_abstr[5]);
  and (_04944_, _04943_, _12782_);
  and (_04945_, _04944_, _04942_);
  or (_04946_, _04945_, _04938_);
  and (_13828_[5], _04946_, _13707_);
  nor (_04947_, _12782_, _03315_);
  and (_04948_, _03164_, \oc8051_golden_model_1.ACC [6]);
  not (_04949_, _04948_);
  nand (_04950_, _04129_, _03986_);
  and (_04951_, _04950_, _04949_);
  nand (_04952_, _04951_, _02758_);
  or (_04953_, _02758_, ACC_abstr[6]);
  and (_04954_, _04953_, _12782_);
  and (_04955_, _04954_, _04952_);
  or (_04956_, _04955_, _04947_);
  and (_13828_[6], _04956_, _13707_);
  or (_04957_, _12782_, \oc8051_golden_model_1.DPL [0]);
  and (_04958_, _04957_, _13707_);
  and (_04959_, _02715_, DPL_abstr[0]);
  or (_04960_, _04959_, _12786_);
  or (_04961_, _03178_, \oc8051_golden_model_1.DPL [0]);
  and (_04962_, _03669_, _02758_);
  and (_04963_, _04962_, _04961_);
  or (_04964_, _04963_, _04960_);
  and (_13831_[0], _04964_, _04958_);
  nand (_04965_, _04072_, _03178_);
  or (_04966_, _03178_, \oc8051_golden_model_1.DPL [1]);
  and (_04967_, _04966_, _02758_);
  and (_04968_, _04967_, _04965_);
  and (_04969_, _02715_, DPL_abstr[1]);
  or (_04970_, _04969_, _12786_);
  or (_04971_, _04970_, _04968_);
  or (_04972_, _12782_, \oc8051_golden_model_1.DPL [1]);
  and (_04973_, _04972_, _13707_);
  and (_13831_[1], _04973_, _04971_);
  or (_04974_, _12782_, \oc8051_golden_model_1.DPL [2]);
  and (_04975_, _04974_, _13707_);
  and (_04976_, _02715_, DPL_abstr[2]);
  or (_04977_, _04976_, _12786_);
  or (_04978_, _04083_, _03975_);
  or (_04979_, _03178_, \oc8051_golden_model_1.DPL [2]);
  and (_04980_, _04979_, _02758_);
  and (_04981_, _04980_, _04978_);
  or (_04982_, _04981_, _04977_);
  and (_13831_[2], _04982_, _04975_);
  or (_04983_, _12782_, \oc8051_golden_model_1.DPL [3]);
  and (_04984_, _04983_, _13707_);
  and (_04985_, _02715_, DPL_abstr[3]);
  or (_04986_, _04985_, _12786_);
  nand (_04987_, _04096_, _03178_);
  or (_04988_, _03178_, \oc8051_golden_model_1.DPL [3]);
  and (_04989_, _04988_, _02758_);
  and (_04990_, _04989_, _04987_);
  or (_04991_, _04990_, _04986_);
  and (_13831_[3], _04991_, _04984_);
  or (_04992_, _12782_, \oc8051_golden_model_1.DPL [4]);
  and (_04993_, _04992_, _13707_);
  and (_04994_, _02715_, DPL_abstr[4]);
  or (_04995_, _04994_, _12786_);
  nand (_04996_, _04107_, _03178_);
  or (_04997_, _03178_, \oc8051_golden_model_1.DPL [4]);
  and (_04998_, _04997_, _02758_);
  and (_04999_, _04998_, _04996_);
  or (_05000_, _04999_, _04995_);
  and (_13831_[4], _05000_, _04993_);
  or (_05001_, _04118_, _03975_);
  or (_05002_, _03178_, \oc8051_golden_model_1.DPL [5]);
  and (_05003_, _05002_, _02758_);
  and (_05004_, _05003_, _05001_);
  and (_05005_, _02715_, DPL_abstr[5]);
  or (_05006_, _05005_, _12786_);
  or (_05007_, _05006_, _05004_);
  or (_05008_, _12782_, \oc8051_golden_model_1.DPL [5]);
  and (_05009_, _05008_, _13707_);
  and (_13831_[5], _05009_, _05007_);
  or (_05010_, _12782_, \oc8051_golden_model_1.DPL [6]);
  and (_05011_, _05010_, _13707_);
  and (_05012_, _02715_, DPL_abstr[6]);
  or (_05013_, _05012_, _12786_);
  or (_05014_, _04129_, _03975_);
  or (_05015_, _03178_, \oc8051_golden_model_1.DPL [6]);
  and (_05016_, _05015_, _02758_);
  and (_05017_, _05016_, _05014_);
  or (_05018_, _05017_, _05013_);
  and (_13831_[6], _05018_, _05011_);
  or (_05019_, _12782_, \oc8051_golden_model_1.DPH [0]);
  and (_05020_, _05019_, _13707_);
  and (_05021_, _03967_, \oc8051_golden_model_1.DPH [0]);
  and (_05022_, _04053_, _03229_);
  or (_05023_, _05022_, _05021_);
  and (_05024_, _05023_, _02758_);
  and (_05025_, _02715_, DPH_abstr[0]);
  or (_05026_, _05025_, _12786_);
  or (_05027_, _05026_, _05024_);
  and (_13830_[0], _05027_, _05020_);
  or (_05028_, _12782_, \oc8051_golden_model_1.DPH [1]);
  and (_05029_, _05028_, _13707_);
  and (_05030_, _03967_, \oc8051_golden_model_1.DPH [1]);
  nor (_05031_, _04072_, _03967_);
  or (_05032_, _05031_, _05030_);
  and (_05033_, _05032_, _02758_);
  and (_05034_, _02715_, DPH_abstr[1]);
  or (_05035_, _05034_, _12786_);
  or (_05036_, _05035_, _05033_);
  and (_13830_[1], _05036_, _05029_);
  or (_05037_, _04083_, _03967_);
  or (_05038_, _03229_, \oc8051_golden_model_1.DPH [2]);
  and (_05039_, _05038_, _02758_);
  and (_05040_, _05039_, _05037_);
  and (_05041_, _02715_, DPH_abstr[2]);
  or (_05042_, _05041_, _12786_);
  or (_05043_, _05042_, _05040_);
  or (_05044_, _12782_, \oc8051_golden_model_1.DPH [2]);
  and (_05045_, _05044_, _13707_);
  and (_13830_[2], _05045_, _05043_);
  or (_05046_, _12782_, \oc8051_golden_model_1.DPH [3]);
  and (_05047_, _05046_, _13707_);
  and (_05048_, _02715_, DPH_abstr[3]);
  or (_05049_, _05048_, _12786_);
  nand (_05050_, _04096_, _03229_);
  or (_05051_, _03229_, \oc8051_golden_model_1.DPH [3]);
  and (_05052_, _05051_, _02758_);
  and (_05053_, _05052_, _05050_);
  or (_05054_, _05053_, _05049_);
  and (_13830_[3], _05054_, _05047_);
  or (_05055_, _12782_, \oc8051_golden_model_1.DPH [4]);
  and (_05056_, _05055_, _13707_);
  and (_05057_, _02715_, DPH_abstr[4]);
  or (_05058_, _05057_, _12786_);
  nand (_05059_, _04107_, _03229_);
  or (_05060_, _03229_, \oc8051_golden_model_1.DPH [4]);
  and (_05061_, _05060_, _02758_);
  and (_05062_, _05061_, _05059_);
  or (_05063_, _05062_, _05058_);
  and (_13830_[4], _05063_, _05056_);
  or (_05064_, _12782_, \oc8051_golden_model_1.DPH [5]);
  and (_05065_, _05064_, _13707_);
  and (_05066_, _02715_, DPH_abstr[5]);
  or (_05067_, _05066_, _12786_);
  or (_05068_, _04118_, _03967_);
  or (_05069_, _03229_, \oc8051_golden_model_1.DPH [5]);
  and (_05070_, _05069_, _02758_);
  and (_05071_, _05070_, _05068_);
  or (_05072_, _05071_, _05067_);
  and (_13830_[5], _05072_, _05065_);
  or (_05073_, _04129_, _03967_);
  or (_05074_, _03229_, \oc8051_golden_model_1.DPH [6]);
  and (_05075_, _05074_, _02758_);
  and (_05076_, _05075_, _05073_);
  and (_05077_, _02715_, DPH_abstr[6]);
  or (_05078_, _05077_, _12786_);
  or (_05079_, _05078_, _05076_);
  or (_05080_, _12782_, \oc8051_golden_model_1.DPH [6]);
  and (_05081_, _05080_, _13707_);
  and (_13830_[6], _05081_, _05079_);
  and (_13832_[0], \oc8051_golden_model_1.IE [0], _13707_);
  and (_13832_[1], \oc8051_golden_model_1.IE [1], _13707_);
  and (_13832_[2], \oc8051_golden_model_1.IE [2], _13707_);
  and (_13832_[3], \oc8051_golden_model_1.IE [3], _13707_);
  and (_13832_[4], \oc8051_golden_model_1.IE [4], _13707_);
  and (_13832_[5], \oc8051_golden_model_1.IE [5], _13707_);
  and (_13832_[6], \oc8051_golden_model_1.IE [6], _13707_);
  and (_13833_[0], \oc8051_golden_model_1.IP [0], _13707_);
  and (_13833_[1], \oc8051_golden_model_1.IP [1], _13707_);
  and (_13833_[2], \oc8051_golden_model_1.IP [2], _13707_);
  and (_13833_[3], \oc8051_golden_model_1.IP [3], _13707_);
  and (_13833_[4], \oc8051_golden_model_1.IP [4], _13707_);
  and (_13833_[5], \oc8051_golden_model_1.IP [5], _13707_);
  and (_13833_[6], \oc8051_golden_model_1.IP [6], _13707_);
  and (_05082_, _02715_, P0_abstr[0]);
  or (_05083_, _03217_, \oc8051_golden_model_1.P0 [0]);
  and (_05084_, _05083_, _02758_);
  and (_05085_, _05084_, _03664_);
  or (_05086_, _05085_, _05082_);
  and (_05087_, _05086_, _12782_);
  nor (_05088_, \oc8051_golden_model_1.P0 [0], rst);
  nor (_05089_, _05088_, _00002_);
  or (_13834_[0], _05089_, _05087_);
  and (_05090_, _02715_, P0_abstr[1]);
  nand (_05091_, _04072_, _03217_);
  or (_05092_, _03217_, \oc8051_golden_model_1.P0 [1]);
  and (_05093_, _05092_, _02758_);
  and (_05094_, _05093_, _05091_);
  or (_05095_, _05094_, _05090_);
  and (_05096_, _05095_, _12782_);
  nor (_05097_, \oc8051_golden_model_1.P0 [1], rst);
  nor (_05098_, _05097_, _00002_);
  or (_13834_[1], _05098_, _05096_);
  and (_05099_, _02715_, P0_abstr[2]);
  or (_05100_, _04083_, _03952_);
  or (_05101_, _03217_, \oc8051_golden_model_1.P0 [2]);
  and (_05102_, _05101_, _02758_);
  and (_05103_, _05102_, _05100_);
  or (_05104_, _05103_, _05099_);
  and (_05105_, _05104_, _12782_);
  nor (_05106_, \oc8051_golden_model_1.P0 [2], rst);
  nor (_05107_, _05106_, _00002_);
  or (_13834_[2], _05107_, _05105_);
  and (_05108_, _02715_, P0_abstr[3]);
  nand (_05109_, _04096_, _03217_);
  or (_05110_, _03217_, \oc8051_golden_model_1.P0 [3]);
  and (_05111_, _05110_, _02758_);
  and (_05112_, _05111_, _05109_);
  or (_05113_, _05112_, _05108_);
  and (_05114_, _05113_, _12782_);
  nor (_05115_, \oc8051_golden_model_1.P0 [3], rst);
  nor (_05116_, _05115_, _00002_);
  or (_13834_[3], _05116_, _05114_);
  and (_05117_, _02715_, P0_abstr[4]);
  nand (_05118_, _04107_, _03217_);
  or (_05119_, _03217_, \oc8051_golden_model_1.P0 [4]);
  and (_05120_, _05119_, _02758_);
  and (_05121_, _05120_, _05118_);
  or (_05122_, _05121_, _05117_);
  and (_05123_, _05122_, _12782_);
  nor (_05124_, \oc8051_golden_model_1.P0 [4], rst);
  nor (_05125_, _05124_, _00002_);
  or (_13834_[4], _05125_, _05123_);
  and (_05126_, _02715_, P0_abstr[5]);
  or (_05127_, _04118_, _03952_);
  or (_05128_, _03217_, \oc8051_golden_model_1.P0 [5]);
  and (_05129_, _05128_, _02758_);
  and (_05130_, _05129_, _05127_);
  or (_05131_, _05130_, _05126_);
  and (_05132_, _05131_, _12782_);
  nor (_05133_, \oc8051_golden_model_1.P0 [5], rst);
  nor (_05134_, _05133_, _00002_);
  or (_13834_[5], _05134_, _05132_);
  and (_05135_, _02715_, P0_abstr[6]);
  or (_05136_, _04129_, _03952_);
  or (_05137_, _03217_, \oc8051_golden_model_1.P0 [6]);
  and (_05138_, _05137_, _02758_);
  and (_05139_, _05138_, _05136_);
  or (_05140_, _05139_, _05135_);
  and (_05141_, _05140_, _12782_);
  nor (_05142_, \oc8051_golden_model_1.P0 [6], rst);
  nor (_05143_, _05142_, _00002_);
  or (_13834_[6], _05143_, _05141_);
  and (_05144_, _02715_, P1_abstr[0]);
  or (_05145_, _03198_, \oc8051_golden_model_1.P1 [0]);
  and (_05146_, _05145_, _02758_);
  and (_05147_, _05146_, _03678_);
  or (_05148_, _05147_, _05144_);
  and (_05149_, _05148_, _12782_);
  nor (_05150_, \oc8051_golden_model_1.P1 [0], rst);
  nor (_05151_, _05150_, _00002_);
  or (_13835_[0], _05151_, _05149_);
  and (_05152_, _02715_, P1_abstr[1]);
  nand (_05153_, _04072_, _03198_);
  or (_05154_, _03198_, \oc8051_golden_model_1.P1 [1]);
  and (_05155_, _05154_, _02758_);
  and (_05156_, _05155_, _05153_);
  or (_05157_, _05156_, _05152_);
  and (_05158_, _05157_, _12782_);
  nor (_05159_, \oc8051_golden_model_1.P1 [1], rst);
  nor (_05160_, _05159_, _00002_);
  or (_13835_[1], _05160_, _05158_);
  and (_05161_, _02715_, P1_abstr[2]);
  or (_05162_, _04083_, _03941_);
  or (_05163_, _03198_, \oc8051_golden_model_1.P1 [2]);
  and (_05164_, _05163_, _02758_);
  and (_05165_, _05164_, _05162_);
  or (_05166_, _05165_, _05161_);
  and (_05167_, _05166_, _12782_);
  nor (_05168_, \oc8051_golden_model_1.P1 [2], rst);
  nor (_05169_, _05168_, _00002_);
  or (_13835_[2], _05169_, _05167_);
  and (_05170_, _02715_, P1_abstr[3]);
  nand (_05171_, _04096_, _03198_);
  or (_05172_, _03198_, \oc8051_golden_model_1.P1 [3]);
  and (_05173_, _05172_, _02758_);
  and (_05174_, _05173_, _05171_);
  or (_05175_, _05174_, _05170_);
  and (_05176_, _05175_, _12782_);
  nor (_05177_, \oc8051_golden_model_1.P1 [3], rst);
  nor (_05178_, _05177_, _00002_);
  or (_13835_[3], _05178_, _05176_);
  and (_05179_, _02715_, P1_abstr[4]);
  nand (_05180_, _04107_, _03198_);
  or (_05181_, _03198_, \oc8051_golden_model_1.P1 [4]);
  and (_05182_, _05181_, _02758_);
  and (_05183_, _05182_, _05180_);
  or (_05184_, _05183_, _05179_);
  and (_05185_, _05184_, _12782_);
  nor (_05186_, \oc8051_golden_model_1.P1 [4], rst);
  nor (_05187_, _05186_, _00002_);
  or (_13835_[4], _05187_, _05185_);
  and (_05188_, _02715_, P1_abstr[5]);
  or (_05189_, _04118_, _03941_);
  or (_05190_, _03198_, \oc8051_golden_model_1.P1 [5]);
  and (_05191_, _05190_, _02758_);
  and (_05192_, _05191_, _05189_);
  or (_05193_, _05192_, _05188_);
  and (_05194_, _05193_, _12782_);
  nor (_05195_, \oc8051_golden_model_1.P1 [5], rst);
  nor (_05196_, _05195_, _00002_);
  or (_13835_[5], _05196_, _05194_);
  and (_05197_, _02715_, P1_abstr[6]);
  or (_05198_, _04129_, _03941_);
  or (_05199_, _03198_, \oc8051_golden_model_1.P1 [6]);
  and (_05200_, _05199_, _02758_);
  and (_05201_, _05200_, _05198_);
  or (_05202_, _05201_, _05197_);
  and (_05203_, _05202_, _12782_);
  nor (_05204_, \oc8051_golden_model_1.P1 [6], rst);
  nor (_05205_, _05204_, _00002_);
  or (_13835_[6], _05205_, _05203_);
  and (_05206_, _02715_, P2_abstr[0]);
  or (_05207_, _03208_, \oc8051_golden_model_1.P2 [0]);
  and (_05208_, _05207_, _02758_);
  and (_05209_, _05208_, _03685_);
  or (_05210_, _05209_, _05206_);
  and (_05211_, _05210_, _12782_);
  nor (_05212_, \oc8051_golden_model_1.P2 [0], rst);
  nor (_05213_, _05212_, _00002_);
  or (_13836_[0], _05213_, _05211_);
  and (_05214_, _02715_, P2_abstr[1]);
  nand (_05215_, _04072_, _03208_);
  or (_05216_, _03208_, \oc8051_golden_model_1.P2 [1]);
  and (_05217_, _05216_, _02758_);
  and (_05218_, _05217_, _05215_);
  or (_05219_, _05218_, _05214_);
  and (_05220_, _05219_, _12782_);
  nor (_05221_, \oc8051_golden_model_1.P2 [1], rst);
  nor (_05222_, _05221_, _00002_);
  or (_13836_[1], _05222_, _05220_);
  and (_05223_, _02715_, P2_abstr[2]);
  or (_05224_, _04083_, _03930_);
  or (_05225_, _03208_, \oc8051_golden_model_1.P2 [2]);
  and (_05226_, _05225_, _02758_);
  and (_05227_, _05226_, _05224_);
  or (_05228_, _05227_, _05223_);
  and (_05229_, _05228_, _12782_);
  nor (_05230_, \oc8051_golden_model_1.P2 [2], rst);
  nor (_05231_, _05230_, _00002_);
  or (_13836_[2], _05231_, _05229_);
  and (_05232_, _02715_, P2_abstr[3]);
  nand (_05233_, _04096_, _03208_);
  or (_05234_, _03208_, \oc8051_golden_model_1.P2 [3]);
  and (_05235_, _05234_, _02758_);
  and (_05236_, _05235_, _05233_);
  or (_05237_, _05236_, _05232_);
  and (_05238_, _05237_, _12782_);
  nor (_05239_, \oc8051_golden_model_1.P2 [3], rst);
  nor (_05240_, _05239_, _00002_);
  or (_13836_[3], _05240_, _05238_);
  and (_05241_, _02715_, P2_abstr[4]);
  nand (_05242_, _04107_, _03208_);
  or (_05243_, _03208_, \oc8051_golden_model_1.P2 [4]);
  and (_05244_, _05243_, _02758_);
  and (_05245_, _05244_, _05242_);
  or (_05246_, _05245_, _05241_);
  and (_05247_, _05246_, _12782_);
  nor (_05248_, \oc8051_golden_model_1.P2 [4], rst);
  nor (_05249_, _05248_, _00002_);
  or (_13836_[4], _05249_, _05247_);
  and (_05250_, _02715_, P2_abstr[5]);
  or (_05251_, _04118_, _03930_);
  or (_05252_, _03208_, \oc8051_golden_model_1.P2 [5]);
  and (_05253_, _05252_, _02758_);
  and (_05254_, _05253_, _05251_);
  or (_05255_, _05254_, _05250_);
  and (_05256_, _05255_, _12782_);
  nor (_05257_, \oc8051_golden_model_1.P2 [5], rst);
  nor (_05258_, _05257_, _00002_);
  or (_13836_[5], _05258_, _05256_);
  and (_05259_, _02715_, P2_abstr[6]);
  or (_05260_, _04129_, _03930_);
  or (_05261_, _03208_, \oc8051_golden_model_1.P2 [6]);
  and (_05262_, _05261_, _02758_);
  and (_05263_, _05262_, _05260_);
  or (_05264_, _05263_, _05259_);
  and (_05265_, _05264_, _12782_);
  nor (_05266_, \oc8051_golden_model_1.P2 [6], rst);
  nor (_05267_, _05266_, _00002_);
  or (_13836_[6], _05267_, _05265_);
  and (_05268_, _02715_, P3_abstr[0]);
  or (_05269_, _03213_, \oc8051_golden_model_1.P3 [0]);
  and (_05270_, _05269_, _02758_);
  and (_05271_, _05270_, _03688_);
  or (_05272_, _05271_, _05268_);
  and (_05273_, _05272_, _12782_);
  nor (_05274_, \oc8051_golden_model_1.P3 [0], rst);
  nor (_05275_, _05274_, _00002_);
  or (_13837_[0], _05275_, _05273_);
  and (_05276_, _02715_, P3_abstr[1]);
  nand (_05277_, _04072_, _03213_);
  or (_05278_, _03213_, \oc8051_golden_model_1.P3 [1]);
  and (_05279_, _05278_, _02758_);
  and (_05280_, _05279_, _05277_);
  or (_05281_, _05280_, _05276_);
  and (_05282_, _05281_, _12782_);
  nor (_05283_, \oc8051_golden_model_1.P3 [1], rst);
  nor (_05284_, _05283_, _00002_);
  or (_13837_[1], _05284_, _05282_);
  and (_05285_, _02715_, P3_abstr[2]);
  or (_05286_, _04083_, _03786_);
  or (_05287_, _03213_, \oc8051_golden_model_1.P3 [2]);
  and (_05288_, _05287_, _02758_);
  and (_05289_, _05288_, _05286_);
  or (_05290_, _05289_, _05285_);
  and (_05291_, _05290_, _12782_);
  nor (_05292_, \oc8051_golden_model_1.P3 [2], rst);
  nor (_05293_, _05292_, _00002_);
  or (_13837_[2], _05293_, _05291_);
  and (_05294_, _02715_, P3_abstr[3]);
  nand (_05295_, _04096_, _03213_);
  or (_05296_, _03213_, \oc8051_golden_model_1.P3 [3]);
  and (_05297_, _05296_, _02758_);
  and (_05298_, _05297_, _05295_);
  or (_05299_, _05298_, _05294_);
  and (_05300_, _05299_, _12782_);
  nor (_05301_, \oc8051_golden_model_1.P3 [3], rst);
  nor (_05302_, _05301_, _00002_);
  or (_13837_[3], _05302_, _05300_);
  and (_05303_, _02715_, P3_abstr[4]);
  nand (_05304_, _04107_, _03213_);
  or (_05305_, _03213_, \oc8051_golden_model_1.P3 [4]);
  and (_05306_, _05305_, _02758_);
  and (_05307_, _05306_, _05304_);
  or (_05308_, _05307_, _05303_);
  and (_05309_, _05308_, _12782_);
  nor (_05310_, \oc8051_golden_model_1.P3 [4], rst);
  nor (_05311_, _05310_, _00002_);
  or (_13837_[4], _05311_, _05309_);
  and (_05312_, _02715_, P3_abstr[5]);
  or (_05313_, _04118_, _03786_);
  or (_05314_, _03213_, \oc8051_golden_model_1.P3 [5]);
  and (_05315_, _05314_, _02758_);
  and (_05316_, _05315_, _05313_);
  or (_05317_, _05316_, _05312_);
  and (_05318_, _05317_, _12782_);
  nor (_05319_, \oc8051_golden_model_1.P3 [5], rst);
  nor (_05320_, _05319_, _00002_);
  or (_13837_[5], _05320_, _05318_);
  and (_05321_, _02715_, P3_abstr[6]);
  or (_05322_, _04129_, _03786_);
  or (_05323_, _03213_, \oc8051_golden_model_1.P3 [6]);
  and (_05324_, _05323_, _02758_);
  and (_05325_, _05324_, _05322_);
  or (_05326_, _05325_, _05321_);
  and (_05327_, _05326_, _12782_);
  nor (_05328_, \oc8051_golden_model_1.P3 [6], rst);
  nor (_05329_, _05328_, _00002_);
  or (_13837_[6], _05329_, _05327_);
  nor (_05330_, _02758_, PSW_abstr[0]);
  and (_05331_, _03987_, _03985_);
  not (_05332_, _04911_);
  or (_05333_, _04901_, _04891_);
  nand (_05334_, _04901_, _04891_);
  and (_05335_, _05334_, _05333_);
  nand (_05336_, _05335_, _05332_);
  or (_05337_, _05335_, _05332_);
  nand (_05338_, _05337_, _05336_);
  nand (_05339_, _04932_, _04922_);
  or (_05340_, _04932_, _04922_);
  and (_05341_, _05340_, _05339_);
  nand (_05342_, _05341_, _05338_);
  or (_05343_, _05341_, _05338_);
  and (_05344_, _05343_, _05342_);
  nand (_05345_, _05344_, _05331_);
  or (_05346_, _05344_, _05331_);
  nand (_05347_, _05346_, _05345_);
  or (_05348_, _04951_, _04941_);
  nand (_05349_, _04951_, _04941_);
  and (_05350_, _05349_, _05348_);
  not (_05351_, _05350_);
  nand (_05352_, _05351_, _05347_);
  or (_05353_, _05351_, _05347_);
  nand (_05354_, _05353_, _05352_);
  and (_05355_, _05354_, _02758_);
  nor (_05356_, _05355_, _05330_);
  or (_05357_, _05356_, _12786_);
  or (_05358_, _12782_, \oc8051_golden_model_1.PSW [0]);
  and (_05359_, _05358_, _13707_);
  and (_13840_[0], _05359_, _05357_);
  and (_05360_, _02715_, PSW_abstr[1]);
  and (_05361_, _03599_, _03597_);
  and (_05362_, _04072_, _03155_);
  or (_05363_, _05362_, _02715_);
  nor (_05364_, _05363_, _05361_);
  nor (_05365_, _05364_, _05360_);
  nand (_05366_, _05365_, _12782_);
  or (_05367_, _12782_, \oc8051_golden_model_1.PSW [1]);
  and (_05368_, _05367_, _13707_);
  and (_13840_[1], _05368_, _05366_);
  and (_05369_, _02715_, PSW_abstr[2]);
  and (_05370_, _03599_, _03760_);
  nor (_05371_, _04083_, _03599_);
  or (_05372_, _05371_, _02715_);
  nor (_05373_, _05372_, _05370_);
  nor (_05374_, _05373_, _05369_);
  nand (_05375_, _05374_, _12782_);
  or (_05376_, _12782_, \oc8051_golden_model_1.PSW [2]);
  and (_05377_, _05376_, _13707_);
  and (_13840_[2], _05377_, _05375_);
  and (_05378_, _02715_, PSW_abstr[3]);
  nor (_05379_, _03155_, \oc8051_golden_model_1.PSW [3]);
  and (_05380_, _04096_, _03155_);
  or (_05381_, _05380_, _02715_);
  nor (_05382_, _05381_, _05379_);
  nor (_05383_, _05382_, _05378_);
  nand (_05384_, _05383_, _12782_);
  or (_05385_, _12782_, \oc8051_golden_model_1.PSW [3]);
  and (_05386_, _05385_, _13707_);
  and (_13840_[3], _05386_, _05384_);
  and (_05387_, _02715_, PSW_abstr[4]);
  not (_05388_, \oc8051_golden_model_1.PSW [4]);
  and (_05389_, _03599_, _05388_);
  and (_05390_, _04107_, _03155_);
  or (_05391_, _05390_, _02715_);
  nor (_05392_, _05391_, _05389_);
  nor (_05393_, _05392_, _05387_);
  nand (_05394_, _05393_, _12782_);
  or (_05395_, _12782_, \oc8051_golden_model_1.PSW [4]);
  and (_05396_, _05395_, _13707_);
  and (_13840_[4], _05396_, _05394_);
  and (_05397_, _02715_, PSW_abstr[5]);
  not (_05398_, \oc8051_golden_model_1.PSW [5]);
  and (_05399_, _03599_, _05398_);
  nor (_05400_, _04118_, _03599_);
  or (_05401_, _05400_, _02715_);
  nor (_05402_, _05401_, _05399_);
  or (_05403_, _05402_, _05397_);
  or (_05404_, _05403_, _12786_);
  or (_05405_, _12782_, \oc8051_golden_model_1.PSW [5]);
  and (_05406_, _05405_, _13707_);
  and (_13840_[5], _05406_, _05404_);
  and (_05407_, _02715_, PSW_abstr[6]);
  or (_05408_, _04129_, _03599_);
  nor (_05409_, _03155_, \oc8051_golden_model_1.PSW [6]);
  nor (_05410_, _05409_, _02715_);
  and (_05411_, _05410_, _05408_);
  or (_05412_, _05411_, _05407_);
  or (_05413_, _05412_, _12786_);
  or (_05414_, _12782_, \oc8051_golden_model_1.PSW [6]);
  and (_05415_, _05414_, _13707_);
  and (_13840_[6], _05415_, _05413_);
  and (_13838_[0], \oc8051_golden_model_1.PCON [0], _13707_);
  and (_13838_[1], \oc8051_golden_model_1.PCON [1], _13707_);
  and (_13838_[2], \oc8051_golden_model_1.PCON [2], _13707_);
  and (_13838_[3], \oc8051_golden_model_1.PCON [3], _13707_);
  and (_13838_[4], \oc8051_golden_model_1.PCON [4], _13707_);
  and (_13838_[5], \oc8051_golden_model_1.PCON [5], _13707_);
  and (_13838_[6], \oc8051_golden_model_1.PCON [6], _13707_);
  and (_13841_[0], \oc8051_golden_model_1.SBUF [0], _13707_);
  and (_13841_[1], \oc8051_golden_model_1.SBUF [1], _13707_);
  and (_13841_[2], \oc8051_golden_model_1.SBUF [2], _13707_);
  and (_13841_[3], \oc8051_golden_model_1.SBUF [3], _13707_);
  and (_13841_[4], \oc8051_golden_model_1.SBUF [4], _13707_);
  and (_13841_[5], \oc8051_golden_model_1.SBUF [5], _13707_);
  and (_13841_[6], \oc8051_golden_model_1.SBUF [6], _13707_);
  and (_13842_[0], \oc8051_golden_model_1.SCON [0], _13707_);
  and (_13842_[1], \oc8051_golden_model_1.SCON [1], _13707_);
  and (_13842_[2], \oc8051_golden_model_1.SCON [2], _13707_);
  and (_13842_[3], \oc8051_golden_model_1.SCON [3], _13707_);
  and (_13842_[4], \oc8051_golden_model_1.SCON [4], _13707_);
  and (_13842_[5], \oc8051_golden_model_1.SCON [5], _13707_);
  and (_13842_[6], \oc8051_golden_model_1.SCON [6], _13707_);
  and (_05416_, _02715_, SP_abstr[0]);
  or (_05417_, _03067_, \oc8051_golden_model_1.SP [0]);
  and (_05418_, _03672_, _02758_);
  and (_05419_, _05418_, _05417_);
  or (_05420_, _05419_, _05416_);
  and (_05421_, _05420_, _12782_);
  nor (_05422_, \oc8051_golden_model_1.SP [0], rst);
  nor (_05423_, _05422_, _00002_);
  or (_13843_[0], _05423_, _05421_);
  and (_05424_, _02715_, SP_abstr[1]);
  nand (_05425_, _04072_, _03067_);
  or (_05426_, _03067_, \oc8051_golden_model_1.SP [1]);
  and (_05427_, _05426_, _02758_);
  and (_05428_, _05427_, _05425_);
  or (_05429_, _05428_, _05424_);
  and (_05430_, _05429_, _12782_);
  nor (_05431_, \oc8051_golden_model_1.SP [1], rst);
  nor (_05432_, _05431_, _00002_);
  or (_13843_[1], _05432_, _05430_);
  and (_05433_, _02715_, SP_abstr[2]);
  or (_05434_, _04083_, _03068_);
  or (_05435_, _03067_, \oc8051_golden_model_1.SP [2]);
  and (_05436_, _05435_, _02758_);
  and (_05437_, _05436_, _05434_);
  or (_05438_, _05437_, _05433_);
  and (_05439_, _05438_, _12782_);
  nor (_05440_, \oc8051_golden_model_1.SP [2], rst);
  nor (_05441_, _05440_, _00002_);
  or (_13843_[2], _05441_, _05439_);
  nand (_05442_, _04096_, _03067_);
  or (_05443_, _03067_, \oc8051_golden_model_1.SP [3]);
  and (_05444_, _05443_, _02758_);
  and (_05445_, _05444_, _05442_);
  and (_05446_, _02715_, SP_abstr[3]);
  or (_05447_, _05446_, _12786_);
  or (_05448_, _05447_, _05445_);
  or (_05449_, _12782_, \oc8051_golden_model_1.SP [3]);
  and (_05450_, _05449_, _13707_);
  and (_13843_[3], _05450_, _05448_);
  nand (_05451_, _04107_, _03067_);
  or (_05452_, _03067_, \oc8051_golden_model_1.SP [4]);
  and (_05453_, _05452_, _02758_);
  and (_05454_, _05453_, _05451_);
  and (_05455_, _02715_, SP_abstr[4]);
  or (_05456_, _05455_, _12786_);
  or (_05457_, _05456_, _05454_);
  or (_05458_, _12782_, \oc8051_golden_model_1.SP [4]);
  and (_05459_, _05458_, _13707_);
  and (_13843_[4], _05459_, _05457_);
  or (_05460_, _04118_, _03068_);
  or (_05461_, _03067_, \oc8051_golden_model_1.SP [5]);
  and (_05462_, _05461_, _02758_);
  and (_05463_, _05462_, _05460_);
  and (_05464_, _02715_, SP_abstr[5]);
  or (_05465_, _05464_, _12786_);
  or (_05466_, _05465_, _05463_);
  or (_05467_, _12782_, \oc8051_golden_model_1.SP [5]);
  and (_05468_, _05467_, _13707_);
  and (_13843_[5], _05468_, _05466_);
  or (_05469_, _12782_, \oc8051_golden_model_1.SP [6]);
  and (_05470_, _05469_, _13707_);
  and (_05471_, _02715_, SP_abstr[6]);
  or (_05472_, _05471_, _12786_);
  or (_05473_, _04129_, _03068_);
  or (_05474_, _03067_, \oc8051_golden_model_1.SP [6]);
  and (_05475_, _05474_, _02758_);
  and (_05476_, _05475_, _05473_);
  or (_05477_, _05476_, _05472_);
  and (_13843_[6], _05477_, _05470_);
  and (_13844_[0], \oc8051_golden_model_1.TCON [0], _13707_);
  and (_13844_[1], \oc8051_golden_model_1.TCON [1], _13707_);
  and (_13844_[2], \oc8051_golden_model_1.TCON [2], _13707_);
  and (_13844_[3], \oc8051_golden_model_1.TCON [3], _13707_);
  and (_13844_[4], \oc8051_golden_model_1.TCON [4], _13707_);
  and (_13844_[5], \oc8051_golden_model_1.TCON [5], _13707_);
  and (_13844_[6], \oc8051_golden_model_1.TCON [6], _13707_);
  and (_13845_[0], \oc8051_golden_model_1.TH0 [0], _13707_);
  and (_13845_[1], \oc8051_golden_model_1.TH0 [1], _13707_);
  and (_13845_[2], \oc8051_golden_model_1.TH0 [2], _13707_);
  and (_13845_[3], \oc8051_golden_model_1.TH0 [3], _13707_);
  and (_13845_[4], \oc8051_golden_model_1.TH0 [4], _13707_);
  and (_13845_[5], \oc8051_golden_model_1.TH0 [5], _13707_);
  and (_13845_[6], \oc8051_golden_model_1.TH0 [6], _13707_);
  and (_13846_[0], \oc8051_golden_model_1.TH1 [0], _13707_);
  and (_13846_[1], \oc8051_golden_model_1.TH1 [1], _13707_);
  and (_13846_[2], \oc8051_golden_model_1.TH1 [2], _13707_);
  and (_13846_[3], \oc8051_golden_model_1.TH1 [3], _13707_);
  and (_13846_[4], \oc8051_golden_model_1.TH1 [4], _13707_);
  and (_13846_[5], \oc8051_golden_model_1.TH1 [5], _13707_);
  and (_13846_[6], \oc8051_golden_model_1.TH1 [6], _13707_);
  and (_13847_[0], \oc8051_golden_model_1.TL0 [0], _13707_);
  and (_13847_[1], \oc8051_golden_model_1.TL0 [1], _13707_);
  and (_13847_[2], \oc8051_golden_model_1.TL0 [2], _13707_);
  and (_13847_[3], \oc8051_golden_model_1.TL0 [3], _13707_);
  and (_13847_[4], \oc8051_golden_model_1.TL0 [4], _13707_);
  and (_13847_[5], \oc8051_golden_model_1.TL0 [5], _13707_);
  and (_13847_[6], \oc8051_golden_model_1.TL0 [6], _13707_);
  and (_13848_[0], \oc8051_golden_model_1.TL1 [0], _13707_);
  and (_13848_[1], \oc8051_golden_model_1.TL1 [1], _13707_);
  and (_13848_[2], \oc8051_golden_model_1.TL1 [2], _13707_);
  and (_13848_[3], \oc8051_golden_model_1.TL1 [3], _13707_);
  and (_13848_[4], \oc8051_golden_model_1.TL1 [4], _13707_);
  and (_13848_[5], \oc8051_golden_model_1.TL1 [5], _13707_);
  and (_13848_[6], \oc8051_golden_model_1.TL1 [6], _13707_);
  and (_13849_[0], \oc8051_golden_model_1.TMOD [0], _13707_);
  and (_13849_[1], \oc8051_golden_model_1.TMOD [1], _13707_);
  and (_13849_[2], \oc8051_golden_model_1.TMOD [2], _13707_);
  and (_13849_[3], \oc8051_golden_model_1.TMOD [3], _13707_);
  and (_13849_[4], \oc8051_golden_model_1.TMOD [4], _13707_);
  and (_13849_[5], \oc8051_golden_model_1.TMOD [5], _13707_);
  and (_13849_[6], \oc8051_golden_model_1.TMOD [6], _13707_);
  and (_05478_, _02715_, XRAM_ADDR_abstr[0]);
  or (_05479_, _05478_, _12786_);
  or (_05480_, _12782_, \oc8051_golden_model_1.XRAM_ADDR [0]);
  and (_05481_, _05480_, _13707_);
  and (_13850_[0], _05481_, _05479_);
  and (_05482_, _02715_, XRAM_ADDR_abstr[1]);
  or (_05483_, _05482_, _12786_);
  or (_05484_, _12782_, \oc8051_golden_model_1.XRAM_ADDR [1]);
  and (_05485_, _05484_, _13707_);
  and (_13850_[1], _05485_, _05483_);
  and (_05486_, _02715_, XRAM_ADDR_abstr[2]);
  or (_05487_, _05486_, _12786_);
  or (_05488_, _12782_, \oc8051_golden_model_1.XRAM_ADDR [2]);
  and (_05489_, _05488_, _13707_);
  and (_13850_[2], _05489_, _05487_);
  and (_05490_, _02715_, XRAM_ADDR_abstr[3]);
  or (_05491_, _05490_, _12786_);
  or (_05492_, _12782_, \oc8051_golden_model_1.XRAM_ADDR [3]);
  and (_05493_, _05492_, _13707_);
  and (_13850_[3], _05493_, _05491_);
  and (_05494_, _02715_, XRAM_ADDR_abstr[4]);
  or (_05495_, _05494_, _12786_);
  or (_05496_, _12782_, \oc8051_golden_model_1.XRAM_ADDR [4]);
  and (_05497_, _05496_, _13707_);
  and (_13850_[4], _05497_, _05495_);
  and (_05498_, _02715_, XRAM_ADDR_abstr[5]);
  or (_05499_, _05498_, _12786_);
  or (_05500_, _12782_, \oc8051_golden_model_1.XRAM_ADDR [5]);
  and (_05501_, _05500_, _13707_);
  and (_13850_[5], _05501_, _05499_);
  and (_05502_, _02715_, XRAM_ADDR_abstr[6]);
  or (_05503_, _05502_, _12786_);
  or (_05504_, _12782_, \oc8051_golden_model_1.XRAM_ADDR [6]);
  and (_05505_, _05504_, _13707_);
  and (_13850_[6], _05505_, _05503_);
  and (_05506_, _02715_, XRAM_ADDR_abstr[7]);
  or (_05507_, _05506_, _12786_);
  or (_05508_, _12782_, \oc8051_golden_model_1.XRAM_ADDR [7]);
  and (_05509_, _05508_, _13707_);
  and (_13850_[7], _05509_, _05507_);
  and (_05510_, _02715_, XRAM_ADDR_abstr[8]);
  or (_05511_, _05510_, _12786_);
  or (_05512_, _12782_, \oc8051_golden_model_1.XRAM_ADDR [8]);
  and (_05513_, _05512_, _13707_);
  and (_13850_[8], _05513_, _05511_);
  and (_05514_, _02715_, XRAM_ADDR_abstr[9]);
  or (_05515_, _05514_, _12786_);
  or (_05516_, _12782_, \oc8051_golden_model_1.XRAM_ADDR [9]);
  and (_05517_, _05516_, _13707_);
  and (_13850_[9], _05517_, _05515_);
  and (_05518_, _02715_, XRAM_ADDR_abstr[10]);
  or (_05519_, _05518_, _12786_);
  or (_05520_, _12782_, \oc8051_golden_model_1.XRAM_ADDR [10]);
  and (_05521_, _05520_, _13707_);
  and (_13850_[10], _05521_, _05519_);
  and (_05522_, _02715_, XRAM_ADDR_abstr[11]);
  or (_05523_, _05522_, _12786_);
  or (_05524_, _12782_, \oc8051_golden_model_1.XRAM_ADDR [11]);
  and (_05525_, _05524_, _13707_);
  and (_13850_[11], _05525_, _05523_);
  and (_05526_, _02715_, XRAM_ADDR_abstr[12]);
  or (_05527_, _05526_, _12786_);
  or (_05528_, _12782_, \oc8051_golden_model_1.XRAM_ADDR [12]);
  and (_05529_, _05528_, _13707_);
  and (_13850_[12], _05529_, _05527_);
  and (_05530_, _02715_, XRAM_ADDR_abstr[13]);
  or (_05531_, _05530_, _12786_);
  or (_05532_, _12782_, \oc8051_golden_model_1.XRAM_ADDR [13]);
  and (_05533_, _05532_, _13707_);
  and (_13850_[13], _05533_, _05531_);
  and (_05534_, _02715_, XRAM_ADDR_abstr[14]);
  or (_05535_, _05534_, _12786_);
  or (_05536_, _12782_, \oc8051_golden_model_1.XRAM_ADDR [14]);
  and (_05537_, _05536_, _13707_);
  and (_13850_[14], _05537_, _05535_);
  and (_05538_, _02715_, PC_abstr[0]);
  not (_05539_, _05538_);
  and (_05540_, _05539_, _02764_);
  nand (_05541_, _05540_, _12782_);
  or (_05542_, _12782_, \oc8051_golden_model_1.PC [0]);
  and (_05543_, _05542_, _13707_);
  and (_13839_[0], _05543_, _05541_);
  and (_05544_, _02758_, \oc8051_golden_model_1.PC [1]);
  nor (_05545_, _02758_, PC_abstr[1]);
  nor (_05546_, _05545_, _05544_);
  or (_05547_, _05546_, _12786_);
  or (_05548_, _12782_, \oc8051_golden_model_1.PC [1]);
  and (_05549_, _05548_, _13707_);
  and (_13839_[1], _05549_, _05547_);
  nor (_05550_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [1]);
  nor (_05551_, _05550_, _02720_);
  nor (_05552_, _05551_, _02715_);
  nor (_05553_, _02758_, PC_abstr[2]);
  nor (_05554_, _05553_, _05552_);
  or (_05555_, _05554_, _12786_);
  or (_05556_, _12782_, \oc8051_golden_model_1.PC [2]);
  and (_05557_, _05556_, _13707_);
  and (_13839_[2], _05557_, _05555_);
  nor (_05558_, _02758_, PC_abstr[3]);
  nor (_05559_, _02720_, \oc8051_golden_model_1.PC [3]);
  nor (_05560_, _05559_, _02721_);
  nor (_05561_, _05560_, _02715_);
  nor (_05562_, _05561_, _05558_);
  or (_05563_, _05562_, _12786_);
  or (_05564_, _12782_, \oc8051_golden_model_1.PC [3]);
  and (_05565_, _05564_, _13707_);
  and (_13839_[3], _05565_, _05563_);
  nor (_05566_, _02721_, \oc8051_golden_model_1.PC [4]);
  nor (_05567_, _05566_, _02722_);
  nor (_05568_, _05567_, _02715_);
  nor (_05569_, _02758_, PC_abstr[4]);
  nor (_05570_, _05569_, _05568_);
  or (_05571_, _05570_, _12786_);
  or (_05572_, _12782_, \oc8051_golden_model_1.PC [4]);
  and (_05573_, _05572_, _13707_);
  and (_13839_[4], _05573_, _05571_);
  nor (_05574_, _02722_, \oc8051_golden_model_1.PC [5]);
  nor (_05575_, _05574_, _02723_);
  nor (_05576_, _05575_, _02715_);
  nor (_05577_, _02758_, PC_abstr[5]);
  nor (_05578_, _05577_, _05576_);
  or (_05579_, _05578_, _12786_);
  or (_05580_, _12782_, \oc8051_golden_model_1.PC [5]);
  and (_05581_, _05580_, _13707_);
  and (_13839_[5], _05581_, _05579_);
  nor (_05582_, _02723_, \oc8051_golden_model_1.PC [6]);
  nor (_05583_, _05582_, _02724_);
  nor (_05584_, _05583_, _02715_);
  nor (_05585_, _02758_, PC_abstr[6]);
  nor (_05586_, _05585_, _05584_);
  or (_05587_, _05586_, _12786_);
  or (_05588_, _12782_, \oc8051_golden_model_1.PC [6]);
  and (_05589_, _05588_, _13707_);
  and (_13839_[6], _05589_, _05587_);
  nor (_05590_, _02724_, \oc8051_golden_model_1.PC [7]);
  nor (_05591_, _05590_, _02725_);
  nor (_05592_, _05591_, _02715_);
  nor (_05593_, _02758_, PC_abstr[7]);
  nor (_05594_, _05593_, _05592_);
  or (_05595_, _05594_, _12786_);
  or (_05596_, _12782_, \oc8051_golden_model_1.PC [7]);
  and (_05597_, _05596_, _13707_);
  and (_13839_[7], _05597_, _05595_);
  nor (_05598_, _02725_, \oc8051_golden_model_1.PC [8]);
  nor (_05599_, _05598_, _02726_);
  nor (_05600_, _05599_, _02715_);
  nor (_05601_, _02758_, PC_abstr[8]);
  nor (_05602_, _05601_, _05600_);
  or (_05603_, _05602_, _12786_);
  or (_05604_, _12782_, \oc8051_golden_model_1.PC [8]);
  and (_05605_, _05604_, _13707_);
  and (_13839_[8], _05605_, _05603_);
  nor (_05606_, _02726_, \oc8051_golden_model_1.PC [9]);
  nor (_05607_, _05606_, _02727_);
  nor (_05608_, _05607_, _02715_);
  nor (_05609_, _02758_, PC_abstr[9]);
  nor (_05610_, _05609_, _05608_);
  or (_05611_, _05610_, _12786_);
  or (_05612_, _12782_, \oc8051_golden_model_1.PC [9]);
  and (_05613_, _05612_, _13707_);
  and (_13839_[9], _05613_, _05611_);
  nor (_05614_, _02727_, \oc8051_golden_model_1.PC [10]);
  nor (_05615_, _05614_, _02728_);
  nor (_05616_, _05615_, _02715_);
  nor (_05617_, _02758_, PC_abstr[10]);
  nor (_05618_, _05617_, _05616_);
  or (_05619_, _05618_, _12786_);
  or (_05620_, _12782_, \oc8051_golden_model_1.PC [10]);
  and (_05621_, _05620_, _13707_);
  and (_13839_[10], _05621_, _05619_);
  nor (_05622_, _02728_, \oc8051_golden_model_1.PC [11]);
  nor (_05623_, _05622_, _02729_);
  nor (_05624_, _05623_, _02715_);
  nor (_05625_, _02758_, PC_abstr[11]);
  nor (_05626_, _05625_, _05624_);
  or (_05627_, _05626_, _12786_);
  or (_05628_, _12782_, \oc8051_golden_model_1.PC [11]);
  and (_05629_, _05628_, _13707_);
  and (_13839_[11], _05629_, _05627_);
  nor (_05630_, _02729_, \oc8051_golden_model_1.PC [12]);
  nor (_05631_, _05630_, _02730_);
  nor (_05632_, _05631_, _02715_);
  nor (_05633_, _02758_, PC_abstr[12]);
  nor (_05634_, _05633_, _05632_);
  or (_05635_, _05634_, _12786_);
  or (_05636_, _12782_, \oc8051_golden_model_1.PC [12]);
  and (_05637_, _05636_, _13707_);
  and (_13839_[12], _05637_, _05635_);
  nor (_05638_, _02730_, \oc8051_golden_model_1.PC [13]);
  nor (_05639_, _05638_, _02731_);
  nor (_05640_, _05639_, _02715_);
  nor (_05641_, _02758_, PC_abstr[13]);
  nor (_05642_, _05641_, _05640_);
  or (_05643_, _05642_, _12786_);
  or (_05644_, _12782_, \oc8051_golden_model_1.PC [13]);
  and (_05645_, _05644_, _13707_);
  and (_13839_[13], _05645_, _05643_);
  nor (_05646_, _02731_, \oc8051_golden_model_1.PC [14]);
  nor (_05647_, _05646_, _02732_);
  nor (_05648_, _05647_, _02715_);
  nor (_05649_, _02758_, PC_abstr[14]);
  nor (_05650_, _05649_, _05648_);
  or (_05651_, _05650_, _12786_);
  or (_05652_, _12782_, \oc8051_golden_model_1.PC [14]);
  and (_05653_, _05652_, _13707_);
  and (_13839_[14], _05653_, _05651_);
  and (_05654_, _02715_, XRAM_DATA_OUT_abstr[0]);
  or (_05655_, _05654_, _12786_);
  or (_05656_, _12782_, \oc8051_golden_model_1.XRAM_DATA_OUT [0]);
  and (_05657_, _05656_, _13707_);
  and (_13851_[0], _05657_, _05655_);
  and (_05658_, _02715_, XRAM_DATA_OUT_abstr[1]);
  or (_05659_, _05658_, _12786_);
  or (_05660_, _12782_, \oc8051_golden_model_1.XRAM_DATA_OUT [1]);
  and (_05661_, _05660_, _13707_);
  and (_13851_[1], _05661_, _05659_);
  and (_05662_, _02715_, XRAM_DATA_OUT_abstr[2]);
  or (_05663_, _05662_, _12786_);
  or (_05664_, _12782_, \oc8051_golden_model_1.XRAM_DATA_OUT [2]);
  and (_05665_, _05664_, _13707_);
  and (_13851_[2], _05665_, _05663_);
  and (_05666_, _02715_, XRAM_DATA_OUT_abstr[3]);
  or (_05667_, _05666_, _12786_);
  or (_05668_, _12782_, \oc8051_golden_model_1.XRAM_DATA_OUT [3]);
  and (_05669_, _05668_, _13707_);
  and (_13851_[3], _05669_, _05667_);
  and (_05670_, _02715_, XRAM_DATA_OUT_abstr[4]);
  or (_05671_, _05670_, _12786_);
  or (_05672_, _12782_, \oc8051_golden_model_1.XRAM_DATA_OUT [4]);
  and (_05673_, _05672_, _13707_);
  and (_13851_[4], _05673_, _05671_);
  and (_05674_, _02715_, XRAM_DATA_OUT_abstr[5]);
  or (_05675_, _05674_, _12786_);
  or (_05676_, _12782_, \oc8051_golden_model_1.XRAM_DATA_OUT [5]);
  and (_05677_, _05676_, _13707_);
  and (_13851_[5], _05677_, _05675_);
  and (_05678_, _02715_, XRAM_DATA_OUT_abstr[6]);
  or (_05679_, _05678_, _12786_);
  or (_05680_, _12782_, \oc8051_golden_model_1.XRAM_DATA_OUT [6]);
  and (_05681_, _05680_, _13707_);
  and (_13851_[6], _05681_, _05679_);
  and (_00007_[6], _00854_, _13707_);
  and (_00007_[5], _00870_, _13707_);
  and (_00007_[4], _00836_, _13707_);
  and (_00007_[3], _00845_, _13707_);
  and (_00007_[2], _00861_, _13707_);
  and (_00007_[1], _00877_, _13707_);
  and (_00007_[0], _00829_, _13707_);
  and (_00006_[6], _00924_, _13707_);
  and (_00006_[5], _00940_, _13707_);
  and (_00006_[4], _00906_, _13707_);
  and (_00006_[3], _00915_, _13707_);
  and (_00006_[2], _00931_, _13707_);
  and (_00006_[1], _00947_, _13707_);
  and (_00006_[0], _00899_, _13707_);
  and (_00005_[6], _00772_, _13707_);
  and (_00005_[5], _00756_, _13707_);
  and (_00005_[4], _00739_, _13707_);
  and (_00005_[3], _00748_, _13707_);
  and (_00005_[2], _00779_, _13707_);
  and (_00005_[1], _00763_, _13707_);
  and (_00005_[0], _00732_, _13707_);
  and (_00004_[6], _00994_, _13707_);
  and (_00004_[5], _01010_, _13707_);
  and (_00004_[4], _00985_, _13707_);
  and (_00004_[3], _00970_, _13707_);
  and (_00004_[2], _01001_, _13707_);
  and (_00004_[1], _01018_, _13707_);
  and (_00004_[0], _00978_, _13707_);
  and (_05682_, _12786_, xram_data_in_reg[6]);
  and (_05683_, _12782_, xram_data_in[6]);
  or (_05684_, _05683_, _05682_);
  and (_00010_[6], _05684_, _13707_);
  and (_05685_, _12786_, xram_data_in_reg[5]);
  and (_05686_, _12782_, xram_data_in[5]);
  or (_05687_, _05686_, _05685_);
  and (_00010_[5], _05687_, _13707_);
  and (_05688_, _12786_, xram_data_in_reg[4]);
  and (_05689_, _12782_, xram_data_in[4]);
  or (_05690_, _05689_, _05688_);
  and (_00010_[4], _05690_, _13707_);
  and (_05691_, _12786_, xram_data_in_reg[3]);
  and (_05692_, _12782_, xram_data_in[3]);
  or (_05693_, _05692_, _05691_);
  and (_00010_[3], _05693_, _13707_);
  and (_05694_, _12786_, xram_data_in_reg[2]);
  and (_05695_, _12782_, xram_data_in[2]);
  or (_05696_, _05695_, _05694_);
  and (_00010_[2], _05696_, _13707_);
  and (_05697_, _12786_, xram_data_in_reg[1]);
  and (_05698_, _12782_, xram_data_in[1]);
  or (_05699_, _05698_, _05697_);
  and (_00010_[1], _05699_, _13707_);
  and (_05700_, _12786_, xram_data_in_reg[0]);
  and (_05701_, _12782_, xram_data_in[0]);
  or (_05702_, _05701_, _05700_);
  and (_00010_[0], _05702_, _13707_);
  not (_05703_, _00684_);
  nand (_05704_, _05356_, _05703_);
  or (_05705_, _05356_, _05703_);
  nand (_05706_, _05393_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  or (_05707_, _05393_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_05708_, _05707_, _05706_);
  or (_05709_, _05383_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  nand (_05710_, _05383_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_05711_, _05710_, _05709_);
  nand (_05712_, _05365_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  or (_05713_, _05365_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_05714_, _05713_, _05712_);
  nand (_05715_, _05374_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_05716_, _05374_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  and (_05717_, _05716_, _05715_);
  and (_05718_, _05717_, _05714_);
  and (_05719_, _05718_, _05711_);
  and (_05720_, _05719_, _05708_);
  nand (_05721_, _03915_, _09391_);
  or (_05722_, _03915_, _09391_);
  and (_05723_, _05722_, _05721_);
  nand (_05724_, _05412_, _08273_);
  or (_05725_, _05412_, _08273_);
  and (_05726_, _05725_, _05724_);
  not (_05727_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  or (_05728_, _05403_, _05727_);
  nand (_05729_, _05403_, _05727_);
  and (_05730_, _05729_, _05728_);
  and (_05731_, _05730_, _05726_);
  and (_05732_, _05731_, _05723_);
  and (_05733_, _05732_, _05720_);
  not (_05734_, \oc8051_golden_model_1.SP [7]);
  nand (_05735_, _08999_, _05734_);
  or (_05736_, _08999_, _05734_);
  and (_05737_, _05736_, _05735_);
  or (_05738_, _09043_, \oc8051_golden_model_1.SP [6]);
  nand (_05739_, _09043_, \oc8051_golden_model_1.SP [6]);
  and (_05740_, _05739_, _05738_);
  nand (_05741_, _09037_, \oc8051_golden_model_1.SP [5]);
  or (_05742_, _09037_, \oc8051_golden_model_1.SP [5]);
  and (_05743_, _05742_, _05741_);
  or (_05744_, _09031_, \oc8051_golden_model_1.SP [4]);
  nand (_05745_, _09031_, \oc8051_golden_model_1.SP [4]);
  and (_05746_, _05745_, _05744_);
  or (_05747_, _09025_, \oc8051_golden_model_1.SP [3]);
  nand (_05748_, _09025_, \oc8051_golden_model_1.SP [3]);
  and (_05749_, _05748_, _05747_);
  nor (_05750_, \oc8051_golden_model_1.IRAM[5] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  and (_05751_, \oc8051_golden_model_1.IRAM[5] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  nor (_05752_, _05751_, _05750_);
  nor (_05753_, \oc8051_golden_model_1.IRAM[5] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  and (_05754_, \oc8051_golden_model_1.IRAM[5] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  nor (_05755_, _05754_, _05753_);
  nor (_05756_, _05755_, _05752_);
  and (_05757_, \oc8051_golden_model_1.IRAM[5] [5], _10756_);
  nor (_05758_, \oc8051_golden_model_1.IRAM[5] [5], _10756_);
  nor (_05759_, _05758_, _05757_);
  nor (_05760_, \oc8051_golden_model_1.IRAM[5] [4], _10753_);
  and (_05761_, \oc8051_golden_model_1.IRAM[5] [4], _10753_);
  nor (_05762_, _05761_, _05760_);
  and (_05763_, _05762_, _05759_);
  and (_05764_, _05763_, _05756_);
  nor (_05765_, \oc8051_golden_model_1.IRAM[4] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  and (_05766_, \oc8051_golden_model_1.IRAM[4] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  nor (_05767_, _05766_, _05765_);
  not (_05768_, _05767_);
  and (_05769_, \oc8051_golden_model_1.IRAM[4] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  nor (_05770_, \oc8051_golden_model_1.IRAM[4] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  or (_05771_, _05770_, _05769_);
  and (_05772_, _05771_, _05768_);
  nor (_05773_, \oc8051_golden_model_1.IRAM[4] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  and (_05774_, \oc8051_golden_model_1.IRAM[4] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  nor (_05775_, _05774_, _05773_);
  nand (_05776_, \oc8051_golden_model_1.IRAM[4] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  or (_05777_, \oc8051_golden_model_1.IRAM[4] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  and (_05778_, _05777_, _05776_);
  nor (_05779_, _05778_, _05775_);
  and (_05780_, _05779_, _05772_);
  and (_05781_, _05780_, _05764_);
  and (_05782_, _03711_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  and (_05783_, \oc8051_golden_model_1.IRAM[7] [2], _10794_);
  nor (_05784_, _05783_, _05782_);
  nand (_05785_, \oc8051_golden_model_1.IRAM[7] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  or (_05786_, \oc8051_golden_model_1.IRAM[7] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  and (_05787_, _05786_, _05785_);
  not (_05788_, _05787_);
  and (_05789_, _05788_, _05784_);
  nor (_05790_, \oc8051_golden_model_1.IRAM[7] [7], _10570_);
  and (_05791_, \oc8051_golden_model_1.IRAM[7] [7], _10570_);
  nor (_05792_, _05791_, _05790_);
  nand (_05793_, \oc8051_golden_model_1.IRAM[7] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  or (_05794_, \oc8051_golden_model_1.IRAM[7] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  and (_05795_, _05794_, _05793_);
  not (_05796_, _05795_);
  and (_05797_, _05796_, _05792_);
  and (_05798_, _05797_, _05789_);
  nor (_05799_, \oc8051_golden_model_1.IRAM[6] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  and (_05800_, \oc8051_golden_model_1.IRAM[6] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  nor (_05801_, _05800_, _05799_);
  nor (_05802_, \oc8051_golden_model_1.IRAM[6] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  and (_05803_, \oc8051_golden_model_1.IRAM[6] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  nor (_05804_, _05803_, _05802_);
  nor (_05805_, _05804_, _05801_);
  nor (_05806_, \oc8051_golden_model_1.IRAM[6] [4], _10775_);
  and (_05807_, \oc8051_golden_model_1.IRAM[6] [4], _10775_);
  nor (_05808_, _05807_, _05806_);
  nor (_05809_, \oc8051_golden_model_1.IRAM[6] [5], _10778_);
  and (_05810_, \oc8051_golden_model_1.IRAM[6] [5], _10778_);
  nor (_05811_, _05810_, _05809_);
  and (_05812_, _05811_, _05808_);
  and (_05813_, _05812_, _05805_);
  and (_05814_, _05813_, _05798_);
  and (_05815_, _05814_, _05781_);
  nor (_05816_, \oc8051_golden_model_1.IRAM[1] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  and (_05817_, \oc8051_golden_model_1.IRAM[1] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  nor (_05818_, _05817_, _05816_);
  not (_05819_, _05818_);
  and (_05820_, \oc8051_golden_model_1.IRAM[1] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  nor (_05821_, \oc8051_golden_model_1.IRAM[1] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  or (_05822_, _05821_, _05820_);
  and (_05823_, _05822_, _05819_);
  nor (_05824_, \oc8051_golden_model_1.IRAM[1] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  and (_05825_, \oc8051_golden_model_1.IRAM[1] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  nor (_05826_, _05825_, _05824_);
  not (_05827_, _05826_);
  and (_05828_, \oc8051_golden_model_1.IRAM[1] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  nor (_05829_, \oc8051_golden_model_1.IRAM[1] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  or (_05830_, _05829_, _05828_);
  and (_05831_, _05830_, _05827_);
  and (_05832_, _05831_, _05823_);
  and (_05833_, _03623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  and (_05834_, \oc8051_golden_model_1.IRAM[0] [0], _10625_);
  nor (_05835_, _05834_, _05833_);
  nor (_05836_, \oc8051_golden_model_1.IRAM[0] [1], _10629_);
  and (_05837_, \oc8051_golden_model_1.IRAM[0] [1], _10629_);
  nor (_05838_, _05837_, _05836_);
  and (_05839_, _05838_, _05835_);
  nor (_05840_, \oc8051_golden_model_1.IRAM[0] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  and (_05841_, \oc8051_golden_model_1.IRAM[0] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  nor (_05842_, _05841_, _05840_);
  nor (_05843_, \oc8051_golden_model_1.IRAM[0] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  and (_05844_, \oc8051_golden_model_1.IRAM[0] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nor (_05845_, _05844_, _05843_);
  nor (_05846_, _05845_, _05842_);
  and (_05847_, _05846_, _05839_);
  and (_05848_, _05847_, _05832_);
  and (_05849_, _03628_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  and (_05850_, \oc8051_golden_model_1.IRAM[3] [0], _10698_);
  nor (_05851_, _05850_, _05849_);
  nor (_05852_, \oc8051_golden_model_1.IRAM[3] [1], _10701_);
  and (_05853_, \oc8051_golden_model_1.IRAM[3] [1], _10701_);
  nor (_05854_, _05853_, _05852_);
  and (_05855_, _05854_, _05851_);
  nor (_05856_, \oc8051_golden_model_1.IRAM[3] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  and (_05857_, \oc8051_golden_model_1.IRAM[3] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  nor (_05858_, _05857_, _05856_);
  nor (_05859_, \oc8051_golden_model_1.IRAM[3] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  and (_05860_, \oc8051_golden_model_1.IRAM[3] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  nor (_05861_, _05860_, _05859_);
  nor (_05862_, _05861_, _05858_);
  and (_05863_, _05862_, _05855_);
  and (_05864_, _03721_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  and (_05865_, \oc8051_golden_model_1.IRAM[2] [2], _10680_);
  nor (_05866_, _05865_, _05864_);
  nand (_05867_, \oc8051_golden_model_1.IRAM[2] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or (_05868_, \oc8051_golden_model_1.IRAM[2] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  and (_05869_, _05868_, _05867_);
  not (_05870_, _05869_);
  and (_05871_, _05870_, _05866_);
  and (_05872_, \oc8051_golden_model_1.IRAM[2] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  nor (_05873_, \oc8051_golden_model_1.IRAM[2] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  or (_05874_, _05873_, _05872_);
  nor (_05875_, \oc8051_golden_model_1.IRAM[2] [7], _10694_);
  and (_05876_, \oc8051_golden_model_1.IRAM[2] [7], _10694_);
  nor (_05877_, _05876_, _05875_);
  and (_05878_, _05877_, _05874_);
  and (_05879_, _05878_, _05871_);
  and (_05880_, _05879_, _05863_);
  and (_05881_, _05880_, _05848_);
  and (_05882_, _05881_, _05815_);
  nor (_05883_, \oc8051_golden_model_1.IRAM[13] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  and (_05884_, \oc8051_golden_model_1.IRAM[13] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  nor (_05885_, _05884_, _05883_);
  not (_05886_, _05885_);
  and (_05887_, \oc8051_golden_model_1.IRAM[13] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  nor (_05888_, \oc8051_golden_model_1.IRAM[13] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  or (_05889_, _05888_, _05887_);
  and (_05890_, _05889_, _05886_);
  nor (_05891_, \oc8051_golden_model_1.IRAM[13] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  and (_05892_, \oc8051_golden_model_1.IRAM[13] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  nor (_05893_, _05892_, _05891_);
  nand (_05894_, \oc8051_golden_model_1.IRAM[13] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  or (_05895_, \oc8051_golden_model_1.IRAM[13] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  and (_05896_, _05895_, _05894_);
  nor (_05897_, _05896_, _05893_);
  and (_05898_, _05897_, _05890_);
  nor (_05899_, \oc8051_golden_model_1.IRAM[12] [0], _10897_);
  and (_05900_, \oc8051_golden_model_1.IRAM[12] [0], _10897_);
  nor (_05901_, _05900_, _05899_);
  nor (_05902_, \oc8051_golden_model_1.IRAM[12] [1], _10900_);
  and (_05903_, \oc8051_golden_model_1.IRAM[12] [1], _10900_);
  nor (_05904_, _05903_, _05902_);
  and (_05905_, _05904_, _05901_);
  nor (_05906_, \oc8051_golden_model_1.IRAM[12] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  and (_05907_, \oc8051_golden_model_1.IRAM[12] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  nor (_05908_, _05907_, _05906_);
  nor (_05909_, \oc8051_golden_model_1.IRAM[12] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  and (_05910_, \oc8051_golden_model_1.IRAM[12] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  nor (_05911_, _05910_, _05909_);
  nor (_05912_, _05911_, _05908_);
  and (_05913_, _05912_, _05905_);
  and (_05914_, _05913_, _05898_);
  nor (_05915_, \oc8051_golden_model_1.IRAM[15] [0], _10960_);
  and (_05916_, \oc8051_golden_model_1.IRAM[15] [0], _10960_);
  nor (_05917_, _05916_, _05915_);
  and (_05918_, \oc8051_golden_model_1.IRAM[15] [1], _10963_);
  nor (_05919_, \oc8051_golden_model_1.IRAM[15] [1], _10963_);
  nor (_05920_, _05919_, _05918_);
  and (_05921_, _05920_, _05917_);
  nor (_05922_, \oc8051_golden_model_1.IRAM[15] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  and (_05923_, \oc8051_golden_model_1.IRAM[15] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  nor (_05924_, _05923_, _05922_);
  nor (_05925_, \oc8051_golden_model_1.IRAM[15] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  and (_05926_, \oc8051_golden_model_1.IRAM[15] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  nor (_05927_, _05926_, _05925_);
  nor (_05928_, _05927_, _05924_);
  and (_05929_, _05928_, _05921_);
  and (_05930_, \oc8051_golden_model_1.IRAM[14] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  nor (_05931_, \oc8051_golden_model_1.IRAM[14] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  or (_05932_, _05931_, _05930_);
  and (_05933_, \oc8051_golden_model_1.IRAM[14] [2], _10944_);
  nor (_05934_, \oc8051_golden_model_1.IRAM[14] [2], _10944_);
  nor (_05935_, _05934_, _05933_);
  and (_05936_, _05935_, _05932_);
  nor (_05937_, \oc8051_golden_model_1.IRAM[14] [7], _10595_);
  and (_05938_, \oc8051_golden_model_1.IRAM[14] [7], _10595_);
  nor (_05939_, _05938_, _05937_);
  nand (_05940_, \oc8051_golden_model_1.IRAM[14] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  or (_05941_, \oc8051_golden_model_1.IRAM[14] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  and (_05942_, _05941_, _05940_);
  not (_05943_, _05942_);
  and (_05944_, _05943_, _05939_);
  and (_05945_, _05944_, _05936_);
  and (_05946_, _05945_, _05929_);
  and (_05947_, _05946_, _05914_);
  nor (_05948_, \oc8051_golden_model_1.IRAM[9] [5], _10844_);
  and (_05949_, \oc8051_golden_model_1.IRAM[9] [5], _10844_);
  nor (_05950_, _05949_, _05948_);
  nor (_05951_, \oc8051_golden_model_1.IRAM[9] [4], _10841_);
  and (_05952_, \oc8051_golden_model_1.IRAM[9] [4], _10841_);
  nor (_05953_, _05952_, _05951_);
  and (_05954_, _05953_, _05950_);
  nor (_05955_, \oc8051_golden_model_1.IRAM[9] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  and (_05956_, \oc8051_golden_model_1.IRAM[9] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  nor (_05957_, _05956_, _05955_);
  nor (_05958_, \oc8051_golden_model_1.IRAM[9] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  and (_05959_, \oc8051_golden_model_1.IRAM[9] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  nor (_05960_, _05959_, _05958_);
  nor (_05961_, _05960_, _05957_);
  and (_05962_, _05961_, _05954_);
  nor (_05963_, \oc8051_golden_model_1.IRAM[8] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  and (_05964_, \oc8051_golden_model_1.IRAM[8] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  nor (_05965_, _05964_, _05963_);
  nor (_05966_, \oc8051_golden_model_1.IRAM[8] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  and (_05967_, \oc8051_golden_model_1.IRAM[8] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  nor (_05968_, _05967_, _05966_);
  nor (_05969_, _05968_, _05965_);
  nor (_05970_, \oc8051_golden_model_1.IRAM[8] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  and (_05971_, \oc8051_golden_model_1.IRAM[8] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  nor (_05972_, _05971_, _05970_);
  nor (_05973_, \oc8051_golden_model_1.IRAM[8] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  and (_05974_, \oc8051_golden_model_1.IRAM[8] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  nor (_05975_, _05974_, _05973_);
  nor (_05976_, _05975_, _05972_);
  and (_05977_, _05976_, _05969_);
  and (_05978_, _05977_, _05962_);
  and (_05979_, \oc8051_golden_model_1.IRAM[11] [2], _10880_);
  nor (_05980_, \oc8051_golden_model_1.IRAM[11] [2], _10880_);
  nor (_05981_, _05980_, _05979_);
  nand (_05982_, \oc8051_golden_model_1.IRAM[11] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  or (_05983_, \oc8051_golden_model_1.IRAM[11] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  and (_05984_, _05983_, _05982_);
  not (_05985_, _05984_);
  and (_05986_, _05985_, _05981_);
  nor (_05987_, \oc8051_golden_model_1.IRAM[11] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  and (_05988_, \oc8051_golden_model_1.IRAM[11] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  nor (_05989_, _05988_, _05987_);
  not (_05990_, _05989_);
  nor (_05991_, \oc8051_golden_model_1.IRAM[11] [7], _10893_);
  and (_05992_, \oc8051_golden_model_1.IRAM[11] [7], _10893_);
  nor (_05993_, _05992_, _05991_);
  and (_05994_, _05993_, _05990_);
  and (_05995_, _05994_, _05986_);
  nor (_05996_, \oc8051_golden_model_1.IRAM[10] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  and (_05997_, \oc8051_golden_model_1.IRAM[10] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  nor (_05998_, _05997_, _05996_);
  nor (_05999_, \oc8051_golden_model_1.IRAM[10] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  and (_06000_, \oc8051_golden_model_1.IRAM[10] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  nor (_06001_, _06000_, _05999_);
  nor (_06002_, _06001_, _05998_);
  and (_06003_, \oc8051_golden_model_1.IRAM[10] [4], _10863_);
  nor (_06004_, \oc8051_golden_model_1.IRAM[10] [4], _10863_);
  nor (_06005_, _06004_, _06003_);
  nor (_06006_, \oc8051_golden_model_1.IRAM[10] [5], _10866_);
  and (_06007_, \oc8051_golden_model_1.IRAM[10] [5], _10866_);
  nor (_06008_, _06007_, _06006_);
  and (_06009_, _06008_, _06005_);
  and (_06010_, _06009_, _06002_);
  and (_06011_, _06010_, _05995_);
  and (_06012_, _06011_, _05978_);
  and (_06013_, _06012_, _05947_);
  and (_06014_, _06013_, _05882_);
  nor (_06015_, \oc8051_golden_model_1.IRAM[5] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  and (_06016_, \oc8051_golden_model_1.IRAM[5] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  nor (_06017_, _06016_, _06015_);
  nand (_06018_, \oc8051_golden_model_1.IRAM[5] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  or (_06019_, \oc8051_golden_model_1.IRAM[5] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  and (_06020_, _06019_, _06018_);
  nor (_06021_, _06020_, _06017_);
  nor (_06022_, \oc8051_golden_model_1.IRAM[5] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  and (_06023_, \oc8051_golden_model_1.IRAM[5] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  nor (_06024_, _06023_, _06022_);
  nand (_06025_, \oc8051_golden_model_1.IRAM[5] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  or (_06026_, \oc8051_golden_model_1.IRAM[5] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  and (_06027_, _06026_, _06025_);
  nor (_06028_, _06027_, _06024_);
  and (_06029_, _06028_, _06021_);
  and (_06030_, _03611_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  and (_06031_, \oc8051_golden_model_1.IRAM[4] [0], _10722_);
  nor (_06032_, _06031_, _06030_);
  nor (_06033_, \oc8051_golden_model_1.IRAM[4] [1], _10725_);
  and (_06034_, \oc8051_golden_model_1.IRAM[4] [1], _10725_);
  nor (_06035_, _06034_, _06033_);
  and (_06036_, _06035_, _06032_);
  nor (_06037_, \oc8051_golden_model_1.IRAM[4] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  and (_06038_, \oc8051_golden_model_1.IRAM[4] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  nor (_06039_, _06038_, _06037_);
  nor (_06040_, \oc8051_golden_model_1.IRAM[4] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  and (_06041_, \oc8051_golden_model_1.IRAM[4] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  nor (_06042_, _06041_, _06040_);
  nor (_06043_, _06042_, _06039_);
  and (_06044_, _06043_, _06036_);
  and (_06045_, _06044_, _06029_);
  nor (_06046_, \oc8051_golden_model_1.IRAM[7] [1], _10791_);
  and (_06047_, \oc8051_golden_model_1.IRAM[7] [1], _10791_);
  nor (_06048_, _06047_, _06046_);
  and (_06049_, _03617_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  and (_06050_, \oc8051_golden_model_1.IRAM[7] [0], _10788_);
  nor (_06051_, _06050_, _06049_);
  and (_06052_, _06051_, _06048_);
  nor (_06053_, \oc8051_golden_model_1.IRAM[7] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  and (_06054_, \oc8051_golden_model_1.IRAM[7] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  nor (_06055_, _06054_, _06053_);
  nor (_06056_, \oc8051_golden_model_1.IRAM[7] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  and (_06057_, \oc8051_golden_model_1.IRAM[7] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  nor (_06058_, _06057_, _06056_);
  nor (_06059_, _06058_, _06055_);
  and (_06060_, _06059_, _06052_);
  and (_06061_, \oc8051_golden_model_1.IRAM[6] [2], _10770_);
  and (_06062_, _03709_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  nor (_06063_, _06062_, _06061_);
  and (_06064_, \oc8051_golden_model_1.IRAM[6] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  nor (_06065_, \oc8051_golden_model_1.IRAM[6] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or (_06066_, _06065_, _06064_);
  and (_06067_, _06066_, _06063_);
  nor (_06068_, \oc8051_golden_model_1.IRAM[6] [7], _10784_);
  and (_06069_, \oc8051_golden_model_1.IRAM[6] [7], _10784_);
  nor (_06070_, _06069_, _06068_);
  nand (_06071_, \oc8051_golden_model_1.IRAM[6] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  or (_06072_, \oc8051_golden_model_1.IRAM[6] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  and (_06073_, _06072_, _06071_);
  not (_06074_, _06073_);
  and (_06075_, _06074_, _06070_);
  and (_06076_, _06075_, _06067_);
  and (_06077_, _06076_, _06060_);
  and (_06078_, _06077_, _06045_);
  nor (_06079_, \oc8051_golden_model_1.IRAM[1] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  and (_06080_, \oc8051_golden_model_1.IRAM[1] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  nor (_06081_, _06080_, _06079_);
  nor (_06082_, \oc8051_golden_model_1.IRAM[1] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  and (_06083_, \oc8051_golden_model_1.IRAM[1] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  nor (_06084_, _06083_, _06082_);
  nor (_06085_, _06084_, _06081_);
  nor (_06086_, \oc8051_golden_model_1.IRAM[1] [4], _10663_);
  and (_06087_, \oc8051_golden_model_1.IRAM[1] [4], _10663_);
  nor (_06088_, _06087_, _06086_);
  nor (_06089_, \oc8051_golden_model_1.IRAM[1] [5], _10666_);
  and (_06090_, \oc8051_golden_model_1.IRAM[1] [5], _10666_);
  nor (_06091_, _06090_, _06089_);
  and (_06092_, _06091_, _06088_);
  and (_06093_, _06092_, _06085_);
  nor (_06094_, \oc8051_golden_model_1.IRAM[0] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  and (_06095_, \oc8051_golden_model_1.IRAM[0] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  nor (_06096_, _06095_, _06094_);
  nand (_06097_, \oc8051_golden_model_1.IRAM[0] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  or (_06098_, \oc8051_golden_model_1.IRAM[0] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  and (_06099_, _06098_, _06097_);
  nor (_06100_, _06099_, _06096_);
  nor (_06101_, \oc8051_golden_model_1.IRAM[0] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  and (_06102_, \oc8051_golden_model_1.IRAM[0] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  nor (_06103_, _06102_, _06101_);
  nand (_06104_, \oc8051_golden_model_1.IRAM[0] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  or (_06105_, \oc8051_golden_model_1.IRAM[0] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  and (_06106_, _06105_, _06104_);
  nor (_06107_, _06106_, _06103_);
  and (_06108_, _06107_, _06100_);
  and (_06109_, _06108_, _06093_);
  and (_06110_, \oc8051_golden_model_1.IRAM[3] [2], _10704_);
  and (_06111_, _03723_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  nor (_06112_, _06111_, _06110_);
  nand (_06113_, \oc8051_golden_model_1.IRAM[3] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  or (_06114_, \oc8051_golden_model_1.IRAM[3] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  and (_06115_, _06114_, _06113_);
  not (_06116_, _06115_);
  and (_06117_, _06116_, _06112_);
  nor (_06118_, \oc8051_golden_model_1.IRAM[3] [7], _10558_);
  and (_06119_, \oc8051_golden_model_1.IRAM[3] [7], _10558_);
  nor (_06120_, _06119_, _06118_);
  nand (_06121_, \oc8051_golden_model_1.IRAM[3] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  or (_06122_, \oc8051_golden_model_1.IRAM[3] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  and (_06123_, _06122_, _06121_);
  not (_06124_, _06123_);
  and (_06125_, _06124_, _06120_);
  and (_06126_, _06125_, _06117_);
  nor (_06127_, \oc8051_golden_model_1.IRAM[2] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  and (_06128_, \oc8051_golden_model_1.IRAM[2] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  nor (_06129_, _06128_, _06127_);
  nor (_06130_, \oc8051_golden_model_1.IRAM[2] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  and (_06131_, \oc8051_golden_model_1.IRAM[2] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  nor (_06132_, _06131_, _06130_);
  nor (_06133_, _06132_, _06129_);
  nor (_06134_, \oc8051_golden_model_1.IRAM[2] [5], _10689_);
  and (_06135_, \oc8051_golden_model_1.IRAM[2] [5], _10689_);
  nor (_06136_, _06135_, _06134_);
  nor (_06137_, \oc8051_golden_model_1.IRAM[2] [4], _10686_);
  and (_06138_, \oc8051_golden_model_1.IRAM[2] [4], _10686_);
  nor (_06139_, _06138_, _06137_);
  and (_06140_, _06139_, _06136_);
  and (_06141_, _06140_, _06133_);
  and (_06142_, _06141_, _06126_);
  and (_06143_, _06142_, _06109_);
  and (_06144_, _06143_, _06078_);
  nor (_06145_, \oc8051_golden_model_1.IRAM[13] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  and (_06146_, \oc8051_golden_model_1.IRAM[13] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  nor (_06147_, _06146_, _06145_);
  nor (_06148_, \oc8051_golden_model_1.IRAM[13] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  and (_06149_, \oc8051_golden_model_1.IRAM[13] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  nor (_06150_, _06149_, _06148_);
  nor (_06151_, _06150_, _06147_);
  and (_06152_, \oc8051_golden_model_1.IRAM[13] [5], _10930_);
  nor (_06153_, \oc8051_golden_model_1.IRAM[13] [5], _10930_);
  nor (_06154_, _06153_, _06152_);
  and (_06155_, \oc8051_golden_model_1.IRAM[13] [4], _10927_);
  nor (_06156_, \oc8051_golden_model_1.IRAM[13] [4], _10927_);
  nor (_06157_, _06156_, _06155_);
  and (_06158_, _06157_, _06154_);
  and (_06159_, _06158_, _06151_);
  nor (_06160_, \oc8051_golden_model_1.IRAM[12] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  and (_06161_, \oc8051_golden_model_1.IRAM[12] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  nor (_06162_, _06161_, _06160_);
  not (_06163_, _06162_);
  and (_06164_, \oc8051_golden_model_1.IRAM[12] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  nor (_06165_, \oc8051_golden_model_1.IRAM[12] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  or (_06166_, _06165_, _06164_);
  and (_06167_, _06166_, _06163_);
  nor (_06168_, \oc8051_golden_model_1.IRAM[12] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  and (_06169_, \oc8051_golden_model_1.IRAM[12] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  nor (_06170_, _06169_, _06168_);
  nand (_06171_, \oc8051_golden_model_1.IRAM[12] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  or (_06172_, \oc8051_golden_model_1.IRAM[12] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  and (_06173_, _06172_, _06171_);
  nor (_06174_, _06173_, _06170_);
  and (_06175_, _06174_, _06167_);
  and (_06176_, _06175_, _06159_);
  nor (_06177_, \oc8051_golden_model_1.IRAM[15] [2], _10966_);
  and (_06178_, \oc8051_golden_model_1.IRAM[15] [2], _10966_);
  nor (_06179_, _06178_, _06177_);
  nand (_06180_, \oc8051_golden_model_1.IRAM[15] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  or (_06181_, \oc8051_golden_model_1.IRAM[15] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  and (_06182_, _06181_, _06180_);
  not (_06183_, _06182_);
  and (_06184_, _06183_, _06179_);
  nor (_06185_, \oc8051_golden_model_1.IRAM[15] [7], _10617_);
  and (_06186_, \oc8051_golden_model_1.IRAM[15] [7], _10617_);
  nor (_06187_, _06186_, _06185_);
  nand (_06188_, \oc8051_golden_model_1.IRAM[15] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  or (_06189_, \oc8051_golden_model_1.IRAM[15] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  and (_06190_, _06189_, _06188_);
  not (_06191_, _06190_);
  and (_06192_, _06191_, _06187_);
  and (_06193_, _06192_, _06184_);
  nor (_06194_, \oc8051_golden_model_1.IRAM[14] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  and (_06195_, \oc8051_golden_model_1.IRAM[14] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  nor (_06196_, _06195_, _06194_);
  nor (_06197_, \oc8051_golden_model_1.IRAM[14] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  and (_06198_, \oc8051_golden_model_1.IRAM[14] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  nor (_06199_, _06198_, _06197_);
  nor (_06200_, _06199_, _06196_);
  and (_06201_, \oc8051_golden_model_1.IRAM[14] [5], _10952_);
  nor (_06202_, \oc8051_golden_model_1.IRAM[14] [5], _10952_);
  nor (_06203_, _06202_, _06201_);
  nor (_06204_, \oc8051_golden_model_1.IRAM[14] [4], _10949_);
  and (_06205_, \oc8051_golden_model_1.IRAM[14] [4], _10949_);
  nor (_06206_, _06205_, _06204_);
  and (_06207_, _06206_, _06203_);
  and (_06208_, _06207_, _06200_);
  and (_06209_, _06208_, _06193_);
  and (_06210_, _06209_, _06176_);
  nor (_06211_, \oc8051_golden_model_1.IRAM[9] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  and (_06212_, \oc8051_golden_model_1.IRAM[9] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  nor (_06213_, _06212_, _06211_);
  nor (_06214_, \oc8051_golden_model_1.IRAM[9] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  and (_06215_, \oc8051_golden_model_1.IRAM[9] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  nor (_06216_, _06215_, _06214_);
  nor (_06217_, _06216_, _06213_);
  nor (_06218_, \oc8051_golden_model_1.IRAM[9] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  and (_06219_, \oc8051_golden_model_1.IRAM[9] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  nor (_06220_, _06219_, _06218_);
  nor (_06221_, \oc8051_golden_model_1.IRAM[9] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  and (_06222_, \oc8051_golden_model_1.IRAM[9] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  nor (_06223_, _06222_, _06221_);
  nor (_06224_, _06223_, _06220_);
  and (_06225_, _06224_, _06217_);
  nor (_06226_, \oc8051_golden_model_1.IRAM[8] [0], _10812_);
  and (_06227_, \oc8051_golden_model_1.IRAM[8] [0], _10812_);
  nor (_06228_, _06227_, _06226_);
  nor (_06229_, \oc8051_golden_model_1.IRAM[8] [1], _10815_);
  and (_06230_, \oc8051_golden_model_1.IRAM[8] [1], _10815_);
  nor (_06231_, _06230_, _06229_);
  and (_06232_, _06231_, _06228_);
  nor (_06233_, \oc8051_golden_model_1.IRAM[8] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  and (_06234_, \oc8051_golden_model_1.IRAM[8] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  nor (_06235_, _06234_, _06233_);
  nor (_06236_, \oc8051_golden_model_1.IRAM[8] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  and (_06237_, \oc8051_golden_model_1.IRAM[8] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  nor (_06238_, _06237_, _06236_);
  nor (_06239_, _06238_, _06235_);
  and (_06240_, _06239_, _06232_);
  and (_06241_, _06240_, _06225_);
  nor (_06242_, \oc8051_golden_model_1.IRAM[11] [0], _10874_);
  and (_06243_, \oc8051_golden_model_1.IRAM[11] [0], _10874_);
  nor (_06244_, _06243_, _06242_);
  and (_06245_, \oc8051_golden_model_1.IRAM[11] [1], _10877_);
  nor (_06246_, \oc8051_golden_model_1.IRAM[11] [1], _10877_);
  nor (_06247_, _06246_, _06245_);
  and (_06248_, _06247_, _06244_);
  nor (_06249_, \oc8051_golden_model_1.IRAM[11] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  and (_06250_, \oc8051_golden_model_1.IRAM[11] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  nor (_06251_, _06250_, _06249_);
  nor (_06252_, \oc8051_golden_model_1.IRAM[11] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  and (_06253_, \oc8051_golden_model_1.IRAM[11] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  nor (_06254_, _06253_, _06252_);
  nor (_06255_, _06254_, _06251_);
  and (_06256_, _06255_, _06248_);
  and (_06257_, \oc8051_golden_model_1.IRAM[10] [2], _10857_);
  nor (_06258_, \oc8051_golden_model_1.IRAM[10] [2], _10857_);
  nor (_06259_, _06258_, _06257_);
  nand (_06260_, \oc8051_golden_model_1.IRAM[10] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  or (_06261_, \oc8051_golden_model_1.IRAM[10] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  and (_06262_, _06261_, _06260_);
  not (_06263_, _06262_);
  and (_06264_, _06263_, _06259_);
  nor (_06265_, \oc8051_golden_model_1.IRAM[10] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  and (_06266_, \oc8051_golden_model_1.IRAM[10] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  nor (_06267_, _06266_, _06265_);
  not (_06268_, _06267_);
  nor (_06269_, \oc8051_golden_model_1.IRAM[10] [7], _10584_);
  and (_06270_, \oc8051_golden_model_1.IRAM[10] [7], _10584_);
  nor (_06271_, _06270_, _06269_);
  and (_06272_, _06271_, _06268_);
  and (_06273_, _06272_, _06264_);
  and (_06274_, _06273_, _06256_);
  and (_06275_, _06274_, _06241_);
  and (_06276_, _06275_, _06210_);
  and (_06277_, _06276_, _06144_);
  and (_06278_, _06277_, _06014_);
  nor (_06279_, \oc8051_golden_model_1.ACC [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_06280_, \oc8051_golden_model_1.ACC [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor (_06281_, _06280_, _06279_);
  nor (_06282_, \oc8051_golden_model_1.ACC [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and (_06283_, \oc8051_golden_model_1.ACC [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_06284_, _06283_, _06282_);
  nor (_06285_, _06284_, _06281_);
  nor (_06286_, \oc8051_golden_model_1.ACC [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_06287_, \oc8051_golden_model_1.ACC [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor (_06288_, _06287_, _06286_);
  nor (_06289_, \oc8051_golden_model_1.ACC [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_06290_, \oc8051_golden_model_1.ACC [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_06291_, _06290_, _06289_);
  nor (_06292_, _06291_, _06288_);
  and (_06293_, _06292_, _06285_);
  and (_06294_, _03758_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_06295_, \oc8051_golden_model_1.ACC [2], _06976_);
  nor (_06296_, _06295_, _06294_);
  and (_06297_, \oc8051_golden_model_1.ACC [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor (_06298_, \oc8051_golden_model_1.ACC [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_06299_, _06298_, _06297_);
  and (_06300_, _06299_, _06296_);
  and (_06301_, _03158_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_06302_, \oc8051_golden_model_1.ACC [7], _06960_);
  nor (_06304_, _06302_, _06301_);
  and (_06305_, \oc8051_golden_model_1.ACC [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor (_06306_, \oc8051_golden_model_1.ACC [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_06307_, _06306_, _06305_);
  and (_06308_, _06307_, _06304_);
  and (_06309_, _06308_, _06300_);
  and (_06310_, _06309_, _06293_);
  nor (_06311_, \oc8051_golden_model_1.B [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_06312_, \oc8051_golden_model_1.B [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  nor (_06313_, _06312_, _06311_);
  nor (_06314_, \oc8051_golden_model_1.B [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  and (_06315_, \oc8051_golden_model_1.B [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nor (_06316_, _06315_, _06314_);
  nor (_06317_, _06316_, _06313_);
  nor (_06318_, \oc8051_golden_model_1.B [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_06319_, \oc8051_golden_model_1.B [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nor (_06320_, _06319_, _06318_);
  nor (_06321_, \oc8051_golden_model_1.B [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_06322_, \oc8051_golden_model_1.B [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nor (_06323_, _06322_, _06321_);
  nor (_06324_, _06323_, _06320_);
  and (_06325_, _06324_, _06317_);
  nor (_06326_, \oc8051_golden_model_1.B [2], _08226_);
  and (_06327_, \oc8051_golden_model_1.B [2], _08226_);
  nor (_06328_, _06327_, _06326_);
  and (_06329_, \oc8051_golden_model_1.B [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nor (_06330_, \oc8051_golden_model_1.B [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  or (_06331_, _06330_, _06329_);
  and (_06332_, _06331_, _06328_);
  nor (_06333_, \oc8051_golden_model_1.B [7], _08009_);
  and (_06334_, \oc8051_golden_model_1.B [7], _08009_);
  nor (_06335_, _06334_, _06333_);
  and (_06336_, \oc8051_golden_model_1.B [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  nor (_06337_, \oc8051_golden_model_1.B [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  or (_06338_, _06337_, _06336_);
  and (_06339_, _06338_, _06335_);
  and (_06340_, _06339_, _06332_);
  and (_06341_, _06340_, _06325_);
  and (_06342_, _06341_, _06310_);
  nor (_06343_, \oc8051_golden_model_1.DPH [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  and (_06344_, \oc8051_golden_model_1.DPH [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  nor (_06345_, _06344_, _06343_);
  nor (_06346_, \oc8051_golden_model_1.DPH [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and (_06347_, \oc8051_golden_model_1.DPH [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  nor (_06348_, _06347_, _06346_);
  nor (_06349_, _06348_, _06345_);
  nor (_06350_, \oc8051_golden_model_1.DPH [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  and (_06351_, \oc8051_golden_model_1.DPH [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  nor (_06352_, _06351_, _06350_);
  nor (_06353_, \oc8051_golden_model_1.DPH [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  and (_06354_, \oc8051_golden_model_1.DPH [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  nor (_06355_, _06354_, _06353_);
  nor (_06356_, _06355_, _06352_);
  and (_06357_, _06356_, _06349_);
  not (_06358_, \oc8051_golden_model_1.DPH [2]);
  and (_06359_, _06358_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  nor (_06360_, _06358_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  nor (_06361_, _06360_, _06359_);
  and (_06362_, \oc8051_golden_model_1.DPH [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  nor (_06363_, \oc8051_golden_model_1.DPH [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_06364_, _06363_, _06362_);
  and (_06365_, _06364_, _06361_);
  not (_06366_, \oc8051_golden_model_1.DPH [7]);
  and (_06367_, _06366_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  nor (_06368_, _06366_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  nor (_06369_, _06368_, _06367_);
  and (_06370_, \oc8051_golden_model_1.DPH [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  nor (_06371_, \oc8051_golden_model_1.DPH [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_06372_, _06371_, _06370_);
  and (_06373_, _06372_, _06369_);
  and (_06374_, _06373_, _06365_);
  and (_06375_, _06374_, _06357_);
  nor (_06376_, \oc8051_golden_model_1.DPL [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_06377_, \oc8051_golden_model_1.DPL [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  nor (_06378_, _06377_, _06376_);
  nor (_06379_, \oc8051_golden_model_1.DPL [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_06380_, \oc8051_golden_model_1.DPL [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  nor (_06381_, _06380_, _06379_);
  nor (_06382_, _06381_, _06378_);
  nor (_06383_, \oc8051_golden_model_1.DPL [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_06384_, \oc8051_golden_model_1.DPL [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  nor (_06385_, _06384_, _06383_);
  nor (_06386_, \oc8051_golden_model_1.DPL [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_06387_, \oc8051_golden_model_1.DPL [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  nor (_06388_, _06387_, _06386_);
  nor (_06389_, _06388_, _06385_);
  and (_06390_, _06389_, _06382_);
  nor (_06391_, \oc8051_golden_model_1.DPL [2], _09363_);
  and (_06392_, \oc8051_golden_model_1.DPL [2], _09363_);
  nor (_06393_, _06392_, _06391_);
  and (_06394_, \oc8051_golden_model_1.DPL [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  nor (_06395_, \oc8051_golden_model_1.DPL [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  or (_06396_, _06395_, _06394_);
  and (_06397_, _06396_, _06393_);
  nor (_06398_, \oc8051_golden_model_1.DPL [7], _09137_);
  and (_06399_, \oc8051_golden_model_1.DPL [7], _09137_);
  nor (_06400_, _06399_, _06398_);
  and (_06401_, \oc8051_golden_model_1.DPL [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  nor (_06402_, \oc8051_golden_model_1.DPL [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  or (_06403_, _06402_, _06401_);
  and (_06404_, _06403_, _06400_);
  and (_06405_, _06404_, _06397_);
  and (_06406_, _06405_, _06390_);
  and (_06407_, _06406_, _06375_);
  and (_06408_, _06407_, _06342_);
  nor (_06409_, \oc8051_golden_model_1.P3 [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_06410_, \oc8051_golden_model_1.P3 [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  nor (_06411_, _06410_, _06409_);
  nor (_06412_, \oc8051_golden_model_1.P3 [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and (_06413_, \oc8051_golden_model_1.P3 [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  nor (_06414_, _06413_, _06412_);
  nor (_06415_, _06414_, _06411_);
  nor (_06416_, \oc8051_golden_model_1.P3 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_06417_, \oc8051_golden_model_1.P3 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  nor (_06418_, _06417_, _06416_);
  nor (_06419_, \oc8051_golden_model_1.P3 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_06420_, \oc8051_golden_model_1.P3 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  nor (_06421_, _06420_, _06419_);
  nor (_06422_, _06421_, _06418_);
  and (_06423_, _06422_, _06415_);
  and (_06424_, _03785_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_06425_, \oc8051_golden_model_1.P3 [2], _09960_);
  nor (_06426_, _06425_, _06424_);
  and (_06427_, \oc8051_golden_model_1.P3 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  nor (_06428_, \oc8051_golden_model_1.P3 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_06429_, _06428_, _06427_);
  and (_06430_, _06429_, _06426_);
  and (_06431_, _03926_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and (_06432_, \oc8051_golden_model_1.P3 [7], _09655_);
  nor (_06433_, _06432_, _06431_);
  and (_06434_, \oc8051_golden_model_1.P3 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  nor (_06435_, \oc8051_golden_model_1.P3 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or (_06436_, _06435_, _06434_);
  and (_06437_, _06436_, _06433_);
  and (_06438_, _06437_, _06430_);
  and (_06439_, _06438_, _06423_);
  nor (_06440_, \oc8051_golden_model_1.P1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_06441_, \oc8051_golden_model_1.P1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  nor (_06442_, _06441_, _06440_);
  nor (_06443_, \oc8051_golden_model_1.P1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and (_06444_, \oc8051_golden_model_1.P1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  nor (_06445_, _06444_, _06443_);
  nor (_06446_, _06445_, _06442_);
  nor (_06447_, \oc8051_golden_model_1.P1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_06448_, \oc8051_golden_model_1.P1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  nor (_06449_, _06448_, _06447_);
  nor (_06450_, \oc8051_golden_model_1.P1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_06451_, \oc8051_golden_model_1.P1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  nor (_06452_, _06451_, _06450_);
  nor (_06453_, _06452_, _06449_);
  and (_06454_, _06453_, _06446_);
  nor (_06455_, \oc8051_golden_model_1.P1 [2], _09792_);
  and (_06456_, \oc8051_golden_model_1.P1 [2], _09792_);
  nor (_06457_, _06456_, _06455_);
  and (_06458_, \oc8051_golden_model_1.P1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  nor (_06459_, \oc8051_golden_model_1.P1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or (_06460_, _06459_, _06458_);
  and (_06461_, _06460_, _06457_);
  and (_06462_, _03948_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_06463_, \oc8051_golden_model_1.P1 [7], _09627_);
  nor (_06464_, _06463_, _06462_);
  and (_06465_, \oc8051_golden_model_1.P1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  nor (_06466_, \oc8051_golden_model_1.P1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  or (_06467_, _06466_, _06465_);
  and (_06468_, _06467_, _06464_);
  and (_06469_, _06468_, _06461_);
  and (_06470_, _06469_, _06454_);
  and (_06471_, _06470_, _06439_);
  nor (_06472_, \oc8051_golden_model_1.P2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_06473_, \oc8051_golden_model_1.P2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  nor (_06474_, _06473_, _06472_);
  nor (_06475_, \oc8051_golden_model_1.P2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and (_06476_, \oc8051_golden_model_1.P2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  nor (_06477_, _06476_, _06475_);
  nor (_06478_, _06477_, _06474_);
  nor (_06479_, \oc8051_golden_model_1.P2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_06480_, \oc8051_golden_model_1.P2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  nor (_06481_, _06480_, _06479_);
  nor (_06482_, \oc8051_golden_model_1.P2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_06483_, \oc8051_golden_model_1.P2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  nor (_06484_, _06483_, _06482_);
  nor (_06485_, _06484_, _06481_);
  and (_06486_, _06485_, _06478_);
  nor (_06487_, \oc8051_golden_model_1.P2 [2], _09877_);
  and (_06488_, \oc8051_golden_model_1.P2 [2], _09877_);
  nor (_06489_, _06488_, _06487_);
  and (_06490_, \oc8051_golden_model_1.P2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  nor (_06491_, \oc8051_golden_model_1.P2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_06492_, _06491_, _06490_);
  and (_06493_, _06492_, _06489_);
  and (_06494_, _03937_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_06495_, \oc8051_golden_model_1.P2 [7], _09647_);
  nor (_06496_, _06495_, _06494_);
  and (_06497_, \oc8051_golden_model_1.P2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  nor (_06498_, \oc8051_golden_model_1.P2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or (_06499_, _06498_, _06497_);
  and (_06500_, _06499_, _06496_);
  and (_06501_, _06500_, _06493_);
  and (_06502_, _06501_, _06486_);
  nor (_06503_, \oc8051_golden_model_1.P0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_06504_, \oc8051_golden_model_1.P0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  nor (_06505_, _06504_, _06503_);
  nor (_06506_, \oc8051_golden_model_1.P0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  and (_06507_, \oc8051_golden_model_1.P0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  nor (_06508_, _06507_, _06506_);
  nor (_06509_, _06508_, _06505_);
  nor (_06510_, \oc8051_golden_model_1.P0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_06511_, \oc8051_golden_model_1.P0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  nor (_06512_, _06511_, _06510_);
  nor (_06513_, \oc8051_golden_model_1.P0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_06514_, \oc8051_golden_model_1.P0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  nor (_06515_, _06514_, _06513_);
  nor (_06516_, _06515_, _06512_);
  and (_06517_, _06516_, _06509_);
  nor (_06518_, \oc8051_golden_model_1.P0 [2], _09707_);
  and (_06519_, \oc8051_golden_model_1.P0 [2], _09707_);
  nor (_06520_, _06519_, _06518_);
  and (_06521_, \oc8051_golden_model_1.P0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  nor (_06522_, \oc8051_golden_model_1.P0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or (_06523_, _06522_, _06521_);
  and (_06524_, _06523_, _06520_);
  and (_06525_, _03960_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_06526_, \oc8051_golden_model_1.P0 [7], _09617_);
  nor (_06527_, _06526_, _06525_);
  and (_06528_, \oc8051_golden_model_1.P0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  nor (_06529_, \oc8051_golden_model_1.P0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  or (_06530_, _06529_, _06528_);
  and (_06531_, _06530_, _06527_);
  and (_06532_, _06531_, _06524_);
  and (_06533_, _06532_, _06517_);
  and (_06534_, _06533_, _06502_);
  and (_06535_, _06534_, _06471_);
  and (_06536_, _06535_, _06408_);
  and (_06537_, _06536_, _06278_);
  or (_06538_, _09007_, \oc8051_golden_model_1.SP [0]);
  nand (_06539_, _09007_, \oc8051_golden_model_1.SP [0]);
  and (_06540_, _06539_, _06538_);
  and (_06541_, _06540_, _06537_);
  nand (_06542_, _09013_, \oc8051_golden_model_1.SP [1]);
  or (_06543_, _09013_, \oc8051_golden_model_1.SP [1]);
  and (_06544_, _06543_, _06542_);
  and (_06545_, _06544_, _06541_);
  nand (_06546_, _09019_, \oc8051_golden_model_1.SP [2]);
  or (_06547_, _09019_, \oc8051_golden_model_1.SP [2]);
  and (_06548_, _06547_, _06546_);
  and (_06549_, _06548_, _06545_);
  and (_06550_, _06549_, _05749_);
  and (_06551_, _06550_, _05746_);
  and (_06552_, _06551_, _05743_);
  and (_06553_, _06552_, _05740_);
  and (_06554_, _06553_, _05737_);
  and (_06555_, _06554_, _05733_);
  and (_06556_, _06555_, _05705_);
  nand (_06557_, _06556_, _05704_);
  nand (_06558_, _06557_, inst_finished_r);
  and (_06559_, _06558_, eq_state_2);
  or (_00001_, _06559_, rst);
  and (_06560_, _02738_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor (_06561_, _05650_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_06562_, _05650_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor (_06563_, _06562_, _06561_);
  nor (_06564_, _02738_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  or (_06565_, _06564_, _06563_);
  nor (_06566_, _06565_, _06560_);
  nor (_06567_, _05634_, _06865_);
  and (_06568_, _05634_, _06865_);
  or (_06569_, _06568_, _06567_);
  nor (_06570_, _05578_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_06571_, _05578_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nor (_06572_, _06571_, _06570_);
  nor (_06573_, _05540_, _07171_);
  and (_06574_, _05540_, _07171_);
  nor (_06575_, _06574_, _06573_);
  nor (_06576_, _05586_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_06577_, _05586_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_06578_, _06577_, _06576_);
  or (_06579_, _06578_, _06575_);
  or (_06580_, _06579_, _06572_);
  nor (_06581_, _05626_, _07021_);
  and (_06582_, _05626_, _07021_);
  nor (_06583_, _06582_, _06581_);
  nor (_06584_, _05546_, _07119_);
  and (_06585_, _05546_, _07119_);
  nor (_06586_, _06585_, _06584_);
  nor (_06587_, _05618_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_06588_, _05618_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  nor (_06589_, _06588_, _06587_);
  not (_06590_, _06589_);
  and (_06591_, _06590_, _06586_);
  nand (_06592_, _06591_, _06583_);
  or (_06593_, _06592_, _06580_);
  nor (_06594_, _06593_, _06569_);
  and (_06595_, _05642_, _07040_);
  nor (_06596_, _05642_, _07040_);
  or (_06597_, _06596_, _06595_);
  nor (_06598_, _05562_, _07019_);
  and (_06599_, _05562_, _07019_);
  nor (_06600_, _06599_, _06598_);
  nor (_06601_, _05610_, _07121_);
  and (_06602_, _05610_, _07121_);
  nor (_06603_, _06602_, _06601_);
  nand (_06604_, _06603_, _06600_);
  nor (_06605_, _05554_, _07138_);
  and (_06606_, _05554_, _07138_);
  nor (_06607_, _06606_, _06605_);
  nor (_06608_, _05602_, _07173_);
  and (_06609_, _05602_, _07173_);
  nor (_06610_, _06609_, _06608_);
  nand (_06611_, _06610_, _06607_);
  nor (_06612_, _05570_, _06859_);
  and (_06613_, _05570_, _06859_);
  nor (_06614_, _06613_, _06612_);
  nor (_06615_, _05594_, _07094_);
  and (_06616_, _05594_, _07094_);
  nor (_06617_, _06616_, _06615_);
  nand (_06618_, _06617_, _06614_);
  or (_06619_, _06618_, _06611_);
  or (_06620_, _06619_, _06604_);
  nor (_06621_, _06620_, _06597_);
  and (_06622_, _06621_, _06594_);
  and (_06623_, _06622_, _06566_);
  nor (_06624_, _06623_, _12786_);
  nor (_06625_, _05658_, _00435_);
  and (_06626_, _05658_, _00435_);
  nor (_06627_, _06626_, _06625_);
  nor (_06628_, _05678_, _00465_);
  and (_06629_, _05678_, _00465_);
  nor (_06630_, _06629_, _06628_);
  and (_06631_, _06630_, _06627_);
  nor (_06632_, _05654_, _00429_);
  and (_06633_, _05654_, _00429_);
  nor (_06634_, _06633_, _06632_);
  nor (_06635_, _02716_, _13332_);
  and (_06636_, _02716_, _13332_);
  nor (_06637_, _06636_, _06635_);
  and (_06638_, _06637_, _06634_);
  and (_06639_, _06638_, _06631_);
  nor (_06640_, _05662_, _00440_);
  and (_06641_, _05662_, _00440_);
  nor (_06642_, _06641_, _06640_);
  nor (_06643_, _05670_, _00451_);
  and (_06644_, _05670_, _00451_);
  nor (_06645_, _06644_, _06643_);
  and (_06646_, _06645_, _06642_);
  nor (_06647_, _05666_, _00445_);
  and (_06648_, _05666_, _00445_);
  nor (_06649_, _06648_, _06647_);
  nor (_06650_, _05674_, _00458_);
  and (_06651_, _05674_, _00458_);
  nor (_06652_, _06651_, _06650_);
  and (_06653_, _06652_, _06649_);
  and (_06654_, _06653_, _06646_);
  and (_06655_, _06654_, _06639_);
  nor (_06656_, _05514_, _00544_);
  and (_06657_, _05514_, _00544_);
  nor (_06658_, _06657_, _06656_);
  nor (_06659_, _05522_, _00555_);
  and (_06660_, _05522_, _00555_);
  or (_06661_, _06660_, _06659_);
  not (_06662_, _06661_);
  and (_06663_, _06662_, _06658_);
  nor (_06664_, _02742_, _13342_);
  and (_06665_, _02742_, _13342_);
  nor (_06666_, _06665_, _06664_);
  nor (_06667_, _05526_, _00560_);
  and (_06668_, _05526_, _00560_);
  nor (_06669_, _06668_, _06667_);
  and (_06670_, _06669_, _06666_);
  and (_06671_, _06670_, _06663_);
  nor (_06672_, _05478_, _00472_);
  and (_06673_, _05478_, _00472_);
  nor (_06674_, _06673_, _06672_);
  nor (_06675_, _05486_, _00488_);
  and (_06676_, _05486_, _00488_);
  nor (_06677_, _06676_, _06675_);
  and (_06678_, _06677_, _06674_);
  nor (_06679_, _05498_, _00515_);
  and (_06680_, _05498_, _00515_);
  nor (_06681_, _06680_, _06679_);
  nor (_06682_, _05506_, _00532_);
  and (_06683_, _05506_, _00532_);
  nor (_06684_, _06683_, _06682_);
  and (_06685_, _06684_, _06681_);
  and (_06686_, _06685_, _06678_);
  and (_06687_, _06686_, _06671_);
  nor (_06688_, _05510_, _00539_);
  and (_06689_, _05510_, _00539_);
  nor (_06690_, _06689_, _06688_);
  and (_06691_, _05518_, _00550_);
  nor (_06692_, _05518_, _00550_);
  nor (_06693_, _06692_, _06691_);
  and (_06694_, _06693_, _06690_);
  nor (_06695_, _05534_, _00570_);
  and (_06696_, _05534_, _00570_);
  nor (_06697_, _06696_, _06695_);
  and (_06698_, _05530_, _00565_);
  nor (_06699_, _05530_, _00565_);
  or (_06700_, _06699_, _06698_);
  not (_06701_, _06700_);
  and (_06702_, _06701_, _06697_);
  and (_06703_, _06702_, _06694_);
  nor (_06704_, _05490_, _00495_);
  and (_06705_, _05490_, _00495_);
  nor (_06706_, _06705_, _06704_);
  nor (_06707_, _05482_, _00481_);
  and (_06708_, _05482_, _00481_);
  or (_06709_, _06708_, _06707_);
  not (_06710_, _06709_);
  and (_06711_, _06710_, _06706_);
  nor (_06712_, _05502_, _00525_);
  and (_06713_, _05502_, _00525_);
  nor (_06714_, _06713_, _06712_);
  nor (_06715_, _05494_, _00505_);
  and (_06716_, _05494_, _00505_);
  nor (_06717_, _06716_, _06715_);
  and (_06718_, _06717_, _06714_);
  and (_06719_, _06718_, _06711_);
  and (_06720_, _06719_, _06703_);
  and (_06721_, _06720_, _06687_);
  and (_06722_, _06721_, _06655_);
  or (_06723_, _06722_, _12786_);
  nand (_06724_, _06723_, eq_state_1);
  nor (_06725_, _06724_, _06624_);
  or (_00000_, _06725_, rst);
  and (_00008_, _05733_, _13707_);
  not (_06726_, _02438_);
  or (_06727_, _06726_, _02393_);
  not (_06728_, _02667_);
  nand (_06729_, _06728_, _02621_);
  or (_06730_, _02576_, _02484_);
  and (_06731_, _06730_, _02529_);
  or (_06732_, _06731_, _06729_);
  or (_06733_, _02576_, _02529_);
  and (_06734_, _06733_, _02484_);
  or (_06735_, _02529_, _02484_);
  and (_06736_, _06735_, _02621_);
  or (_06737_, _06736_, _06728_);
  or (_06738_, _06737_, _06734_);
  and (_06739_, _06738_, _06732_);
  or (_06740_, _06739_, _02712_);
  not (_06741_, _02712_);
  or (_06742_, _02667_, _02621_);
  or (_06743_, _06742_, _06741_);
  or (_06744_, _06743_, _06733_);
  nand (_06745_, _02713_, _02529_);
  or (_06746_, _06745_, _02622_);
  and (_06747_, _06746_, _06744_);
  or (_06748_, _06747_, _02484_);
  and (_06749_, _06748_, _06740_);
  or (_06750_, _06749_, _06727_);
  and (_06751_, _06741_, _02529_);
  and (_06752_, _06751_, _02439_);
  nor (_06753_, _06730_, _06729_);
  nand (_06754_, _06753_, _06752_);
  and (_06755_, _06754_, op0_cnst);
  and (_06756_, _06755_, _06750_);
  or (_00003_, _06756_, rst);
  and (_00009_, _02758_, _13707_);
  and (_00007_[7], _00822_, _13707_);
  and (_00006_[7], _00892_, _13707_);
  and (_00005_[7], _00788_, _13707_);
  and (_00004_[7], _00963_, _13707_);
  and (_06757_, _12786_, xram_data_in_reg[7]);
  and (_06758_, _12782_, xram_data_in[7]);
  or (_06759_, _06758_, _06757_);
  and (_00010_[7], _06759_, _13707_);
  not (_06760_, _06655_);
  and (_06761_, _02758_, eq_state_1);
  and (_06762_, _06761_, _06756_);
  and (_06763_, _06762_, _06559_);
  and (_06764_, _06763_, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  and (property_invalid_xram_data_out, _06764_, _06760_);
  not (_06765_, _06721_);
  and (property_invalid_xram_addr, _06764_, _06765_);
  and (_06766_, inst_finished_r, eq_state_2);
  and (_06767_, _06766_, this_op_cnst_r);
  and (_06768_, _06767_, _06756_);
  and (_06769_, _06768_, _06725_);
  and (_06770_, _03597_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  nor (_06771_, _03597_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  or (_06772_, _06771_, _06770_);
  and (_06773_, _03760_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  and (_06774_, \oc8051_golden_model_1.PSW [2], _09434_);
  or (_06775_, _06774_, _06773_);
  or (_06776_, _06775_, _06772_);
  and (_06777_, _05388_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_06778_, \oc8051_golden_model_1.PSW [4], _09455_);
  or (_06779_, _06778_, _06777_);
  nand (_06780_, \oc8051_golden_model_1.PSW [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  or (_06781_, \oc8051_golden_model_1.PSW [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_06782_, _06781_, _06780_);
  or (_06783_, _06782_, _06779_);
  or (_06784_, _06783_, _06776_);
  and (_06785_, _03911_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  and (_06786_, \oc8051_golden_model_1.PSW [7], _09391_);
  or (_06787_, _06786_, _06785_);
  and (_06788_, _05398_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_06789_, \oc8051_golden_model_1.PSW [5], _05727_);
  or (_06790_, _06789_, _06788_);
  nand (_06791_, \oc8051_golden_model_1.PSW [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  or (_06792_, \oc8051_golden_model_1.PSW [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_06793_, _06792_, _06791_);
  or (_06794_, _06793_, _06790_);
  or (_06795_, _06794_, _06787_);
  nor (_06796_, _06795_, _06784_);
  nor (_06797_, _06796_, property_valid_psw_1_r);
  and (property_invalid_psw, _06797_, _06769_);
  not (_06798_, _06439_);
  and (property_invalid_p3, _06769_, _06798_);
  not (_06799_, _06502_);
  and (property_invalid_p2, _06769_, _06799_);
  not (_06800_, _06470_);
  and (property_invalid_p1, _06769_, _06800_);
  not (_06801_, _06533_);
  and (property_invalid_p0, _06769_, _06801_);
  not (_06802_, _06278_);
  and (property_invalid_iram, _06769_, _06802_);
  not (_06803_, _06375_);
  and (property_invalid_dph, _06769_, _06803_);
  not (_06804_, _06406_);
  and (property_invalid_dpl, _06769_, _06804_);
  not (_06805_, _06341_);
  and (property_invalid_b_reg, _06769_, _06805_);
  not (_06806_, _06310_);
  and (property_invalid_acc, _06769_, _06806_);
  and (property_invalid_pc, _06763_, _06624_);
  buf (_13759_, _13707_);
  buf (_13810_, _13707_);
  buf (_00048_, _13707_);
  buf (_00099_, _13707_);
  buf (_00149_, _13707_);
  buf (_00197_, _13707_);
  buf (_00244_, _13707_);
  buf (_00284_, _13707_);
  buf (_00324_, _13707_);
  buf (_00366_, _13707_);
  buf (_00408_, _13707_);
  buf (_00452_, _13707_);
  buf (_00499_, _13707_);
  buf (_00545_, _13707_);
  buf (_13827_, _13707_);
  buf (_13933_[7], _13911_[7]);
  buf (_13934_[7], _13912_[7]);
  buf (_13945_[7], _13911_[7]);
  buf (_13946_[7], _13912_[7]);
  buf (_13933_[0], _13911_[0]);
  buf (_13933_[1], _13911_[1]);
  buf (_13933_[2], _13911_[2]);
  buf (_13933_[3], _13911_[3]);
  buf (_13933_[4], _13911_[4]);
  buf (_13933_[5], _13911_[5]);
  buf (_13933_[6], _13911_[6]);
  buf (_13934_[0], _13912_[0]);
  buf (_13934_[1], _13912_[1]);
  buf (_13934_[2], _13912_[2]);
  buf (_13934_[3], _13912_[3]);
  buf (_13934_[4], _13912_[4]);
  buf (_13934_[5], _13912_[5]);
  buf (_13934_[6], _13912_[6]);
  buf (_13945_[0], _13911_[0]);
  buf (_13945_[1], _13911_[1]);
  buf (_13945_[2], _13911_[2]);
  buf (_13945_[3], _13911_[3]);
  buf (_13945_[4], _13911_[4]);
  buf (_13945_[5], _13911_[5]);
  buf (_13945_[6], _13911_[6]);
  buf (_13946_[0], _13912_[0]);
  buf (_13946_[1], _13912_[1]);
  buf (_13946_[2], _13912_[2]);
  buf (_13946_[3], _13912_[3]);
  buf (_13946_[4], _13912_[4]);
  buf (_13946_[5], _13912_[5]);
  buf (_13946_[6], _13912_[6]);
  buf (_13970_, _13926_);
  buf (_13965_, _13926_);
  dff (xram_data_in_reg[0], _00010_[0]);
  dff (xram_data_in_reg[1], _00010_[1]);
  dff (xram_data_in_reg[2], _00010_[2]);
  dff (xram_data_in_reg[3], _00010_[3]);
  dff (xram_data_in_reg[4], _00010_[4]);
  dff (xram_data_in_reg[5], _00010_[5]);
  dff (xram_data_in_reg[6], _00010_[6]);
  dff (xram_data_in_reg[7], _00010_[7]);
  dff (p0in_reg[0], _00004_[0]);
  dff (p0in_reg[1], _00004_[1]);
  dff (p0in_reg[2], _00004_[2]);
  dff (p0in_reg[3], _00004_[3]);
  dff (p0in_reg[4], _00004_[4]);
  dff (p0in_reg[5], _00004_[5]);
  dff (p0in_reg[6], _00004_[6]);
  dff (p0in_reg[7], _00004_[7]);
  dff (p1in_reg[0], _00005_[0]);
  dff (p1in_reg[1], _00005_[1]);
  dff (p1in_reg[2], _00005_[2]);
  dff (p1in_reg[3], _00005_[3]);
  dff (p1in_reg[4], _00005_[4]);
  dff (p1in_reg[5], _00005_[5]);
  dff (p1in_reg[6], _00005_[6]);
  dff (p1in_reg[7], _00005_[7]);
  dff (p2in_reg[0], _00006_[0]);
  dff (p2in_reg[1], _00006_[1]);
  dff (p2in_reg[2], _00006_[2]);
  dff (p2in_reg[3], _00006_[3]);
  dff (p2in_reg[4], _00006_[4]);
  dff (p2in_reg[5], _00006_[5]);
  dff (p2in_reg[6], _00006_[6]);
  dff (p2in_reg[7], _00006_[7]);
  dff (p3in_reg[0], _00007_[0]);
  dff (p3in_reg[1], _00007_[1]);
  dff (p3in_reg[2], _00007_[2]);
  dff (p3in_reg[3], _00007_[3]);
  dff (p3in_reg[4], _00007_[4]);
  dff (p3in_reg[5], _00007_[5]);
  dff (p3in_reg[6], _00007_[6]);
  dff (p3in_reg[7], _00007_[7]);
  dff (inst_finished_r, _00002_);
  dff (this_op_cnst_r, _00009_);
  dff (op0_cnst, _00003_);
  dff (property_valid_psw_1_r, _00008_);
  dff (eq_state_1, _00000_);
  dff (eq_state_2, _00001_);
  dff (\oc8051_gm_cxrom_1.cell0.data [0], _13711_);
  dff (\oc8051_gm_cxrom_1.cell0.data [1], _13715_);
  dff (\oc8051_gm_cxrom_1.cell0.data [2], _13718_);
  dff (\oc8051_gm_cxrom_1.cell0.data [3], _13722_);
  dff (\oc8051_gm_cxrom_1.cell0.data [4], _13726_);
  dff (\oc8051_gm_cxrom_1.cell0.data [5], _13730_);
  dff (\oc8051_gm_cxrom_1.cell0.data [6], _13734_);
  dff (\oc8051_gm_cxrom_1.cell0.data [7], _13704_);
  dff (\oc8051_gm_cxrom_1.cell0.valid , _13707_);
  dff (\oc8051_gm_cxrom_1.cell1.data [0], _13763_);
  dff (\oc8051_gm_cxrom_1.cell1.data [1], _13767_);
  dff (\oc8051_gm_cxrom_1.cell1.data [2], _13771_);
  dff (\oc8051_gm_cxrom_1.cell1.data [3], _13775_);
  dff (\oc8051_gm_cxrom_1.cell1.data [4], _13779_);
  dff (\oc8051_gm_cxrom_1.cell1.data [5], _13782_);
  dff (\oc8051_gm_cxrom_1.cell1.data [6], _13786_);
  dff (\oc8051_gm_cxrom_1.cell1.data [7], _13756_);
  dff (\oc8051_gm_cxrom_1.cell1.valid , _13759_);
  dff (\oc8051_gm_cxrom_1.cell10.data [0], _00369_);
  dff (\oc8051_gm_cxrom_1.cell10.data [1], _00373_);
  dff (\oc8051_gm_cxrom_1.cell10.data [2], _00376_);
  dff (\oc8051_gm_cxrom_1.cell10.data [3], _00379_);
  dff (\oc8051_gm_cxrom_1.cell10.data [4], _00382_);
  dff (\oc8051_gm_cxrom_1.cell10.data [5], _00386_);
  dff (\oc8051_gm_cxrom_1.cell10.data [6], _00389_);
  dff (\oc8051_gm_cxrom_1.cell10.data [7], _00364_);
  dff (\oc8051_gm_cxrom_1.cell10.valid , _00366_);
  dff (\oc8051_gm_cxrom_1.cell11.data [0], _00411_);
  dff (\oc8051_gm_cxrom_1.cell11.data [1], _00415_);
  dff (\oc8051_gm_cxrom_1.cell11.data [2], _00418_);
  dff (\oc8051_gm_cxrom_1.cell11.data [3], _00421_);
  dff (\oc8051_gm_cxrom_1.cell11.data [4], _00424_);
  dff (\oc8051_gm_cxrom_1.cell11.data [5], _00428_);
  dff (\oc8051_gm_cxrom_1.cell11.data [6], _00431_);
  dff (\oc8051_gm_cxrom_1.cell11.data [7], _00406_);
  dff (\oc8051_gm_cxrom_1.cell11.valid , _00408_);
  dff (\oc8051_gm_cxrom_1.cell12.data [0], _00456_);
  dff (\oc8051_gm_cxrom_1.cell12.data [1], _00459_);
  dff (\oc8051_gm_cxrom_1.cell12.data [2], _00463_);
  dff (\oc8051_gm_cxrom_1.cell12.data [3], _00466_);
  dff (\oc8051_gm_cxrom_1.cell12.data [4], _00470_);
  dff (\oc8051_gm_cxrom_1.cell12.data [5], _00473_);
  dff (\oc8051_gm_cxrom_1.cell12.data [6], _00477_);
  dff (\oc8051_gm_cxrom_1.cell12.data [7], _00450_);
  dff (\oc8051_gm_cxrom_1.cell12.valid , _00452_);
  dff (\oc8051_gm_cxrom_1.cell13.data [0], _00503_);
  dff (\oc8051_gm_cxrom_1.cell13.data [1], _00506_);
  dff (\oc8051_gm_cxrom_1.cell13.data [2], _00510_);
  dff (\oc8051_gm_cxrom_1.cell13.data [3], _00514_);
  dff (\oc8051_gm_cxrom_1.cell13.data [4], _00517_);
  dff (\oc8051_gm_cxrom_1.cell13.data [5], _00521_);
  dff (\oc8051_gm_cxrom_1.cell13.data [6], _00524_);
  dff (\oc8051_gm_cxrom_1.cell13.data [7], _00496_);
  dff (\oc8051_gm_cxrom_1.cell13.valid , _00499_);
  dff (\oc8051_gm_cxrom_1.cell14.data [0], _13825_[0]);
  dff (\oc8051_gm_cxrom_1.cell14.data [1], _13825_[1]);
  dff (\oc8051_gm_cxrom_1.cell14.data [2], _13825_[2]);
  dff (\oc8051_gm_cxrom_1.cell14.data [3], _13825_[3]);
  dff (\oc8051_gm_cxrom_1.cell14.data [4], _13825_[4]);
  dff (\oc8051_gm_cxrom_1.cell14.data [5], _13825_[5]);
  dff (\oc8051_gm_cxrom_1.cell14.data [6], _13825_[6]);
  dff (\oc8051_gm_cxrom_1.cell14.data [7], _13825_[7]);
  dff (\oc8051_gm_cxrom_1.cell14.valid , _00545_);
  dff (\oc8051_gm_cxrom_1.cell15.data [0], _13826_[0]);
  dff (\oc8051_gm_cxrom_1.cell15.data [1], _13826_[1]);
  dff (\oc8051_gm_cxrom_1.cell15.data [2], _13826_[2]);
  dff (\oc8051_gm_cxrom_1.cell15.data [3], _13826_[3]);
  dff (\oc8051_gm_cxrom_1.cell15.data [4], _13826_[4]);
  dff (\oc8051_gm_cxrom_1.cell15.data [5], _13826_[5]);
  dff (\oc8051_gm_cxrom_1.cell15.data [6], _13826_[6]);
  dff (\oc8051_gm_cxrom_1.cell15.data [7], _13826_[7]);
  dff (\oc8051_gm_cxrom_1.cell15.valid , _13827_);
  dff (\oc8051_gm_cxrom_1.cell2.data [0], _13814_);
  dff (\oc8051_gm_cxrom_1.cell2.data [1], _13818_);
  dff (\oc8051_gm_cxrom_1.cell2.data [2], _13822_);
  dff (\oc8051_gm_cxrom_1.cell2.data [3], _00012_);
  dff (\oc8051_gm_cxrom_1.cell2.data [4], _00016_);
  dff (\oc8051_gm_cxrom_1.cell2.data [5], _00020_);
  dff (\oc8051_gm_cxrom_1.cell2.data [6], _00024_);
  dff (\oc8051_gm_cxrom_1.cell2.data [7], _13808_);
  dff (\oc8051_gm_cxrom_1.cell2.valid , _13810_);
  dff (\oc8051_gm_cxrom_1.cell3.data [0], _00052_);
  dff (\oc8051_gm_cxrom_1.cell3.data [1], _00056_);
  dff (\oc8051_gm_cxrom_1.cell3.data [2], _00059_);
  dff (\oc8051_gm_cxrom_1.cell3.data [3], _00063_);
  dff (\oc8051_gm_cxrom_1.cell3.data [4], _00067_);
  dff (\oc8051_gm_cxrom_1.cell3.data [5], _00071_);
  dff (\oc8051_gm_cxrom_1.cell3.data [6], _00075_);
  dff (\oc8051_gm_cxrom_1.cell3.data [7], _00045_);
  dff (\oc8051_gm_cxrom_1.cell3.valid , _00048_);
  dff (\oc8051_gm_cxrom_1.cell4.data [0], _00103_);
  dff (\oc8051_gm_cxrom_1.cell4.data [1], _00107_);
  dff (\oc8051_gm_cxrom_1.cell4.data [2], _00111_);
  dff (\oc8051_gm_cxrom_1.cell4.data [3], _00114_);
  dff (\oc8051_gm_cxrom_1.cell4.data [4], _00118_);
  dff (\oc8051_gm_cxrom_1.cell4.data [5], _00122_);
  dff (\oc8051_gm_cxrom_1.cell4.data [6], _00126_);
  dff (\oc8051_gm_cxrom_1.cell4.data [7], _00096_);
  dff (\oc8051_gm_cxrom_1.cell4.valid , _00099_);
  dff (\oc8051_gm_cxrom_1.cell5.data [0], _00153_);
  dff (\oc8051_gm_cxrom_1.cell5.data [1], _00156_);
  dff (\oc8051_gm_cxrom_1.cell5.data [2], _00160_);
  dff (\oc8051_gm_cxrom_1.cell5.data [3], _00163_);
  dff (\oc8051_gm_cxrom_1.cell5.data [4], _00167_);
  dff (\oc8051_gm_cxrom_1.cell5.data [5], _00171_);
  dff (\oc8051_gm_cxrom_1.cell5.data [6], _00174_);
  dff (\oc8051_gm_cxrom_1.cell5.data [7], _00146_);
  dff (\oc8051_gm_cxrom_1.cell5.valid , _00149_);
  dff (\oc8051_gm_cxrom_1.cell6.data [0], _00200_);
  dff (\oc8051_gm_cxrom_1.cell6.data [1], _00204_);
  dff (\oc8051_gm_cxrom_1.cell6.data [2], _00207_);
  dff (\oc8051_gm_cxrom_1.cell6.data [3], _00211_);
  dff (\oc8051_gm_cxrom_1.cell6.data [4], _00215_);
  dff (\oc8051_gm_cxrom_1.cell6.data [5], _00218_);
  dff (\oc8051_gm_cxrom_1.cell6.data [6], _00222_);
  dff (\oc8051_gm_cxrom_1.cell6.data [7], _00194_);
  dff (\oc8051_gm_cxrom_1.cell6.valid , _00197_);
  dff (\oc8051_gm_cxrom_1.cell7.data [0], _00248_);
  dff (\oc8051_gm_cxrom_1.cell7.data [1], _00251_);
  dff (\oc8051_gm_cxrom_1.cell7.data [2], _00255_);
  dff (\oc8051_gm_cxrom_1.cell7.data [3], _00259_);
  dff (\oc8051_gm_cxrom_1.cell7.data [4], _00262_);
  dff (\oc8051_gm_cxrom_1.cell7.data [5], _00266_);
  dff (\oc8051_gm_cxrom_1.cell7.data [6], _00269_);
  dff (\oc8051_gm_cxrom_1.cell7.data [7], _00241_);
  dff (\oc8051_gm_cxrom_1.cell7.valid , _00244_);
  dff (\oc8051_gm_cxrom_1.cell8.data [0], _00287_);
  dff (\oc8051_gm_cxrom_1.cell8.data [1], _00291_);
  dff (\oc8051_gm_cxrom_1.cell8.data [2], _00294_);
  dff (\oc8051_gm_cxrom_1.cell8.data [3], _00297_);
  dff (\oc8051_gm_cxrom_1.cell8.data [4], _00300_);
  dff (\oc8051_gm_cxrom_1.cell8.data [5], _00304_);
  dff (\oc8051_gm_cxrom_1.cell8.data [6], _00307_);
  dff (\oc8051_gm_cxrom_1.cell8.data [7], _00282_);
  dff (\oc8051_gm_cxrom_1.cell8.valid , _00284_);
  dff (\oc8051_gm_cxrom_1.cell9.data [0], _00327_);
  dff (\oc8051_gm_cxrom_1.cell9.data [1], _00331_);
  dff (\oc8051_gm_cxrom_1.cell9.data [2], _00334_);
  dff (\oc8051_gm_cxrom_1.cell9.data [3], _00337_);
  dff (\oc8051_gm_cxrom_1.cell9.data [4], _00340_);
  dff (\oc8051_gm_cxrom_1.cell9.data [5], _00344_);
  dff (\oc8051_gm_cxrom_1.cell9.data [6], _00347_);
  dff (\oc8051_gm_cxrom_1.cell9.data [7], _00322_);
  dff (\oc8051_gm_cxrom_1.cell9.valid , _00324_);
  dff (\oc8051_golden_model_1.IRAM[15] [0], _13905_[0]);
  dff (\oc8051_golden_model_1.IRAM[15] [1], _13905_[1]);
  dff (\oc8051_golden_model_1.IRAM[15] [2], _13905_[2]);
  dff (\oc8051_golden_model_1.IRAM[15] [3], _13905_[3]);
  dff (\oc8051_golden_model_1.IRAM[15] [4], _13905_[4]);
  dff (\oc8051_golden_model_1.IRAM[15] [5], _13905_[5]);
  dff (\oc8051_golden_model_1.IRAM[15] [6], _13905_[6]);
  dff (\oc8051_golden_model_1.IRAM[15] [7], _13905_[7]);
  dff (\oc8051_golden_model_1.IRAM[14] [0], _13904_[0]);
  dff (\oc8051_golden_model_1.IRAM[14] [1], _13904_[1]);
  dff (\oc8051_golden_model_1.IRAM[14] [2], _13904_[2]);
  dff (\oc8051_golden_model_1.IRAM[14] [3], _13904_[3]);
  dff (\oc8051_golden_model_1.IRAM[14] [4], _13904_[4]);
  dff (\oc8051_golden_model_1.IRAM[14] [5], _13904_[5]);
  dff (\oc8051_golden_model_1.IRAM[14] [6], _13904_[6]);
  dff (\oc8051_golden_model_1.IRAM[14] [7], _13904_[7]);
  dff (\oc8051_golden_model_1.IRAM[13] [0], _13903_[0]);
  dff (\oc8051_golden_model_1.IRAM[13] [1], _13903_[1]);
  dff (\oc8051_golden_model_1.IRAM[13] [2], _13903_[2]);
  dff (\oc8051_golden_model_1.IRAM[13] [3], _13903_[3]);
  dff (\oc8051_golden_model_1.IRAM[13] [4], _13903_[4]);
  dff (\oc8051_golden_model_1.IRAM[13] [5], _13903_[5]);
  dff (\oc8051_golden_model_1.IRAM[13] [6], _13903_[6]);
  dff (\oc8051_golden_model_1.IRAM[13] [7], _13903_[7]);
  dff (\oc8051_golden_model_1.IRAM[12] [0], _13902_[0]);
  dff (\oc8051_golden_model_1.IRAM[12] [1], _13902_[1]);
  dff (\oc8051_golden_model_1.IRAM[12] [2], _13902_[2]);
  dff (\oc8051_golden_model_1.IRAM[12] [3], _13902_[3]);
  dff (\oc8051_golden_model_1.IRAM[12] [4], _13902_[4]);
  dff (\oc8051_golden_model_1.IRAM[12] [5], _13902_[5]);
  dff (\oc8051_golden_model_1.IRAM[12] [6], _13902_[6]);
  dff (\oc8051_golden_model_1.IRAM[12] [7], _13902_[7]);
  dff (\oc8051_golden_model_1.IRAM[11] [0], _13901_[0]);
  dff (\oc8051_golden_model_1.IRAM[11] [1], _13901_[1]);
  dff (\oc8051_golden_model_1.IRAM[11] [2], _13901_[2]);
  dff (\oc8051_golden_model_1.IRAM[11] [3], _13901_[3]);
  dff (\oc8051_golden_model_1.IRAM[11] [4], _13901_[4]);
  dff (\oc8051_golden_model_1.IRAM[11] [5], _13901_[5]);
  dff (\oc8051_golden_model_1.IRAM[11] [6], _13901_[6]);
  dff (\oc8051_golden_model_1.IRAM[11] [7], _13901_[7]);
  dff (\oc8051_golden_model_1.IRAM[10] [0], _13900_[0]);
  dff (\oc8051_golden_model_1.IRAM[10] [1], _13900_[1]);
  dff (\oc8051_golden_model_1.IRAM[10] [2], _13900_[2]);
  dff (\oc8051_golden_model_1.IRAM[10] [3], _13900_[3]);
  dff (\oc8051_golden_model_1.IRAM[10] [4], _13900_[4]);
  dff (\oc8051_golden_model_1.IRAM[10] [5], _13900_[5]);
  dff (\oc8051_golden_model_1.IRAM[10] [6], _13900_[6]);
  dff (\oc8051_golden_model_1.IRAM[10] [7], _13900_[7]);
  dff (\oc8051_golden_model_1.IRAM[9] [0], _13892_);
  dff (\oc8051_golden_model_1.IRAM[9] [1], _13893_);
  dff (\oc8051_golden_model_1.IRAM[9] [2], _13894_);
  dff (\oc8051_golden_model_1.IRAM[9] [3], _13895_);
  dff (\oc8051_golden_model_1.IRAM[9] [4], _13896_);
  dff (\oc8051_golden_model_1.IRAM[9] [5], _13897_);
  dff (\oc8051_golden_model_1.IRAM[9] [6], _13898_);
  dff (\oc8051_golden_model_1.IRAM[9] [7], _13899_);
  dff (\oc8051_golden_model_1.IRAM[8] [0], _13909_[0]);
  dff (\oc8051_golden_model_1.IRAM[8] [1], _13909_[1]);
  dff (\oc8051_golden_model_1.IRAM[8] [2], _13909_[2]);
  dff (\oc8051_golden_model_1.IRAM[8] [3], _13909_[3]);
  dff (\oc8051_golden_model_1.IRAM[8] [4], _13909_[4]);
  dff (\oc8051_golden_model_1.IRAM[8] [5], _13909_[5]);
  dff (\oc8051_golden_model_1.IRAM[8] [6], _13909_[6]);
  dff (\oc8051_golden_model_1.IRAM[8] [7], _13909_[7]);
  dff (\oc8051_golden_model_1.IRAM[7] [0], _13884_);
  dff (\oc8051_golden_model_1.IRAM[7] [1], _13885_);
  dff (\oc8051_golden_model_1.IRAM[7] [2], _13886_);
  dff (\oc8051_golden_model_1.IRAM[7] [3], _13887_);
  dff (\oc8051_golden_model_1.IRAM[7] [4], _13888_);
  dff (\oc8051_golden_model_1.IRAM[7] [5], _13889_);
  dff (\oc8051_golden_model_1.IRAM[7] [6], _13890_);
  dff (\oc8051_golden_model_1.IRAM[7] [7], _13891_);
  dff (\oc8051_golden_model_1.IRAM[6] [0], _13908_[0]);
  dff (\oc8051_golden_model_1.IRAM[6] [1], _13908_[1]);
  dff (\oc8051_golden_model_1.IRAM[6] [2], _13908_[2]);
  dff (\oc8051_golden_model_1.IRAM[6] [3], _13908_[3]);
  dff (\oc8051_golden_model_1.IRAM[6] [4], _13908_[4]);
  dff (\oc8051_golden_model_1.IRAM[6] [5], _13908_[5]);
  dff (\oc8051_golden_model_1.IRAM[6] [6], _13908_[6]);
  dff (\oc8051_golden_model_1.IRAM[6] [7], _13908_[7]);
  dff (\oc8051_golden_model_1.IRAM[5] [0], _13907_[0]);
  dff (\oc8051_golden_model_1.IRAM[5] [1], _13907_[1]);
  dff (\oc8051_golden_model_1.IRAM[5] [2], _13907_[2]);
  dff (\oc8051_golden_model_1.IRAM[5] [3], _13907_[3]);
  dff (\oc8051_golden_model_1.IRAM[5] [4], _13907_[4]);
  dff (\oc8051_golden_model_1.IRAM[5] [5], _13907_[5]);
  dff (\oc8051_golden_model_1.IRAM[5] [6], _13907_[6]);
  dff (\oc8051_golden_model_1.IRAM[5] [7], _13907_[7]);
  dff (\oc8051_golden_model_1.IRAM[4] [0], _13906_[0]);
  dff (\oc8051_golden_model_1.IRAM[4] [1], _13906_[1]);
  dff (\oc8051_golden_model_1.IRAM[4] [2], _13906_[2]);
  dff (\oc8051_golden_model_1.IRAM[4] [3], _13906_[3]);
  dff (\oc8051_golden_model_1.IRAM[4] [4], _13906_[4]);
  dff (\oc8051_golden_model_1.IRAM[4] [5], _13906_[5]);
  dff (\oc8051_golden_model_1.IRAM[4] [6], _13906_[6]);
  dff (\oc8051_golden_model_1.IRAM[4] [7], _13906_[7]);
  dff (\oc8051_golden_model_1.IRAM[3] [0], _13876_);
  dff (\oc8051_golden_model_1.IRAM[3] [1], _13877_);
  dff (\oc8051_golden_model_1.IRAM[3] [2], _13878_);
  dff (\oc8051_golden_model_1.IRAM[3] [3], _13879_);
  dff (\oc8051_golden_model_1.IRAM[3] [4], _13880_);
  dff (\oc8051_golden_model_1.IRAM[3] [5], _13881_);
  dff (\oc8051_golden_model_1.IRAM[3] [6], _13882_);
  dff (\oc8051_golden_model_1.IRAM[3] [7], _13883_);
  dff (\oc8051_golden_model_1.IRAM[2] [0], _13868_);
  dff (\oc8051_golden_model_1.IRAM[2] [1], _13869_);
  dff (\oc8051_golden_model_1.IRAM[2] [2], _13870_);
  dff (\oc8051_golden_model_1.IRAM[2] [3], _13871_);
  dff (\oc8051_golden_model_1.IRAM[2] [4], _13872_);
  dff (\oc8051_golden_model_1.IRAM[2] [5], _13873_);
  dff (\oc8051_golden_model_1.IRAM[2] [6], _13874_);
  dff (\oc8051_golden_model_1.IRAM[2] [7], _13875_);
  dff (\oc8051_golden_model_1.IRAM[1] [0], _13860_);
  dff (\oc8051_golden_model_1.IRAM[1] [1], _13861_);
  dff (\oc8051_golden_model_1.IRAM[1] [2], _13862_);
  dff (\oc8051_golden_model_1.IRAM[1] [3], _13863_);
  dff (\oc8051_golden_model_1.IRAM[1] [4], _13864_);
  dff (\oc8051_golden_model_1.IRAM[1] [5], _13865_);
  dff (\oc8051_golden_model_1.IRAM[1] [6], _13866_);
  dff (\oc8051_golden_model_1.IRAM[1] [7], _13867_);
  dff (\oc8051_golden_model_1.IRAM[0] [0], _13852_);
  dff (\oc8051_golden_model_1.IRAM[0] [1], _13853_);
  dff (\oc8051_golden_model_1.IRAM[0] [2], _13854_);
  dff (\oc8051_golden_model_1.IRAM[0] [3], _13855_);
  dff (\oc8051_golden_model_1.IRAM[0] [4], _13856_);
  dff (\oc8051_golden_model_1.IRAM[0] [5], _13857_);
  dff (\oc8051_golden_model_1.IRAM[0] [6], _13858_);
  dff (\oc8051_golden_model_1.IRAM[0] [7], _13859_);
  dff (\oc8051_golden_model_1.B [0], _13829_[0]);
  dff (\oc8051_golden_model_1.B [1], _13829_[1]);
  dff (\oc8051_golden_model_1.B [2], _13829_[2]);
  dff (\oc8051_golden_model_1.B [3], _13829_[3]);
  dff (\oc8051_golden_model_1.B [4], _13829_[4]);
  dff (\oc8051_golden_model_1.B [5], _13829_[5]);
  dff (\oc8051_golden_model_1.B [6], _13829_[6]);
  dff (\oc8051_golden_model_1.B [7], _13829_[7]);
  dff (\oc8051_golden_model_1.ACC [0], _13828_[0]);
  dff (\oc8051_golden_model_1.ACC [1], _13828_[1]);
  dff (\oc8051_golden_model_1.ACC [2], _13828_[2]);
  dff (\oc8051_golden_model_1.ACC [3], _13828_[3]);
  dff (\oc8051_golden_model_1.ACC [4], _13828_[4]);
  dff (\oc8051_golden_model_1.ACC [5], _13828_[5]);
  dff (\oc8051_golden_model_1.ACC [6], _13828_[6]);
  dff (\oc8051_golden_model_1.ACC [7], _13828_[7]);
  dff (\oc8051_golden_model_1.DPL [0], _13831_[0]);
  dff (\oc8051_golden_model_1.DPL [1], _13831_[1]);
  dff (\oc8051_golden_model_1.DPL [2], _13831_[2]);
  dff (\oc8051_golden_model_1.DPL [3], _13831_[3]);
  dff (\oc8051_golden_model_1.DPL [4], _13831_[4]);
  dff (\oc8051_golden_model_1.DPL [5], _13831_[5]);
  dff (\oc8051_golden_model_1.DPL [6], _13831_[6]);
  dff (\oc8051_golden_model_1.DPL [7], _13831_[7]);
  dff (\oc8051_golden_model_1.DPH [0], _13830_[0]);
  dff (\oc8051_golden_model_1.DPH [1], _13830_[1]);
  dff (\oc8051_golden_model_1.DPH [2], _13830_[2]);
  dff (\oc8051_golden_model_1.DPH [3], _13830_[3]);
  dff (\oc8051_golden_model_1.DPH [4], _13830_[4]);
  dff (\oc8051_golden_model_1.DPH [5], _13830_[5]);
  dff (\oc8051_golden_model_1.DPH [6], _13830_[6]);
  dff (\oc8051_golden_model_1.DPH [7], _13830_[7]);
  dff (\oc8051_golden_model_1.IE [0], _13832_[0]);
  dff (\oc8051_golden_model_1.IE [1], _13832_[1]);
  dff (\oc8051_golden_model_1.IE [2], _13832_[2]);
  dff (\oc8051_golden_model_1.IE [3], _13832_[3]);
  dff (\oc8051_golden_model_1.IE [4], _13832_[4]);
  dff (\oc8051_golden_model_1.IE [5], _13832_[5]);
  dff (\oc8051_golden_model_1.IE [6], _13832_[6]);
  dff (\oc8051_golden_model_1.IE [7], _13832_[7]);
  dff (\oc8051_golden_model_1.IP [0], _13833_[0]);
  dff (\oc8051_golden_model_1.IP [1], _13833_[1]);
  dff (\oc8051_golden_model_1.IP [2], _13833_[2]);
  dff (\oc8051_golden_model_1.IP [3], _13833_[3]);
  dff (\oc8051_golden_model_1.IP [4], _13833_[4]);
  dff (\oc8051_golden_model_1.IP [5], _13833_[5]);
  dff (\oc8051_golden_model_1.IP [6], _13833_[6]);
  dff (\oc8051_golden_model_1.IP [7], _13833_[7]);
  dff (\oc8051_golden_model_1.P0 [0], _13834_[0]);
  dff (\oc8051_golden_model_1.P0 [1], _13834_[1]);
  dff (\oc8051_golden_model_1.P0 [2], _13834_[2]);
  dff (\oc8051_golden_model_1.P0 [3], _13834_[3]);
  dff (\oc8051_golden_model_1.P0 [4], _13834_[4]);
  dff (\oc8051_golden_model_1.P0 [5], _13834_[5]);
  dff (\oc8051_golden_model_1.P0 [6], _13834_[6]);
  dff (\oc8051_golden_model_1.P0 [7], _13834_[7]);
  dff (\oc8051_golden_model_1.P1 [0], _13835_[0]);
  dff (\oc8051_golden_model_1.P1 [1], _13835_[1]);
  dff (\oc8051_golden_model_1.P1 [2], _13835_[2]);
  dff (\oc8051_golden_model_1.P1 [3], _13835_[3]);
  dff (\oc8051_golden_model_1.P1 [4], _13835_[4]);
  dff (\oc8051_golden_model_1.P1 [5], _13835_[5]);
  dff (\oc8051_golden_model_1.P1 [6], _13835_[6]);
  dff (\oc8051_golden_model_1.P1 [7], _13835_[7]);
  dff (\oc8051_golden_model_1.P2 [0], _13836_[0]);
  dff (\oc8051_golden_model_1.P2 [1], _13836_[1]);
  dff (\oc8051_golden_model_1.P2 [2], _13836_[2]);
  dff (\oc8051_golden_model_1.P2 [3], _13836_[3]);
  dff (\oc8051_golden_model_1.P2 [4], _13836_[4]);
  dff (\oc8051_golden_model_1.P2 [5], _13836_[5]);
  dff (\oc8051_golden_model_1.P2 [6], _13836_[6]);
  dff (\oc8051_golden_model_1.P2 [7], _13836_[7]);
  dff (\oc8051_golden_model_1.P3 [0], _13837_[0]);
  dff (\oc8051_golden_model_1.P3 [1], _13837_[1]);
  dff (\oc8051_golden_model_1.P3 [2], _13837_[2]);
  dff (\oc8051_golden_model_1.P3 [3], _13837_[3]);
  dff (\oc8051_golden_model_1.P3 [4], _13837_[4]);
  dff (\oc8051_golden_model_1.P3 [5], _13837_[5]);
  dff (\oc8051_golden_model_1.P3 [6], _13837_[6]);
  dff (\oc8051_golden_model_1.P3 [7], _13837_[7]);
  dff (\oc8051_golden_model_1.PSW [0], _13840_[0]);
  dff (\oc8051_golden_model_1.PSW [1], _13840_[1]);
  dff (\oc8051_golden_model_1.PSW [2], _13840_[2]);
  dff (\oc8051_golden_model_1.PSW [3], _13840_[3]);
  dff (\oc8051_golden_model_1.PSW [4], _13840_[4]);
  dff (\oc8051_golden_model_1.PSW [5], _13840_[5]);
  dff (\oc8051_golden_model_1.PSW [6], _13840_[6]);
  dff (\oc8051_golden_model_1.PSW [7], _13840_[7]);
  dff (\oc8051_golden_model_1.PCON [0], _13838_[0]);
  dff (\oc8051_golden_model_1.PCON [1], _13838_[1]);
  dff (\oc8051_golden_model_1.PCON [2], _13838_[2]);
  dff (\oc8051_golden_model_1.PCON [3], _13838_[3]);
  dff (\oc8051_golden_model_1.PCON [4], _13838_[4]);
  dff (\oc8051_golden_model_1.PCON [5], _13838_[5]);
  dff (\oc8051_golden_model_1.PCON [6], _13838_[6]);
  dff (\oc8051_golden_model_1.PCON [7], _13838_[7]);
  dff (\oc8051_golden_model_1.SBUF [0], _13841_[0]);
  dff (\oc8051_golden_model_1.SBUF [1], _13841_[1]);
  dff (\oc8051_golden_model_1.SBUF [2], _13841_[2]);
  dff (\oc8051_golden_model_1.SBUF [3], _13841_[3]);
  dff (\oc8051_golden_model_1.SBUF [4], _13841_[4]);
  dff (\oc8051_golden_model_1.SBUF [5], _13841_[5]);
  dff (\oc8051_golden_model_1.SBUF [6], _13841_[6]);
  dff (\oc8051_golden_model_1.SBUF [7], _13841_[7]);
  dff (\oc8051_golden_model_1.SCON [0], _13842_[0]);
  dff (\oc8051_golden_model_1.SCON [1], _13842_[1]);
  dff (\oc8051_golden_model_1.SCON [2], _13842_[2]);
  dff (\oc8051_golden_model_1.SCON [3], _13842_[3]);
  dff (\oc8051_golden_model_1.SCON [4], _13842_[4]);
  dff (\oc8051_golden_model_1.SCON [5], _13842_[5]);
  dff (\oc8051_golden_model_1.SCON [6], _13842_[6]);
  dff (\oc8051_golden_model_1.SCON [7], _13842_[7]);
  dff (\oc8051_golden_model_1.SP [0], _13843_[0]);
  dff (\oc8051_golden_model_1.SP [1], _13843_[1]);
  dff (\oc8051_golden_model_1.SP [2], _13843_[2]);
  dff (\oc8051_golden_model_1.SP [3], _13843_[3]);
  dff (\oc8051_golden_model_1.SP [4], _13843_[4]);
  dff (\oc8051_golden_model_1.SP [5], _13843_[5]);
  dff (\oc8051_golden_model_1.SP [6], _13843_[6]);
  dff (\oc8051_golden_model_1.SP [7], _13843_[7]);
  dff (\oc8051_golden_model_1.TCON [0], _13844_[0]);
  dff (\oc8051_golden_model_1.TCON [1], _13844_[1]);
  dff (\oc8051_golden_model_1.TCON [2], _13844_[2]);
  dff (\oc8051_golden_model_1.TCON [3], _13844_[3]);
  dff (\oc8051_golden_model_1.TCON [4], _13844_[4]);
  dff (\oc8051_golden_model_1.TCON [5], _13844_[5]);
  dff (\oc8051_golden_model_1.TCON [6], _13844_[6]);
  dff (\oc8051_golden_model_1.TCON [7], _13844_[7]);
  dff (\oc8051_golden_model_1.TH0 [0], _13845_[0]);
  dff (\oc8051_golden_model_1.TH0 [1], _13845_[1]);
  dff (\oc8051_golden_model_1.TH0 [2], _13845_[2]);
  dff (\oc8051_golden_model_1.TH0 [3], _13845_[3]);
  dff (\oc8051_golden_model_1.TH0 [4], _13845_[4]);
  dff (\oc8051_golden_model_1.TH0 [5], _13845_[5]);
  dff (\oc8051_golden_model_1.TH0 [6], _13845_[6]);
  dff (\oc8051_golden_model_1.TH0 [7], _13845_[7]);
  dff (\oc8051_golden_model_1.TH1 [0], _13846_[0]);
  dff (\oc8051_golden_model_1.TH1 [1], _13846_[1]);
  dff (\oc8051_golden_model_1.TH1 [2], _13846_[2]);
  dff (\oc8051_golden_model_1.TH1 [3], _13846_[3]);
  dff (\oc8051_golden_model_1.TH1 [4], _13846_[4]);
  dff (\oc8051_golden_model_1.TH1 [5], _13846_[5]);
  dff (\oc8051_golden_model_1.TH1 [6], _13846_[6]);
  dff (\oc8051_golden_model_1.TH1 [7], _13846_[7]);
  dff (\oc8051_golden_model_1.TL0 [0], _13847_[0]);
  dff (\oc8051_golden_model_1.TL0 [1], _13847_[1]);
  dff (\oc8051_golden_model_1.TL0 [2], _13847_[2]);
  dff (\oc8051_golden_model_1.TL0 [3], _13847_[3]);
  dff (\oc8051_golden_model_1.TL0 [4], _13847_[4]);
  dff (\oc8051_golden_model_1.TL0 [5], _13847_[5]);
  dff (\oc8051_golden_model_1.TL0 [6], _13847_[6]);
  dff (\oc8051_golden_model_1.TL0 [7], _13847_[7]);
  dff (\oc8051_golden_model_1.TL1 [0], _13848_[0]);
  dff (\oc8051_golden_model_1.TL1 [1], _13848_[1]);
  dff (\oc8051_golden_model_1.TL1 [2], _13848_[2]);
  dff (\oc8051_golden_model_1.TL1 [3], _13848_[3]);
  dff (\oc8051_golden_model_1.TL1 [4], _13848_[4]);
  dff (\oc8051_golden_model_1.TL1 [5], _13848_[5]);
  dff (\oc8051_golden_model_1.TL1 [6], _13848_[6]);
  dff (\oc8051_golden_model_1.TL1 [7], _13848_[7]);
  dff (\oc8051_golden_model_1.TMOD [0], _13849_[0]);
  dff (\oc8051_golden_model_1.TMOD [1], _13849_[1]);
  dff (\oc8051_golden_model_1.TMOD [2], _13849_[2]);
  dff (\oc8051_golden_model_1.TMOD [3], _13849_[3]);
  dff (\oc8051_golden_model_1.TMOD [4], _13849_[4]);
  dff (\oc8051_golden_model_1.TMOD [5], _13849_[5]);
  dff (\oc8051_golden_model_1.TMOD [6], _13849_[6]);
  dff (\oc8051_golden_model_1.TMOD [7], _13849_[7]);
  dff (\oc8051_golden_model_1.XRAM_ADDR [0], _13850_[0]);
  dff (\oc8051_golden_model_1.XRAM_ADDR [1], _13850_[1]);
  dff (\oc8051_golden_model_1.XRAM_ADDR [2], _13850_[2]);
  dff (\oc8051_golden_model_1.XRAM_ADDR [3], _13850_[3]);
  dff (\oc8051_golden_model_1.XRAM_ADDR [4], _13850_[4]);
  dff (\oc8051_golden_model_1.XRAM_ADDR [5], _13850_[5]);
  dff (\oc8051_golden_model_1.XRAM_ADDR [6], _13850_[6]);
  dff (\oc8051_golden_model_1.XRAM_ADDR [7], _13850_[7]);
  dff (\oc8051_golden_model_1.XRAM_ADDR [8], _13850_[8]);
  dff (\oc8051_golden_model_1.XRAM_ADDR [9], _13850_[9]);
  dff (\oc8051_golden_model_1.XRAM_ADDR [10], _13850_[10]);
  dff (\oc8051_golden_model_1.XRAM_ADDR [11], _13850_[11]);
  dff (\oc8051_golden_model_1.XRAM_ADDR [12], _13850_[12]);
  dff (\oc8051_golden_model_1.XRAM_ADDR [13], _13850_[13]);
  dff (\oc8051_golden_model_1.XRAM_ADDR [14], _13850_[14]);
  dff (\oc8051_golden_model_1.XRAM_ADDR [15], _13850_[15]);
  dff (\oc8051_golden_model_1.PC [0], _13839_[0]);
  dff (\oc8051_golden_model_1.PC [1], _13839_[1]);
  dff (\oc8051_golden_model_1.PC [2], _13839_[2]);
  dff (\oc8051_golden_model_1.PC [3], _13839_[3]);
  dff (\oc8051_golden_model_1.PC [4], _13839_[4]);
  dff (\oc8051_golden_model_1.PC [5], _13839_[5]);
  dff (\oc8051_golden_model_1.PC [6], _13839_[6]);
  dff (\oc8051_golden_model_1.PC [7], _13839_[7]);
  dff (\oc8051_golden_model_1.PC [8], _13839_[8]);
  dff (\oc8051_golden_model_1.PC [9], _13839_[9]);
  dff (\oc8051_golden_model_1.PC [10], _13839_[10]);
  dff (\oc8051_golden_model_1.PC [11], _13839_[11]);
  dff (\oc8051_golden_model_1.PC [12], _13839_[12]);
  dff (\oc8051_golden_model_1.PC [13], _13839_[13]);
  dff (\oc8051_golden_model_1.PC [14], _13839_[14]);
  dff (\oc8051_golden_model_1.PC [15], _13839_[15]);
  dff (\oc8051_golden_model_1.XRAM_DATA_OUT [0], _13851_[0]);
  dff (\oc8051_golden_model_1.XRAM_DATA_OUT [1], _13851_[1]);
  dff (\oc8051_golden_model_1.XRAM_DATA_OUT [2], _13851_[2]);
  dff (\oc8051_golden_model_1.XRAM_DATA_OUT [3], _13851_[3]);
  dff (\oc8051_golden_model_1.XRAM_DATA_OUT [4], _13851_[4]);
  dff (\oc8051_golden_model_1.XRAM_DATA_OUT [5], _13851_[5]);
  dff (\oc8051_golden_model_1.XRAM_DATA_OUT [6], _13851_[6]);
  dff (\oc8051_golden_model_1.XRAM_DATA_OUT [7], _13851_[7]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _03008_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _03019_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _03040_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _03061_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4], _03082_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5], _01048_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], _03093_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1], _01017_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0], _03104_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1], _03115_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2], _03126_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3], _03137_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4], _03148_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5], _03160_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6], _03171_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7], _01069_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], _02746_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _07572_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0], _02947_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1], _03159_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2], _03362_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3], _03563_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4], _03764_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5], _03957_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6], _04143_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7], _04316_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8], _04402_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9], _04488_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10], _04574_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11], _04659_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12], _04745_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13], _04830_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [14], _04921_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [15], _07759_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [0], _13910_[0]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [1], _13910_[1]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [2], _13910_[2]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [3], _13910_[3]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [4], _13910_[4]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [5], _13910_[5]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [6], _13910_[6]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [7], _13910_[7]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [0], _13911_[0]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [1], _13911_[1]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [2], _13911_[2]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [3], _13911_[3]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [4], _13911_[4]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [5], _13911_[5]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [6], _13911_[6]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [7], _13911_[7]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [0], _13912_[0]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [1], _13912_[1]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [2], _13912_[2]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [3], _13912_[3]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [4], _13912_[4]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [5], _13912_[5]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [6], _13912_[6]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [7], _13912_[7]);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], _13913_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], _13913_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], _13913_[2]);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [0], _13914_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [1], _13914_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [2], _13914_[2]);
  dff (\oc8051_top_1.oc8051_decoder1.state [0], _13915_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.state [1], _13915_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.op [0], _13916_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.op [1], _13916_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.op [2], _13916_[2]);
  dff (\oc8051_top_1.oc8051_decoder1.op [3], _13916_[3]);
  dff (\oc8051_top_1.oc8051_decoder1.op [4], _13916_[4]);
  dff (\oc8051_top_1.oc8051_decoder1.op [5], _13916_[5]);
  dff (\oc8051_top_1.oc8051_decoder1.op [6], _13916_[6]);
  dff (\oc8051_top_1.oc8051_decoder1.op [7], _13916_[7]);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel3 , _13917_);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [0], _13918_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [1], _13918_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [0], _13919_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [1], _13919_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _13920_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _13920_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], _13920_[2]);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [0], _13921_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [1], _13921_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [2], _13921_[2]);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [0], _13922_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [1], _13922_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [0], _13923_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [1], _13923_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [2], _13923_[2]);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [3], _13923_[3]);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [0], _13924_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [1], _13924_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.wr , _13925_);
  dff (\oc8051_top_1.oc8051_indi_addr1.wr_bit_r , _13926_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [0], _13927_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [1], _13927_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [2], _13927_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [3], _13927_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [4], _13927_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [5], _13927_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [6], _13927_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [7], _13927_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [8], _13927_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [9], _13927_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [10], _13927_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [11], _13927_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [12], _13927_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [13], _13927_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [14], _13927_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [15], _13927_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _13928_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _13928_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _13928_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _13928_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _13928_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _13928_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _13928_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _13928_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _13928_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _13928_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _13928_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _13928_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _13928_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _13928_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _13928_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _13928_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [0], _13952_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [1], _13952_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [2], _13952_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [3], _13952_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [4], _13952_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [5], _13952_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [6], _13952_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [7], _13952_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [8], _13952_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [9], _13952_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [10], _13952_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [11], _13952_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [12], _13952_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [13], _13952_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [14], _13952_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [15], _13952_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [16], _13952_[16]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [17], _13952_[17]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [18], _13952_[18]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [19], _13952_[19]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [20], _13952_[20]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [21], _13952_[21]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [22], _13952_[22]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [23], _13952_[23]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [24], _13952_[24]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [25], _13952_[25]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [26], _13952_[26]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [27], _13952_[27]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [28], _13952_[28]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [29], _13952_[29]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [30], _13952_[30]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [31], _13952_[31]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _13929_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dack_ir , _13930_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [0], _13931_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [1], _13931_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [2], _13931_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [3], _13931_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [4], _13931_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [0], _13932_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [1], _13932_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [2], _13932_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [3], _13932_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [4], _13932_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [5], _13932_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [6], _13932_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [7], _13932_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [0], _13933_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [1], _13933_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [2], _13933_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [3], _13933_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [4], _13933_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [5], _13933_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [6], _13933_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [7], _13933_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [0], _13934_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [1], _13934_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [2], _13934_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [3], _13934_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [4], _13934_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [5], _13934_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [6], _13934_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [7], _13934_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _13935_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _13936_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], _13937_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _13937_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], _13937_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], _13937_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _13937_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], _13937_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], _13937_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [7], _13937_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [0], _13938_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [1], _13938_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _13938_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [3], _13938_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [4], _13938_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [5], _13938_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [6], _13938_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [7], _13938_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [8], _13938_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [9], _13938_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [10], _13938_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [11], _13938_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [12], _13938_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [13], _13938_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [14], _13938_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [15], _13938_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [0], _13939_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [1], _13939_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [2], _13939_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [3], _13939_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [4], _13939_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [5], _13939_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [6], _13939_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [7], _13939_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [8], _13939_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [9], _13939_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [10], _13939_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [11], _13939_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [12], _13939_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [13], _13939_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [14], _13939_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [15], _13939_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack , _13940_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_t , _13942_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_buff , _13941_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], _13943_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], _13943_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _13943_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], _13943_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _13943_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], _13943_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _13943_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _13943_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [0], _13944_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [1], _13944_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [2], _13944_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [0], _13945_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [1], _13945_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [2], _13945_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [3], _13945_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [4], _13945_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [5], _13945_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [6], _13945_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [7], _13945_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [0], _13946_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [1], _13946_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [2], _13946_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [3], _13946_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [4], _13946_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [5], _13946_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [6], _13946_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [7], _13946_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.reti , _13947_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [0], _13948_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [1], _13948_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [2], _13948_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [3], _13948_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [4], _13948_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [5], _13948_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [6], _13948_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [7], _13948_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdone , _13949_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst , _13950_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], _13951_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], _13951_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], _13951_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], _13951_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [0], _13953_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [1], _13953_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [2], _13953_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [3], _13953_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [4], _13953_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [5], _13953_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [6], _13953_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [7], _13953_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [8], _13953_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [9], _13953_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [10], _13953_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [11], _13953_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [12], _13953_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [13], _13953_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [14], _13953_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [15], _13953_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [16], _13953_[16]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [17], _13953_[17]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [18], _13953_[18]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [19], _13953_[19]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [20], _13953_[20]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [21], _13953_[21]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [22], _13953_[22]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [23], _13953_[23]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [24], _13953_[24]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [25], _13953_[25]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [26], _13953_[26]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [27], _13953_[27]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [28], _13953_[28]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [29], _13953_[29]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [30], _13953_[30]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [31], _13953_[31]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [0], _13954_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [1], _13954_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [2], _13954_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [3], _13954_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [4], _13954_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [5], _13954_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [6], _13954_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [7], _13954_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dwe_o , _13955_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dstb_o , _13956_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [0], _13957_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [1], _13957_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [2], _13957_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [3], _13957_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [4], _13957_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [5], _13957_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [6], _13957_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [7], _13957_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [8], _13957_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [9], _13957_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [10], _13957_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [11], _13957_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [12], _13957_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [13], _13957_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [14], _13957_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [15], _13957_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dmem_wait , _13958_);
  dff (\oc8051_top_1.oc8051_memory_interface1.istb_t , _13959_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imem_wait , _13960_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _13961_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _13961_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _13961_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _13961_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [4], _13961_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [5], _13961_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [6], _13961_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [7], _13961_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [8], _13961_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [9], _13961_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [10], _13961_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [11], _13961_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [12], _13961_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [13], _13961_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [14], _13961_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [15], _13961_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_ind , _13962_);
  dff (\oc8051_top_1.oc8051_ram_top1.rd_en_r , _13963_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _13964_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _13964_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _13964_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _13964_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _13964_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _13964_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _13964_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [7], _13964_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_addr_r , _13965_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [0], _13966_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [1], _13966_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [2], _13966_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0], _11586_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1], _11591_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2], _11596_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3], _11601_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4], _11606_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5], _11612_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6], _11617_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7], _11619_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0], _11626_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1], _11630_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2], _11633_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3], _11637_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4], _11640_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5], _11644_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6], _11647_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7], _11650_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0], _11801_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1], _11804_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2], _11808_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3], _11811_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4], _11815_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5], _11818_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6], _11822_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7], _11824_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0], _11773_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1], _11776_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2], _11780_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3], _11783_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4], _11787_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5], _11790_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6], _11794_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7], _11796_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0], _11744_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1], _11748_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2], _11751_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3], _11755_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4], _11758_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5], _11762_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6], _11766_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7], _11768_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0], _11716_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1], _11720_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2], _11723_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3], _11727_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4], _11730_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5], _11734_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6], _11737_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7], _11740_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0], _11686_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1], _11689_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2], _11693_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3], _11696_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4], _11700_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5], _11703_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6], _11707_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7], _11710_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0], _11657_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1], _11660_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2], _11664_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3], _11667_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4], _11671_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5], _11674_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6], _11678_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7], _11681_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0], _11831_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1], _11835_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2], _11838_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3], _11842_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4], _11845_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5], _11849_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6], _11852_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7], _11855_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0], _12001_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1], _12004_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2], _12008_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3], _12011_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4], _12015_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5], _12018_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6], _12022_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7], _12024_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0], _11972_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1], _11976_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2], _11979_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3], _11983_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4], _11986_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5], _11990_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6], _11994_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7], _11996_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0], _11944_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1], _11948_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2], _11951_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3], _11955_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4], _11958_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5], _11962_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6], _11965_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7], _11968_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0], _11915_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1], _11919_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2], _11922_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3], _11926_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4], _11929_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5], _11933_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6], _11937_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7], _11939_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0], _11887_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1], _11891_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2], _11894_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3], _11898_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4], _11901_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5], _11905_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6], _11908_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7], _11911_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0], _11859_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1], _11863_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2], _11866_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3], _11870_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4], _11873_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5], _11877_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6], _11880_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7], _11883_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0], _12029_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1], _12032_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2], _12036_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3], _12039_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4], _12043_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5], _12046_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6], _12050_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7], _11343_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0], _13685_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1], _13687_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2], _13688_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3], _13690_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4], _13692_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5], _13694_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6], _13696_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7], _11331_);
  dff (\oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  dff (\oc8051_top_1.oc8051_rom1.ea_int , 1'b1);
  dff (\oc8051_top_1.oc8051_sfr1.bit_out , _13967_);
  dff (\oc8051_top_1.oc8051_sfr1.wait_data , _13968_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [0], _13969_[0]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [1], _13969_[1]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [2], _13969_[2]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [3], _13969_[3]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [4], _13969_[4]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [5], _13969_[5]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [6], _13969_[6]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [7], _13969_[7]);
  dff (\oc8051_top_1.oc8051_sfr1.wr_bit_r , _13970_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], _07525_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], _07527_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], _07529_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3], _07531_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4], _07533_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], _07535_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], _07537_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], _07355_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0], _06807_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1], _06808_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2], _06809_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3], _06810_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4], _06811_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5], _06812_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6], _06813_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7], _06303_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], _06825_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], _06826_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], _06827_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], _06828_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], _06829_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], _06830_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], _06831_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7], _06823_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0], _06832_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1], _06833_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2], _06834_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3], _06835_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4], _06836_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5], _06837_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6], _06838_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7], _06824_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0], _11189_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1], _11191_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2], _11193_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3], _11195_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4], _11197_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5], _11199_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6], _11201_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7], _08547_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0], _11203_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1], _11205_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2], _11207_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3], _11209_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4], _11211_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5], _11213_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6], _11215_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7], _08550_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0], _11217_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1], _11219_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2], _11221_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3], _11223_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4], _11225_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5], _11227_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6], _11229_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7], _08553_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0], _11231_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1], _11233_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2], _11235_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3], _11237_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4], _11239_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5], _11241_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6], _11243_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7], _08556_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1], _07290_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], _07292_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3], _07294_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4], _07296_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5], _07298_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6], _07300_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], _06839_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop , _06814_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], _06816_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], _06817_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2], _06818_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3], _06819_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4], _06820_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5], _06821_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6], _06822_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7], _06815_);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div0 , \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div1 , \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [0], psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [0], psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [1], \oc8051_top_1.oc8051_sfr1.psw_next [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [2], \oc8051_top_1.oc8051_sfr1.psw_next [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [3], \oc8051_top_1.oc8051_sfr1.psw_next [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [4], \oc8051_top_1.oc8051_sfr1.psw_next [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [5], \oc8051_top_1.oc8051_sfr1.psw_next [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [6], \oc8051_top_1.oc8051_sfr1.psw_next [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [7], \oc8051_top_1.oc8051_sfr1.psw_next [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [1], \oc8051_top_1.oc8051_sfr1.psw_next [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [2], \oc8051_top_1.oc8051_sfr1.psw_next [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [3], \oc8051_top_1.oc8051_sfr1.psw_next [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [4], \oc8051_top_1.oc8051_sfr1.psw_next [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [5], \oc8051_top_1.oc8051_sfr1.psw_next [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [6], \oc8051_top_1.oc8051_sfr1.psw_next [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [7], \oc8051_top_1.oc8051_sfr1.psw_next [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.p , psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell0.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell0.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell0.word [0], word_in[0]);
  buf(\oc8051_gm_cxrom_1.cell0.word [1], word_in[1]);
  buf(\oc8051_gm_cxrom_1.cell0.word [2], word_in[2]);
  buf(\oc8051_gm_cxrom_1.cell0.word [3], word_in[3]);
  buf(\oc8051_gm_cxrom_1.cell0.word [4], word_in[4]);
  buf(\oc8051_gm_cxrom_1.cell0.word [5], word_in[5]);
  buf(\oc8051_gm_cxrom_1.cell0.word [6], word_in[6]);
  buf(\oc8051_gm_cxrom_1.cell0.word [7], word_in[7]);
  buf(\oc8051_gm_cxrom_1.cell1.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell1.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell1.word [0], word_in[8]);
  buf(\oc8051_gm_cxrom_1.cell1.word [1], word_in[9]);
  buf(\oc8051_gm_cxrom_1.cell1.word [2], word_in[10]);
  buf(\oc8051_gm_cxrom_1.cell1.word [3], word_in[11]);
  buf(\oc8051_gm_cxrom_1.cell1.word [4], word_in[12]);
  buf(\oc8051_gm_cxrom_1.cell1.word [5], word_in[13]);
  buf(\oc8051_gm_cxrom_1.cell1.word [6], word_in[14]);
  buf(\oc8051_gm_cxrom_1.cell1.word [7], word_in[15]);
  buf(\oc8051_gm_cxrom_1.cell2.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell2.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell2.word [0], word_in[16]);
  buf(\oc8051_gm_cxrom_1.cell2.word [1], word_in[17]);
  buf(\oc8051_gm_cxrom_1.cell2.word [2], word_in[18]);
  buf(\oc8051_gm_cxrom_1.cell2.word [3], word_in[19]);
  buf(\oc8051_gm_cxrom_1.cell2.word [4], word_in[20]);
  buf(\oc8051_gm_cxrom_1.cell2.word [5], word_in[21]);
  buf(\oc8051_gm_cxrom_1.cell2.word [6], word_in[22]);
  buf(\oc8051_gm_cxrom_1.cell2.word [7], word_in[23]);
  buf(\oc8051_gm_cxrom_1.cell3.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell3.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell3.word [0], word_in[24]);
  buf(\oc8051_gm_cxrom_1.cell3.word [1], word_in[25]);
  buf(\oc8051_gm_cxrom_1.cell3.word [2], word_in[26]);
  buf(\oc8051_gm_cxrom_1.cell3.word [3], word_in[27]);
  buf(\oc8051_gm_cxrom_1.cell3.word [4], word_in[28]);
  buf(\oc8051_gm_cxrom_1.cell3.word [5], word_in[29]);
  buf(\oc8051_gm_cxrom_1.cell3.word [6], word_in[30]);
  buf(\oc8051_gm_cxrom_1.cell3.word [7], word_in[31]);
  buf(\oc8051_gm_cxrom_1.cell4.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell4.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell4.word [0], word_in[32]);
  buf(\oc8051_gm_cxrom_1.cell4.word [1], word_in[33]);
  buf(\oc8051_gm_cxrom_1.cell4.word [2], word_in[34]);
  buf(\oc8051_gm_cxrom_1.cell4.word [3], word_in[35]);
  buf(\oc8051_gm_cxrom_1.cell4.word [4], word_in[36]);
  buf(\oc8051_gm_cxrom_1.cell4.word [5], word_in[37]);
  buf(\oc8051_gm_cxrom_1.cell4.word [6], word_in[38]);
  buf(\oc8051_gm_cxrom_1.cell4.word [7], word_in[39]);
  buf(\oc8051_gm_cxrom_1.cell5.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell5.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell5.word [0], word_in[40]);
  buf(\oc8051_gm_cxrom_1.cell5.word [1], word_in[41]);
  buf(\oc8051_gm_cxrom_1.cell5.word [2], word_in[42]);
  buf(\oc8051_gm_cxrom_1.cell5.word [3], word_in[43]);
  buf(\oc8051_gm_cxrom_1.cell5.word [4], word_in[44]);
  buf(\oc8051_gm_cxrom_1.cell5.word [5], word_in[45]);
  buf(\oc8051_gm_cxrom_1.cell5.word [6], word_in[46]);
  buf(\oc8051_gm_cxrom_1.cell5.word [7], word_in[47]);
  buf(\oc8051_gm_cxrom_1.cell6.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell6.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell6.word [0], word_in[48]);
  buf(\oc8051_gm_cxrom_1.cell6.word [1], word_in[49]);
  buf(\oc8051_gm_cxrom_1.cell6.word [2], word_in[50]);
  buf(\oc8051_gm_cxrom_1.cell6.word [3], word_in[51]);
  buf(\oc8051_gm_cxrom_1.cell6.word [4], word_in[52]);
  buf(\oc8051_gm_cxrom_1.cell6.word [5], word_in[53]);
  buf(\oc8051_gm_cxrom_1.cell6.word [6], word_in[54]);
  buf(\oc8051_gm_cxrom_1.cell6.word [7], word_in[55]);
  buf(\oc8051_gm_cxrom_1.cell7.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell7.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell7.word [0], word_in[56]);
  buf(\oc8051_gm_cxrom_1.cell7.word [1], word_in[57]);
  buf(\oc8051_gm_cxrom_1.cell7.word [2], word_in[58]);
  buf(\oc8051_gm_cxrom_1.cell7.word [3], word_in[59]);
  buf(\oc8051_gm_cxrom_1.cell7.word [4], word_in[60]);
  buf(\oc8051_gm_cxrom_1.cell7.word [5], word_in[61]);
  buf(\oc8051_gm_cxrom_1.cell7.word [6], word_in[62]);
  buf(\oc8051_gm_cxrom_1.cell7.word [7], word_in[63]);
  buf(\oc8051_gm_cxrom_1.cell8.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell8.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell8.word [0], word_in[64]);
  buf(\oc8051_gm_cxrom_1.cell8.word [1], word_in[65]);
  buf(\oc8051_gm_cxrom_1.cell8.word [2], word_in[66]);
  buf(\oc8051_gm_cxrom_1.cell8.word [3], word_in[67]);
  buf(\oc8051_gm_cxrom_1.cell8.word [4], word_in[68]);
  buf(\oc8051_gm_cxrom_1.cell8.word [5], word_in[69]);
  buf(\oc8051_gm_cxrom_1.cell8.word [6], word_in[70]);
  buf(\oc8051_gm_cxrom_1.cell8.word [7], word_in[71]);
  buf(\oc8051_gm_cxrom_1.cell9.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell9.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell9.word [0], word_in[72]);
  buf(\oc8051_gm_cxrom_1.cell9.word [1], word_in[73]);
  buf(\oc8051_gm_cxrom_1.cell9.word [2], word_in[74]);
  buf(\oc8051_gm_cxrom_1.cell9.word [3], word_in[75]);
  buf(\oc8051_gm_cxrom_1.cell9.word [4], word_in[76]);
  buf(\oc8051_gm_cxrom_1.cell9.word [5], word_in[77]);
  buf(\oc8051_gm_cxrom_1.cell9.word [6], word_in[78]);
  buf(\oc8051_gm_cxrom_1.cell9.word [7], word_in[79]);
  buf(\oc8051_gm_cxrom_1.cell10.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell10.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell10.word [0], word_in[80]);
  buf(\oc8051_gm_cxrom_1.cell10.word [1], word_in[81]);
  buf(\oc8051_gm_cxrom_1.cell10.word [2], word_in[82]);
  buf(\oc8051_gm_cxrom_1.cell10.word [3], word_in[83]);
  buf(\oc8051_gm_cxrom_1.cell10.word [4], word_in[84]);
  buf(\oc8051_gm_cxrom_1.cell10.word [5], word_in[85]);
  buf(\oc8051_gm_cxrom_1.cell10.word [6], word_in[86]);
  buf(\oc8051_gm_cxrom_1.cell10.word [7], word_in[87]);
  buf(\oc8051_gm_cxrom_1.cell11.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell11.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell11.word [0], word_in[88]);
  buf(\oc8051_gm_cxrom_1.cell11.word [1], word_in[89]);
  buf(\oc8051_gm_cxrom_1.cell11.word [2], word_in[90]);
  buf(\oc8051_gm_cxrom_1.cell11.word [3], word_in[91]);
  buf(\oc8051_gm_cxrom_1.cell11.word [4], word_in[92]);
  buf(\oc8051_gm_cxrom_1.cell11.word [5], word_in[93]);
  buf(\oc8051_gm_cxrom_1.cell11.word [6], word_in[94]);
  buf(\oc8051_gm_cxrom_1.cell11.word [7], word_in[95]);
  buf(\oc8051_gm_cxrom_1.cell12.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell12.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell12.word [0], word_in[96]);
  buf(\oc8051_gm_cxrom_1.cell12.word [1], word_in[97]);
  buf(\oc8051_gm_cxrom_1.cell12.word [2], word_in[98]);
  buf(\oc8051_gm_cxrom_1.cell12.word [3], word_in[99]);
  buf(\oc8051_gm_cxrom_1.cell12.word [4], word_in[100]);
  buf(\oc8051_gm_cxrom_1.cell12.word [5], word_in[101]);
  buf(\oc8051_gm_cxrom_1.cell12.word [6], word_in[102]);
  buf(\oc8051_gm_cxrom_1.cell12.word [7], word_in[103]);
  buf(\oc8051_gm_cxrom_1.cell13.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell13.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell13.word [0], word_in[104]);
  buf(\oc8051_gm_cxrom_1.cell13.word [1], word_in[105]);
  buf(\oc8051_gm_cxrom_1.cell13.word [2], word_in[106]);
  buf(\oc8051_gm_cxrom_1.cell13.word [3], word_in[107]);
  buf(\oc8051_gm_cxrom_1.cell13.word [4], word_in[108]);
  buf(\oc8051_gm_cxrom_1.cell13.word [5], word_in[109]);
  buf(\oc8051_gm_cxrom_1.cell13.word [6], word_in[110]);
  buf(\oc8051_gm_cxrom_1.cell13.word [7], word_in[111]);
  buf(\oc8051_gm_cxrom_1.cell14.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell14.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell14.word [0], word_in[112]);
  buf(\oc8051_gm_cxrom_1.cell14.word [1], word_in[113]);
  buf(\oc8051_gm_cxrom_1.cell14.word [2], word_in[114]);
  buf(\oc8051_gm_cxrom_1.cell14.word [3], word_in[115]);
  buf(\oc8051_gm_cxrom_1.cell14.word [4], word_in[116]);
  buf(\oc8051_gm_cxrom_1.cell14.word [5], word_in[117]);
  buf(\oc8051_gm_cxrom_1.cell14.word [6], word_in[118]);
  buf(\oc8051_gm_cxrom_1.cell14.word [7], word_in[119]);
  buf(\oc8051_gm_cxrom_1.cell15.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell15.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell15.word [0], word_in[120]);
  buf(\oc8051_gm_cxrom_1.cell15.word [1], word_in[121]);
  buf(\oc8051_gm_cxrom_1.cell15.word [2], word_in[122]);
  buf(\oc8051_gm_cxrom_1.cell15.word [3], word_in[123]);
  buf(\oc8051_gm_cxrom_1.cell15.word [4], word_in[124]);
  buf(\oc8051_gm_cxrom_1.cell15.word [5], word_in[125]);
  buf(\oc8051_gm_cxrom_1.cell15.word [6], word_in[126]);
  buf(\oc8051_gm_cxrom_1.cell15.word [7], word_in[127]);
  buf(\oc8051_top_1.oc8051_decoder1.clk , clk);
  buf(\oc8051_top_1.oc8051_decoder1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.oc8051_decoder1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.oc8051_comp1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_comp1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_comp1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_comp1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_comp1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_comp1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_comp1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_comp1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_comp1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_alu1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_in , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.rst , rst);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.oc8051_memory_interface1.dack_i , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.ddat_i [0], xram_data_in_reg[0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.ddat_i [1], xram_data_in_reg[1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.ddat_i [2], xram_data_in_reg[2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.ddat_i [3], xram_data_in_reg[3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.ddat_i [4], xram_data_in_reg[4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.ddat_i [5], xram_data_in_reg[5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.ddat_i [6], xram_data_in_reg[6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.ddat_i [7], xram_data_in_reg[7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.oc8051_indi_addr1.clk , clk);
  buf(\oc8051_top_1.oc8051_indi_addr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [0], psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p , psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_next [0], psw_impl[0]);
  buf(\oc8051_top_1.oc8051_rom1.rst , rst);
  buf(\oc8051_top_1.oc8051_rom1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.rst , rst);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  buf(\oc8051_gm_cxrom_1.clk , clk);
  buf(\oc8051_gm_cxrom_1.rst , rst);
  buf(\oc8051_gm_cxrom_1.word_in [0], word_in[0]);
  buf(\oc8051_gm_cxrom_1.word_in [1], word_in[1]);
  buf(\oc8051_gm_cxrom_1.word_in [2], word_in[2]);
  buf(\oc8051_gm_cxrom_1.word_in [3], word_in[3]);
  buf(\oc8051_gm_cxrom_1.word_in [4], word_in[4]);
  buf(\oc8051_gm_cxrom_1.word_in [5], word_in[5]);
  buf(\oc8051_gm_cxrom_1.word_in [6], word_in[6]);
  buf(\oc8051_gm_cxrom_1.word_in [7], word_in[7]);
  buf(\oc8051_gm_cxrom_1.word_in [8], word_in[8]);
  buf(\oc8051_gm_cxrom_1.word_in [9], word_in[9]);
  buf(\oc8051_gm_cxrom_1.word_in [10], word_in[10]);
  buf(\oc8051_gm_cxrom_1.word_in [11], word_in[11]);
  buf(\oc8051_gm_cxrom_1.word_in [12], word_in[12]);
  buf(\oc8051_gm_cxrom_1.word_in [13], word_in[13]);
  buf(\oc8051_gm_cxrom_1.word_in [14], word_in[14]);
  buf(\oc8051_gm_cxrom_1.word_in [15], word_in[15]);
  buf(\oc8051_gm_cxrom_1.word_in [16], word_in[16]);
  buf(\oc8051_gm_cxrom_1.word_in [17], word_in[17]);
  buf(\oc8051_gm_cxrom_1.word_in [18], word_in[18]);
  buf(\oc8051_gm_cxrom_1.word_in [19], word_in[19]);
  buf(\oc8051_gm_cxrom_1.word_in [20], word_in[20]);
  buf(\oc8051_gm_cxrom_1.word_in [21], word_in[21]);
  buf(\oc8051_gm_cxrom_1.word_in [22], word_in[22]);
  buf(\oc8051_gm_cxrom_1.word_in [23], word_in[23]);
  buf(\oc8051_gm_cxrom_1.word_in [24], word_in[24]);
  buf(\oc8051_gm_cxrom_1.word_in [25], word_in[25]);
  buf(\oc8051_gm_cxrom_1.word_in [26], word_in[26]);
  buf(\oc8051_gm_cxrom_1.word_in [27], word_in[27]);
  buf(\oc8051_gm_cxrom_1.word_in [28], word_in[28]);
  buf(\oc8051_gm_cxrom_1.word_in [29], word_in[29]);
  buf(\oc8051_gm_cxrom_1.word_in [30], word_in[30]);
  buf(\oc8051_gm_cxrom_1.word_in [31], word_in[31]);
  buf(\oc8051_gm_cxrom_1.word_in [32], word_in[32]);
  buf(\oc8051_gm_cxrom_1.word_in [33], word_in[33]);
  buf(\oc8051_gm_cxrom_1.word_in [34], word_in[34]);
  buf(\oc8051_gm_cxrom_1.word_in [35], word_in[35]);
  buf(\oc8051_gm_cxrom_1.word_in [36], word_in[36]);
  buf(\oc8051_gm_cxrom_1.word_in [37], word_in[37]);
  buf(\oc8051_gm_cxrom_1.word_in [38], word_in[38]);
  buf(\oc8051_gm_cxrom_1.word_in [39], word_in[39]);
  buf(\oc8051_gm_cxrom_1.word_in [40], word_in[40]);
  buf(\oc8051_gm_cxrom_1.word_in [41], word_in[41]);
  buf(\oc8051_gm_cxrom_1.word_in [42], word_in[42]);
  buf(\oc8051_gm_cxrom_1.word_in [43], word_in[43]);
  buf(\oc8051_gm_cxrom_1.word_in [44], word_in[44]);
  buf(\oc8051_gm_cxrom_1.word_in [45], word_in[45]);
  buf(\oc8051_gm_cxrom_1.word_in [46], word_in[46]);
  buf(\oc8051_gm_cxrom_1.word_in [47], word_in[47]);
  buf(\oc8051_gm_cxrom_1.word_in [48], word_in[48]);
  buf(\oc8051_gm_cxrom_1.word_in [49], word_in[49]);
  buf(\oc8051_gm_cxrom_1.word_in [50], word_in[50]);
  buf(\oc8051_gm_cxrom_1.word_in [51], word_in[51]);
  buf(\oc8051_gm_cxrom_1.word_in [52], word_in[52]);
  buf(\oc8051_gm_cxrom_1.word_in [53], word_in[53]);
  buf(\oc8051_gm_cxrom_1.word_in [54], word_in[54]);
  buf(\oc8051_gm_cxrom_1.word_in [55], word_in[55]);
  buf(\oc8051_gm_cxrom_1.word_in [56], word_in[56]);
  buf(\oc8051_gm_cxrom_1.word_in [57], word_in[57]);
  buf(\oc8051_gm_cxrom_1.word_in [58], word_in[58]);
  buf(\oc8051_gm_cxrom_1.word_in [59], word_in[59]);
  buf(\oc8051_gm_cxrom_1.word_in [60], word_in[60]);
  buf(\oc8051_gm_cxrom_1.word_in [61], word_in[61]);
  buf(\oc8051_gm_cxrom_1.word_in [62], word_in[62]);
  buf(\oc8051_gm_cxrom_1.word_in [63], word_in[63]);
  buf(\oc8051_gm_cxrom_1.word_in [64], word_in[64]);
  buf(\oc8051_gm_cxrom_1.word_in [65], word_in[65]);
  buf(\oc8051_gm_cxrom_1.word_in [66], word_in[66]);
  buf(\oc8051_gm_cxrom_1.word_in [67], word_in[67]);
  buf(\oc8051_gm_cxrom_1.word_in [68], word_in[68]);
  buf(\oc8051_gm_cxrom_1.word_in [69], word_in[69]);
  buf(\oc8051_gm_cxrom_1.word_in [70], word_in[70]);
  buf(\oc8051_gm_cxrom_1.word_in [71], word_in[71]);
  buf(\oc8051_gm_cxrom_1.word_in [72], word_in[72]);
  buf(\oc8051_gm_cxrom_1.word_in [73], word_in[73]);
  buf(\oc8051_gm_cxrom_1.word_in [74], word_in[74]);
  buf(\oc8051_gm_cxrom_1.word_in [75], word_in[75]);
  buf(\oc8051_gm_cxrom_1.word_in [76], word_in[76]);
  buf(\oc8051_gm_cxrom_1.word_in [77], word_in[77]);
  buf(\oc8051_gm_cxrom_1.word_in [78], word_in[78]);
  buf(\oc8051_gm_cxrom_1.word_in [79], word_in[79]);
  buf(\oc8051_gm_cxrom_1.word_in [80], word_in[80]);
  buf(\oc8051_gm_cxrom_1.word_in [81], word_in[81]);
  buf(\oc8051_gm_cxrom_1.word_in [82], word_in[82]);
  buf(\oc8051_gm_cxrom_1.word_in [83], word_in[83]);
  buf(\oc8051_gm_cxrom_1.word_in [84], word_in[84]);
  buf(\oc8051_gm_cxrom_1.word_in [85], word_in[85]);
  buf(\oc8051_gm_cxrom_1.word_in [86], word_in[86]);
  buf(\oc8051_gm_cxrom_1.word_in [87], word_in[87]);
  buf(\oc8051_gm_cxrom_1.word_in [88], word_in[88]);
  buf(\oc8051_gm_cxrom_1.word_in [89], word_in[89]);
  buf(\oc8051_gm_cxrom_1.word_in [90], word_in[90]);
  buf(\oc8051_gm_cxrom_1.word_in [91], word_in[91]);
  buf(\oc8051_gm_cxrom_1.word_in [92], word_in[92]);
  buf(\oc8051_gm_cxrom_1.word_in [93], word_in[93]);
  buf(\oc8051_gm_cxrom_1.word_in [94], word_in[94]);
  buf(\oc8051_gm_cxrom_1.word_in [95], word_in[95]);
  buf(\oc8051_gm_cxrom_1.word_in [96], word_in[96]);
  buf(\oc8051_gm_cxrom_1.word_in [97], word_in[97]);
  buf(\oc8051_gm_cxrom_1.word_in [98], word_in[98]);
  buf(\oc8051_gm_cxrom_1.word_in [99], word_in[99]);
  buf(\oc8051_gm_cxrom_1.word_in [100], word_in[100]);
  buf(\oc8051_gm_cxrom_1.word_in [101], word_in[101]);
  buf(\oc8051_gm_cxrom_1.word_in [102], word_in[102]);
  buf(\oc8051_gm_cxrom_1.word_in [103], word_in[103]);
  buf(\oc8051_gm_cxrom_1.word_in [104], word_in[104]);
  buf(\oc8051_gm_cxrom_1.word_in [105], word_in[105]);
  buf(\oc8051_gm_cxrom_1.word_in [106], word_in[106]);
  buf(\oc8051_gm_cxrom_1.word_in [107], word_in[107]);
  buf(\oc8051_gm_cxrom_1.word_in [108], word_in[108]);
  buf(\oc8051_gm_cxrom_1.word_in [109], word_in[109]);
  buf(\oc8051_gm_cxrom_1.word_in [110], word_in[110]);
  buf(\oc8051_gm_cxrom_1.word_in [111], word_in[111]);
  buf(\oc8051_gm_cxrom_1.word_in [112], word_in[112]);
  buf(\oc8051_gm_cxrom_1.word_in [113], word_in[113]);
  buf(\oc8051_gm_cxrom_1.word_in [114], word_in[114]);
  buf(\oc8051_gm_cxrom_1.word_in [115], word_in[115]);
  buf(\oc8051_gm_cxrom_1.word_in [116], word_in[116]);
  buf(\oc8051_gm_cxrom_1.word_in [117], word_in[117]);
  buf(\oc8051_gm_cxrom_1.word_in [118], word_in[118]);
  buf(\oc8051_gm_cxrom_1.word_in [119], word_in[119]);
  buf(\oc8051_gm_cxrom_1.word_in [120], word_in[120]);
  buf(\oc8051_gm_cxrom_1.word_in [121], word_in[121]);
  buf(\oc8051_gm_cxrom_1.word_in [122], word_in[122]);
  buf(\oc8051_gm_cxrom_1.word_in [123], word_in[123]);
  buf(\oc8051_gm_cxrom_1.word_in [124], word_in[124]);
  buf(\oc8051_gm_cxrom_1.word_in [125], word_in[125]);
  buf(\oc8051_gm_cxrom_1.word_in [126], word_in[126]);
  buf(\oc8051_gm_cxrom_1.word_in [127], word_in[127]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [0], \oc8051_golden_model_1.PC [0]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [1], \oc8051_golden_model_1.PC [1]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [2], \oc8051_golden_model_1.PC [2]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [3], \oc8051_golden_model_1.PC [3]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [4], \oc8051_golden_model_1.PC [4]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [5], \oc8051_golden_model_1.PC [5]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [6], \oc8051_golden_model_1.PC [6]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [7], \oc8051_golden_model_1.PC [7]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [8], \oc8051_golden_model_1.PC [8]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [9], \oc8051_golden_model_1.PC [9]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [10], \oc8051_golden_model_1.PC [10]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [11], \oc8051_golden_model_1.PC [11]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [12], \oc8051_golden_model_1.PC [12]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [13], \oc8051_golden_model_1.PC [13]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [14], \oc8051_golden_model_1.PC [14]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [15], \oc8051_golden_model_1.PC [15]);
  buf(\oc8051_gm_cxrom_1.rd_addr_2 [0], RD_ROM_2_ABSTR_ADDR[0]);
  buf(\oc8051_gm_cxrom_1.rd_addr_2 [1], RD_ROM_2_ABSTR_ADDR[1]);
  buf(\oc8051_gm_cxrom_1.rd_addr_2 [2], RD_ROM_2_ABSTR_ADDR[2]);
  buf(\oc8051_gm_cxrom_1.rd_addr_2 [3], RD_ROM_2_ABSTR_ADDR[3]);
  buf(\oc8051_gm_cxrom_1.rd_addr_2 [4], RD_ROM_2_ABSTR_ADDR[4]);
  buf(\oc8051_gm_cxrom_1.rd_addr_2 [5], RD_ROM_2_ABSTR_ADDR[5]);
  buf(\oc8051_gm_cxrom_1.rd_addr_2 [6], RD_ROM_2_ABSTR_ADDR[6]);
  buf(\oc8051_gm_cxrom_1.rd_addr_2 [7], RD_ROM_2_ABSTR_ADDR[7]);
  buf(\oc8051_gm_cxrom_1.rd_addr_2 [8], RD_ROM_2_ABSTR_ADDR[8]);
  buf(\oc8051_gm_cxrom_1.rd_addr_2 [9], RD_ROM_2_ABSTR_ADDR[9]);
  buf(\oc8051_gm_cxrom_1.rd_addr_2 [10], RD_ROM_2_ABSTR_ADDR[10]);
  buf(\oc8051_gm_cxrom_1.rd_addr_2 [11], RD_ROM_2_ABSTR_ADDR[11]);
  buf(\oc8051_gm_cxrom_1.rd_addr_2 [12], RD_ROM_2_ABSTR_ADDR[12]);
  buf(\oc8051_gm_cxrom_1.rd_addr_2 [13], RD_ROM_2_ABSTR_ADDR[13]);
  buf(\oc8051_gm_cxrom_1.rd_addr_2 [14], RD_ROM_2_ABSTR_ADDR[14]);
  buf(\oc8051_gm_cxrom_1.rd_addr_2 [15], RD_ROM_2_ABSTR_ADDR[15]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [0], \oc8051_golden_model_1.PC [0]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [1], \oc8051_golden_model_1.PC [1]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [2], \oc8051_golden_model_1.PC [2]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [3], \oc8051_golden_model_1.PC [3]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [4], \oc8051_golden_model_1.PC [4]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [5], \oc8051_golden_model_1.PC [5]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [6], \oc8051_golden_model_1.PC [6]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [7], \oc8051_golden_model_1.PC [7]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [8], \oc8051_golden_model_1.PC [8]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [9], \oc8051_golden_model_1.PC [9]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [10], \oc8051_golden_model_1.PC [10]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [11], \oc8051_golden_model_1.PC [11]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [12], \oc8051_golden_model_1.PC [12]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [13], \oc8051_golden_model_1.PC [13]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [14], \oc8051_golden_model_1.PC [14]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [15], \oc8051_golden_model_1.PC [15]);
  buf(\oc8051_golden_model_1.RD_ROM_2_ADDR [0], RD_ROM_2_ABSTR_ADDR[0]);
  buf(\oc8051_golden_model_1.RD_ROM_2_ADDR [1], RD_ROM_2_ABSTR_ADDR[1]);
  buf(\oc8051_golden_model_1.RD_ROM_2_ADDR [2], RD_ROM_2_ABSTR_ADDR[2]);
  buf(\oc8051_golden_model_1.RD_ROM_2_ADDR [3], RD_ROM_2_ABSTR_ADDR[3]);
  buf(\oc8051_golden_model_1.RD_ROM_2_ADDR [4], RD_ROM_2_ABSTR_ADDR[4]);
  buf(\oc8051_golden_model_1.RD_ROM_2_ADDR [5], RD_ROM_2_ABSTR_ADDR[5]);
  buf(\oc8051_golden_model_1.RD_ROM_2_ADDR [6], RD_ROM_2_ABSTR_ADDR[6]);
  buf(\oc8051_golden_model_1.RD_ROM_2_ADDR [7], RD_ROM_2_ABSTR_ADDR[7]);
  buf(\oc8051_golden_model_1.RD_ROM_2_ADDR [8], RD_ROM_2_ABSTR_ADDR[8]);
  buf(\oc8051_golden_model_1.RD_ROM_2_ADDR [9], RD_ROM_2_ABSTR_ADDR[9]);
  buf(\oc8051_golden_model_1.RD_ROM_2_ADDR [10], RD_ROM_2_ABSTR_ADDR[10]);
  buf(\oc8051_golden_model_1.RD_ROM_2_ADDR [11], RD_ROM_2_ABSTR_ADDR[11]);
  buf(\oc8051_golden_model_1.RD_ROM_2_ADDR [12], RD_ROM_2_ABSTR_ADDR[12]);
  buf(\oc8051_golden_model_1.RD_ROM_2_ADDR [13], RD_ROM_2_ABSTR_ADDR[13]);
  buf(\oc8051_golden_model_1.RD_ROM_2_ADDR [14], RD_ROM_2_ABSTR_ADDR[14]);
  buf(\oc8051_golden_model_1.RD_ROM_2_ADDR [15], RD_ROM_2_ABSTR_ADDR[15]);
  buf(\oc8051_golden_model_1.SBUF_next [0], \oc8051_golden_model_1.SBUF [0]);
  buf(\oc8051_golden_model_1.SBUF_next [1], \oc8051_golden_model_1.SBUF [1]);
  buf(\oc8051_golden_model_1.SBUF_next [2], \oc8051_golden_model_1.SBUF [2]);
  buf(\oc8051_golden_model_1.SBUF_next [3], \oc8051_golden_model_1.SBUF [3]);
  buf(\oc8051_golden_model_1.SBUF_next [4], \oc8051_golden_model_1.SBUF [4]);
  buf(\oc8051_golden_model_1.SBUF_next [5], \oc8051_golden_model_1.SBUF [5]);
  buf(\oc8051_golden_model_1.SBUF_next [6], \oc8051_golden_model_1.SBUF [6]);
  buf(\oc8051_golden_model_1.SBUF_next [7], \oc8051_golden_model_1.SBUF [7]);
  buf(\oc8051_golden_model_1.SCON_next [0], \oc8051_golden_model_1.SCON [0]);
  buf(\oc8051_golden_model_1.SCON_next [1], \oc8051_golden_model_1.SCON [1]);
  buf(\oc8051_golden_model_1.SCON_next [2], \oc8051_golden_model_1.SCON [2]);
  buf(\oc8051_golden_model_1.SCON_next [3], \oc8051_golden_model_1.SCON [3]);
  buf(\oc8051_golden_model_1.SCON_next [4], \oc8051_golden_model_1.SCON [4]);
  buf(\oc8051_golden_model_1.SCON_next [5], \oc8051_golden_model_1.SCON [5]);
  buf(\oc8051_golden_model_1.SCON_next [6], \oc8051_golden_model_1.SCON [6]);
  buf(\oc8051_golden_model_1.SCON_next [7], \oc8051_golden_model_1.SCON [7]);
  buf(\oc8051_golden_model_1.PCON_next [0], \oc8051_golden_model_1.PCON [0]);
  buf(\oc8051_golden_model_1.PCON_next [1], \oc8051_golden_model_1.PCON [1]);
  buf(\oc8051_golden_model_1.PCON_next [2], \oc8051_golden_model_1.PCON [2]);
  buf(\oc8051_golden_model_1.PCON_next [3], \oc8051_golden_model_1.PCON [3]);
  buf(\oc8051_golden_model_1.PCON_next [4], \oc8051_golden_model_1.PCON [4]);
  buf(\oc8051_golden_model_1.PCON_next [5], \oc8051_golden_model_1.PCON [5]);
  buf(\oc8051_golden_model_1.PCON_next [6], \oc8051_golden_model_1.PCON [6]);
  buf(\oc8051_golden_model_1.PCON_next [7], \oc8051_golden_model_1.PCON [7]);
  buf(\oc8051_golden_model_1.TCON_next [0], \oc8051_golden_model_1.TCON [0]);
  buf(\oc8051_golden_model_1.TCON_next [1], \oc8051_golden_model_1.TCON [1]);
  buf(\oc8051_golden_model_1.TCON_next [2], \oc8051_golden_model_1.TCON [2]);
  buf(\oc8051_golden_model_1.TCON_next [3], \oc8051_golden_model_1.TCON [3]);
  buf(\oc8051_golden_model_1.TCON_next [4], \oc8051_golden_model_1.TCON [4]);
  buf(\oc8051_golden_model_1.TCON_next [5], \oc8051_golden_model_1.TCON [5]);
  buf(\oc8051_golden_model_1.TCON_next [6], \oc8051_golden_model_1.TCON [6]);
  buf(\oc8051_golden_model_1.TCON_next [7], \oc8051_golden_model_1.TCON [7]);
  buf(\oc8051_golden_model_1.TL0_next [0], \oc8051_golden_model_1.TL0 [0]);
  buf(\oc8051_golden_model_1.TL0_next [1], \oc8051_golden_model_1.TL0 [1]);
  buf(\oc8051_golden_model_1.TL0_next [2], \oc8051_golden_model_1.TL0 [2]);
  buf(\oc8051_golden_model_1.TL0_next [3], \oc8051_golden_model_1.TL0 [3]);
  buf(\oc8051_golden_model_1.TL0_next [4], \oc8051_golden_model_1.TL0 [4]);
  buf(\oc8051_golden_model_1.TL0_next [5], \oc8051_golden_model_1.TL0 [5]);
  buf(\oc8051_golden_model_1.TL0_next [6], \oc8051_golden_model_1.TL0 [6]);
  buf(\oc8051_golden_model_1.TL0_next [7], \oc8051_golden_model_1.TL0 [7]);
  buf(\oc8051_golden_model_1.TL1_next [0], \oc8051_golden_model_1.TL1 [0]);
  buf(\oc8051_golden_model_1.TL1_next [1], \oc8051_golden_model_1.TL1 [1]);
  buf(\oc8051_golden_model_1.TL1_next [2], \oc8051_golden_model_1.TL1 [2]);
  buf(\oc8051_golden_model_1.TL1_next [3], \oc8051_golden_model_1.TL1 [3]);
  buf(\oc8051_golden_model_1.TL1_next [4], \oc8051_golden_model_1.TL1 [4]);
  buf(\oc8051_golden_model_1.TL1_next [5], \oc8051_golden_model_1.TL1 [5]);
  buf(\oc8051_golden_model_1.TL1_next [6], \oc8051_golden_model_1.TL1 [6]);
  buf(\oc8051_golden_model_1.TL1_next [7], \oc8051_golden_model_1.TL1 [7]);
  buf(\oc8051_golden_model_1.TH0_next [0], \oc8051_golden_model_1.TH0 [0]);
  buf(\oc8051_golden_model_1.TH0_next [1], \oc8051_golden_model_1.TH0 [1]);
  buf(\oc8051_golden_model_1.TH0_next [2], \oc8051_golden_model_1.TH0 [2]);
  buf(\oc8051_golden_model_1.TH0_next [3], \oc8051_golden_model_1.TH0 [3]);
  buf(\oc8051_golden_model_1.TH0_next [4], \oc8051_golden_model_1.TH0 [4]);
  buf(\oc8051_golden_model_1.TH0_next [5], \oc8051_golden_model_1.TH0 [5]);
  buf(\oc8051_golden_model_1.TH0_next [6], \oc8051_golden_model_1.TH0 [6]);
  buf(\oc8051_golden_model_1.TH0_next [7], \oc8051_golden_model_1.TH0 [7]);
  buf(\oc8051_golden_model_1.TH1_next [0], \oc8051_golden_model_1.TH1 [0]);
  buf(\oc8051_golden_model_1.TH1_next [1], \oc8051_golden_model_1.TH1 [1]);
  buf(\oc8051_golden_model_1.TH1_next [2], \oc8051_golden_model_1.TH1 [2]);
  buf(\oc8051_golden_model_1.TH1_next [3], \oc8051_golden_model_1.TH1 [3]);
  buf(\oc8051_golden_model_1.TH1_next [4], \oc8051_golden_model_1.TH1 [4]);
  buf(\oc8051_golden_model_1.TH1_next [5], \oc8051_golden_model_1.TH1 [5]);
  buf(\oc8051_golden_model_1.TH1_next [6], \oc8051_golden_model_1.TH1 [6]);
  buf(\oc8051_golden_model_1.TH1_next [7], \oc8051_golden_model_1.TH1 [7]);
  buf(\oc8051_golden_model_1.TMOD_next [0], \oc8051_golden_model_1.TMOD [0]);
  buf(\oc8051_golden_model_1.TMOD_next [1], \oc8051_golden_model_1.TMOD [1]);
  buf(\oc8051_golden_model_1.TMOD_next [2], \oc8051_golden_model_1.TMOD [2]);
  buf(\oc8051_golden_model_1.TMOD_next [3], \oc8051_golden_model_1.TMOD [3]);
  buf(\oc8051_golden_model_1.TMOD_next [4], \oc8051_golden_model_1.TMOD [4]);
  buf(\oc8051_golden_model_1.TMOD_next [5], \oc8051_golden_model_1.TMOD [5]);
  buf(\oc8051_golden_model_1.TMOD_next [6], \oc8051_golden_model_1.TMOD [6]);
  buf(\oc8051_golden_model_1.TMOD_next [7], \oc8051_golden_model_1.TMOD [7]);
  buf(\oc8051_golden_model_1.IE_next [0], \oc8051_golden_model_1.IE [0]);
  buf(\oc8051_golden_model_1.IE_next [1], \oc8051_golden_model_1.IE [1]);
  buf(\oc8051_golden_model_1.IE_next [2], \oc8051_golden_model_1.IE [2]);
  buf(\oc8051_golden_model_1.IE_next [3], \oc8051_golden_model_1.IE [3]);
  buf(\oc8051_golden_model_1.IE_next [4], \oc8051_golden_model_1.IE [4]);
  buf(\oc8051_golden_model_1.IE_next [5], \oc8051_golden_model_1.IE [5]);
  buf(\oc8051_golden_model_1.IE_next [6], \oc8051_golden_model_1.IE [6]);
  buf(\oc8051_golden_model_1.IE_next [7], \oc8051_golden_model_1.IE [7]);
  buf(\oc8051_golden_model_1.IP_next [0], \oc8051_golden_model_1.IP [0]);
  buf(\oc8051_golden_model_1.IP_next [1], \oc8051_golden_model_1.IP [1]);
  buf(\oc8051_golden_model_1.IP_next [2], \oc8051_golden_model_1.IP [2]);
  buf(\oc8051_golden_model_1.IP_next [3], \oc8051_golden_model_1.IP [3]);
  buf(\oc8051_golden_model_1.IP_next [4], \oc8051_golden_model_1.IP [4]);
  buf(\oc8051_golden_model_1.IP_next [5], \oc8051_golden_model_1.IP [5]);
  buf(\oc8051_golden_model_1.IP_next [6], \oc8051_golden_model_1.IP [6]);
  buf(\oc8051_golden_model_1.IP_next [7], \oc8051_golden_model_1.IP [7]);
  buf(\oc8051_golden_model_1.clk , clk);
  buf(\oc8051_golden_model_1.rst , rst);
  buf(\oc8051_golden_model_1.XRAM_DATA_IN [0], xram_data_in_reg[0]);
  buf(\oc8051_golden_model_1.XRAM_DATA_IN [1], xram_data_in_reg[1]);
  buf(\oc8051_golden_model_1.XRAM_DATA_IN [2], xram_data_in_reg[2]);
  buf(\oc8051_golden_model_1.XRAM_DATA_IN [3], xram_data_in_reg[3]);
  buf(\oc8051_golden_model_1.XRAM_DATA_IN [4], xram_data_in_reg[4]);
  buf(\oc8051_golden_model_1.XRAM_DATA_IN [5], xram_data_in_reg[5]);
  buf(\oc8051_golden_model_1.XRAM_DATA_IN [6], xram_data_in_reg[6]);
  buf(\oc8051_golden_model_1.XRAM_DATA_IN [7], xram_data_in_reg[7]);
  buf(\oc8051_golden_model_1.RD_IRAM_0_ABSTR_ADDR [0], RD_IRAM_0_ABSTR_ADDR[0]);
  buf(\oc8051_golden_model_1.RD_IRAM_0_ABSTR_ADDR [1], RD_IRAM_0_ABSTR_ADDR[1]);
  buf(\oc8051_golden_model_1.RD_IRAM_0_ABSTR_ADDR [2], RD_IRAM_0_ABSTR_ADDR[2]);
  buf(\oc8051_golden_model_1.RD_IRAM_0_ABSTR_ADDR [3], RD_IRAM_0_ABSTR_ADDR[3]);
  buf(\oc8051_golden_model_1.RD_IRAM_0_ABSTR_ADDR [4], RD_IRAM_0_ABSTR_ADDR[4]);
  buf(\oc8051_golden_model_1.RD_IRAM_0_ABSTR_ADDR [5], RD_IRAM_0_ABSTR_ADDR[5]);
  buf(\oc8051_golden_model_1.RD_IRAM_0_ABSTR_ADDR [6], RD_IRAM_0_ABSTR_ADDR[6]);
  buf(\oc8051_golden_model_1.RD_IRAM_0_ABSTR_ADDR [7], RD_IRAM_0_ABSTR_ADDR[7]);
  buf(\oc8051_golden_model_1.RD_IRAM_1_ABSTR_ADDR [0], RD_IRAM_1_ABSTR_ADDR[0]);
  buf(\oc8051_golden_model_1.RD_IRAM_1_ABSTR_ADDR [1], RD_IRAM_1_ABSTR_ADDR[1]);
  buf(\oc8051_golden_model_1.RD_IRAM_1_ABSTR_ADDR [2], RD_IRAM_1_ABSTR_ADDR[2]);
  buf(\oc8051_golden_model_1.RD_IRAM_1_ABSTR_ADDR [3], RD_IRAM_1_ABSTR_ADDR[3]);
  buf(\oc8051_golden_model_1.RD_IRAM_1_ABSTR_ADDR [4], RD_IRAM_1_ABSTR_ADDR[4]);
  buf(\oc8051_golden_model_1.RD_IRAM_1_ABSTR_ADDR [5], RD_IRAM_1_ABSTR_ADDR[5]);
  buf(\oc8051_golden_model_1.RD_IRAM_1_ABSTR_ADDR [6], RD_IRAM_1_ABSTR_ADDR[6]);
  buf(\oc8051_golden_model_1.RD_IRAM_1_ABSTR_ADDR [7], RD_IRAM_1_ABSTR_ADDR[7]);
  buf(\oc8051_golden_model_1.RD_ROM_1_ABSTR_ADDR [0], RD_ROM_1_ABSTR_ADDR[0]);
  buf(\oc8051_golden_model_1.RD_ROM_1_ABSTR_ADDR [1], RD_ROM_1_ABSTR_ADDR[1]);
  buf(\oc8051_golden_model_1.RD_ROM_1_ABSTR_ADDR [2], RD_ROM_1_ABSTR_ADDR[2]);
  buf(\oc8051_golden_model_1.RD_ROM_1_ABSTR_ADDR [3], RD_ROM_1_ABSTR_ADDR[3]);
  buf(\oc8051_golden_model_1.RD_ROM_1_ABSTR_ADDR [4], RD_ROM_1_ABSTR_ADDR[4]);
  buf(\oc8051_golden_model_1.RD_ROM_1_ABSTR_ADDR [5], RD_ROM_1_ABSTR_ADDR[5]);
  buf(\oc8051_golden_model_1.RD_ROM_1_ABSTR_ADDR [6], RD_ROM_1_ABSTR_ADDR[6]);
  buf(\oc8051_golden_model_1.RD_ROM_1_ABSTR_ADDR [7], RD_ROM_1_ABSTR_ADDR[7]);
  buf(\oc8051_golden_model_1.RD_ROM_1_ABSTR_ADDR [8], RD_ROM_1_ABSTR_ADDR[8]);
  buf(\oc8051_golden_model_1.RD_ROM_1_ABSTR_ADDR [9], RD_ROM_1_ABSTR_ADDR[9]);
  buf(\oc8051_golden_model_1.RD_ROM_1_ABSTR_ADDR [10], RD_ROM_1_ABSTR_ADDR[10]);
  buf(\oc8051_golden_model_1.RD_ROM_1_ABSTR_ADDR [11], RD_ROM_1_ABSTR_ADDR[11]);
  buf(\oc8051_golden_model_1.RD_ROM_1_ABSTR_ADDR [12], RD_ROM_1_ABSTR_ADDR[12]);
  buf(\oc8051_golden_model_1.RD_ROM_1_ABSTR_ADDR [13], RD_ROM_1_ABSTR_ADDR[13]);
  buf(\oc8051_golden_model_1.RD_ROM_1_ABSTR_ADDR [14], RD_ROM_1_ABSTR_ADDR[14]);
  buf(\oc8051_golden_model_1.RD_ROM_1_ABSTR_ADDR [15], RD_ROM_1_ABSTR_ADDR[15]);
  buf(\oc8051_golden_model_1.RD_ROM_2_ABSTR_ADDR [0], RD_ROM_2_ABSTR_ADDR[0]);
  buf(\oc8051_golden_model_1.RD_ROM_2_ABSTR_ADDR [1], RD_ROM_2_ABSTR_ADDR[1]);
  buf(\oc8051_golden_model_1.RD_ROM_2_ABSTR_ADDR [2], RD_ROM_2_ABSTR_ADDR[2]);
  buf(\oc8051_golden_model_1.RD_ROM_2_ABSTR_ADDR [3], RD_ROM_2_ABSTR_ADDR[3]);
  buf(\oc8051_golden_model_1.RD_ROM_2_ABSTR_ADDR [4], RD_ROM_2_ABSTR_ADDR[4]);
  buf(\oc8051_golden_model_1.RD_ROM_2_ABSTR_ADDR [5], RD_ROM_2_ABSTR_ADDR[5]);
  buf(\oc8051_golden_model_1.RD_ROM_2_ABSTR_ADDR [6], RD_ROM_2_ABSTR_ADDR[6]);
  buf(\oc8051_golden_model_1.RD_ROM_2_ABSTR_ADDR [7], RD_ROM_2_ABSTR_ADDR[7]);
  buf(\oc8051_golden_model_1.RD_ROM_2_ABSTR_ADDR [8], RD_ROM_2_ABSTR_ADDR[8]);
  buf(\oc8051_golden_model_1.RD_ROM_2_ABSTR_ADDR [9], RD_ROM_2_ABSTR_ADDR[9]);
  buf(\oc8051_golden_model_1.RD_ROM_2_ABSTR_ADDR [10], RD_ROM_2_ABSTR_ADDR[10]);
  buf(\oc8051_golden_model_1.RD_ROM_2_ABSTR_ADDR [11], RD_ROM_2_ABSTR_ADDR[11]);
  buf(\oc8051_golden_model_1.RD_ROM_2_ABSTR_ADDR [12], RD_ROM_2_ABSTR_ADDR[12]);
  buf(\oc8051_golden_model_1.RD_ROM_2_ABSTR_ADDR [13], RD_ROM_2_ABSTR_ADDR[13]);
  buf(\oc8051_golden_model_1.RD_ROM_2_ABSTR_ADDR [14], RD_ROM_2_ABSTR_ADDR[14]);
  buf(\oc8051_golden_model_1.RD_ROM_2_ABSTR_ADDR [15], RD_ROM_2_ABSTR_ADDR[15]);
  buf(\oc8051_golden_model_1.ACC_abstr [0], ACC_abstr[0]);
  buf(\oc8051_golden_model_1.ACC_abstr [1], ACC_abstr[1]);
  buf(\oc8051_golden_model_1.ACC_abstr [2], ACC_abstr[2]);
  buf(\oc8051_golden_model_1.ACC_abstr [3], ACC_abstr[3]);
  buf(\oc8051_golden_model_1.ACC_abstr [4], ACC_abstr[4]);
  buf(\oc8051_golden_model_1.ACC_abstr [5], ACC_abstr[5]);
  buf(\oc8051_golden_model_1.ACC_abstr [6], ACC_abstr[6]);
  buf(\oc8051_golden_model_1.ACC_abstr [7], ACC_abstr[7]);
  buf(\oc8051_golden_model_1.P2_abstr [0], P2_abstr[0]);
  buf(\oc8051_golden_model_1.P2_abstr [1], P2_abstr[1]);
  buf(\oc8051_golden_model_1.P2_abstr [2], P2_abstr[2]);
  buf(\oc8051_golden_model_1.P2_abstr [3], P2_abstr[3]);
  buf(\oc8051_golden_model_1.P2_abstr [4], P2_abstr[4]);
  buf(\oc8051_golden_model_1.P2_abstr [5], P2_abstr[5]);
  buf(\oc8051_golden_model_1.P2_abstr [6], P2_abstr[6]);
  buf(\oc8051_golden_model_1.P2_abstr [7], P2_abstr[7]);
  buf(\oc8051_golden_model_1.P0_abstr [0], P0_abstr[0]);
  buf(\oc8051_golden_model_1.P0_abstr [1], P0_abstr[1]);
  buf(\oc8051_golden_model_1.P0_abstr [2], P0_abstr[2]);
  buf(\oc8051_golden_model_1.P0_abstr [3], P0_abstr[3]);
  buf(\oc8051_golden_model_1.P0_abstr [4], P0_abstr[4]);
  buf(\oc8051_golden_model_1.P0_abstr [5], P0_abstr[5]);
  buf(\oc8051_golden_model_1.P0_abstr [6], P0_abstr[6]);
  buf(\oc8051_golden_model_1.P0_abstr [7], P0_abstr[7]);
  buf(\oc8051_golden_model_1.B_abstr [0], B_abstr[0]);
  buf(\oc8051_golden_model_1.B_abstr [1], B_abstr[1]);
  buf(\oc8051_golden_model_1.B_abstr [2], B_abstr[2]);
  buf(\oc8051_golden_model_1.B_abstr [3], B_abstr[3]);
  buf(\oc8051_golden_model_1.B_abstr [4], B_abstr[4]);
  buf(\oc8051_golden_model_1.B_abstr [5], B_abstr[5]);
  buf(\oc8051_golden_model_1.B_abstr [6], B_abstr[6]);
  buf(\oc8051_golden_model_1.B_abstr [7], B_abstr[7]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_abstr [0], XRAM_ADDR_abstr[0]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_abstr [1], XRAM_ADDR_abstr[1]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_abstr [2], XRAM_ADDR_abstr[2]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_abstr [3], XRAM_ADDR_abstr[3]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_abstr [4], XRAM_ADDR_abstr[4]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_abstr [5], XRAM_ADDR_abstr[5]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_abstr [6], XRAM_ADDR_abstr[6]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_abstr [7], XRAM_ADDR_abstr[7]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_abstr [8], XRAM_ADDR_abstr[8]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_abstr [9], XRAM_ADDR_abstr[9]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_abstr [10], XRAM_ADDR_abstr[10]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_abstr [11], XRAM_ADDR_abstr[11]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_abstr [12], XRAM_ADDR_abstr[12]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_abstr [13], XRAM_ADDR_abstr[13]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_abstr [14], XRAM_ADDR_abstr[14]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_abstr [15], XRAM_ADDR_abstr[15]);
  buf(\oc8051_golden_model_1.P3_abstr [0], P3_abstr[0]);
  buf(\oc8051_golden_model_1.P3_abstr [1], P3_abstr[1]);
  buf(\oc8051_golden_model_1.P3_abstr [2], P3_abstr[2]);
  buf(\oc8051_golden_model_1.P3_abstr [3], P3_abstr[3]);
  buf(\oc8051_golden_model_1.P3_abstr [4], P3_abstr[4]);
  buf(\oc8051_golden_model_1.P3_abstr [5], P3_abstr[5]);
  buf(\oc8051_golden_model_1.P3_abstr [6], P3_abstr[6]);
  buf(\oc8051_golden_model_1.P3_abstr [7], P3_abstr[7]);
  buf(\oc8051_golden_model_1.SP_abstr [0], SP_abstr[0]);
  buf(\oc8051_golden_model_1.SP_abstr [1], SP_abstr[1]);
  buf(\oc8051_golden_model_1.SP_abstr [2], SP_abstr[2]);
  buf(\oc8051_golden_model_1.SP_abstr [3], SP_abstr[3]);
  buf(\oc8051_golden_model_1.SP_abstr [4], SP_abstr[4]);
  buf(\oc8051_golden_model_1.SP_abstr [5], SP_abstr[5]);
  buf(\oc8051_golden_model_1.SP_abstr [6], SP_abstr[6]);
  buf(\oc8051_golden_model_1.SP_abstr [7], SP_abstr[7]);
  buf(\oc8051_golden_model_1.PC_abstr [0], PC_abstr[0]);
  buf(\oc8051_golden_model_1.PC_abstr [1], PC_abstr[1]);
  buf(\oc8051_golden_model_1.PC_abstr [2], PC_abstr[2]);
  buf(\oc8051_golden_model_1.PC_abstr [3], PC_abstr[3]);
  buf(\oc8051_golden_model_1.PC_abstr [4], PC_abstr[4]);
  buf(\oc8051_golden_model_1.PC_abstr [5], PC_abstr[5]);
  buf(\oc8051_golden_model_1.PC_abstr [6], PC_abstr[6]);
  buf(\oc8051_golden_model_1.PC_abstr [7], PC_abstr[7]);
  buf(\oc8051_golden_model_1.PC_abstr [8], PC_abstr[8]);
  buf(\oc8051_golden_model_1.PC_abstr [9], PC_abstr[9]);
  buf(\oc8051_golden_model_1.PC_abstr [10], PC_abstr[10]);
  buf(\oc8051_golden_model_1.PC_abstr [11], PC_abstr[11]);
  buf(\oc8051_golden_model_1.PC_abstr [12], PC_abstr[12]);
  buf(\oc8051_golden_model_1.PC_abstr [13], PC_abstr[13]);
  buf(\oc8051_golden_model_1.PC_abstr [14], PC_abstr[14]);
  buf(\oc8051_golden_model_1.PC_abstr [15], PC_abstr[15]);
  buf(\oc8051_golden_model_1.P1_abstr [0], P1_abstr[0]);
  buf(\oc8051_golden_model_1.P1_abstr [1], P1_abstr[1]);
  buf(\oc8051_golden_model_1.P1_abstr [2], P1_abstr[2]);
  buf(\oc8051_golden_model_1.P1_abstr [3], P1_abstr[3]);
  buf(\oc8051_golden_model_1.P1_abstr [4], P1_abstr[4]);
  buf(\oc8051_golden_model_1.P1_abstr [5], P1_abstr[5]);
  buf(\oc8051_golden_model_1.P1_abstr [6], P1_abstr[6]);
  buf(\oc8051_golden_model_1.P1_abstr [7], P1_abstr[7]);
  buf(\oc8051_golden_model_1.XRAM_DATA_OUT_abstr [0], XRAM_DATA_OUT_abstr[0]);
  buf(\oc8051_golden_model_1.XRAM_DATA_OUT_abstr [1], XRAM_DATA_OUT_abstr[1]);
  buf(\oc8051_golden_model_1.XRAM_DATA_OUT_abstr [2], XRAM_DATA_OUT_abstr[2]);
  buf(\oc8051_golden_model_1.XRAM_DATA_OUT_abstr [3], XRAM_DATA_OUT_abstr[3]);
  buf(\oc8051_golden_model_1.XRAM_DATA_OUT_abstr [4], XRAM_DATA_OUT_abstr[4]);
  buf(\oc8051_golden_model_1.XRAM_DATA_OUT_abstr [5], XRAM_DATA_OUT_abstr[5]);
  buf(\oc8051_golden_model_1.XRAM_DATA_OUT_abstr [6], XRAM_DATA_OUT_abstr[6]);
  buf(\oc8051_golden_model_1.XRAM_DATA_OUT_abstr [7], XRAM_DATA_OUT_abstr[7]);
  buf(\oc8051_golden_model_1.DPL_abstr [0], DPL_abstr[0]);
  buf(\oc8051_golden_model_1.DPL_abstr [1], DPL_abstr[1]);
  buf(\oc8051_golden_model_1.DPL_abstr [2], DPL_abstr[2]);
  buf(\oc8051_golden_model_1.DPL_abstr [3], DPL_abstr[3]);
  buf(\oc8051_golden_model_1.DPL_abstr [4], DPL_abstr[4]);
  buf(\oc8051_golden_model_1.DPL_abstr [5], DPL_abstr[5]);
  buf(\oc8051_golden_model_1.DPL_abstr [6], DPL_abstr[6]);
  buf(\oc8051_golden_model_1.DPL_abstr [7], DPL_abstr[7]);
  buf(\oc8051_golden_model_1.PSW_abstr [0], PSW_abstr[0]);
  buf(\oc8051_golden_model_1.PSW_abstr [1], PSW_abstr[1]);
  buf(\oc8051_golden_model_1.PSW_abstr [2], PSW_abstr[2]);
  buf(\oc8051_golden_model_1.PSW_abstr [3], PSW_abstr[3]);
  buf(\oc8051_golden_model_1.PSW_abstr [4], PSW_abstr[4]);
  buf(\oc8051_golden_model_1.PSW_abstr [5], PSW_abstr[5]);
  buf(\oc8051_golden_model_1.PSW_abstr [6], PSW_abstr[6]);
  buf(\oc8051_golden_model_1.PSW_abstr [7], PSW_abstr[7]);
  buf(\oc8051_golden_model_1.DPH_abstr [0], DPH_abstr[0]);
  buf(\oc8051_golden_model_1.DPH_abstr [1], DPH_abstr[1]);
  buf(\oc8051_golden_model_1.DPH_abstr [2], DPH_abstr[2]);
  buf(\oc8051_golden_model_1.DPH_abstr [3], DPH_abstr[3]);
  buf(\oc8051_golden_model_1.DPH_abstr [4], DPH_abstr[4]);
  buf(\oc8051_golden_model_1.DPH_abstr [5], DPH_abstr[5]);
  buf(\oc8051_golden_model_1.DPH_abstr [6], DPH_abstr[6]);
  buf(\oc8051_golden_model_1.DPH_abstr [7], DPH_abstr[7]);
  buf(\oc8051_golden_model_1.WR_COND_ABSTR_IRAM_0 , WR_COND_ABSTR_IRAM_0);
  buf(\oc8051_golden_model_1.WR_ADDR_ABSTR_IRAM_0 [0], WR_ADDR_ABSTR_IRAM_0[0]);
  buf(\oc8051_golden_model_1.WR_ADDR_ABSTR_IRAM_0 [1], WR_ADDR_ABSTR_IRAM_0[1]);
  buf(\oc8051_golden_model_1.WR_ADDR_ABSTR_IRAM_0 [2], WR_ADDR_ABSTR_IRAM_0[2]);
  buf(\oc8051_golden_model_1.WR_ADDR_ABSTR_IRAM_0 [3], WR_ADDR_ABSTR_IRAM_0[3]);
  buf(\oc8051_golden_model_1.WR_DATA_ABSTR_IRAM_0 [0], WR_DATA_ABSTR_IRAM_0[0]);
  buf(\oc8051_golden_model_1.WR_DATA_ABSTR_IRAM_0 [1], WR_DATA_ABSTR_IRAM_0[1]);
  buf(\oc8051_golden_model_1.WR_DATA_ABSTR_IRAM_0 [2], WR_DATA_ABSTR_IRAM_0[2]);
  buf(\oc8051_golden_model_1.WR_DATA_ABSTR_IRAM_0 [3], WR_DATA_ABSTR_IRAM_0[3]);
  buf(\oc8051_golden_model_1.WR_DATA_ABSTR_IRAM_0 [4], WR_DATA_ABSTR_IRAM_0[4]);
  buf(\oc8051_golden_model_1.WR_DATA_ABSTR_IRAM_0 [5], WR_DATA_ABSTR_IRAM_0[5]);
  buf(\oc8051_golden_model_1.WR_DATA_ABSTR_IRAM_0 [6], WR_DATA_ABSTR_IRAM_0[6]);
  buf(\oc8051_golden_model_1.WR_DATA_ABSTR_IRAM_0 [7], WR_DATA_ABSTR_IRAM_0[7]);
  buf(\oc8051_golden_model_1.WR_COND_ABSTR_IRAM_1 , WR_COND_ABSTR_IRAM_1);
  buf(\oc8051_golden_model_1.WR_ADDR_ABSTR_IRAM_1 [0], WR_ADDR_ABSTR_IRAM_1[0]);
  buf(\oc8051_golden_model_1.WR_ADDR_ABSTR_IRAM_1 [1], WR_ADDR_ABSTR_IRAM_1[1]);
  buf(\oc8051_golden_model_1.WR_ADDR_ABSTR_IRAM_1 [2], WR_ADDR_ABSTR_IRAM_1[2]);
  buf(\oc8051_golden_model_1.WR_ADDR_ABSTR_IRAM_1 [3], WR_ADDR_ABSTR_IRAM_1[3]);
  buf(\oc8051_golden_model_1.WR_DATA_ABSTR_IRAM_1 [0], WR_DATA_ABSTR_IRAM_1[0]);
  buf(\oc8051_golden_model_1.WR_DATA_ABSTR_IRAM_1 [1], WR_DATA_ABSTR_IRAM_1[1]);
  buf(\oc8051_golden_model_1.WR_DATA_ABSTR_IRAM_1 [2], WR_DATA_ABSTR_IRAM_1[2]);
  buf(\oc8051_golden_model_1.WR_DATA_ABSTR_IRAM_1 [3], WR_DATA_ABSTR_IRAM_1[3]);
  buf(\oc8051_golden_model_1.WR_DATA_ABSTR_IRAM_1 [4], WR_DATA_ABSTR_IRAM_1[4]);
  buf(\oc8051_golden_model_1.WR_DATA_ABSTR_IRAM_1 [5], WR_DATA_ABSTR_IRAM_1[5]);
  buf(\oc8051_golden_model_1.WR_DATA_ABSTR_IRAM_1 [6], WR_DATA_ABSTR_IRAM_1[6]);
  buf(\oc8051_golden_model_1.WR_DATA_ABSTR_IRAM_1 [7], WR_DATA_ABSTR_IRAM_1[7]);
  buf(\oc8051_golden_model_1.RD_IRAM_1_ADDR [0], RD_IRAM_1_ABSTR_ADDR[0]);
  buf(\oc8051_golden_model_1.RD_IRAM_1_ADDR [1], RD_IRAM_1_ABSTR_ADDR[1]);
  buf(\oc8051_golden_model_1.RD_IRAM_1_ADDR [2], RD_IRAM_1_ABSTR_ADDR[2]);
  buf(\oc8051_golden_model_1.RD_IRAM_1_ADDR [3], RD_IRAM_1_ABSTR_ADDR[3]);
  buf(\oc8051_golden_model_1.RD_IRAM_1_ADDR [4], RD_IRAM_1_ABSTR_ADDR[4]);
  buf(\oc8051_golden_model_1.RD_IRAM_1_ADDR [5], RD_IRAM_1_ABSTR_ADDR[5]);
  buf(\oc8051_golden_model_1.RD_IRAM_1_ADDR [6], RD_IRAM_1_ABSTR_ADDR[6]);
  buf(\oc8051_golden_model_1.RD_IRAM_1_ADDR [7], RD_IRAM_1_ABSTR_ADDR[7]);
  buf(\oc8051_golden_model_1.WR_ADDR_1_IRAM [0], WR_ADDR_ABSTR_IRAM_1[0]);
  buf(\oc8051_golden_model_1.WR_ADDR_1_IRAM [1], WR_ADDR_ABSTR_IRAM_1[1]);
  buf(\oc8051_golden_model_1.WR_ADDR_1_IRAM [2], WR_ADDR_ABSTR_IRAM_1[2]);
  buf(\oc8051_golden_model_1.WR_ADDR_1_IRAM [3], WR_ADDR_ABSTR_IRAM_1[3]);
  buf(\oc8051_golden_model_1.WR_DATA_1_IRAM [0], WR_DATA_ABSTR_IRAM_1[0]);
  buf(\oc8051_golden_model_1.WR_DATA_1_IRAM [1], WR_DATA_ABSTR_IRAM_1[1]);
  buf(\oc8051_golden_model_1.WR_DATA_1_IRAM [2], WR_DATA_ABSTR_IRAM_1[2]);
  buf(\oc8051_golden_model_1.WR_DATA_1_IRAM [3], WR_DATA_ABSTR_IRAM_1[3]);
  buf(\oc8051_golden_model_1.WR_DATA_1_IRAM [4], WR_DATA_ABSTR_IRAM_1[4]);
  buf(\oc8051_golden_model_1.WR_DATA_1_IRAM [5], WR_DATA_ABSTR_IRAM_1[5]);
  buf(\oc8051_golden_model_1.WR_DATA_1_IRAM [6], WR_DATA_ABSTR_IRAM_1[6]);
  buf(\oc8051_golden_model_1.WR_DATA_1_IRAM [7], WR_DATA_ABSTR_IRAM_1[7]);
  buf(\oc8051_golden_model_1.n0006 [0], RD_IRAM_1_ABSTR_ADDR[0]);
  buf(\oc8051_golden_model_1.n0006 [1], RD_IRAM_1_ABSTR_ADDR[1]);
  buf(\oc8051_golden_model_1.n0006 [2], RD_IRAM_1_ABSTR_ADDR[2]);
  buf(\oc8051_golden_model_1.n0006 [3], RD_IRAM_1_ABSTR_ADDR[3]);
  buf(\oc8051_golden_model_1.n0288 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n0288 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n0288 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n0288 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n0289 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n0289 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n0289 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n0289 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n0289 [4], \oc8051_golden_model_1.RD_IRAM_1 [4]);
  buf(\oc8051_golden_model_1.n0289 [5], \oc8051_golden_model_1.RD_IRAM_1 [5]);
  buf(\oc8051_golden_model_1.n0289 [6], \oc8051_golden_model_1.RD_IRAM_1 [6]);
  buf(\oc8051_golden_model_1.n0289 [7], \oc8051_golden_model_1.RD_IRAM_1 [7]);
  buf(\oc8051_golden_model_1.n0115 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0115 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0116 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0116 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0116 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0116 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0116 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0116 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0116 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0116 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0117 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0117 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0117 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0117 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0120 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0120 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0120 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0120 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0120 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0120 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0120 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0120 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0121 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0121 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0121 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0121 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0123 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0123 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0123 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0123 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0123 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0123 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0123 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0123 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0124 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0124 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0124 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0124 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0246 , \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n0126 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0126 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0126 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0126 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0126 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0126 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0126 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0126 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0127 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0127 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0127 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0127 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0247 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n0247 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0247 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0247 [3], 1'b0);
  buf(\oc8051_golden_model_1.n0247 [4], 1'b0);
  buf(\oc8051_golden_model_1.n0247 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0247 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0247 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0129 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0129 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0129 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0129 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0129 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0129 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0129 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0129 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0130 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0130 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0130 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0130 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0132 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0132 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0132 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0132 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0132 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0132 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0132 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0132 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0133 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0133 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0133 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0133 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0135 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0135 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0135 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0135 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0135 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0135 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0135 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0135 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0136 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0136 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0136 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0136 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0138 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0138 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0138 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0138 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0138 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0138 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0138 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0138 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0139 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0139 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0139 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0139 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_top_1.wb_rst_i , rst);
  buf(\oc8051_top_1.wb_clk_i , clk);
  buf(\oc8051_top_1.wbd_ack_i , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_top_1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_top_1.pc_log [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_top_1.pc_log [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_top_1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_top_1.pc_log [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_top_1.pc_log [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_top_1.pc_log [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_top_1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_top_1.pc_log [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_top_1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_top_1.pc_log [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_top_1.pc_log [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_top_1.pc_log [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_top_1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_top_1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_top_1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_top_1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_top_1.pc_log_prev [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_top_1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_top_1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_top_1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_top_1.pc_log_prev [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_top_1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_top_1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_top_1.pc_log_prev [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_top_1.pc_log_prev [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_top_1.pc_log_prev [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_top_1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_top_1.pc_log_prev [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_top_1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_top_1.psw [0], psw_impl[0]);
  buf(\oc8051_top_1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.wbd_dat_i [0], xram_data_in_reg[0]);
  buf(\oc8051_top_1.wbd_dat_i [1], xram_data_in_reg[1]);
  buf(\oc8051_top_1.wbd_dat_i [2], xram_data_in_reg[2]);
  buf(\oc8051_top_1.wbd_dat_i [3], xram_data_in_reg[3]);
  buf(\oc8051_top_1.wbd_dat_i [4], xram_data_in_reg[4]);
  buf(\oc8051_top_1.wbd_dat_i [5], xram_data_in_reg[5]);
  buf(\oc8051_top_1.wbd_dat_i [6], xram_data_in_reg[6]);
  buf(\oc8051_top_1.wbd_dat_i [7], xram_data_in_reg[7]);
  buf(\oc8051_top_1.wbd_we_o , \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  buf(\oc8051_top_1.wbd_stb_o , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.wbd_cyc_o , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.wbd_dat_o [0], \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  buf(\oc8051_top_1.wbd_dat_o [1], \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  buf(\oc8051_top_1.wbd_dat_o [2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  buf(\oc8051_top_1.wbd_dat_o [3], \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  buf(\oc8051_top_1.wbd_dat_o [4], \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  buf(\oc8051_top_1.wbd_dat_o [5], \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  buf(\oc8051_top_1.wbd_dat_o [6], \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  buf(\oc8051_top_1.wbd_dat_o [7], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  buf(\oc8051_top_1.wbd_adr_o [0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(\oc8051_top_1.wbd_adr_o [1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(\oc8051_top_1.wbd_adr_o [2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(\oc8051_top_1.wbd_adr_o [3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(\oc8051_top_1.wbd_adr_o [4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(\oc8051_top_1.wbd_adr_o [5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(\oc8051_top_1.wbd_adr_o [6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(\oc8051_top_1.wbd_adr_o [7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(\oc8051_top_1.wbd_adr_o [8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(\oc8051_top_1.wbd_adr_o [9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(\oc8051_top_1.wbd_adr_o [10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(\oc8051_top_1.wbd_adr_o [11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(\oc8051_top_1.wbd_adr_o [12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(\oc8051_top_1.wbd_adr_o [13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(\oc8051_top_1.wbd_adr_o [14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(\oc8051_top_1.wbd_adr_o [15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(\oc8051_top_1.cxrom_data_out [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.cxrom_data_out [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.cxrom_data_out [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.cxrom_data_out [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.cxrom_data_out [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.cxrom_data_out [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.cxrom_data_out [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.cxrom_data_out [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.cxrom_data_out [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.cxrom_data_out [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.cxrom_data_out [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.cxrom_data_out [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.cxrom_data_out [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.cxrom_data_out [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.cxrom_data_out [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.cxrom_data_out [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.cxrom_data_out [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.cxrom_data_out [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.cxrom_data_out [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.cxrom_data_out [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.cxrom_data_out [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.cxrom_data_out [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.cxrom_data_out [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.cxrom_data_out [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.cxrom_data_out [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.cxrom_data_out [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.cxrom_data_out [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.cxrom_data_out [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.cxrom_data_out [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.cxrom_data_out [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.cxrom_data_out [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.cxrom_data_out [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.p0_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.p0_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.p0_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.p0_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.p0_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.p0_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.p0_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.p0_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.p1_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.p1_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.p1_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.p1_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.p1_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.p1_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.p1_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.p1_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.p2_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.p2_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.p2_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.p2_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.p2_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.p2_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.p2_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.p2_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.p3_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.p3_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.p3_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.p3_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.p3_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.p3_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.p3_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.p3_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.src_sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.src_sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.sfr_out [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.sfr_out [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.sfr_out [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.sfr_out [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.sfr_out [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.sfr_out [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.sfr_out [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.sfr_out [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.rd_ind , \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  buf(\oc8051_top_1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(xram_data_in_model[0], xram_data_in_reg[0]);
  buf(xram_data_in_model[1], xram_data_in_reg[1]);
  buf(xram_data_in_model[2], xram_data_in_reg[2]);
  buf(xram_data_in_model[3], xram_data_in_reg[3]);
  buf(xram_data_in_model[4], xram_data_in_reg[4]);
  buf(xram_data_in_model[5], xram_data_in_reg[5]);
  buf(xram_data_in_model[6], xram_data_in_reg[6]);
  buf(xram_data_in_model[7], xram_data_in_reg[7]);
  buf(rd_rom_2_addr[0], RD_ROM_2_ABSTR_ADDR[0]);
  buf(rd_rom_2_addr[1], RD_ROM_2_ABSTR_ADDR[1]);
  buf(rd_rom_2_addr[2], RD_ROM_2_ABSTR_ADDR[2]);
  buf(rd_rom_2_addr[3], RD_ROM_2_ABSTR_ADDR[3]);
  buf(rd_rom_2_addr[4], RD_ROM_2_ABSTR_ADDR[4]);
  buf(rd_rom_2_addr[5], RD_ROM_2_ABSTR_ADDR[5]);
  buf(rd_rom_2_addr[6], RD_ROM_2_ABSTR_ADDR[6]);
  buf(rd_rom_2_addr[7], RD_ROM_2_ABSTR_ADDR[7]);
  buf(rd_rom_2_addr[8], RD_ROM_2_ABSTR_ADDR[8]);
  buf(rd_rom_2_addr[9], RD_ROM_2_ABSTR_ADDR[9]);
  buf(rd_rom_2_addr[10], RD_ROM_2_ABSTR_ADDR[10]);
  buf(rd_rom_2_addr[11], RD_ROM_2_ABSTR_ADDR[11]);
  buf(rd_rom_2_addr[12], RD_ROM_2_ABSTR_ADDR[12]);
  buf(rd_rom_2_addr[13], RD_ROM_2_ABSTR_ADDR[13]);
  buf(rd_rom_2_addr[14], RD_ROM_2_ABSTR_ADDR[14]);
  buf(rd_rom_2_addr[15], RD_ROM_2_ABSTR_ADDR[15]);
  buf(rd_rom_0_addr[0], \oc8051_golden_model_1.PC [0]);
  buf(rd_rom_0_addr[1], \oc8051_golden_model_1.PC [1]);
  buf(rd_rom_0_addr[2], \oc8051_golden_model_1.PC [2]);
  buf(rd_rom_0_addr[3], \oc8051_golden_model_1.PC [3]);
  buf(rd_rom_0_addr[4], \oc8051_golden_model_1.PC [4]);
  buf(rd_rom_0_addr[5], \oc8051_golden_model_1.PC [5]);
  buf(rd_rom_0_addr[6], \oc8051_golden_model_1.PC [6]);
  buf(rd_rom_0_addr[7], \oc8051_golden_model_1.PC [7]);
  buf(rd_rom_0_addr[8], \oc8051_golden_model_1.PC [8]);
  buf(rd_rom_0_addr[9], \oc8051_golden_model_1.PC [9]);
  buf(rd_rom_0_addr[10], \oc8051_golden_model_1.PC [10]);
  buf(rd_rom_0_addr[11], \oc8051_golden_model_1.PC [11]);
  buf(rd_rom_0_addr[12], \oc8051_golden_model_1.PC [12]);
  buf(rd_rom_0_addr[13], \oc8051_golden_model_1.PC [13]);
  buf(rd_rom_0_addr[14], \oc8051_golden_model_1.PC [14]);
  buf(rd_rom_0_addr[15], \oc8051_golden_model_1.PC [15]);
  buf(TMOD_gm_next[0], \oc8051_golden_model_1.TMOD [0]);
  buf(TMOD_gm_next[1], \oc8051_golden_model_1.TMOD [1]);
  buf(TMOD_gm_next[2], \oc8051_golden_model_1.TMOD [2]);
  buf(TMOD_gm_next[3], \oc8051_golden_model_1.TMOD [3]);
  buf(TMOD_gm_next[4], \oc8051_golden_model_1.TMOD [4]);
  buf(TMOD_gm_next[5], \oc8051_golden_model_1.TMOD [5]);
  buf(TMOD_gm_next[6], \oc8051_golden_model_1.TMOD [6]);
  buf(TMOD_gm_next[7], \oc8051_golden_model_1.TMOD [7]);
  buf(TMOD_gm[0], \oc8051_golden_model_1.TMOD [0]);
  buf(TMOD_gm[1], \oc8051_golden_model_1.TMOD [1]);
  buf(TMOD_gm[2], \oc8051_golden_model_1.TMOD [2]);
  buf(TMOD_gm[3], \oc8051_golden_model_1.TMOD [3]);
  buf(TMOD_gm[4], \oc8051_golden_model_1.TMOD [4]);
  buf(TMOD_gm[5], \oc8051_golden_model_1.TMOD [5]);
  buf(TMOD_gm[6], \oc8051_golden_model_1.TMOD [6]);
  buf(TMOD_gm[7], \oc8051_golden_model_1.TMOD [7]);
  buf(TL1_gm_next[0], \oc8051_golden_model_1.TL1 [0]);
  buf(TL1_gm_next[1], \oc8051_golden_model_1.TL1 [1]);
  buf(TL1_gm_next[2], \oc8051_golden_model_1.TL1 [2]);
  buf(TL1_gm_next[3], \oc8051_golden_model_1.TL1 [3]);
  buf(TL1_gm_next[4], \oc8051_golden_model_1.TL1 [4]);
  buf(TL1_gm_next[5], \oc8051_golden_model_1.TL1 [5]);
  buf(TL1_gm_next[6], \oc8051_golden_model_1.TL1 [6]);
  buf(TL1_gm_next[7], \oc8051_golden_model_1.TL1 [7]);
  buf(TL1_gm[0], \oc8051_golden_model_1.TL1 [0]);
  buf(TL1_gm[1], \oc8051_golden_model_1.TL1 [1]);
  buf(TL1_gm[2], \oc8051_golden_model_1.TL1 [2]);
  buf(TL1_gm[3], \oc8051_golden_model_1.TL1 [3]);
  buf(TL1_gm[4], \oc8051_golden_model_1.TL1 [4]);
  buf(TL1_gm[5], \oc8051_golden_model_1.TL1 [5]);
  buf(TL1_gm[6], \oc8051_golden_model_1.TL1 [6]);
  buf(TL1_gm[7], \oc8051_golden_model_1.TL1 [7]);
  buf(TL0_gm_next[0], \oc8051_golden_model_1.TL0 [0]);
  buf(TL0_gm_next[1], \oc8051_golden_model_1.TL0 [1]);
  buf(TL0_gm_next[2], \oc8051_golden_model_1.TL0 [2]);
  buf(TL0_gm_next[3], \oc8051_golden_model_1.TL0 [3]);
  buf(TL0_gm_next[4], \oc8051_golden_model_1.TL0 [4]);
  buf(TL0_gm_next[5], \oc8051_golden_model_1.TL0 [5]);
  buf(TL0_gm_next[6], \oc8051_golden_model_1.TL0 [6]);
  buf(TL0_gm_next[7], \oc8051_golden_model_1.TL0 [7]);
  buf(TL0_gm[0], \oc8051_golden_model_1.TL0 [0]);
  buf(TL0_gm[1], \oc8051_golden_model_1.TL0 [1]);
  buf(TL0_gm[2], \oc8051_golden_model_1.TL0 [2]);
  buf(TL0_gm[3], \oc8051_golden_model_1.TL0 [3]);
  buf(TL0_gm[4], \oc8051_golden_model_1.TL0 [4]);
  buf(TL0_gm[5], \oc8051_golden_model_1.TL0 [5]);
  buf(TL0_gm[6], \oc8051_golden_model_1.TL0 [6]);
  buf(TL0_gm[7], \oc8051_golden_model_1.TL0 [7]);
  buf(TH1_gm_next[0], \oc8051_golden_model_1.TH1 [0]);
  buf(TH1_gm_next[1], \oc8051_golden_model_1.TH1 [1]);
  buf(TH1_gm_next[2], \oc8051_golden_model_1.TH1 [2]);
  buf(TH1_gm_next[3], \oc8051_golden_model_1.TH1 [3]);
  buf(TH1_gm_next[4], \oc8051_golden_model_1.TH1 [4]);
  buf(TH1_gm_next[5], \oc8051_golden_model_1.TH1 [5]);
  buf(TH1_gm_next[6], \oc8051_golden_model_1.TH1 [6]);
  buf(TH1_gm_next[7], \oc8051_golden_model_1.TH1 [7]);
  buf(TH1_gm[0], \oc8051_golden_model_1.TH1 [0]);
  buf(TH1_gm[1], \oc8051_golden_model_1.TH1 [1]);
  buf(TH1_gm[2], \oc8051_golden_model_1.TH1 [2]);
  buf(TH1_gm[3], \oc8051_golden_model_1.TH1 [3]);
  buf(TH1_gm[4], \oc8051_golden_model_1.TH1 [4]);
  buf(TH1_gm[5], \oc8051_golden_model_1.TH1 [5]);
  buf(TH1_gm[6], \oc8051_golden_model_1.TH1 [6]);
  buf(TH1_gm[7], \oc8051_golden_model_1.TH1 [7]);
  buf(TH0_gm_next[0], \oc8051_golden_model_1.TH0 [0]);
  buf(TH0_gm_next[1], \oc8051_golden_model_1.TH0 [1]);
  buf(TH0_gm_next[2], \oc8051_golden_model_1.TH0 [2]);
  buf(TH0_gm_next[3], \oc8051_golden_model_1.TH0 [3]);
  buf(TH0_gm_next[4], \oc8051_golden_model_1.TH0 [4]);
  buf(TH0_gm_next[5], \oc8051_golden_model_1.TH0 [5]);
  buf(TH0_gm_next[6], \oc8051_golden_model_1.TH0 [6]);
  buf(TH0_gm_next[7], \oc8051_golden_model_1.TH0 [7]);
  buf(TH0_gm[0], \oc8051_golden_model_1.TH0 [0]);
  buf(TH0_gm[1], \oc8051_golden_model_1.TH0 [1]);
  buf(TH0_gm[2], \oc8051_golden_model_1.TH0 [2]);
  buf(TH0_gm[3], \oc8051_golden_model_1.TH0 [3]);
  buf(TH0_gm[4], \oc8051_golden_model_1.TH0 [4]);
  buf(TH0_gm[5], \oc8051_golden_model_1.TH0 [5]);
  buf(TH0_gm[6], \oc8051_golden_model_1.TH0 [6]);
  buf(TH0_gm[7], \oc8051_golden_model_1.TH0 [7]);
  buf(TCON_gm_next[0], \oc8051_golden_model_1.TCON [0]);
  buf(TCON_gm_next[1], \oc8051_golden_model_1.TCON [1]);
  buf(TCON_gm_next[2], \oc8051_golden_model_1.TCON [2]);
  buf(TCON_gm_next[3], \oc8051_golden_model_1.TCON [3]);
  buf(TCON_gm_next[4], \oc8051_golden_model_1.TCON [4]);
  buf(TCON_gm_next[5], \oc8051_golden_model_1.TCON [5]);
  buf(TCON_gm_next[6], \oc8051_golden_model_1.TCON [6]);
  buf(TCON_gm_next[7], \oc8051_golden_model_1.TCON [7]);
  buf(TCON_gm[0], \oc8051_golden_model_1.TCON [0]);
  buf(TCON_gm[1], \oc8051_golden_model_1.TCON [1]);
  buf(TCON_gm[2], \oc8051_golden_model_1.TCON [2]);
  buf(TCON_gm[3], \oc8051_golden_model_1.TCON [3]);
  buf(TCON_gm[4], \oc8051_golden_model_1.TCON [4]);
  buf(TCON_gm[5], \oc8051_golden_model_1.TCON [5]);
  buf(TCON_gm[6], \oc8051_golden_model_1.TCON [6]);
  buf(TCON_gm[7], \oc8051_golden_model_1.TCON [7]);
  buf(SP_gm[0], \oc8051_golden_model_1.SP [0]);
  buf(SP_gm[1], \oc8051_golden_model_1.SP [1]);
  buf(SP_gm[2], \oc8051_golden_model_1.SP [2]);
  buf(SP_gm[3], \oc8051_golden_model_1.SP [3]);
  buf(SP_gm[4], \oc8051_golden_model_1.SP [4]);
  buf(SP_gm[5], \oc8051_golden_model_1.SP [5]);
  buf(SP_gm[6], \oc8051_golden_model_1.SP [6]);
  buf(SP_gm[7], \oc8051_golden_model_1.SP [7]);
  buf(SCON_gm_next[0], \oc8051_golden_model_1.SCON [0]);
  buf(SCON_gm_next[1], \oc8051_golden_model_1.SCON [1]);
  buf(SCON_gm_next[2], \oc8051_golden_model_1.SCON [2]);
  buf(SCON_gm_next[3], \oc8051_golden_model_1.SCON [3]);
  buf(SCON_gm_next[4], \oc8051_golden_model_1.SCON [4]);
  buf(SCON_gm_next[5], \oc8051_golden_model_1.SCON [5]);
  buf(SCON_gm_next[6], \oc8051_golden_model_1.SCON [6]);
  buf(SCON_gm_next[7], \oc8051_golden_model_1.SCON [7]);
  buf(SCON_gm[0], \oc8051_golden_model_1.SCON [0]);
  buf(SCON_gm[1], \oc8051_golden_model_1.SCON [1]);
  buf(SCON_gm[2], \oc8051_golden_model_1.SCON [2]);
  buf(SCON_gm[3], \oc8051_golden_model_1.SCON [3]);
  buf(SCON_gm[4], \oc8051_golden_model_1.SCON [4]);
  buf(SCON_gm[5], \oc8051_golden_model_1.SCON [5]);
  buf(SCON_gm[6], \oc8051_golden_model_1.SCON [6]);
  buf(SCON_gm[7], \oc8051_golden_model_1.SCON [7]);
  buf(SBUF_gm_next[0], \oc8051_golden_model_1.SBUF [0]);
  buf(SBUF_gm_next[1], \oc8051_golden_model_1.SBUF [1]);
  buf(SBUF_gm_next[2], \oc8051_golden_model_1.SBUF [2]);
  buf(SBUF_gm_next[3], \oc8051_golden_model_1.SBUF [3]);
  buf(SBUF_gm_next[4], \oc8051_golden_model_1.SBUF [4]);
  buf(SBUF_gm_next[5], \oc8051_golden_model_1.SBUF [5]);
  buf(SBUF_gm_next[6], \oc8051_golden_model_1.SBUF [6]);
  buf(SBUF_gm_next[7], \oc8051_golden_model_1.SBUF [7]);
  buf(SBUF_gm[0], \oc8051_golden_model_1.SBUF [0]);
  buf(SBUF_gm[1], \oc8051_golden_model_1.SBUF [1]);
  buf(SBUF_gm[2], \oc8051_golden_model_1.SBUF [2]);
  buf(SBUF_gm[3], \oc8051_golden_model_1.SBUF [3]);
  buf(SBUF_gm[4], \oc8051_golden_model_1.SBUF [4]);
  buf(SBUF_gm[5], \oc8051_golden_model_1.SBUF [5]);
  buf(SBUF_gm[6], \oc8051_golden_model_1.SBUF [6]);
  buf(SBUF_gm[7], \oc8051_golden_model_1.SBUF [7]);
  buf(PSW_gm[0], \oc8051_golden_model_1.PSW [0]);
  buf(PSW_gm[1], \oc8051_golden_model_1.PSW [1]);
  buf(PSW_gm[2], \oc8051_golden_model_1.PSW [2]);
  buf(PSW_gm[3], \oc8051_golden_model_1.PSW [3]);
  buf(PSW_gm[4], \oc8051_golden_model_1.PSW [4]);
  buf(PSW_gm[5], \oc8051_golden_model_1.PSW [5]);
  buf(PSW_gm[6], \oc8051_golden_model_1.PSW [6]);
  buf(PSW_gm[7], \oc8051_golden_model_1.PSW [7]);
  buf(PCON_gm_next[0], \oc8051_golden_model_1.PCON [0]);
  buf(PCON_gm_next[1], \oc8051_golden_model_1.PCON [1]);
  buf(PCON_gm_next[2], \oc8051_golden_model_1.PCON [2]);
  buf(PCON_gm_next[3], \oc8051_golden_model_1.PCON [3]);
  buf(PCON_gm_next[4], \oc8051_golden_model_1.PCON [4]);
  buf(PCON_gm_next[5], \oc8051_golden_model_1.PCON [5]);
  buf(PCON_gm_next[6], \oc8051_golden_model_1.PCON [6]);
  buf(PCON_gm_next[7], \oc8051_golden_model_1.PCON [7]);
  buf(PCON_gm[0], \oc8051_golden_model_1.PCON [0]);
  buf(PCON_gm[1], \oc8051_golden_model_1.PCON [1]);
  buf(PCON_gm[2], \oc8051_golden_model_1.PCON [2]);
  buf(PCON_gm[3], \oc8051_golden_model_1.PCON [3]);
  buf(PCON_gm[4], \oc8051_golden_model_1.PCON [4]);
  buf(PCON_gm[5], \oc8051_golden_model_1.PCON [5]);
  buf(PCON_gm[6], \oc8051_golden_model_1.PCON [6]);
  buf(PCON_gm[7], \oc8051_golden_model_1.PCON [7]);
  buf(P3_gm[0], \oc8051_golden_model_1.P3 [0]);
  buf(P3_gm[1], \oc8051_golden_model_1.P3 [1]);
  buf(P3_gm[2], \oc8051_golden_model_1.P3 [2]);
  buf(P3_gm[3], \oc8051_golden_model_1.P3 [3]);
  buf(P3_gm[4], \oc8051_golden_model_1.P3 [4]);
  buf(P3_gm[5], \oc8051_golden_model_1.P3 [5]);
  buf(P3_gm[6], \oc8051_golden_model_1.P3 [6]);
  buf(P3_gm[7], \oc8051_golden_model_1.P3 [7]);
  buf(P2_gm[0], \oc8051_golden_model_1.P2 [0]);
  buf(P2_gm[1], \oc8051_golden_model_1.P2 [1]);
  buf(P2_gm[2], \oc8051_golden_model_1.P2 [2]);
  buf(P2_gm[3], \oc8051_golden_model_1.P2 [3]);
  buf(P2_gm[4], \oc8051_golden_model_1.P2 [4]);
  buf(P2_gm[5], \oc8051_golden_model_1.P2 [5]);
  buf(P2_gm[6], \oc8051_golden_model_1.P2 [6]);
  buf(P2_gm[7], \oc8051_golden_model_1.P2 [7]);
  buf(P1_gm[0], \oc8051_golden_model_1.P1 [0]);
  buf(P1_gm[1], \oc8051_golden_model_1.P1 [1]);
  buf(P1_gm[2], \oc8051_golden_model_1.P1 [2]);
  buf(P1_gm[3], \oc8051_golden_model_1.P1 [3]);
  buf(P1_gm[4], \oc8051_golden_model_1.P1 [4]);
  buf(P1_gm[5], \oc8051_golden_model_1.P1 [5]);
  buf(P1_gm[6], \oc8051_golden_model_1.P1 [6]);
  buf(P1_gm[7], \oc8051_golden_model_1.P1 [7]);
  buf(P0_gm[0], \oc8051_golden_model_1.P0 [0]);
  buf(P0_gm[1], \oc8051_golden_model_1.P0 [1]);
  buf(P0_gm[2], \oc8051_golden_model_1.P0 [2]);
  buf(P0_gm[3], \oc8051_golden_model_1.P0 [3]);
  buf(P0_gm[4], \oc8051_golden_model_1.P0 [4]);
  buf(P0_gm[5], \oc8051_golden_model_1.P0 [5]);
  buf(P0_gm[6], \oc8051_golden_model_1.P0 [6]);
  buf(P0_gm[7], \oc8051_golden_model_1.P0 [7]);
  buf(IP_gm_next[0], \oc8051_golden_model_1.IP [0]);
  buf(IP_gm_next[1], \oc8051_golden_model_1.IP [1]);
  buf(IP_gm_next[2], \oc8051_golden_model_1.IP [2]);
  buf(IP_gm_next[3], \oc8051_golden_model_1.IP [3]);
  buf(IP_gm_next[4], \oc8051_golden_model_1.IP [4]);
  buf(IP_gm_next[5], \oc8051_golden_model_1.IP [5]);
  buf(IP_gm_next[6], \oc8051_golden_model_1.IP [6]);
  buf(IP_gm_next[7], \oc8051_golden_model_1.IP [7]);
  buf(IP_gm[0], \oc8051_golden_model_1.IP [0]);
  buf(IP_gm[1], \oc8051_golden_model_1.IP [1]);
  buf(IP_gm[2], \oc8051_golden_model_1.IP [2]);
  buf(IP_gm[3], \oc8051_golden_model_1.IP [3]);
  buf(IP_gm[4], \oc8051_golden_model_1.IP [4]);
  buf(IP_gm[5], \oc8051_golden_model_1.IP [5]);
  buf(IP_gm[6], \oc8051_golden_model_1.IP [6]);
  buf(IP_gm[7], \oc8051_golden_model_1.IP [7]);
  buf(IE_gm_next[0], \oc8051_golden_model_1.IE [0]);
  buf(IE_gm_next[1], \oc8051_golden_model_1.IE [1]);
  buf(IE_gm_next[2], \oc8051_golden_model_1.IE [2]);
  buf(IE_gm_next[3], \oc8051_golden_model_1.IE [3]);
  buf(IE_gm_next[4], \oc8051_golden_model_1.IE [4]);
  buf(IE_gm_next[5], \oc8051_golden_model_1.IE [5]);
  buf(IE_gm_next[6], \oc8051_golden_model_1.IE [6]);
  buf(IE_gm_next[7], \oc8051_golden_model_1.IE [7]);
  buf(IE_gm[0], \oc8051_golden_model_1.IE [0]);
  buf(IE_gm[1], \oc8051_golden_model_1.IE [1]);
  buf(IE_gm[2], \oc8051_golden_model_1.IE [2]);
  buf(IE_gm[3], \oc8051_golden_model_1.IE [3]);
  buf(IE_gm[4], \oc8051_golden_model_1.IE [4]);
  buf(IE_gm[5], \oc8051_golden_model_1.IE [5]);
  buf(IE_gm[6], \oc8051_golden_model_1.IE [6]);
  buf(IE_gm[7], \oc8051_golden_model_1.IE [7]);
  buf(DPH_gm[0], \oc8051_golden_model_1.DPH [0]);
  buf(DPH_gm[1], \oc8051_golden_model_1.DPH [1]);
  buf(DPH_gm[2], \oc8051_golden_model_1.DPH [2]);
  buf(DPH_gm[3], \oc8051_golden_model_1.DPH [3]);
  buf(DPH_gm[4], \oc8051_golden_model_1.DPH [4]);
  buf(DPH_gm[5], \oc8051_golden_model_1.DPH [5]);
  buf(DPH_gm[6], \oc8051_golden_model_1.DPH [6]);
  buf(DPH_gm[7], \oc8051_golden_model_1.DPH [7]);
  buf(DPL_gm[0], \oc8051_golden_model_1.DPL [0]);
  buf(DPL_gm[1], \oc8051_golden_model_1.DPL [1]);
  buf(DPL_gm[2], \oc8051_golden_model_1.DPL [2]);
  buf(DPL_gm[3], \oc8051_golden_model_1.DPL [3]);
  buf(DPL_gm[4], \oc8051_golden_model_1.DPL [4]);
  buf(DPL_gm[5], \oc8051_golden_model_1.DPL [5]);
  buf(DPL_gm[6], \oc8051_golden_model_1.DPL [6]);
  buf(DPL_gm[7], \oc8051_golden_model_1.DPL [7]);
  buf(B_gm[0], \oc8051_golden_model_1.B [0]);
  buf(B_gm[1], \oc8051_golden_model_1.B [1]);
  buf(B_gm[2], \oc8051_golden_model_1.B [2]);
  buf(B_gm[3], \oc8051_golden_model_1.B [3]);
  buf(B_gm[4], \oc8051_golden_model_1.B [4]);
  buf(B_gm[5], \oc8051_golden_model_1.B [5]);
  buf(B_gm[6], \oc8051_golden_model_1.B [6]);
  buf(B_gm[7], \oc8051_golden_model_1.B [7]);
  buf(ACC_gm[0], \oc8051_golden_model_1.ACC [0]);
  buf(ACC_gm[1], \oc8051_golden_model_1.ACC [1]);
  buf(ACC_gm[2], \oc8051_golden_model_1.ACC [2]);
  buf(ACC_gm[3], \oc8051_golden_model_1.ACC [3]);
  buf(ACC_gm[4], \oc8051_golden_model_1.ACC [4]);
  buf(ACC_gm[5], \oc8051_golden_model_1.ACC [5]);
  buf(ACC_gm[6], \oc8051_golden_model_1.ACC [6]);
  buf(ACC_gm[7], \oc8051_golden_model_1.ACC [7]);
  buf(dptr_impl[0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(dptr_impl[1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(dptr_impl[2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(dptr_impl[3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(dptr_impl[4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(dptr_impl[5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(dptr_impl[6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(dptr_impl[7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(dptr_impl[8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(dptr_impl[9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(dptr_impl[10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(dptr_impl[11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(dptr_impl[12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(dptr_impl[13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(dptr_impl[14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(dptr_impl[15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(b_reg_impl[0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(b_reg_impl[1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(b_reg_impl[2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(b_reg_impl[3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(b_reg_impl[4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(b_reg_impl[5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(b_reg_impl[6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(b_reg_impl[7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(acc_impl[0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(acc_impl[1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(acc_impl[2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(acc_impl[3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(acc_impl[4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(acc_impl[5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(acc_impl[6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(acc_impl[7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(psw_impl[1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(psw_impl[2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(psw_impl[3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(psw_impl[4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(psw_impl[5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(psw_impl[6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(psw_impl[7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(pc1[0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(pc1[1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(pc1[2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(pc1[3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(pc1[4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(pc1[5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(pc1[6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(pc1[7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(pc1[8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(pc1[9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(pc1[10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(pc1[11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(pc1[12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(pc1[13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(pc1[14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(pc1[15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(pc2[0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(pc2[1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(pc2[2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(pc2[3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(pc2[4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(pc2[5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(pc2[6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(pc2[7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(pc2[8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(pc2[9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(pc2[10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(pc2[11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(pc2[12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(pc2[13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(pc2[14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(pc2[15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(cxrom_data_out[0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(cxrom_data_out[1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(cxrom_data_out[2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(cxrom_data_out[3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(cxrom_data_out[4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(cxrom_data_out[5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(cxrom_data_out[6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(cxrom_data_out[7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(cxrom_data_out[8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(cxrom_data_out[9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(cxrom_data_out[10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(cxrom_data_out[11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(cxrom_data_out[12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(cxrom_data_out[13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(cxrom_data_out[14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(cxrom_data_out[15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(cxrom_data_out[16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(cxrom_data_out[17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(cxrom_data_out[18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(cxrom_data_out[19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(cxrom_data_out[20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(cxrom_data_out[21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(cxrom_data_out[22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(cxrom_data_out[23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(cxrom_data_out[24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(cxrom_data_out[25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(cxrom_data_out[26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(cxrom_data_out[27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(cxrom_data_out[28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(cxrom_data_out[29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(cxrom_data_out[30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(cxrom_data_out[31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(wbd_dat_o[0], \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  buf(wbd_dat_o[1], \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  buf(wbd_dat_o[2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  buf(wbd_dat_o[3], \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  buf(wbd_dat_o[4], \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  buf(wbd_dat_o[5], \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  buf(wbd_dat_o[6], \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  buf(wbd_dat_o[7], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  buf(wbd_cyc_o, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_we_o, \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  buf(wbd_ack_i, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_stb_o, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_adr_o[0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(wbd_adr_o[1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(wbd_adr_o[2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(wbd_adr_o[3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(wbd_adr_o[4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(wbd_adr_o[5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(wbd_adr_o[6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(wbd_adr_o[7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(wbd_adr_o[8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(wbd_adr_o[9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(wbd_adr_o[10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(wbd_adr_o[11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(wbd_adr_o[12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(wbd_adr_o[13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(wbd_adr_o[14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(wbd_adr_o[15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(wbd_dat_i[0], xram_data_in_reg[0]);
  buf(wbd_dat_i[1], xram_data_in_reg[1]);
  buf(wbd_dat_i[2], xram_data_in_reg[2]);
  buf(wbd_dat_i[3], xram_data_in_reg[3]);
  buf(wbd_dat_i[4], xram_data_in_reg[4]);
  buf(wbd_dat_i[5], xram_data_in_reg[5]);
  buf(wbd_dat_i[6], xram_data_in_reg[6]);
  buf(wbd_dat_i[7], xram_data_in_reg[7]);
  buf(p3_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(p3_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(p3_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(p3_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(p3_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(p3_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(p3_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(p3_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(p2_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(p2_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(p2_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(p2_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(p2_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(p2_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(p2_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(p2_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(p1_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(p1_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(p1_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(p1_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(p1_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(p1_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(p1_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(p1_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(p0_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(p0_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(p0_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(p0_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(p0_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(p0_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(p0_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(p0_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
endmodule
