
module oc8051_fv_top(clk, rst, word_in, p0_in, p1_in, p2_in, p3_in, rxd_i, t0_i, t1_i, t2_i, t2ex_i, property_invalid_ajmp, ABINPUT, ABINPUT000, ABINPUT001);
  wire _00000_;
  wire _00001_;
  wire _00002_;
  wire _00003_;
  wire _00004_;
  wire _00005_;
  wire _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  wire _08001_;
  wire _08002_;
  wire _08003_;
  wire _08004_;
  wire _08005_;
  wire _08006_;
  wire _08007_;
  wire _08008_;
  wire _08009_;
  wire _08010_;
  wire _08011_;
  wire _08012_;
  wire _08013_;
  wire _08014_;
  wire _08015_;
  wire _08016_;
  wire _08017_;
  wire _08018_;
  wire _08019_;
  wire _08020_;
  wire _08021_;
  wire _08022_;
  wire _08023_;
  wire _08024_;
  wire _08025_;
  wire _08026_;
  wire _08027_;
  wire _08028_;
  wire _08029_;
  wire _08030_;
  wire _08031_;
  wire _08032_;
  wire _08033_;
  wire _08034_;
  wire _08035_;
  wire _08036_;
  wire _08037_;
  wire _08038_;
  wire _08039_;
  wire _08040_;
  wire _08041_;
  wire _08042_;
  wire _08043_;
  wire _08044_;
  wire _08045_;
  wire _08046_;
  wire _08047_;
  wire _08048_;
  wire _08049_;
  wire _08050_;
  wire _08051_;
  wire _08052_;
  wire _08053_;
  wire _08054_;
  wire _08055_;
  wire _08056_;
  wire _08057_;
  wire _08058_;
  wire _08059_;
  wire _08060_;
  wire _08061_;
  wire _08062_;
  wire _08063_;
  wire _08064_;
  wire _08065_;
  wire _08066_;
  wire _08067_;
  wire _08068_;
  wire _08069_;
  wire _08070_;
  wire _08071_;
  wire _08072_;
  wire _08073_;
  wire _08074_;
  wire _08075_;
  wire _08076_;
  wire _08077_;
  wire _08078_;
  wire _08079_;
  wire _08080_;
  wire _08081_;
  wire _08082_;
  wire _08083_;
  wire _08084_;
  wire _08085_;
  wire _08086_;
  wire _08087_;
  wire _08088_;
  wire _08089_;
  wire _08090_;
  wire _08091_;
  wire _08092_;
  wire _08093_;
  wire _08094_;
  wire _08095_;
  wire _08096_;
  wire _08097_;
  wire _08098_;
  wire _08099_;
  wire _08100_;
  wire _08101_;
  wire _08102_;
  wire _08103_;
  wire _08104_;
  wire _08105_;
  wire _08106_;
  wire _08107_;
  wire _08108_;
  wire _08109_;
  wire _08110_;
  wire _08111_;
  wire _08112_;
  wire _08113_;
  wire _08114_;
  wire _08115_;
  wire _08116_;
  wire _08117_;
  wire _08118_;
  wire _08119_;
  wire _08120_;
  wire _08121_;
  wire _08122_;
  wire _08123_;
  wire _08124_;
  wire _08125_;
  wire _08126_;
  wire _08127_;
  wire _08128_;
  wire _08129_;
  wire _08130_;
  wire _08131_;
  wire _08132_;
  wire _08133_;
  wire _08134_;
  wire _08135_;
  wire _08136_;
  wire _08137_;
  wire _08138_;
  wire _08139_;
  wire _08140_;
  wire _08141_;
  wire _08142_;
  wire _08143_;
  wire _08144_;
  wire _08145_;
  wire _08146_;
  wire _08147_;
  wire _08148_;
  wire _08149_;
  wire _08150_;
  wire _08151_;
  wire _08152_;
  wire _08153_;
  wire _08154_;
  wire _08155_;
  wire _08156_;
  wire _08157_;
  wire _08158_;
  wire _08159_;
  wire _08160_;
  wire _08161_;
  wire _08162_;
  wire _08163_;
  wire _08164_;
  wire _08165_;
  wire _08166_;
  wire _08167_;
  wire _08168_;
  wire _08169_;
  wire _08170_;
  wire _08171_;
  wire _08172_;
  wire _08173_;
  wire _08174_;
  wire _08175_;
  wire _08176_;
  wire _08177_;
  wire _08178_;
  wire _08179_;
  wire _08180_;
  wire _08181_;
  wire _08182_;
  wire _08183_;
  wire _08184_;
  wire _08185_;
  wire _08186_;
  wire _08187_;
  wire _08188_;
  wire _08189_;
  wire _08190_;
  wire _08191_;
  wire _08192_;
  wire _08193_;
  wire _08194_;
  wire _08195_;
  wire _08196_;
  wire _08197_;
  wire _08198_;
  wire _08199_;
  wire _08200_;
  wire _08201_;
  wire _08202_;
  wire _08203_;
  wire _08204_;
  wire _08205_;
  wire _08206_;
  wire _08207_;
  wire _08208_;
  wire _08209_;
  wire _08210_;
  wire _08211_;
  wire _08212_;
  wire _08213_;
  wire _08214_;
  wire _08215_;
  wire _08216_;
  wire _08217_;
  wire _08218_;
  wire _08219_;
  wire _08220_;
  wire _08221_;
  wire _08222_;
  wire _08223_;
  wire _08224_;
  wire _08225_;
  wire _08226_;
  wire _08227_;
  wire _08228_;
  wire _08229_;
  wire _08230_;
  wire _08231_;
  wire _08232_;
  wire _08233_;
  wire _08234_;
  wire _08235_;
  wire _08236_;
  wire _08237_;
  wire _08238_;
  wire _08239_;
  wire _08240_;
  wire _08241_;
  wire _08242_;
  wire _08243_;
  wire _08244_;
  wire _08245_;
  wire _08246_;
  wire _08247_;
  wire _08248_;
  wire _08249_;
  wire _08250_;
  wire _08251_;
  wire _08252_;
  wire _08253_;
  wire _08254_;
  wire _08255_;
  wire _08256_;
  wire _08257_;
  wire _08258_;
  wire _08259_;
  wire _08260_;
  wire _08261_;
  wire _08262_;
  wire _08263_;
  wire _08264_;
  wire _08265_;
  wire _08266_;
  wire _08267_;
  wire _08268_;
  wire _08269_;
  wire _08270_;
  wire _08271_;
  wire _08272_;
  wire _08273_;
  wire _08274_;
  wire _08275_;
  wire _08276_;
  wire _08277_;
  wire _08278_;
  wire _08279_;
  wire _08280_;
  wire _08281_;
  wire _08282_;
  wire _08283_;
  wire _08284_;
  wire _08285_;
  wire _08286_;
  wire _08287_;
  wire _08288_;
  wire _08289_;
  wire _08290_;
  wire _08291_;
  wire _08292_;
  wire _08293_;
  wire _08294_;
  wire _08295_;
  wire _08296_;
  wire _08297_;
  wire _08298_;
  wire _08299_;
  wire _08300_;
  wire _08301_;
  wire _08302_;
  wire _08303_;
  wire _08304_;
  wire _08305_;
  wire _08306_;
  wire _08307_;
  wire _08308_;
  wire _08309_;
  wire _08310_;
  wire _08311_;
  wire _08312_;
  wire _08313_;
  wire _08314_;
  wire _08315_;
  wire _08316_;
  wire _08317_;
  wire _08318_;
  wire _08319_;
  wire _08320_;
  wire _08321_;
  wire _08322_;
  wire _08323_;
  wire _08324_;
  wire _08325_;
  wire _08326_;
  wire _08327_;
  wire _08328_;
  wire _08329_;
  wire _08330_;
  wire _08331_;
  wire _08332_;
  wire _08333_;
  wire _08334_;
  wire _08335_;
  wire _08336_;
  wire _08337_;
  wire _08338_;
  wire _08339_;
  wire _08340_;
  wire _08341_;
  wire _08342_;
  wire _08343_;
  wire _08344_;
  wire _08345_;
  wire _08346_;
  wire _08347_;
  wire _08348_;
  wire _08349_;
  wire _08350_;
  wire _08351_;
  wire _08352_;
  wire _08353_;
  wire _08354_;
  wire _08355_;
  wire _08356_;
  wire _08357_;
  wire _08358_;
  wire _08359_;
  wire _08360_;
  wire _08361_;
  wire _08362_;
  wire _08363_;
  wire _08364_;
  wire _08365_;
  wire _08366_;
  wire _08367_;
  wire _08368_;
  wire _08369_;
  wire _08370_;
  wire _08371_;
  wire _08372_;
  wire _08373_;
  wire _08374_;
  wire _08375_;
  wire _08376_;
  wire _08377_;
  wire _08378_;
  wire _08379_;
  wire _08380_;
  wire _08381_;
  wire _08382_;
  wire _08383_;
  wire _08384_;
  wire _08385_;
  wire _08386_;
  wire _08387_;
  wire _08388_;
  wire _08389_;
  wire _08390_;
  wire _08391_;
  wire _08392_;
  wire _08393_;
  wire _08394_;
  wire _08395_;
  wire _08396_;
  wire _08397_;
  wire _08398_;
  wire _08399_;
  wire _08400_;
  wire _08401_;
  wire _08402_;
  wire _08403_;
  wire _08404_;
  wire _08405_;
  wire _08406_;
  wire _08407_;
  wire _08408_;
  wire _08409_;
  wire _08410_;
  wire _08411_;
  wire _08412_;
  wire _08413_;
  wire _08414_;
  wire _08415_;
  wire _08416_;
  wire _08417_;
  wire _08418_;
  wire _08419_;
  wire _08420_;
  wire _08421_;
  wire _08422_;
  wire _08423_;
  wire _08424_;
  wire _08425_;
  wire _08426_;
  wire _08427_;
  wire _08428_;
  wire _08429_;
  wire _08430_;
  wire _08431_;
  wire _08432_;
  wire _08433_;
  wire _08434_;
  wire _08435_;
  wire _08436_;
  wire _08437_;
  wire _08438_;
  wire _08439_;
  wire _08440_;
  wire _08441_;
  wire _08442_;
  wire _08443_;
  wire _08444_;
  wire _08445_;
  wire _08446_;
  wire _08447_;
  wire _08448_;
  wire _08449_;
  wire _08450_;
  wire _08451_;
  wire _08452_;
  wire _08453_;
  wire _08454_;
  wire _08455_;
  wire _08456_;
  wire _08457_;
  wire _08458_;
  wire _08459_;
  wire _08460_;
  wire _08461_;
  wire _08462_;
  wire _08463_;
  wire _08464_;
  wire _08465_;
  wire _08466_;
  wire _08467_;
  wire _08468_;
  wire _08469_;
  wire _08470_;
  wire _08471_;
  wire _08472_;
  wire _08473_;
  wire _08474_;
  wire _08475_;
  wire _08476_;
  wire _08477_;
  wire _08478_;
  wire _08479_;
  wire _08480_;
  wire _08481_;
  wire _08482_;
  wire _08483_;
  wire _08484_;
  wire _08485_;
  wire _08486_;
  wire _08487_;
  wire _08488_;
  wire _08489_;
  wire _08490_;
  wire _08491_;
  wire _08492_;
  wire _08493_;
  wire _08494_;
  wire _08495_;
  wire _08496_;
  wire _08497_;
  wire _08498_;
  wire _08499_;
  wire _08500_;
  wire _08501_;
  wire _08502_;
  wire _08503_;
  wire _08504_;
  wire _08505_;
  wire _08506_;
  wire _08507_;
  wire _08508_;
  wire _08509_;
  wire _08510_;
  wire _08511_;
  wire _08512_;
  wire _08513_;
  wire _08514_;
  wire _08515_;
  wire _08516_;
  wire _08517_;
  wire _08518_;
  wire _08519_;
  wire _08520_;
  wire _08521_;
  wire _08522_;
  wire _08523_;
  wire _08524_;
  wire _08525_;
  wire _08526_;
  wire _08527_;
  wire _08528_;
  wire _08529_;
  wire _08530_;
  wire _08531_;
  wire _08532_;
  wire _08533_;
  wire _08534_;
  wire _08535_;
  wire _08536_;
  wire _08537_;
  wire _08538_;
  wire _08539_;
  wire _08540_;
  wire _08541_;
  wire _08542_;
  wire _08543_;
  wire _08544_;
  wire _08545_;
  wire _08546_;
  wire _08547_;
  wire _08548_;
  wire _08549_;
  wire _08550_;
  wire _08551_;
  wire _08552_;
  wire _08553_;
  wire _08554_;
  wire _08555_;
  wire _08556_;
  wire _08557_;
  wire _08558_;
  wire _08559_;
  wire _08560_;
  wire _08561_;
  wire _08562_;
  wire _08563_;
  wire _08564_;
  wire _08565_;
  wire _08566_;
  wire _08567_;
  wire _08568_;
  wire _08569_;
  wire _08570_;
  wire _08571_;
  wire _08572_;
  wire _08573_;
  wire _08574_;
  wire _08575_;
  wire _08576_;
  wire _08577_;
  wire _08578_;
  wire _08579_;
  wire _08580_;
  wire _08581_;
  wire _08582_;
  wire _08583_;
  wire _08584_;
  wire _08585_;
  wire _08586_;
  wire _08587_;
  wire _08588_;
  wire _08589_;
  wire _08590_;
  wire _08591_;
  wire _08592_;
  wire _08593_;
  wire _08594_;
  wire _08595_;
  wire _08596_;
  wire _08597_;
  wire _08598_;
  wire _08599_;
  wire _08600_;
  wire _08601_;
  wire _08602_;
  wire _08603_;
  wire _08604_;
  wire _08605_;
  wire _08606_;
  wire _08607_;
  wire _08608_;
  wire _08609_;
  wire _08610_;
  wire _08611_;
  wire _08612_;
  wire _08613_;
  wire _08614_;
  wire _08615_;
  wire _08616_;
  wire _08617_;
  wire _08618_;
  wire _08619_;
  wire _08620_;
  wire _08621_;
  wire _08622_;
  wire _08623_;
  wire _08624_;
  wire _08625_;
  wire _08626_;
  wire _08627_;
  wire _08628_;
  wire _08629_;
  wire _08630_;
  wire _08631_;
  wire _08632_;
  wire _08633_;
  wire _08634_;
  wire _08635_;
  wire _08636_;
  wire _08637_;
  wire _08638_;
  wire _08639_;
  wire _08640_;
  wire _08641_;
  wire _08642_;
  wire _08643_;
  wire _08644_;
  wire _08645_;
  wire _08646_;
  wire _08647_;
  wire _08648_;
  wire _08649_;
  wire _08650_;
  wire _08651_;
  wire _08652_;
  wire _08653_;
  wire _08654_;
  wire _08655_;
  wire _08656_;
  wire _08657_;
  wire _08658_;
  wire _08659_;
  wire _08660_;
  wire _08661_;
  wire _08662_;
  wire _08663_;
  wire _08664_;
  wire _08665_;
  wire _08666_;
  wire _08667_;
  wire _08668_;
  wire _08669_;
  wire _08670_;
  wire _08671_;
  wire _08672_;
  wire _08673_;
  wire _08674_;
  wire _08675_;
  wire _08676_;
  wire _08677_;
  wire _08678_;
  wire _08679_;
  wire _08680_;
  wire _08681_;
  wire _08682_;
  wire _08683_;
  wire _08684_;
  wire _08685_;
  wire _08686_;
  wire _08687_;
  wire _08688_;
  wire _08689_;
  wire _08690_;
  wire _08691_;
  wire _08692_;
  wire _08693_;
  wire _08694_;
  wire _08695_;
  wire _08696_;
  wire _08697_;
  wire _08698_;
  wire _08699_;
  wire _08700_;
  wire _08701_;
  wire _08702_;
  wire _08703_;
  wire _08704_;
  wire _08705_;
  wire _08706_;
  wire _08707_;
  wire _08708_;
  wire _08709_;
  wire _08710_;
  wire _08711_;
  wire _08712_;
  wire _08713_;
  wire _08714_;
  wire _08715_;
  wire _08716_;
  wire _08717_;
  wire _08718_;
  wire _08719_;
  wire _08720_;
  wire _08721_;
  wire _08722_;
  wire _08723_;
  wire _08724_;
  wire _08725_;
  wire _08726_;
  wire _08727_;
  wire _08728_;
  wire _08729_;
  wire _08730_;
  wire _08731_;
  wire _08732_;
  wire _08733_;
  wire _08734_;
  wire _08735_;
  wire _08736_;
  wire _08737_;
  wire _08738_;
  wire _08739_;
  wire _08740_;
  wire _08741_;
  wire _08742_;
  wire _08743_;
  wire _08744_;
  wire _08745_;
  wire _08746_;
  wire _08747_;
  wire _08748_;
  wire _08749_;
  wire _08750_;
  wire _08751_;
  wire _08752_;
  wire _08753_;
  wire _08754_;
  wire _08755_;
  wire _08756_;
  wire _08757_;
  wire _08758_;
  wire _08759_;
  wire _08760_;
  wire _08761_;
  wire _08762_;
  wire _08763_;
  wire _08764_;
  wire _08765_;
  wire _08766_;
  wire _08767_;
  wire _08768_;
  wire _08769_;
  wire _08770_;
  wire _08771_;
  wire _08772_;
  wire _08773_;
  wire _08774_;
  wire _08775_;
  wire _08776_;
  wire _08777_;
  wire _08778_;
  wire _08779_;
  wire _08780_;
  wire _08781_;
  wire _08782_;
  wire _08783_;
  wire _08784_;
  wire _08785_;
  wire _08786_;
  wire _08787_;
  wire _08788_;
  wire _08789_;
  wire _08790_;
  wire _08791_;
  wire _08792_;
  wire _08793_;
  wire _08794_;
  wire _08795_;
  wire _08796_;
  wire _08797_;
  wire _08798_;
  wire _08799_;
  wire _08800_;
  wire _08801_;
  wire _08802_;
  wire _08803_;
  wire _08804_;
  wire _08805_;
  wire _08806_;
  wire _08807_;
  wire _08808_;
  wire _08809_;
  wire _08810_;
  wire _08811_;
  wire _08812_;
  wire _08813_;
  wire _08814_;
  wire _08815_;
  wire _08816_;
  wire _08817_;
  wire _08818_;
  wire _08819_;
  wire _08820_;
  wire _08821_;
  wire _08822_;
  wire _08823_;
  wire _08824_;
  wire _08825_;
  wire _08826_;
  wire _08827_;
  wire _08828_;
  wire _08829_;
  wire _08830_;
  wire _08831_;
  wire _08832_;
  wire _08833_;
  wire _08834_;
  wire _08835_;
  wire _08836_;
  wire _08837_;
  wire _08838_;
  wire _08839_;
  wire _08840_;
  wire _08841_;
  wire _08842_;
  wire _08843_;
  wire _08844_;
  wire _08845_;
  wire _08846_;
  wire _08847_;
  wire _08848_;
  wire _08849_;
  wire _08850_;
  wire _08851_;
  wire _08852_;
  wire _08853_;
  wire _08854_;
  wire _08855_;
  wire _08856_;
  wire _08857_;
  wire _08858_;
  wire _08859_;
  wire _08860_;
  wire _08861_;
  wire _08862_;
  wire _08863_;
  wire _08864_;
  wire _08865_;
  wire _08866_;
  wire _08867_;
  wire _08868_;
  wire _08869_;
  wire _08870_;
  wire _08871_;
  wire _08872_;
  wire _08873_;
  wire _08874_;
  wire _08875_;
  wire _08876_;
  wire _08877_;
  wire _08878_;
  wire _08879_;
  wire _08880_;
  wire _08881_;
  wire _08882_;
  wire _08883_;
  wire _08884_;
  wire _08885_;
  wire _08886_;
  wire _08887_;
  wire _08888_;
  wire _08889_;
  wire _08890_;
  wire _08891_;
  wire _08892_;
  wire _08893_;
  wire _08894_;
  wire _08895_;
  wire _08896_;
  wire _08897_;
  wire _08898_;
  wire _08899_;
  wire _08900_;
  wire _08901_;
  wire _08902_;
  wire _08903_;
  wire _08904_;
  wire _08905_;
  wire _08906_;
  wire _08907_;
  wire _08908_;
  wire _08909_;
  wire _08910_;
  wire _08911_;
  wire _08912_;
  wire _08913_;
  wire _08914_;
  wire _08915_;
  wire _08916_;
  wire _08917_;
  wire _08918_;
  wire _08919_;
  wire _08920_;
  wire _08921_;
  wire _08922_;
  wire _08923_;
  wire _08924_;
  wire _08925_;
  wire _08926_;
  wire _08927_;
  wire _08928_;
  wire _08929_;
  wire _08930_;
  wire _08931_;
  wire _08932_;
  wire _08933_;
  wire _08934_;
  wire _08935_;
  wire _08936_;
  wire _08937_;
  wire _08938_;
  wire _08939_;
  wire _08940_;
  wire _08941_;
  wire _08942_;
  wire _08943_;
  wire _08944_;
  wire _08945_;
  wire _08946_;
  wire _08947_;
  wire _08948_;
  wire _08949_;
  wire _08950_;
  wire _08951_;
  wire _08952_;
  wire _08953_;
  wire _08954_;
  wire _08955_;
  wire _08956_;
  wire _08957_;
  wire _08958_;
  wire _08959_;
  wire _08960_;
  wire _08961_;
  wire _08962_;
  wire _08963_;
  wire _08964_;
  wire _08965_;
  wire _08966_;
  wire _08967_;
  wire _08968_;
  wire _08969_;
  wire _08970_;
  wire _08971_;
  wire _08972_;
  wire _08973_;
  wire _08974_;
  wire _08975_;
  wire _08976_;
  wire _08977_;
  wire _08978_;
  wire _08979_;
  wire _08980_;
  wire _08981_;
  wire _08982_;
  wire _08983_;
  wire _08984_;
  wire _08985_;
  wire _08986_;
  wire _08987_;
  wire _08988_;
  wire _08989_;
  wire _08990_;
  wire _08991_;
  wire _08992_;
  wire _08993_;
  wire _08994_;
  wire _08995_;
  wire _08996_;
  wire _08997_;
  wire _08998_;
  wire _08999_;
  wire _09000_;
  wire _09001_;
  wire _09002_;
  wire _09003_;
  wire _09004_;
  wire _09005_;
  wire _09006_;
  wire _09007_;
  wire _09008_;
  wire _09009_;
  wire _09010_;
  wire _09011_;
  wire _09012_;
  wire _09013_;
  wire _09014_;
  wire _09015_;
  wire _09016_;
  wire _09017_;
  wire _09018_;
  wire _09019_;
  wire _09020_;
  wire _09021_;
  wire _09022_;
  wire _09023_;
  wire _09024_;
  wire _09025_;
  wire _09026_;
  wire _09027_;
  wire _09028_;
  wire _09029_;
  wire _09030_;
  wire _09031_;
  wire _09032_;
  wire _09033_;
  wire _09034_;
  wire _09035_;
  wire _09036_;
  wire _09037_;
  wire _09038_;
  wire _09039_;
  wire _09040_;
  wire _09041_;
  wire _09042_;
  wire _09043_;
  wire _09044_;
  wire _09045_;
  wire _09046_;
  wire _09047_;
  wire _09048_;
  wire _09049_;
  wire _09050_;
  wire _09051_;
  wire _09052_;
  wire _09053_;
  wire _09054_;
  wire _09055_;
  wire _09056_;
  wire _09057_;
  wire _09058_;
  wire _09059_;
  wire _09060_;
  wire _09061_;
  wire _09062_;
  wire _09063_;
  wire _09064_;
  wire _09065_;
  wire _09066_;
  wire _09067_;
  wire _09068_;
  wire _09069_;
  wire _09070_;
  wire _09071_;
  wire _09072_;
  wire _09073_;
  wire _09074_;
  wire _09075_;
  wire _09076_;
  wire _09077_;
  wire _09078_;
  wire _09079_;
  wire _09080_;
  wire _09081_;
  wire _09082_;
  wire _09083_;
  wire _09084_;
  wire _09085_;
  wire _09086_;
  wire _09087_;
  wire _09088_;
  wire _09089_;
  wire _09090_;
  wire _09091_;
  wire _09092_;
  wire _09093_;
  wire _09094_;
  wire _09095_;
  wire _09096_;
  wire _09097_;
  wire _09098_;
  wire _09099_;
  wire _09100_;
  wire _09101_;
  wire _09102_;
  wire _09103_;
  wire _09104_;
  wire _09105_;
  wire _09106_;
  wire _09107_;
  wire _09108_;
  wire _09109_;
  wire _09110_;
  wire _09111_;
  wire _09112_;
  wire _09113_;
  wire _09114_;
  wire _09115_;
  wire _09116_;
  wire _09117_;
  wire _09118_;
  wire _09119_;
  wire _09120_;
  wire _09121_;
  wire _09122_;
  wire _09123_;
  wire _09124_;
  wire _09125_;
  wire _09126_;
  wire _09127_;
  wire _09128_;
  wire _09129_;
  wire _09130_;
  wire _09131_;
  wire _09132_;
  wire _09133_;
  wire _09134_;
  wire _09135_;
  wire _09136_;
  wire _09137_;
  wire _09138_;
  wire _09139_;
  wire _09140_;
  wire _09141_;
  wire _09142_;
  wire _09143_;
  wire _09144_;
  wire _09145_;
  wire _09146_;
  wire _09147_;
  wire _09148_;
  wire _09149_;
  wire _09150_;
  wire _09151_;
  wire _09152_;
  wire _09153_;
  wire _09154_;
  wire _09155_;
  wire _09156_;
  wire _09157_;
  wire _09158_;
  wire _09159_;
  wire _09160_;
  wire _09161_;
  wire _09162_;
  wire _09163_;
  wire _09164_;
  wire _09165_;
  wire _09166_;
  wire _09167_;
  wire _09168_;
  wire _09169_;
  wire _09170_;
  wire _09171_;
  wire _09172_;
  wire _09173_;
  wire _09174_;
  wire _09175_;
  wire _09176_;
  wire _09177_;
  wire _09178_;
  wire _09179_;
  wire _09180_;
  wire _09181_;
  wire _09182_;
  wire _09183_;
  wire _09184_;
  wire _09185_;
  wire _09186_;
  wire _09187_;
  wire _09188_;
  wire _09189_;
  wire _09190_;
  wire _09191_;
  wire _09192_;
  wire _09193_;
  wire _09194_;
  wire _09195_;
  wire _09196_;
  wire _09197_;
  wire _09198_;
  wire _09199_;
  wire _09200_;
  wire _09201_;
  wire _09202_;
  wire _09203_;
  wire _09204_;
  wire _09205_;
  wire _09206_;
  wire _09207_;
  wire _09208_;
  wire _09209_;
  wire _09210_;
  wire _09211_;
  wire _09212_;
  wire _09213_;
  wire _09214_;
  wire _09215_;
  wire _09216_;
  wire _09217_;
  wire _09218_;
  wire _09219_;
  wire _09220_;
  wire _09221_;
  wire _09222_;
  wire _09223_;
  wire _09224_;
  wire _09225_;
  wire _09226_;
  wire _09227_;
  wire _09228_;
  wire _09229_;
  wire _09230_;
  wire _09231_;
  wire _09232_;
  wire _09233_;
  wire _09234_;
  wire _09235_;
  wire _09236_;
  wire _09237_;
  wire _09238_;
  wire _09239_;
  wire _09240_;
  wire _09241_;
  wire _09242_;
  wire _09243_;
  wire _09244_;
  wire _09245_;
  wire _09246_;
  wire _09247_;
  wire _09248_;
  wire _09249_;
  wire _09250_;
  wire _09251_;
  wire _09252_;
  wire _09253_;
  wire _09254_;
  wire _09255_;
  wire _09256_;
  wire _09257_;
  wire _09258_;
  wire _09259_;
  wire _09260_;
  wire _09261_;
  wire _09262_;
  wire _09263_;
  wire _09264_;
  wire _09265_;
  wire _09266_;
  wire _09267_;
  wire _09268_;
  wire _09269_;
  wire _09270_;
  wire _09271_;
  wire _09272_;
  wire _09273_;
  wire _09274_;
  wire _09275_;
  wire _09276_;
  wire _09277_;
  wire _09278_;
  wire _09279_;
  wire _09280_;
  wire _09281_;
  wire _09282_;
  wire _09283_;
  wire _09284_;
  wire _09285_;
  wire _09286_;
  wire _09287_;
  wire _09288_;
  wire _09289_;
  wire _09290_;
  wire _09291_;
  wire _09292_;
  wire _09293_;
  wire _09294_;
  wire _09295_;
  wire _09296_;
  wire _09297_;
  wire _09298_;
  wire _09299_;
  wire _09300_;
  wire _09301_;
  wire _09302_;
  wire _09303_;
  wire _09304_;
  wire _09305_;
  wire _09306_;
  wire _09307_;
  wire _09308_;
  wire _09309_;
  wire _09310_;
  wire _09311_;
  wire _09312_;
  wire _09313_;
  wire _09314_;
  wire _09315_;
  wire _09316_;
  wire _09317_;
  wire _09318_;
  wire _09319_;
  wire _09320_;
  wire _09321_;
  wire _09322_;
  wire _09323_;
  wire _09324_;
  wire _09325_;
  wire _09326_;
  wire _09327_;
  wire _09328_;
  wire _09329_;
  wire _09330_;
  wire _09331_;
  wire _09332_;
  wire _09333_;
  wire _09334_;
  wire _09335_;
  wire _09336_;
  wire _09337_;
  wire _09338_;
  wire _09339_;
  wire _09340_;
  wire _09341_;
  wire _09342_;
  wire _09343_;
  wire _09344_;
  wire _09345_;
  wire _09346_;
  wire _09347_;
  wire _09348_;
  wire _09349_;
  wire _09350_;
  wire _09351_;
  wire _09352_;
  wire _09353_;
  wire _09354_;
  wire _09355_;
  wire _09356_;
  wire _09357_;
  wire _09358_;
  wire _09359_;
  wire _09360_;
  wire _09361_;
  wire _09362_;
  wire _09363_;
  wire _09364_;
  wire _09365_;
  wire _09366_;
  wire _09367_;
  wire _09368_;
  wire _09369_;
  wire _09370_;
  wire _09371_;
  wire _09372_;
  wire _09373_;
  wire _09374_;
  wire _09375_;
  wire _09376_;
  wire _09377_;
  wire _09378_;
  wire _09379_;
  wire _09380_;
  wire _09381_;
  wire _09382_;
  wire _09383_;
  wire _09384_;
  wire _09385_;
  wire _09386_;
  wire _09387_;
  wire _09388_;
  wire _09389_;
  wire _09390_;
  wire _09391_;
  wire _09392_;
  wire _09393_;
  wire _09394_;
  wire _09395_;
  wire _09396_;
  wire _09397_;
  wire _09398_;
  wire _09399_;
  wire _09400_;
  wire _09401_;
  wire _09402_;
  wire _09403_;
  wire _09404_;
  wire _09405_;
  wire _09406_;
  wire _09407_;
  wire _09408_;
  wire _09409_;
  wire _09410_;
  wire _09411_;
  wire _09412_;
  wire _09413_;
  wire _09414_;
  wire _09415_;
  wire _09416_;
  wire _09417_;
  wire _09418_;
  wire _09419_;
  wire _09420_;
  wire _09421_;
  wire _09422_;
  wire _09423_;
  wire _09424_;
  wire _09425_;
  wire _09426_;
  wire _09427_;
  wire _09428_;
  wire _09429_;
  wire _09430_;
  wire _09431_;
  wire _09432_;
  wire _09433_;
  wire _09434_;
  wire _09435_;
  wire _09436_;
  wire _09437_;
  wire _09438_;
  wire _09439_;
  wire _09440_;
  wire _09441_;
  wire _09442_;
  wire _09443_;
  wire _09444_;
  wire _09445_;
  wire _09446_;
  wire _09447_;
  wire _09448_;
  wire _09449_;
  wire _09450_;
  wire _09451_;
  wire _09452_;
  wire _09453_;
  wire _09454_;
  wire _09455_;
  wire _09456_;
  wire _09457_;
  wire _09458_;
  wire _09459_;
  wire _09460_;
  wire _09461_;
  wire _09462_;
  wire _09463_;
  wire _09464_;
  wire _09465_;
  wire _09466_;
  wire _09467_;
  wire _09468_;
  wire _09469_;
  wire _09470_;
  wire _09471_;
  wire _09472_;
  wire _09473_;
  wire _09474_;
  wire _09475_;
  wire _09476_;
  wire _09477_;
  wire _09478_;
  wire _09479_;
  wire _09480_;
  wire _09481_;
  wire _09482_;
  wire _09483_;
  wire _09484_;
  wire _09485_;
  wire _09486_;
  wire _09487_;
  wire _09488_;
  wire _09489_;
  wire _09490_;
  wire _09491_;
  wire _09492_;
  wire _09493_;
  wire _09494_;
  wire _09495_;
  wire _09496_;
  wire _09497_;
  wire _09498_;
  wire _09499_;
  wire _09500_;
  wire _09501_;
  wire _09502_;
  wire _09503_;
  wire _09504_;
  wire _09505_;
  wire _09506_;
  wire _09507_;
  wire _09508_;
  wire _09509_;
  wire _09510_;
  wire _09511_;
  wire _09512_;
  wire _09513_;
  wire _09514_;
  wire _09515_;
  wire _09516_;
  wire _09517_;
  wire _09518_;
  wire _09519_;
  wire _09520_;
  wire _09521_;
  wire _09522_;
  wire _09523_;
  wire _09524_;
  wire _09525_;
  wire _09526_;
  wire _09527_;
  wire _09528_;
  wire _09529_;
  wire _09530_;
  wire _09531_;
  wire _09532_;
  wire _09533_;
  wire _09534_;
  wire _09535_;
  wire _09536_;
  wire _09537_;
  wire _09538_;
  wire _09539_;
  wire _09540_;
  wire _09541_;
  wire _09542_;
  wire _09543_;
  wire _09544_;
  wire _09545_;
  wire _09546_;
  wire _09547_;
  wire _09548_;
  wire _09549_;
  wire _09550_;
  wire _09551_;
  wire _09552_;
  wire _09553_;
  wire _09554_;
  wire _09555_;
  wire _09556_;
  wire _09557_;
  wire _09558_;
  wire _09559_;
  wire _09560_;
  wire _09561_;
  wire _09562_;
  wire _09563_;
  wire _09564_;
  wire _09565_;
  wire _09566_;
  wire _09567_;
  wire _09568_;
  wire _09569_;
  wire _09570_;
  wire _09571_;
  wire _09572_;
  wire _09573_;
  wire _09574_;
  wire _09575_;
  wire _09576_;
  wire _09577_;
  wire _09578_;
  wire _09579_;
  wire _09580_;
  wire _09581_;
  wire _09582_;
  wire _09583_;
  wire _09584_;
  wire _09585_;
  wire _09586_;
  wire _09587_;
  wire _09588_;
  wire _09589_;
  wire _09590_;
  wire _09591_;
  wire _09592_;
  wire _09593_;
  wire _09594_;
  wire _09595_;
  wire _09596_;
  wire _09597_;
  wire _09598_;
  wire _09599_;
  wire _09600_;
  wire _09601_;
  wire _09602_;
  wire _09603_;
  wire _09604_;
  wire _09605_;
  wire _09606_;
  wire _09607_;
  wire _09608_;
  wire _09609_;
  wire _09610_;
  wire _09611_;
  wire _09612_;
  wire _09613_;
  wire _09614_;
  wire _09615_;
  wire _09616_;
  wire _09617_;
  wire _09618_;
  wire _09619_;
  wire _09620_;
  wire _09621_;
  wire _09622_;
  wire _09623_;
  wire _09624_;
  wire _09625_;
  wire _09626_;
  wire _09627_;
  wire _09628_;
  wire _09629_;
  wire _09630_;
  wire _09631_;
  wire _09632_;
  wire _09633_;
  wire _09634_;
  wire _09635_;
  wire _09636_;
  wire _09637_;
  wire _09638_;
  wire _09639_;
  wire _09640_;
  wire _09641_;
  wire _09642_;
  wire _09643_;
  wire _09644_;
  wire _09645_;
  wire _09646_;
  wire _09647_;
  wire _09648_;
  wire _09649_;
  wire _09650_;
  wire _09651_;
  wire _09652_;
  wire _09653_;
  wire _09654_;
  wire _09655_;
  wire _09656_;
  wire _09657_;
  wire _09658_;
  wire _09659_;
  wire _09660_;
  wire _09661_;
  wire _09662_;
  wire _09663_;
  wire _09664_;
  wire _09665_;
  wire _09666_;
  wire _09667_;
  wire _09668_;
  wire _09669_;
  wire _09670_;
  wire _09671_;
  wire _09672_;
  wire _09673_;
  wire _09674_;
  wire _09675_;
  wire _09676_;
  wire _09677_;
  wire _09678_;
  wire _09679_;
  wire _09680_;
  wire _09681_;
  wire _09682_;
  wire _09683_;
  wire _09684_;
  wire _09685_;
  wire _09686_;
  wire _09687_;
  wire _09688_;
  wire _09689_;
  wire _09690_;
  wire _09691_;
  wire _09692_;
  wire _09693_;
  wire _09694_;
  wire _09695_;
  wire _09696_;
  wire _09697_;
  wire _09698_;
  wire _09699_;
  wire _09700_;
  wire _09701_;
  wire _09702_;
  wire _09703_;
  wire _09704_;
  wire _09705_;
  wire _09706_;
  wire _09707_;
  wire _09708_;
  wire _09709_;
  wire _09710_;
  wire _09711_;
  wire _09712_;
  wire _09713_;
  wire _09714_;
  wire _09715_;
  wire _09716_;
  wire _09717_;
  wire _09718_;
  wire _09719_;
  wire _09720_;
  wire _09721_;
  wire _09722_;
  wire _09723_;
  wire _09724_;
  wire _09725_;
  wire _09726_;
  wire _09727_;
  wire _09728_;
  wire _09729_;
  wire _09730_;
  wire _09731_;
  wire _09732_;
  wire _09733_;
  wire _09734_;
  wire _09735_;
  wire _09736_;
  wire _09737_;
  wire _09738_;
  wire _09739_;
  wire _09740_;
  wire _09741_;
  wire _09742_;
  wire _09743_;
  wire _09744_;
  wire _09745_;
  wire _09746_;
  wire _09747_;
  wire _09748_;
  wire _09749_;
  wire _09750_;
  wire _09751_;
  wire _09752_;
  wire _09753_;
  wire _09754_;
  wire _09755_;
  wire _09756_;
  wire _09757_;
  wire _09758_;
  wire _09759_;
  wire _09760_;
  wire _09761_;
  wire _09762_;
  wire _09763_;
  wire _09764_;
  wire _09765_;
  wire _09766_;
  wire _09767_;
  wire _09768_;
  wire _09769_;
  wire _09770_;
  wire _09771_;
  wire _09772_;
  wire _09773_;
  wire _09774_;
  wire _09775_;
  wire _09776_;
  wire _09777_;
  wire _09778_;
  wire _09779_;
  wire _09780_;
  wire _09781_;
  wire _09782_;
  wire _09783_;
  wire _09784_;
  wire _09785_;
  wire _09786_;
  wire _09787_;
  wire _09788_;
  wire _09789_;
  wire _09790_;
  wire _09791_;
  wire _09792_;
  wire _09793_;
  wire _09794_;
  wire _09795_;
  wire _09796_;
  wire _09797_;
  wire _09798_;
  wire _09799_;
  wire _09800_;
  wire _09801_;
  wire _09802_;
  wire _09803_;
  wire _09804_;
  wire _09805_;
  wire _09806_;
  wire _09807_;
  wire _09808_;
  wire _09809_;
  wire _09810_;
  wire _09811_;
  wire _09812_;
  wire _09813_;
  wire _09814_;
  wire _09815_;
  wire _09816_;
  wire _09817_;
  wire _09818_;
  wire _09819_;
  wire _09820_;
  wire _09821_;
  wire _09822_;
  wire _09823_;
  wire _09824_;
  wire _09825_;
  wire _09826_;
  wire _09827_;
  wire _09828_;
  wire _09829_;
  wire _09830_;
  wire _09831_;
  wire _09832_;
  wire _09833_;
  wire _09834_;
  wire _09835_;
  wire _09836_;
  wire _09837_;
  wire _09838_;
  wire _09839_;
  wire _09840_;
  wire _09841_;
  wire _09842_;
  wire _09843_;
  wire _09844_;
  wire _09845_;
  wire _09846_;
  wire _09847_;
  wire _09848_;
  wire _09849_;
  wire _09850_;
  wire _09851_;
  wire _09852_;
  wire _09853_;
  wire _09854_;
  wire _09855_;
  wire _09856_;
  wire _09857_;
  wire _09858_;
  wire _09859_;
  wire _09860_;
  wire _09861_;
  wire _09862_;
  wire _09863_;
  wire _09864_;
  wire _09865_;
  wire _09866_;
  wire _09867_;
  wire _09868_;
  wire _09869_;
  wire _09870_;
  wire _09871_;
  wire _09872_;
  wire _09873_;
  wire _09874_;
  wire _09875_;
  wire _09876_;
  wire _09877_;
  wire _09878_;
  wire _09879_;
  wire _09880_;
  wire _09881_;
  wire _09882_;
  wire _09883_;
  wire _09884_;
  wire _09885_;
  wire _09886_;
  wire _09887_;
  wire _09888_;
  wire _09889_;
  wire _09890_;
  wire _09891_;
  wire _09892_;
  wire _09893_;
  wire _09894_;
  wire _09895_;
  wire _09896_;
  wire _09897_;
  wire _09898_;
  wire _09899_;
  wire _09900_;
  wire _09901_;
  wire _09902_;
  wire _09903_;
  wire _09904_;
  wire _09905_;
  wire _09906_;
  wire _09907_;
  wire _09908_;
  wire _09909_;
  wire _09910_;
  wire _09911_;
  wire _09912_;
  wire _09913_;
  wire _09914_;
  wire _09915_;
  wire _09916_;
  wire _09917_;
  wire _09918_;
  wire _09919_;
  wire _09920_;
  wire _09921_;
  wire _09922_;
  wire _09923_;
  wire _09924_;
  wire _09925_;
  wire _09926_;
  wire _09927_;
  wire _09928_;
  wire _09929_;
  wire _09930_;
  wire _09931_;
  wire _09932_;
  wire _09933_;
  wire _09934_;
  wire _09935_;
  wire _09936_;
  wire _09937_;
  wire _09938_;
  wire _09939_;
  wire _09940_;
  wire _09941_;
  wire _09942_;
  wire _09943_;
  wire _09944_;
  wire _09945_;
  wire _09946_;
  wire _09947_;
  wire _09948_;
  wire _09949_;
  wire _09950_;
  wire _09951_;
  wire _09952_;
  wire _09953_;
  wire _09954_;
  wire _09955_;
  wire _09956_;
  wire _09957_;
  wire _09958_;
  wire _09959_;
  wire _09960_;
  wire _09961_;
  wire _09962_;
  wire _09963_;
  wire _09964_;
  wire _09965_;
  wire _09966_;
  wire _09967_;
  wire _09968_;
  wire _09969_;
  wire _09970_;
  wire _09971_;
  wire _09972_;
  wire _09973_;
  wire _09974_;
  wire _09975_;
  wire _09976_;
  wire _09977_;
  wire _09978_;
  wire _09979_;
  wire _09980_;
  wire _09981_;
  wire _09982_;
  wire _09983_;
  wire _09984_;
  wire _09985_;
  wire _09986_;
  wire _09987_;
  wire _09988_;
  wire _09989_;
  wire _09990_;
  wire _09991_;
  wire _09992_;
  wire _09993_;
  wire _09994_;
  wire _09995_;
  wire _09996_;
  wire _09997_;
  wire _09998_;
  wire _09999_;
  wire _10000_;
  wire _10001_;
  wire _10002_;
  wire _10003_;
  wire _10004_;
  wire _10005_;
  wire _10006_;
  wire _10007_;
  wire _10008_;
  wire _10009_;
  wire _10010_;
  wire _10011_;
  wire _10012_;
  wire _10013_;
  wire _10014_;
  wire _10015_;
  wire _10016_;
  wire _10017_;
  wire _10018_;
  wire _10019_;
  wire _10020_;
  wire _10021_;
  wire _10022_;
  wire _10023_;
  wire _10024_;
  wire _10025_;
  wire _10026_;
  wire _10027_;
  wire _10028_;
  wire _10029_;
  wire _10030_;
  wire _10031_;
  wire _10032_;
  wire _10033_;
  wire _10034_;
  wire _10035_;
  wire _10036_;
  wire _10037_;
  wire _10038_;
  wire _10039_;
  wire _10040_;
  wire _10041_;
  wire _10042_;
  wire _10043_;
  wire _10044_;
  wire _10045_;
  wire _10046_;
  wire _10047_;
  wire _10048_;
  wire _10049_;
  wire _10050_;
  wire _10051_;
  wire _10052_;
  wire _10053_;
  wire _10054_;
  wire _10055_;
  wire _10056_;
  wire _10057_;
  wire _10058_;
  wire _10059_;
  wire _10060_;
  wire _10061_;
  wire _10062_;
  wire _10063_;
  wire _10064_;
  wire _10065_;
  wire _10066_;
  wire _10067_;
  wire _10068_;
  wire _10069_;
  wire _10070_;
  wire _10071_;
  wire _10072_;
  wire _10073_;
  wire _10074_;
  wire _10075_;
  wire _10076_;
  wire _10077_;
  wire _10078_;
  wire _10079_;
  wire _10080_;
  wire _10081_;
  wire _10082_;
  wire _10083_;
  wire _10084_;
  wire _10085_;
  wire _10086_;
  wire _10087_;
  wire _10088_;
  wire _10089_;
  wire _10090_;
  wire _10091_;
  wire _10092_;
  wire _10093_;
  wire _10094_;
  wire _10095_;
  wire _10096_;
  wire _10097_;
  wire _10098_;
  wire _10099_;
  wire _10100_;
  wire _10101_;
  wire _10102_;
  wire _10103_;
  wire _10104_;
  wire _10105_;
  wire _10106_;
  wire _10107_;
  wire _10108_;
  wire _10109_;
  wire _10110_;
  wire _10111_;
  wire _10112_;
  wire _10113_;
  wire _10114_;
  wire _10115_;
  wire _10116_;
  wire _10117_;
  wire _10118_;
  wire _10119_;
  wire _10120_;
  wire _10121_;
  wire _10122_;
  wire _10123_;
  wire _10124_;
  wire _10125_;
  wire _10126_;
  wire _10127_;
  wire _10128_;
  wire _10129_;
  wire _10130_;
  wire _10131_;
  wire _10132_;
  wire _10133_;
  wire _10134_;
  wire _10135_;
  wire _10136_;
  wire _10137_;
  wire _10138_;
  wire _10139_;
  wire _10140_;
  wire _10141_;
  wire _10142_;
  wire _10143_;
  wire _10144_;
  wire _10145_;
  wire _10146_;
  wire _10147_;
  wire _10148_;
  wire _10149_;
  wire _10150_;
  wire _10151_;
  wire _10152_;
  wire _10153_;
  wire _10154_;
  wire _10155_;
  wire _10156_;
  wire _10157_;
  wire _10158_;
  wire _10159_;
  wire _10160_;
  wire _10161_;
  wire _10162_;
  wire _10163_;
  wire _10164_;
  wire _10165_;
  wire _10166_;
  wire _10167_;
  wire _10168_;
  wire _10169_;
  wire _10170_;
  wire _10171_;
  wire _10172_;
  wire _10173_;
  wire _10174_;
  wire _10175_;
  wire _10176_;
  wire _10177_;
  wire _10178_;
  wire _10179_;
  wire _10180_;
  wire _10181_;
  wire _10182_;
  wire _10183_;
  wire _10184_;
  wire _10185_;
  wire _10186_;
  wire _10187_;
  wire _10188_;
  wire _10189_;
  wire _10190_;
  wire _10191_;
  wire _10192_;
  wire _10193_;
  wire _10194_;
  wire _10195_;
  wire _10196_;
  wire _10197_;
  wire _10198_;
  wire _10199_;
  wire _10200_;
  wire _10201_;
  wire _10202_;
  wire _10203_;
  wire _10204_;
  wire _10205_;
  wire _10206_;
  wire _10207_;
  wire _10208_;
  wire _10209_;
  wire _10210_;
  wire _10211_;
  wire _10212_;
  wire _10213_;
  wire _10214_;
  wire _10215_;
  wire _10216_;
  wire _10217_;
  wire _10218_;
  wire _10219_;
  wire _10220_;
  wire _10221_;
  wire _10222_;
  wire _10223_;
  wire _10224_;
  wire _10225_;
  wire _10226_;
  wire _10227_;
  wire _10228_;
  wire _10229_;
  wire _10230_;
  wire _10231_;
  wire _10232_;
  wire _10233_;
  wire _10234_;
  wire _10235_;
  wire _10236_;
  wire _10237_;
  wire _10238_;
  wire _10239_;
  wire _10240_;
  wire _10241_;
  wire _10242_;
  wire _10243_;
  wire _10244_;
  wire _10245_;
  wire _10246_;
  wire _10247_;
  wire _10248_;
  wire _10249_;
  wire _10250_;
  wire _10251_;
  wire _10252_;
  wire _10253_;
  wire _10254_;
  wire _10255_;
  wire _10256_;
  wire _10257_;
  wire _10258_;
  wire _10259_;
  wire _10260_;
  wire _10261_;
  wire _10262_;
  wire _10263_;
  wire _10264_;
  wire _10265_;
  wire _10266_;
  wire _10267_;
  wire _10268_;
  wire _10269_;
  wire _10270_;
  wire _10271_;
  wire _10272_;
  wire _10273_;
  wire _10274_;
  wire _10275_;
  wire _10276_;
  wire _10277_;
  wire _10278_;
  wire _10279_;
  wire _10280_;
  wire _10281_;
  wire _10282_;
  wire _10283_;
  wire _10284_;
  wire _10285_;
  wire _10286_;
  wire _10287_;
  wire _10288_;
  wire _10289_;
  wire _10290_;
  wire _10291_;
  wire _10292_;
  wire _10293_;
  wire _10294_;
  wire _10295_;
  wire _10296_;
  wire _10297_;
  wire _10298_;
  wire _10299_;
  wire _10300_;
  wire _10301_;
  wire _10302_;
  wire _10303_;
  wire _10304_;
  wire _10305_;
  wire _10306_;
  wire _10307_;
  wire _10308_;
  wire _10309_;
  wire _10310_;
  wire _10311_;
  wire _10312_;
  wire _10313_;
  wire _10314_;
  wire _10315_;
  wire _10316_;
  wire _10317_;
  wire _10318_;
  wire _10319_;
  wire _10320_;
  wire _10321_;
  wire _10322_;
  wire _10323_;
  wire _10324_;
  wire _10325_;
  wire _10326_;
  wire _10327_;
  wire _10328_;
  wire _10329_;
  wire _10330_;
  wire _10331_;
  wire _10332_;
  wire _10333_;
  wire _10334_;
  wire _10335_;
  wire _10336_;
  wire _10337_;
  wire _10338_;
  wire _10339_;
  wire _10340_;
  wire _10341_;
  wire _10342_;
  wire _10343_;
  wire _10344_;
  wire _10345_;
  wire _10346_;
  wire _10347_;
  wire _10348_;
  wire _10349_;
  wire _10350_;
  wire _10351_;
  wire _10352_;
  wire _10353_;
  wire _10354_;
  wire _10355_;
  wire _10356_;
  wire _10357_;
  wire _10358_;
  wire _10359_;
  wire _10360_;
  wire _10361_;
  wire _10362_;
  wire _10363_;
  wire _10364_;
  wire _10365_;
  wire _10366_;
  wire _10367_;
  wire _10368_;
  wire _10369_;
  wire _10370_;
  wire _10371_;
  wire _10372_;
  wire _10373_;
  wire _10374_;
  wire _10375_;
  wire _10376_;
  wire _10377_;
  wire _10378_;
  wire _10379_;
  wire _10380_;
  wire _10381_;
  wire _10382_;
  wire _10383_;
  wire _10384_;
  wire _10385_;
  wire _10386_;
  wire _10387_;
  wire _10388_;
  wire _10389_;
  wire _10390_;
  wire _10391_;
  wire _10392_;
  wire _10393_;
  wire _10394_;
  wire _10395_;
  wire _10396_;
  wire _10397_;
  wire _10398_;
  wire _10399_;
  wire _10400_;
  wire _10401_;
  wire _10402_;
  wire _10403_;
  wire _10404_;
  wire _10405_;
  wire _10406_;
  wire _10407_;
  wire _10408_;
  wire _10409_;
  wire _10410_;
  wire _10411_;
  wire _10412_;
  wire _10413_;
  wire _10414_;
  wire _10415_;
  wire _10416_;
  wire _10417_;
  wire _10418_;
  wire _10419_;
  wire _10420_;
  wire _10421_;
  wire _10422_;
  wire _10423_;
  wire _10424_;
  wire _10425_;
  wire _10426_;
  wire _10427_;
  wire _10428_;
  wire _10429_;
  wire _10430_;
  wire _10431_;
  wire _10432_;
  wire _10433_;
  wire _10434_;
  wire _10435_;
  wire _10436_;
  wire _10437_;
  wire _10438_;
  wire _10439_;
  wire _10440_;
  wire _10441_;
  wire _10442_;
  wire _10443_;
  wire _10444_;
  wire _10445_;
  wire _10446_;
  wire _10447_;
  wire _10448_;
  wire _10449_;
  wire _10450_;
  wire _10451_;
  wire _10452_;
  wire _10453_;
  wire _10454_;
  wire _10455_;
  wire _10456_;
  wire _10457_;
  wire _10458_;
  wire _10459_;
  wire _10460_;
  wire _10461_;
  wire _10462_;
  wire _10463_;
  wire _10464_;
  wire _10465_;
  wire _10466_;
  wire _10467_;
  wire _10468_;
  wire _10469_;
  wire _10470_;
  wire _10471_;
  wire _10472_;
  wire _10473_;
  wire _10474_;
  wire _10475_;
  wire _10476_;
  wire _10477_;
  wire _10478_;
  wire _10479_;
  wire _10480_;
  wire _10481_;
  wire _10482_;
  wire _10483_;
  wire _10484_;
  wire _10485_;
  wire _10486_;
  wire _10487_;
  wire _10488_;
  wire _10489_;
  wire _10490_;
  wire _10491_;
  wire _10492_;
  wire _10493_;
  wire _10494_;
  wire _10495_;
  wire _10496_;
  wire _10497_;
  wire _10498_;
  wire _10499_;
  wire _10500_;
  wire _10501_;
  wire _10502_;
  wire _10503_;
  wire _10504_;
  wire _10505_;
  wire _10506_;
  wire _10507_;
  wire _10508_;
  wire _10509_;
  wire _10510_;
  wire _10511_;
  wire _10512_;
  wire _10513_;
  wire _10514_;
  wire _10515_;
  wire _10516_;
  wire _10517_;
  wire _10518_;
  wire _10519_;
  wire _10520_;
  wire _10521_;
  wire _10522_;
  wire _10523_;
  wire _10524_;
  wire _10525_;
  wire _10526_;
  wire _10527_;
  wire _10528_;
  wire _10529_;
  wire _10530_;
  wire _10531_;
  wire _10532_;
  wire _10533_;
  wire _10534_;
  wire _10535_;
  wire _10536_;
  wire _10537_;
  wire _10538_;
  wire _10539_;
  wire _10540_;
  wire _10541_;
  wire _10542_;
  wire _10543_;
  wire _10544_;
  wire _10545_;
  wire _10546_;
  wire _10547_;
  wire _10548_;
  wire _10549_;
  wire _10550_;
  wire _10551_;
  wire _10552_;
  wire _10553_;
  wire _10554_;
  wire _10555_;
  wire _10556_;
  wire _10557_;
  wire _10558_;
  wire _10559_;
  wire _10560_;
  wire _10561_;
  wire _10562_;
  wire _10563_;
  wire _10564_;
  wire _10565_;
  wire _10566_;
  wire _10567_;
  wire _10568_;
  wire _10569_;
  wire _10570_;
  wire _10571_;
  wire _10572_;
  wire _10573_;
  wire _10574_;
  wire _10575_;
  wire _10576_;
  wire _10577_;
  wire _10578_;
  wire _10579_;
  wire _10580_;
  wire _10581_;
  wire _10582_;
  wire _10583_;
  wire _10584_;
  wire _10585_;
  wire _10586_;
  wire _10587_;
  wire _10588_;
  wire _10589_;
  wire _10590_;
  wire _10591_;
  wire _10592_;
  wire _10593_;
  wire _10594_;
  wire _10595_;
  wire _10596_;
  wire _10597_;
  wire _10598_;
  wire _10599_;
  wire _10600_;
  wire _10601_;
  wire _10602_;
  wire _10603_;
  wire _10604_;
  wire _10605_;
  wire _10606_;
  wire _10607_;
  wire _10608_;
  wire _10609_;
  wire _10610_;
  wire _10611_;
  wire _10612_;
  wire _10613_;
  wire _10614_;
  wire _10615_;
  wire _10616_;
  wire _10617_;
  wire _10618_;
  wire _10619_;
  wire _10620_;
  wire _10621_;
  wire _10622_;
  wire _10623_;
  wire _10624_;
  wire _10625_;
  wire _10626_;
  wire _10627_;
  wire _10628_;
  wire _10629_;
  wire _10630_;
  wire _10631_;
  wire _10632_;
  wire _10633_;
  wire _10634_;
  wire _10635_;
  wire _10636_;
  wire _10637_;
  wire _10638_;
  wire _10639_;
  wire _10640_;
  wire _10641_;
  wire _10642_;
  wire _10643_;
  wire _10644_;
  wire _10645_;
  wire _10646_;
  wire _10647_;
  wire _10648_;
  wire _10649_;
  wire _10650_;
  wire _10651_;
  wire _10652_;
  wire _10653_;
  wire _10654_;
  wire _10655_;
  wire _10656_;
  wire _10657_;
  wire _10658_;
  wire _10659_;
  wire _10660_;
  wire _10661_;
  wire _10662_;
  wire _10663_;
  wire _10664_;
  wire _10665_;
  wire _10666_;
  wire _10667_;
  wire _10668_;
  wire _10669_;
  wire _10670_;
  wire _10671_;
  wire _10672_;
  wire _10673_;
  wire _10674_;
  wire _10675_;
  wire _10676_;
  wire _10677_;
  wire _10678_;
  wire _10679_;
  wire _10680_;
  wire _10681_;
  wire _10682_;
  wire _10683_;
  wire _10684_;
  wire _10685_;
  wire _10686_;
  wire _10687_;
  wire _10688_;
  wire _10689_;
  wire _10690_;
  wire _10691_;
  wire _10692_;
  wire _10693_;
  wire _10694_;
  wire _10695_;
  wire _10696_;
  wire _10697_;
  wire _10698_;
  wire _10699_;
  wire _10700_;
  wire _10701_;
  wire _10702_;
  wire _10703_;
  wire _10704_;
  wire _10705_;
  wire _10706_;
  wire _10707_;
  wire _10708_;
  wire _10709_;
  wire _10710_;
  wire _10711_;
  wire _10712_;
  wire _10713_;
  wire _10714_;
  wire _10715_;
  wire _10716_;
  wire _10717_;
  wire _10718_;
  wire _10719_;
  wire _10720_;
  wire _10721_;
  wire _10722_;
  wire _10723_;
  wire _10724_;
  wire _10725_;
  wire _10726_;
  wire _10727_;
  wire _10728_;
  wire _10729_;
  wire _10730_;
  wire _10731_;
  wire _10732_;
  wire _10733_;
  wire _10734_;
  wire _10735_;
  wire _10736_;
  wire _10737_;
  wire _10738_;
  wire _10739_;
  wire _10740_;
  wire _10741_;
  wire _10742_;
  wire _10743_;
  wire _10744_;
  wire _10745_;
  wire _10746_;
  wire _10747_;
  wire _10748_;
  wire _10749_;
  wire _10750_;
  wire _10751_;
  wire _10752_;
  wire _10753_;
  wire _10754_;
  wire _10755_;
  wire _10756_;
  wire _10757_;
  wire _10758_;
  wire _10759_;
  wire _10760_;
  wire _10761_;
  wire _10762_;
  wire _10763_;
  wire _10764_;
  wire _10765_;
  wire _10766_;
  wire _10767_;
  wire _10768_;
  wire _10769_;
  wire _10770_;
  wire _10771_;
  wire _10772_;
  wire _10773_;
  wire _10774_;
  wire _10775_;
  wire _10776_;
  wire _10777_;
  wire _10778_;
  wire _10779_;
  wire _10780_;
  wire _10781_;
  wire _10782_;
  wire _10783_;
  wire _10784_;
  wire _10785_;
  wire _10786_;
  wire _10787_;
  wire _10788_;
  wire _10789_;
  wire _10790_;
  wire _10791_;
  wire _10792_;
  wire _10793_;
  wire _10794_;
  wire _10795_;
  wire _10796_;
  wire _10797_;
  wire _10798_;
  wire _10799_;
  wire _10800_;
  wire _10801_;
  wire _10802_;
  wire _10803_;
  wire _10804_;
  wire _10805_;
  wire _10806_;
  wire _10807_;
  wire _10808_;
  wire _10809_;
  wire _10810_;
  wire _10811_;
  wire _10812_;
  wire _10813_;
  wire _10814_;
  wire _10815_;
  wire _10816_;
  wire _10817_;
  wire _10818_;
  wire _10819_;
  wire _10820_;
  wire _10821_;
  wire _10822_;
  wire _10823_;
  wire _10824_;
  wire _10825_;
  wire _10826_;
  wire _10827_;
  wire _10828_;
  wire _10829_;
  wire _10830_;
  wire _10831_;
  wire _10832_;
  wire _10833_;
  wire _10834_;
  wire _10835_;
  wire _10836_;
  wire _10837_;
  wire _10838_;
  wire _10839_;
  wire _10840_;
  wire _10841_;
  wire _10842_;
  wire _10843_;
  wire _10844_;
  wire _10845_;
  wire _10846_;
  wire _10847_;
  wire _10848_;
  wire _10849_;
  wire _10850_;
  wire _10851_;
  wire _10852_;
  wire _10853_;
  wire _10854_;
  wire _10855_;
  wire _10856_;
  wire _10857_;
  wire _10858_;
  wire _10859_;
  wire _10860_;
  wire _10861_;
  wire _10862_;
  wire _10863_;
  wire _10864_;
  wire _10865_;
  wire _10866_;
  wire _10867_;
  wire _10868_;
  wire _10869_;
  wire _10870_;
  wire _10871_;
  wire _10872_;
  wire _10873_;
  wire _10874_;
  wire _10875_;
  wire _10876_;
  wire _10877_;
  wire _10878_;
  wire _10879_;
  wire _10880_;
  wire _10881_;
  wire _10882_;
  wire _10883_;
  wire _10884_;
  wire _10885_;
  wire _10886_;
  wire _10887_;
  wire _10888_;
  wire _10889_;
  wire _10890_;
  wire _10891_;
  wire _10892_;
  wire _10893_;
  wire _10894_;
  wire _10895_;
  wire _10896_;
  wire _10897_;
  wire _10898_;
  wire _10899_;
  wire _10900_;
  wire _10901_;
  wire _10902_;
  wire _10903_;
  wire _10904_;
  wire _10905_;
  wire _10906_;
  wire _10907_;
  wire _10908_;
  wire _10909_;
  wire _10910_;
  wire _10911_;
  wire _10912_;
  wire _10913_;
  wire _10914_;
  wire _10915_;
  wire _10916_;
  wire _10917_;
  wire _10918_;
  wire _10919_;
  wire _10920_;
  wire _10921_;
  wire _10922_;
  wire _10923_;
  wire _10924_;
  wire _10925_;
  wire _10926_;
  wire _10927_;
  wire _10928_;
  wire _10929_;
  wire _10930_;
  wire _10931_;
  wire _10932_;
  wire _10933_;
  wire _10934_;
  wire _10935_;
  wire _10936_;
  wire _10937_;
  wire _10938_;
  wire _10939_;
  wire _10940_;
  wire _10941_;
  wire _10942_;
  wire _10943_;
  wire _10944_;
  wire _10945_;
  wire _10946_;
  wire _10947_;
  wire _10948_;
  wire _10949_;
  wire _10950_;
  wire _10951_;
  wire _10952_;
  wire _10953_;
  wire _10954_;
  wire _10955_;
  wire _10956_;
  wire _10957_;
  wire _10958_;
  wire _10959_;
  wire _10960_;
  wire _10961_;
  wire _10962_;
  wire _10963_;
  wire _10964_;
  wire _10965_;
  wire _10966_;
  wire _10967_;
  wire _10968_;
  wire _10969_;
  wire _10970_;
  wire _10971_;
  wire _10972_;
  wire _10973_;
  wire _10974_;
  wire _10975_;
  wire _10976_;
  wire _10977_;
  wire _10978_;
  wire _10979_;
  wire _10980_;
  wire _10981_;
  wire _10982_;
  wire _10983_;
  wire _10984_;
  wire _10985_;
  wire _10986_;
  wire _10987_;
  wire _10988_;
  wire _10989_;
  wire _10990_;
  wire _10991_;
  wire _10992_;
  wire _10993_;
  wire _10994_;
  wire _10995_;
  wire _10996_;
  wire _10997_;
  wire _10998_;
  wire _10999_;
  wire _11000_;
  wire _11001_;
  wire _11002_;
  wire _11003_;
  wire _11004_;
  wire _11005_;
  wire _11006_;
  wire _11007_;
  wire _11008_;
  wire _11009_;
  wire _11010_;
  wire _11011_;
  wire _11012_;
  wire _11013_;
  wire _11014_;
  wire _11015_;
  wire _11016_;
  wire _11017_;
  wire _11018_;
  wire _11019_;
  wire _11020_;
  wire _11021_;
  wire _11022_;
  wire _11023_;
  wire _11024_;
  wire _11025_;
  wire _11026_;
  wire _11027_;
  wire _11028_;
  wire _11029_;
  wire _11030_;
  wire _11031_;
  wire _11032_;
  wire _11033_;
  wire _11034_;
  wire _11035_;
  wire _11036_;
  wire _11037_;
  wire _11038_;
  wire _11039_;
  wire _11040_;
  wire _11041_;
  wire _11042_;
  wire _11043_;
  wire _11044_;
  wire _11045_;
  wire _11046_;
  wire _11047_;
  wire _11048_;
  wire _11049_;
  wire _11050_;
  wire _11051_;
  wire _11052_;
  wire _11053_;
  wire _11054_;
  wire _11055_;
  wire _11056_;
  wire _11057_;
  wire _11058_;
  wire _11059_;
  wire _11060_;
  wire _11061_;
  wire _11062_;
  wire _11063_;
  wire _11064_;
  wire _11065_;
  wire _11066_;
  wire _11067_;
  wire _11068_;
  wire _11069_;
  wire _11070_;
  wire _11071_;
  wire _11072_;
  wire _11073_;
  wire _11074_;
  wire _11075_;
  wire _11076_;
  wire _11077_;
  wire _11078_;
  wire _11079_;
  wire _11080_;
  wire _11081_;
  wire _11082_;
  wire _11083_;
  wire _11084_;
  wire _11085_;
  wire _11086_;
  wire _11087_;
  wire _11088_;
  wire _11089_;
  wire _11090_;
  wire _11091_;
  wire _11092_;
  wire _11093_;
  wire _11094_;
  wire _11095_;
  wire _11096_;
  wire _11097_;
  wire _11098_;
  wire _11099_;
  wire _11100_;
  wire _11101_;
  wire _11102_;
  wire _11103_;
  wire _11104_;
  wire _11105_;
  wire _11106_;
  wire _11107_;
  wire _11108_;
  wire _11109_;
  wire _11110_;
  wire _11111_;
  wire _11112_;
  wire _11113_;
  wire _11114_;
  wire _11115_;
  wire _11116_;
  wire _11117_;
  wire _11118_;
  wire _11119_;
  wire _11120_;
  wire _11121_;
  wire _11122_;
  wire _11123_;
  wire _11124_;
  wire _11125_;
  wire _11126_;
  wire _11127_;
  wire _11128_;
  wire _11129_;
  wire _11130_;
  wire _11131_;
  wire _11132_;
  wire _11133_;
  wire _11134_;
  wire _11135_;
  wire _11136_;
  wire _11137_;
  wire _11138_;
  wire _11139_;
  wire _11140_;
  wire _11141_;
  wire _11142_;
  wire _11143_;
  wire _11144_;
  wire _11145_;
  wire _11146_;
  wire _11147_;
  wire _11148_;
  wire _11149_;
  wire _11150_;
  wire _11151_;
  wire _11152_;
  wire _11153_;
  wire _11154_;
  wire _11155_;
  wire _11156_;
  wire _11157_;
  wire _11158_;
  wire _11159_;
  wire _11160_;
  wire _11161_;
  wire _11162_;
  wire _11163_;
  wire _11164_;
  wire _11165_;
  wire _11166_;
  wire _11167_;
  wire _11168_;
  wire _11169_;
  wire _11170_;
  wire _11171_;
  wire _11172_;
  wire _11173_;
  wire _11174_;
  wire _11175_;
  wire _11176_;
  wire _11177_;
  wire _11178_;
  wire _11179_;
  wire _11180_;
  wire _11181_;
  wire _11182_;
  wire _11183_;
  wire _11184_;
  wire _11185_;
  wire _11186_;
  wire _11187_;
  wire _11188_;
  wire _11189_;
  wire _11190_;
  wire _11191_;
  wire _11192_;
  wire _11193_;
  wire _11194_;
  wire _11195_;
  wire _11196_;
  wire _11197_;
  wire _11198_;
  wire _11199_;
  wire _11200_;
  wire _11201_;
  wire _11202_;
  wire _11203_;
  wire _11204_;
  wire _11205_;
  wire _11206_;
  wire _11207_;
  wire _11208_;
  wire _11209_;
  wire _11210_;
  wire _11211_;
  wire _11212_;
  wire _11213_;
  wire _11214_;
  wire _11215_;
  wire _11216_;
  wire _11217_;
  wire _11218_;
  wire _11219_;
  wire _11220_;
  wire _11221_;
  wire _11222_;
  wire _11223_;
  wire _11224_;
  wire _11225_;
  wire _11226_;
  wire _11227_;
  wire _11228_;
  wire _11229_;
  wire _11230_;
  wire _11231_;
  wire _11232_;
  wire _11233_;
  wire _11234_;
  wire _11235_;
  wire _11236_;
  wire _11237_;
  wire _11238_;
  wire _11239_;
  wire _11240_;
  wire _11241_;
  wire _11242_;
  wire _11243_;
  wire _11244_;
  wire _11245_;
  wire _11246_;
  wire _11247_;
  wire _11248_;
  wire _11249_;
  wire _11250_;
  wire _11251_;
  wire _11252_;
  wire _11253_;
  wire _11254_;
  wire _11255_;
  wire _11256_;
  wire _11257_;
  wire _11258_;
  wire _11259_;
  wire _11260_;
  wire _11261_;
  wire _11262_;
  wire _11263_;
  wire _11264_;
  wire _11265_;
  wire _11266_;
  wire _11267_;
  wire _11268_;
  wire _11269_;
  wire _11270_;
  wire _11271_;
  wire _11272_;
  wire _11273_;
  wire _11274_;
  wire _11275_;
  wire _11276_;
  wire _11277_;
  wire _11278_;
  wire _11279_;
  wire _11280_;
  wire _11281_;
  wire _11282_;
  wire _11283_;
  wire _11284_;
  wire _11285_;
  wire _11286_;
  wire _11287_;
  wire _11288_;
  wire _11289_;
  wire _11290_;
  wire _11291_;
  wire _11292_;
  wire _11293_;
  wire _11294_;
  wire _11295_;
  wire _11296_;
  wire _11297_;
  wire _11298_;
  wire _11299_;
  wire _11300_;
  wire _11301_;
  wire _11302_;
  wire _11303_;
  wire _11304_;
  wire _11305_;
  wire _11306_;
  wire _11307_;
  wire _11308_;
  wire _11309_;
  wire _11310_;
  wire _11311_;
  wire _11312_;
  wire _11313_;
  wire _11314_;
  wire _11315_;
  wire _11316_;
  wire _11317_;
  wire _11318_;
  wire _11319_;
  wire _11320_;
  wire _11321_;
  wire _11322_;
  wire _11323_;
  wire _11324_;
  wire _11325_;
  wire _11326_;
  wire _11327_;
  wire _11328_;
  wire _11329_;
  wire _11330_;
  wire _11331_;
  wire _11332_;
  wire _11333_;
  wire _11334_;
  wire _11335_;
  wire _11336_;
  wire _11337_;
  wire _11338_;
  wire _11339_;
  wire _11340_;
  wire _11341_;
  wire _11342_;
  wire _11343_;
  wire _11344_;
  wire _11345_;
  wire _11346_;
  wire _11347_;
  wire _11348_;
  wire _11349_;
  wire _11350_;
  wire _11351_;
  wire _11352_;
  wire _11353_;
  wire _11354_;
  wire _11355_;
  wire _11356_;
  wire _11357_;
  wire _11358_;
  wire _11359_;
  wire _11360_;
  wire _11361_;
  wire _11362_;
  wire _11363_;
  wire _11364_;
  wire _11365_;
  wire _11366_;
  wire _11367_;
  wire _11368_;
  wire _11369_;
  wire _11370_;
  wire _11371_;
  wire _11372_;
  wire _11373_;
  wire _11374_;
  wire _11375_;
  wire _11376_;
  wire _11377_;
  wire _11378_;
  wire _11379_;
  wire _11380_;
  wire _11381_;
  wire _11382_;
  wire _11383_;
  wire _11384_;
  wire _11385_;
  wire _11386_;
  wire _11387_;
  wire _11388_;
  wire _11389_;
  wire _11390_;
  wire _11391_;
  wire _11392_;
  wire _11393_;
  wire _11394_;
  wire _11395_;
  wire _11396_;
  wire _11397_;
  wire _11398_;
  wire _11399_;
  wire _11400_;
  wire _11401_;
  wire _11402_;
  wire _11403_;
  wire _11404_;
  wire _11405_;
  wire _11406_;
  wire _11407_;
  wire _11408_;
  wire _11409_;
  wire _11410_;
  wire _11411_;
  wire _11412_;
  wire _11413_;
  wire _11414_;
  wire _11415_;
  wire _11416_;
  wire _11417_;
  wire _11418_;
  wire _11419_;
  wire _11420_;
  wire _11421_;
  wire _11422_;
  wire _11423_;
  wire _11424_;
  wire _11425_;
  wire _11426_;
  wire _11427_;
  wire _11428_;
  wire _11429_;
  wire _11430_;
  wire _11431_;
  wire _11432_;
  wire _11433_;
  wire _11434_;
  wire _11435_;
  wire _11436_;
  wire _11437_;
  wire _11438_;
  wire _11439_;
  wire _11440_;
  wire _11441_;
  wire _11442_;
  wire _11443_;
  wire _11444_;
  wire _11445_;
  wire _11446_;
  wire _11447_;
  wire _11448_;
  wire _11449_;
  wire _11450_;
  wire _11451_;
  wire _11452_;
  wire _11453_;
  wire _11454_;
  wire _11455_;
  wire _11456_;
  wire _11457_;
  wire _11458_;
  wire _11459_;
  wire _11460_;
  wire _11461_;
  wire _11462_;
  wire _11463_;
  wire _11464_;
  wire _11465_;
  wire _11466_;
  wire _11467_;
  wire _11468_;
  wire _11469_;
  wire _11470_;
  wire _11471_;
  wire _11472_;
  wire _11473_;
  wire _11474_;
  wire _11475_;
  wire _11476_;
  wire _11477_;
  wire _11478_;
  wire _11479_;
  wire _11480_;
  wire _11481_;
  wire _11482_;
  wire _11483_;
  wire _11484_;
  wire _11485_;
  wire _11486_;
  wire _11487_;
  wire _11488_;
  wire _11489_;
  wire _11490_;
  wire _11491_;
  wire _11492_;
  wire _11493_;
  wire _11494_;
  wire _11495_;
  wire _11496_;
  wire _11497_;
  wire _11498_;
  wire _11499_;
  wire _11500_;
  wire _11501_;
  wire _11502_;
  wire _11503_;
  wire _11504_;
  wire _11505_;
  wire _11506_;
  wire _11507_;
  wire _11508_;
  wire _11509_;
  wire _11510_;
  wire _11511_;
  wire _11512_;
  wire _11513_;
  wire _11514_;
  wire _11515_;
  wire _11516_;
  wire _11517_;
  wire _11518_;
  wire _11519_;
  wire _11520_;
  wire _11521_;
  wire _11522_;
  wire _11523_;
  wire _11524_;
  wire _11525_;
  wire _11526_;
  wire _11527_;
  wire _11528_;
  wire _11529_;
  wire _11530_;
  wire _11531_;
  wire _11532_;
  wire _11533_;
  wire _11534_;
  wire _11535_;
  wire _11536_;
  wire _11537_;
  wire _11538_;
  wire _11539_;
  wire _11540_;
  wire _11541_;
  wire _11542_;
  wire _11543_;
  wire _11544_;
  wire _11545_;
  wire _11546_;
  wire _11547_;
  wire _11548_;
  wire _11549_;
  wire _11550_;
  wire _11551_;
  wire _11552_;
  wire _11553_;
  wire _11554_;
  wire _11555_;
  wire _11556_;
  wire _11557_;
  wire _11558_;
  wire _11559_;
  wire _11560_;
  wire _11561_;
  wire _11562_;
  wire _11563_;
  wire _11564_;
  wire _11565_;
  wire _11566_;
  wire _11567_;
  wire _11568_;
  wire _11569_;
  wire _11570_;
  wire _11571_;
  wire _11572_;
  wire _11573_;
  wire _11574_;
  wire _11575_;
  wire _11576_;
  wire _11577_;
  wire _11578_;
  wire _11579_;
  wire _11580_;
  wire _11581_;
  wire _11582_;
  wire _11583_;
  wire _11584_;
  wire _11585_;
  wire _11586_;
  wire _11587_;
  wire _11588_;
  wire _11589_;
  wire _11590_;
  wire _11591_;
  wire _11592_;
  wire _11593_;
  wire _11594_;
  wire _11595_;
  wire _11596_;
  wire _11597_;
  wire _11598_;
  wire _11599_;
  wire _11600_;
  wire _11601_;
  wire _11602_;
  wire _11603_;
  wire _11604_;
  wire _11605_;
  wire _11606_;
  wire _11607_;
  wire _11608_;
  wire _11609_;
  wire _11610_;
  wire _11611_;
  wire _11612_;
  wire _11613_;
  wire _11614_;
  wire _11615_;
  wire _11616_;
  wire _11617_;
  wire _11618_;
  wire _11619_;
  wire _11620_;
  wire _11621_;
  wire _11622_;
  wire _11623_;
  wire _11624_;
  wire _11625_;
  wire _11626_;
  wire _11627_;
  wire _11628_;
  wire _11629_;
  wire _11630_;
  wire _11631_;
  wire _11632_;
  wire _11633_;
  wire _11634_;
  wire _11635_;
  wire _11636_;
  wire _11637_;
  wire _11638_;
  wire _11639_;
  wire _11640_;
  wire _11641_;
  wire _11642_;
  wire _11643_;
  wire _11644_;
  wire _11645_;
  wire _11646_;
  wire _11647_;
  wire _11648_;
  wire _11649_;
  wire _11650_;
  wire _11651_;
  wire _11652_;
  wire _11653_;
  wire _11654_;
  wire _11655_;
  wire _11656_;
  wire _11657_;
  wire _11658_;
  wire _11659_;
  wire _11660_;
  wire _11661_;
  wire _11662_;
  wire _11663_;
  wire _11664_;
  wire _11665_;
  wire _11666_;
  wire _11667_;
  wire _11668_;
  wire _11669_;
  wire _11670_;
  wire _11671_;
  wire _11672_;
  wire _11673_;
  wire _11674_;
  wire _11675_;
  wire _11676_;
  wire _11677_;
  wire _11678_;
  wire _11679_;
  wire _11680_;
  wire _11681_;
  wire _11682_;
  wire _11683_;
  wire _11684_;
  wire _11685_;
  wire _11686_;
  wire _11687_;
  wire _11688_;
  wire _11689_;
  wire _11690_;
  wire _11691_;
  wire _11692_;
  wire _11693_;
  wire _11694_;
  wire _11695_;
  wire _11696_;
  wire _11697_;
  wire _11698_;
  wire _11699_;
  wire _11700_;
  wire _11701_;
  wire _11702_;
  wire _11703_;
  wire _11704_;
  wire _11705_;
  wire _11706_;
  wire _11707_;
  wire _11708_;
  wire _11709_;
  wire _11710_;
  wire _11711_;
  wire _11712_;
  wire _11713_;
  wire _11714_;
  wire _11715_;
  wire _11716_;
  wire _11717_;
  wire _11718_;
  wire _11719_;
  wire _11720_;
  wire _11721_;
  wire _11722_;
  wire _11723_;
  wire _11724_;
  wire _11725_;
  wire _11726_;
  wire _11727_;
  wire _11728_;
  wire _11729_;
  wire _11730_;
  wire _11731_;
  wire _11732_;
  wire _11733_;
  wire _11734_;
  wire _11735_;
  wire _11736_;
  wire _11737_;
  wire _11738_;
  wire _11739_;
  wire _11740_;
  wire _11741_;
  wire _11742_;
  wire _11743_;
  wire _11744_;
  wire _11745_;
  wire _11746_;
  wire _11747_;
  wire _11748_;
  wire _11749_;
  wire _11750_;
  wire _11751_;
  wire _11752_;
  wire _11753_;
  wire _11754_;
  wire _11755_;
  wire _11756_;
  wire _11757_;
  wire _11758_;
  wire _11759_;
  wire _11760_;
  wire _11761_;
  wire _11762_;
  wire _11763_;
  wire _11764_;
  wire _11765_;
  wire _11766_;
  wire _11767_;
  wire _11768_;
  wire _11769_;
  wire _11770_;
  wire _11771_;
  wire _11772_;
  wire _11773_;
  wire _11774_;
  wire _11775_;
  wire _11776_;
  wire _11777_;
  wire _11778_;
  wire _11779_;
  wire _11780_;
  wire _11781_;
  wire _11782_;
  wire _11783_;
  wire _11784_;
  wire _11785_;
  wire _11786_;
  wire _11787_;
  wire _11788_;
  wire _11789_;
  wire _11790_;
  wire _11791_;
  wire _11792_;
  wire _11793_;
  wire _11794_;
  wire _11795_;
  wire _11796_;
  wire _11797_;
  wire _11798_;
  wire _11799_;
  wire _11800_;
  wire _11801_;
  wire _11802_;
  wire _11803_;
  wire _11804_;
  wire _11805_;
  wire _11806_;
  wire _11807_;
  wire _11808_;
  wire _11809_;
  wire _11810_;
  wire _11811_;
  wire _11812_;
  wire _11813_;
  wire _11814_;
  wire _11815_;
  wire _11816_;
  wire _11817_;
  wire _11818_;
  wire _11819_;
  wire _11820_;
  wire _11821_;
  wire _11822_;
  wire _11823_;
  wire _11824_;
  wire _11825_;
  wire _11826_;
  wire _11827_;
  wire _11828_;
  wire _11829_;
  wire _11830_;
  wire _11831_;
  wire _11832_;
  wire _11833_;
  wire _11834_;
  wire _11835_;
  wire _11836_;
  wire _11837_;
  wire _11838_;
  wire _11839_;
  wire _11840_;
  wire _11841_;
  wire _11842_;
  wire _11843_;
  wire _11844_;
  wire _11845_;
  wire _11846_;
  wire _11847_;
  wire _11848_;
  wire _11849_;
  wire _11850_;
  wire _11851_;
  wire _11852_;
  wire _11853_;
  wire _11854_;
  wire _11855_;
  wire _11856_;
  wire _11857_;
  wire _11858_;
  wire _11859_;
  wire _11860_;
  wire _11861_;
  wire _11862_;
  wire _11863_;
  wire _11864_;
  wire _11865_;
  wire _11866_;
  wire _11867_;
  wire _11868_;
  wire _11869_;
  wire _11870_;
  wire _11871_;
  wire _11872_;
  wire _11873_;
  wire _11874_;
  wire _11875_;
  wire _11876_;
  wire _11877_;
  wire _11878_;
  wire _11879_;
  wire _11880_;
  wire _11881_;
  wire _11882_;
  wire _11883_;
  wire _11884_;
  wire _11885_;
  wire _11886_;
  wire _11887_;
  wire _11888_;
  wire _11889_;
  wire _11890_;
  wire _11891_;
  wire _11892_;
  wire _11893_;
  wire _11894_;
  wire _11895_;
  wire _11896_;
  wire _11897_;
  wire _11898_;
  wire _11899_;
  wire _11900_;
  wire _11901_;
  wire _11902_;
  wire _11903_;
  wire _11904_;
  wire _11905_;
  wire _11906_;
  wire _11907_;
  wire _11908_;
  wire _11909_;
  wire _11910_;
  wire _11911_;
  wire _11912_;
  wire _11913_;
  wire _11914_;
  wire _11915_;
  wire _11916_;
  wire _11917_;
  wire _11918_;
  wire _11919_;
  wire _11920_;
  wire _11921_;
  wire _11922_;
  wire _11923_;
  wire _11924_;
  wire _11925_;
  wire _11926_;
  wire _11927_;
  wire _11928_;
  wire _11929_;
  wire _11930_;
  wire _11931_;
  wire _11932_;
  wire _11933_;
  wire _11934_;
  wire _11935_;
  wire _11936_;
  wire _11937_;
  wire _11938_;
  wire _11939_;
  wire _11940_;
  wire _11941_;
  wire _11942_;
  wire _11943_;
  wire _11944_;
  wire _11945_;
  wire _11946_;
  wire _11947_;
  wire _11948_;
  wire _11949_;
  wire _11950_;
  wire _11951_;
  wire _11952_;
  wire _11953_;
  wire _11954_;
  wire _11955_;
  wire _11956_;
  wire _11957_;
  wire _11958_;
  wire _11959_;
  wire _11960_;
  wire _11961_;
  wire _11962_;
  wire _11963_;
  wire _11964_;
  wire _11965_;
  wire _11966_;
  wire _11967_;
  wire _11968_;
  wire _11969_;
  wire _11970_;
  wire _11971_;
  wire _11972_;
  wire _11973_;
  wire _11974_;
  wire _11975_;
  wire _11976_;
  wire _11977_;
  wire _11978_;
  wire _11979_;
  wire _11980_;
  wire _11981_;
  wire _11982_;
  wire _11983_;
  wire _11984_;
  wire _11985_;
  wire _11986_;
  wire _11987_;
  wire _11988_;
  wire _11989_;
  wire _11990_;
  wire _11991_;
  wire _11992_;
  wire _11993_;
  wire _11994_;
  wire _11995_;
  wire _11996_;
  wire _11997_;
  wire _11998_;
  wire _11999_;
  wire _12000_;
  wire _12001_;
  wire _12002_;
  wire _12003_;
  wire _12004_;
  wire _12005_;
  wire _12006_;
  wire _12007_;
  wire _12008_;
  wire _12009_;
  wire _12010_;
  wire _12011_;
  wire _12012_;
  wire _12013_;
  wire _12014_;
  wire _12015_;
  wire _12016_;
  wire _12017_;
  wire _12018_;
  wire _12019_;
  wire _12020_;
  wire _12021_;
  wire _12022_;
  wire _12023_;
  wire _12024_;
  wire _12025_;
  wire _12026_;
  wire _12027_;
  wire _12028_;
  wire _12029_;
  wire _12030_;
  wire _12031_;
  wire _12032_;
  wire _12033_;
  wire _12034_;
  wire _12035_;
  wire _12036_;
  wire _12037_;
  wire _12038_;
  wire _12039_;
  wire _12040_;
  wire _12041_;
  wire _12042_;
  wire _12043_;
  wire _12044_;
  wire _12045_;
  wire _12046_;
  wire _12047_;
  wire _12048_;
  wire _12049_;
  wire _12050_;
  wire _12051_;
  wire _12052_;
  wire _12053_;
  wire _12054_;
  wire _12055_;
  wire _12056_;
  wire _12057_;
  wire _12058_;
  wire _12059_;
  wire _12060_;
  wire _12061_;
  wire _12062_;
  wire _12063_;
  wire _12064_;
  wire _12065_;
  wire _12066_;
  wire _12067_;
  wire _12068_;
  wire _12069_;
  wire _12070_;
  wire _12071_;
  wire _12072_;
  wire _12073_;
  wire _12074_;
  wire _12075_;
  wire _12076_;
  wire _12077_;
  wire _12078_;
  wire _12079_;
  wire _12080_;
  wire _12081_;
  wire _12082_;
  wire _12083_;
  wire _12084_;
  wire _12085_;
  wire _12086_;
  wire _12087_;
  wire _12088_;
  wire _12089_;
  wire _12090_;
  wire _12091_;
  wire _12092_;
  wire _12093_;
  wire _12094_;
  wire _12095_;
  wire _12096_;
  wire _12097_;
  wire _12098_;
  wire _12099_;
  wire _12100_;
  wire _12101_;
  wire _12102_;
  wire _12103_;
  wire _12104_;
  wire _12105_;
  wire _12106_;
  wire _12107_;
  wire _12108_;
  wire _12109_;
  wire _12110_;
  wire _12111_;
  wire _12112_;
  wire _12113_;
  wire _12114_;
  wire _12115_;
  wire _12116_;
  wire _12117_;
  wire _12118_;
  wire _12119_;
  wire _12120_;
  wire _12121_;
  wire _12122_;
  wire _12123_;
  wire _12124_;
  wire _12125_;
  wire _12126_;
  wire _12127_;
  wire _12128_;
  wire _12129_;
  wire _12130_;
  wire _12131_;
  wire _12132_;
  wire _12133_;
  wire _12134_;
  wire _12135_;
  wire _12136_;
  wire _12137_;
  wire _12138_;
  wire _12139_;
  wire _12140_;
  wire _12141_;
  wire _12142_;
  wire _12143_;
  wire _12144_;
  wire _12145_;
  wire _12146_;
  wire _12147_;
  wire _12148_;
  wire _12149_;
  wire _12150_;
  wire _12151_;
  wire _12152_;
  wire _12153_;
  wire _12154_;
  wire _12155_;
  wire _12156_;
  wire _12157_;
  wire _12158_;
  wire _12159_;
  wire _12160_;
  wire _12161_;
  wire _12162_;
  wire _12163_;
  wire _12164_;
  wire _12165_;
  wire _12166_;
  wire _12167_;
  wire _12168_;
  wire _12169_;
  wire _12170_;
  wire _12171_;
  wire _12172_;
  wire _12173_;
  wire _12174_;
  wire _12175_;
  wire _12176_;
  wire _12177_;
  wire _12178_;
  wire _12179_;
  wire _12180_;
  wire _12181_;
  wire _12182_;
  wire _12183_;
  wire _12184_;
  wire _12185_;
  wire _12186_;
  wire _12187_;
  wire _12188_;
  wire _12189_;
  wire _12190_;
  wire _12191_;
  wire _12192_;
  wire _12193_;
  wire _12194_;
  wire _12195_;
  wire _12196_;
  wire _12197_;
  wire _12198_;
  wire _12199_;
  wire _12200_;
  wire _12201_;
  wire _12202_;
  wire _12203_;
  wire _12204_;
  wire _12205_;
  wire _12206_;
  wire _12207_;
  wire _12208_;
  wire _12209_;
  wire _12210_;
  wire _12211_;
  wire _12212_;
  wire _12213_;
  wire _12214_;
  wire _12215_;
  wire _12216_;
  wire _12217_;
  wire _12218_;
  wire _12219_;
  wire _12220_;
  wire _12221_;
  wire _12222_;
  wire _12223_;
  wire _12224_;
  wire _12225_;
  wire _12226_;
  wire _12227_;
  wire _12228_;
  wire _12229_;
  wire _12230_;
  wire _12231_;
  wire _12232_;
  wire _12233_;
  wire _12234_;
  wire _12235_;
  wire _12236_;
  wire _12237_;
  wire _12238_;
  wire _12239_;
  wire _12240_;
  wire _12241_;
  wire _12242_;
  wire _12243_;
  wire _12244_;
  wire _12245_;
  wire _12246_;
  wire _12247_;
  wire _12248_;
  wire _12249_;
  wire _12250_;
  wire _12251_;
  wire _12252_;
  wire _12253_;
  wire _12254_;
  wire _12255_;
  wire _12256_;
  wire _12257_;
  wire _12258_;
  wire _12259_;
  wire _12260_;
  wire _12261_;
  wire _12262_;
  wire _12263_;
  wire _12264_;
  wire _12265_;
  wire _12266_;
  wire _12267_;
  wire _12268_;
  wire _12269_;
  wire _12270_;
  wire _12271_;
  wire _12272_;
  wire _12273_;
  wire _12274_;
  wire _12275_;
  wire _12276_;
  wire _12277_;
  wire _12278_;
  wire _12279_;
  wire _12280_;
  wire _12281_;
  wire _12282_;
  wire _12283_;
  wire _12284_;
  wire _12285_;
  wire _12286_;
  wire _12287_;
  wire _12288_;
  wire _12289_;
  wire _12290_;
  wire _12291_;
  wire _12292_;
  wire _12293_;
  wire _12294_;
  wire _12295_;
  wire _12296_;
  wire _12297_;
  wire _12298_;
  wire _12299_;
  wire _12300_;
  wire _12301_;
  wire _12302_;
  wire _12303_;
  wire _12304_;
  wire _12305_;
  wire _12306_;
  wire _12307_;
  wire _12308_;
  wire _12309_;
  wire _12310_;
  wire _12311_;
  wire _12312_;
  wire _12313_;
  wire _12314_;
  wire _12315_;
  wire _12316_;
  wire _12317_;
  wire _12318_;
  wire _12319_;
  wire _12320_;
  wire _12321_;
  wire _12322_;
  wire _12323_;
  wire _12324_;
  wire _12325_;
  wire _12326_;
  wire _12327_;
  wire _12328_;
  wire _12329_;
  wire _12330_;
  wire _12331_;
  wire _12332_;
  wire _12333_;
  wire _12334_;
  wire _12335_;
  wire _12336_;
  wire _12337_;
  wire _12338_;
  wire _12339_;
  wire _12340_;
  wire _12341_;
  wire _12342_;
  wire _12343_;
  wire _12344_;
  wire _12345_;
  wire _12346_;
  wire _12347_;
  wire _12348_;
  wire _12349_;
  wire _12350_;
  wire _12351_;
  wire _12352_;
  wire _12353_;
  wire _12354_;
  wire _12355_;
  wire _12356_;
  wire _12357_;
  wire _12358_;
  wire _12359_;
  wire _12360_;
  wire _12361_;
  wire _12362_;
  wire _12363_;
  wire _12364_;
  wire _12365_;
  wire _12366_;
  wire _12367_;
  wire _12368_;
  wire _12369_;
  wire _12370_;
  wire _12371_;
  wire _12372_;
  wire _12373_;
  wire _12374_;
  wire _12375_;
  wire _12376_;
  wire _12377_;
  wire _12378_;
  wire _12379_;
  wire _12380_;
  wire _12381_;
  wire _12382_;
  wire _12383_;
  wire _12384_;
  wire _12385_;
  wire _12386_;
  wire _12387_;
  wire _12388_;
  wire _12389_;
  wire _12390_;
  wire _12391_;
  wire _12392_;
  wire _12393_;
  wire _12394_;
  wire _12395_;
  wire _12396_;
  wire _12397_;
  wire _12398_;
  wire _12399_;
  wire _12400_;
  wire _12401_;
  wire _12402_;
  wire _12403_;
  wire _12404_;
  wire _12405_;
  wire _12406_;
  wire _12407_;
  wire _12408_;
  wire _12409_;
  wire _12410_;
  wire _12411_;
  wire _12412_;
  wire _12413_;
  wire _12414_;
  wire _12415_;
  wire _12416_;
  wire _12417_;
  wire _12418_;
  wire _12419_;
  wire _12420_;
  wire _12421_;
  wire _12422_;
  wire _12423_;
  wire _12424_;
  wire _12425_;
  wire _12426_;
  wire _12427_;
  wire _12428_;
  wire _12429_;
  wire _12430_;
  wire _12431_;
  wire _12432_;
  wire _12433_;
  wire _12434_;
  wire _12435_;
  wire _12436_;
  wire _12437_;
  wire _12438_;
  wire _12439_;
  wire _12440_;
  wire _12441_;
  wire _12442_;
  wire _12443_;
  wire _12444_;
  wire _12445_;
  wire _12446_;
  wire _12447_;
  wire _12448_;
  wire _12449_;
  wire _12450_;
  wire _12451_;
  wire _12452_;
  wire _12453_;
  wire _12454_;
  wire _12455_;
  wire _12456_;
  wire _12457_;
  wire _12458_;
  wire _12459_;
  wire _12460_;
  wire _12461_;
  wire _12462_;
  wire _12463_;
  wire _12464_;
  wire _12465_;
  wire _12466_;
  wire _12467_;
  wire _12468_;
  wire _12469_;
  wire _12470_;
  wire _12471_;
  wire _12472_;
  wire _12473_;
  wire _12474_;
  wire _12475_;
  wire _12476_;
  wire _12477_;
  wire _12478_;
  wire _12479_;
  wire _12480_;
  wire _12481_;
  wire _12482_;
  wire _12483_;
  wire _12484_;
  wire _12485_;
  wire _12486_;
  wire _12487_;
  wire _12488_;
  wire _12489_;
  wire _12490_;
  wire _12491_;
  wire _12492_;
  wire _12493_;
  wire _12494_;
  wire _12495_;
  wire _12496_;
  wire _12497_;
  wire _12498_;
  wire _12499_;
  wire _12500_;
  wire _12501_;
  wire _12502_;
  wire _12503_;
  wire _12504_;
  wire _12505_;
  wire _12506_;
  wire _12507_;
  wire _12508_;
  wire _12509_;
  wire _12510_;
  wire _12511_;
  wire _12512_;
  wire _12513_;
  wire _12514_;
  wire _12515_;
  wire _12516_;
  wire _12517_;
  wire _12518_;
  wire _12519_;
  wire _12520_;
  wire _12521_;
  wire _12522_;
  wire _12523_;
  wire _12524_;
  wire _12525_;
  wire _12526_;
  wire _12527_;
  wire _12528_;
  wire _12529_;
  wire _12530_;
  wire _12531_;
  wire _12532_;
  wire _12533_;
  wire _12534_;
  wire _12535_;
  wire _12536_;
  wire _12537_;
  wire _12538_;
  wire _12539_;
  wire _12540_;
  wire _12541_;
  wire _12542_;
  wire _12543_;
  wire _12544_;
  wire _12545_;
  wire _12546_;
  wire _12547_;
  wire _12548_;
  wire _12549_;
  wire _12550_;
  wire _12551_;
  wire _12552_;
  wire _12553_;
  wire _12554_;
  wire _12555_;
  wire _12556_;
  wire _12557_;
  wire _12558_;
  wire _12559_;
  wire _12560_;
  wire _12561_;
  wire _12562_;
  wire _12563_;
  wire _12564_;
  wire _12565_;
  wire _12566_;
  wire _12567_;
  wire _12568_;
  wire _12569_;
  wire _12570_;
  wire _12571_;
  wire _12572_;
  wire _12573_;
  wire _12574_;
  wire _12575_;
  wire _12576_;
  wire _12577_;
  wire _12578_;
  wire _12579_;
  wire _12580_;
  wire _12581_;
  wire _12582_;
  wire _12583_;
  wire _12584_;
  wire _12585_;
  wire _12586_;
  wire _12587_;
  wire _12588_;
  wire _12589_;
  wire _12590_;
  wire _12591_;
  wire _12592_;
  wire _12593_;
  wire _12594_;
  wire _12595_;
  wire _12596_;
  wire _12597_;
  wire _12598_;
  wire _12599_;
  wire _12600_;
  wire _12601_;
  wire _12602_;
  wire _12603_;
  wire _12604_;
  wire _12605_;
  wire _12606_;
  wire _12607_;
  wire _12608_;
  wire _12609_;
  wire _12610_;
  wire _12611_;
  wire _12612_;
  wire _12613_;
  wire _12614_;
  wire _12615_;
  wire _12616_;
  wire _12617_;
  wire _12618_;
  wire _12619_;
  wire _12620_;
  wire _12621_;
  wire _12622_;
  wire _12623_;
  wire _12624_;
  wire _12625_;
  wire _12626_;
  wire _12627_;
  wire _12628_;
  wire _12629_;
  wire _12630_;
  wire _12631_;
  wire _12632_;
  wire _12633_;
  wire _12634_;
  wire _12635_;
  wire _12636_;
  wire _12637_;
  wire _12638_;
  wire _12639_;
  wire _12640_;
  wire _12641_;
  wire _12642_;
  wire _12643_;
  wire _12644_;
  wire _12645_;
  wire _12646_;
  wire _12647_;
  wire _12648_;
  wire _12649_;
  wire _12650_;
  wire _12651_;
  wire _12652_;
  wire _12653_;
  wire _12654_;
  wire _12655_;
  wire _12656_;
  wire _12657_;
  wire _12658_;
  wire _12659_;
  wire _12660_;
  wire _12661_;
  wire _12662_;
  wire _12663_;
  wire _12664_;
  wire _12665_;
  wire _12666_;
  wire _12667_;
  wire _12668_;
  wire _12669_;
  wire _12670_;
  wire _12671_;
  wire _12672_;
  wire _12673_;
  wire _12674_;
  wire _12675_;
  wire _12676_;
  wire _12677_;
  wire _12678_;
  wire _12679_;
  wire _12680_;
  wire _12681_;
  wire _12682_;
  wire _12683_;
  wire _12684_;
  wire _12685_;
  wire _12686_;
  wire _12687_;
  wire _12688_;
  wire _12689_;
  wire _12690_;
  wire _12691_;
  wire _12692_;
  wire _12693_;
  wire _12694_;
  wire _12695_;
  wire _12696_;
  wire _12697_;
  wire _12698_;
  wire _12699_;
  wire _12700_;
  wire _12701_;
  wire _12702_;
  wire _12703_;
  wire _12704_;
  wire _12705_;
  wire _12706_;
  wire _12707_;
  wire _12708_;
  wire _12709_;
  wire _12710_;
  wire _12711_;
  wire _12712_;
  wire _12713_;
  wire _12714_;
  wire _12715_;
  wire _12716_;
  wire _12717_;
  wire _12718_;
  wire _12719_;
  wire _12720_;
  wire _12721_;
  wire _12722_;
  wire _12723_;
  wire _12724_;
  wire _12725_;
  wire _12726_;
  wire _12727_;
  wire _12728_;
  wire _12729_;
  wire _12730_;
  wire _12731_;
  wire _12732_;
  wire _12733_;
  wire _12734_;
  wire _12735_;
  wire _12736_;
  wire _12737_;
  wire _12738_;
  wire _12739_;
  wire _12740_;
  wire _12741_;
  wire _12742_;
  wire _12743_;
  wire _12744_;
  wire _12745_;
  wire _12746_;
  wire _12747_;
  wire _12748_;
  wire _12749_;
  wire _12750_;
  wire _12751_;
  wire _12752_;
  wire _12753_;
  wire _12754_;
  wire _12755_;
  wire _12756_;
  wire _12757_;
  wire _12758_;
  wire _12759_;
  wire _12760_;
  wire _12761_;
  wire _12762_;
  wire _12763_;
  wire _12764_;
  wire _12765_;
  wire _12766_;
  wire _12767_;
  wire _12768_;
  wire _12769_;
  wire _12770_;
  wire _12771_;
  wire _12772_;
  wire _12773_;
  wire _12774_;
  wire _12775_;
  wire _12776_;
  wire _12777_;
  wire _12778_;
  wire _12779_;
  wire _12780_;
  wire _12781_;
  wire _12782_;
  wire _12783_;
  wire _12784_;
  wire _12785_;
  wire _12786_;
  wire _12787_;
  wire _12788_;
  wire _12789_;
  wire _12790_;
  wire _12791_;
  wire _12792_;
  wire _12793_;
  wire _12794_;
  wire _12795_;
  wire _12796_;
  wire _12797_;
  wire _12798_;
  wire _12799_;
  wire _12800_;
  wire _12801_;
  wire _12802_;
  wire _12803_;
  wire _12804_;
  wire _12805_;
  wire _12806_;
  wire _12807_;
  wire _12808_;
  wire _12809_;
  wire _12810_;
  wire _12811_;
  wire _12812_;
  wire _12813_;
  wire _12814_;
  wire _12815_;
  wire _12816_;
  wire _12817_;
  wire _12818_;
  wire _12819_;
  wire _12820_;
  wire _12821_;
  wire _12822_;
  wire _12823_;
  wire _12824_;
  wire _12825_;
  wire _12826_;
  wire _12827_;
  wire _12828_;
  wire _12829_;
  wire _12830_;
  wire _12831_;
  wire _12832_;
  wire _12833_;
  wire _12834_;
  wire _12835_;
  wire _12836_;
  wire _12837_;
  wire _12838_;
  wire _12839_;
  wire _12840_;
  wire _12841_;
  wire _12842_;
  wire _12843_;
  wire _12844_;
  wire _12845_;
  wire _12846_;
  wire _12847_;
  wire _12848_;
  wire _12849_;
  wire _12850_;
  wire _12851_;
  wire _12852_;
  wire _12853_;
  wire _12854_;
  wire _12855_;
  wire _12856_;
  wire _12857_;
  wire _12858_;
  wire _12859_;
  wire _12860_;
  wire _12861_;
  wire _12862_;
  wire _12863_;
  wire _12864_;
  wire _12865_;
  wire _12866_;
  wire _12867_;
  wire _12868_;
  wire _12869_;
  wire _12870_;
  wire _12871_;
  wire _12872_;
  wire _12873_;
  wire _12874_;
  wire _12875_;
  wire _12876_;
  wire _12877_;
  wire _12878_;
  wire _12879_;
  wire _12880_;
  wire _12881_;
  wire _12882_;
  wire _12883_;
  wire _12884_;
  wire _12885_;
  wire _12886_;
  wire _12887_;
  wire _12888_;
  wire _12889_;
  wire _12890_;
  wire _12891_;
  wire _12892_;
  wire _12893_;
  wire _12894_;
  wire _12895_;
  wire _12896_;
  wire _12897_;
  wire _12898_;
  wire _12899_;
  wire _12900_;
  wire _12901_;
  wire _12902_;
  wire _12903_;
  wire _12904_;
  wire _12905_;
  wire _12906_;
  wire _12907_;
  wire _12908_;
  wire _12909_;
  wire _12910_;
  wire _12911_;
  wire _12912_;
  wire _12913_;
  wire _12914_;
  wire _12915_;
  wire _12916_;
  wire _12917_;
  wire _12918_;
  wire _12919_;
  wire _12920_;
  wire _12921_;
  wire _12922_;
  wire _12923_;
  wire _12924_;
  wire _12925_;
  wire _12926_;
  wire _12927_;
  wire _12928_;
  wire _12929_;
  wire _12930_;
  wire _12931_;
  wire _12932_;
  wire _12933_;
  wire _12934_;
  wire _12935_;
  wire _12936_;
  wire _12937_;
  wire _12938_;
  wire _12939_;
  wire _12940_;
  wire _12941_;
  wire _12942_;
  wire _12943_;
  wire _12944_;
  wire _12945_;
  wire _12946_;
  wire _12947_;
  wire _12948_;
  wire _12949_;
  wire _12950_;
  wire _12951_;
  wire _12952_;
  wire _12953_;
  wire _12954_;
  wire _12955_;
  wire _12956_;
  wire _12957_;
  wire _12958_;
  wire _12959_;
  wire _12960_;
  wire _12961_;
  wire _12962_;
  wire _12963_;
  wire _12964_;
  wire _12965_;
  wire _12966_;
  wire _12967_;
  wire _12968_;
  wire _12969_;
  wire _12970_;
  wire _12971_;
  wire _12972_;
  wire _12973_;
  wire _12974_;
  wire _12975_;
  wire _12976_;
  wire _12977_;
  wire _12978_;
  wire _12979_;
  wire _12980_;
  wire _12981_;
  wire _12982_;
  wire _12983_;
  wire _12984_;
  wire _12985_;
  wire _12986_;
  wire _12987_;
  wire _12988_;
  wire _12989_;
  wire _12990_;
  wire _12991_;
  wire _12992_;
  wire _12993_;
  wire _12994_;
  wire _12995_;
  wire _12996_;
  wire _12997_;
  wire _12998_;
  wire _12999_;
  wire _13000_;
  wire _13001_;
  wire _13002_;
  wire _13003_;
  wire _13004_;
  wire _13005_;
  wire _13006_;
  wire _13007_;
  wire _13008_;
  wire _13009_;
  wire _13010_;
  wire _13011_;
  wire _13012_;
  wire _13013_;
  wire _13014_;
  wire _13015_;
  wire _13016_;
  wire _13017_;
  wire _13018_;
  wire _13019_;
  wire _13020_;
  wire _13021_;
  wire _13022_;
  wire _13023_;
  wire _13024_;
  wire _13025_;
  wire _13026_;
  wire _13027_;
  wire _13028_;
  wire _13029_;
  wire _13030_;
  wire _13031_;
  wire _13032_;
  wire _13033_;
  wire _13034_;
  wire _13035_;
  wire _13036_;
  wire _13037_;
  wire _13038_;
  wire _13039_;
  wire _13040_;
  wire _13041_;
  wire _13042_;
  wire _13043_;
  wire _13044_;
  wire _13045_;
  wire _13046_;
  wire _13047_;
  wire _13048_;
  wire _13049_;
  wire _13050_;
  wire _13051_;
  wire _13052_;
  wire _13053_;
  wire _13054_;
  wire _13055_;
  wire _13056_;
  wire _13057_;
  wire _13058_;
  wire _13059_;
  wire _13060_;
  wire _13061_;
  wire _13062_;
  wire _13063_;
  wire _13064_;
  wire _13065_;
  wire _13066_;
  wire _13067_;
  wire _13068_;
  wire _13069_;
  wire _13070_;
  wire _13071_;
  wire _13072_;
  wire _13073_;
  wire _13074_;
  wire _13075_;
  wire _13076_;
  wire _13077_;
  wire _13078_;
  wire _13079_;
  wire _13080_;
  wire _13081_;
  wire _13082_;
  wire _13083_;
  wire _13084_;
  wire _13085_;
  wire _13086_;
  wire _13087_;
  wire _13088_;
  wire _13089_;
  wire _13090_;
  wire _13091_;
  wire _13092_;
  wire _13093_;
  wire _13094_;
  wire _13095_;
  wire _13096_;
  wire _13097_;
  wire _13098_;
  wire _13099_;
  wire _13100_;
  wire _13101_;
  wire _13102_;
  wire _13103_;
  wire _13104_;
  wire _13105_;
  wire _13106_;
  wire _13107_;
  wire _13108_;
  wire _13109_;
  wire _13110_;
  wire _13111_;
  wire _13112_;
  wire _13113_;
  wire _13114_;
  wire _13115_;
  wire _13116_;
  wire _13117_;
  wire _13118_;
  wire _13119_;
  wire _13120_;
  wire _13121_;
  wire _13122_;
  wire _13123_;
  wire _13124_;
  wire _13125_;
  wire _13126_;
  wire _13127_;
  wire _13128_;
  wire _13129_;
  wire _13130_;
  wire _13131_;
  wire _13132_;
  wire _13133_;
  wire _13134_;
  wire _13135_;
  wire _13136_;
  wire _13137_;
  wire _13138_;
  wire _13139_;
  wire _13140_;
  wire _13141_;
  wire _13142_;
  wire _13143_;
  wire _13144_;
  wire _13145_;
  wire _13146_;
  wire _13147_;
  wire _13148_;
  wire _13149_;
  wire _13150_;
  wire _13151_;
  wire _13152_;
  wire _13153_;
  wire _13154_;
  wire _13155_;
  wire _13156_;
  wire _13157_;
  wire _13158_;
  wire _13159_;
  wire _13160_;
  wire _13161_;
  wire _13162_;
  wire _13163_;
  wire _13164_;
  wire _13165_;
  wire _13166_;
  wire _13167_;
  wire _13168_;
  wire _13169_;
  wire _13170_;
  wire _13171_;
  wire _13172_;
  wire _13173_;
  wire _13174_;
  wire _13175_;
  wire _13176_;
  wire _13177_;
  wire _13178_;
  wire _13179_;
  wire _13180_;
  wire _13181_;
  wire _13182_;
  wire _13183_;
  wire _13184_;
  wire _13185_;
  wire _13186_;
  wire _13187_;
  wire _13188_;
  wire _13189_;
  wire _13190_;
  wire _13191_;
  wire _13192_;
  wire _13193_;
  wire _13194_;
  wire _13195_;
  wire _13196_;
  wire _13197_;
  wire _13198_;
  wire _13199_;
  wire _13200_;
  wire _13201_;
  wire _13202_;
  wire _13203_;
  wire _13204_;
  wire _13205_;
  wire _13206_;
  wire _13207_;
  wire _13208_;
  wire _13209_;
  wire _13210_;
  wire _13211_;
  wire _13212_;
  wire _13213_;
  wire _13214_;
  wire _13215_;
  wire _13216_;
  wire _13217_;
  wire _13218_;
  wire _13219_;
  wire _13220_;
  wire _13221_;
  wire _13222_;
  wire _13223_;
  wire _13224_;
  wire _13225_;
  wire _13226_;
  wire _13227_;
  wire _13228_;
  wire _13229_;
  wire _13230_;
  wire _13231_;
  wire _13232_;
  wire _13233_;
  wire _13234_;
  wire _13235_;
  wire _13236_;
  wire _13237_;
  wire _13238_;
  wire _13239_;
  wire _13240_;
  wire _13241_;
  wire _13242_;
  wire _13243_;
  wire _13244_;
  wire _13245_;
  wire _13246_;
  wire _13247_;
  wire _13248_;
  wire _13249_;
  wire _13250_;
  wire _13251_;
  wire _13252_;
  wire _13253_;
  wire _13254_;
  wire _13255_;
  wire _13256_;
  wire _13257_;
  wire _13258_;
  wire _13259_;
  wire _13260_;
  wire _13261_;
  wire _13262_;
  wire _13263_;
  wire _13264_;
  wire _13265_;
  input [8:0] ABINPUT;
  input [16:0] ABINPUT000;
  input [16:0] ABINPUT001;
  input clk;
  wire [31:0] cxrom_data_out;
  wire cy;
  wire first_instr;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein0 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein1 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein2 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein3 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout0 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout1 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout2 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout3 ;
  wire \oc8051_symbolic_cxrom1.clk ;
  wire [31:0] \oc8051_symbolic_cxrom1.cxrom_data_out ;
  wire [15:0] \oc8051_symbolic_cxrom1.pc1 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc10 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc12 ;
  wire [15:0] \oc8051_symbolic_cxrom1.pc2 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc20 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc22 ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[0] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[10] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[11] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[12] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[13] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[14] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[15] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[1] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[2] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[3] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[4] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[5] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[6] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[7] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[8] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[9] ;
  wire [15:0] \oc8051_symbolic_cxrom1.regvalid ;
  wire \oc8051_symbolic_cxrom1.rst ;
  wire [31:0] \oc8051_symbolic_cxrom1.word_in ;
  wire [8:0] \oc8051_top_1.ABINPUT ;
  wire [16:0] \oc8051_top_1.ABINPUT000 ;
  wire [16:0] \oc8051_top_1.ABINPUT001 ;
  wire [7:0] \oc8051_top_1.acc ;
  wire \oc8051_top_1.bit_data ;
  wire [31:0] \oc8051_top_1.cxrom_data_out ;
  wire \oc8051_top_1.cy ;
  wire [1:0] \oc8051_top_1.cy_sel ;
  wire [7:0] \oc8051_top_1.dptr_hi ;
  wire [7:0] \oc8051_top_1.dptr_lo ;
  wire [31:0] \oc8051_top_1.idat_onchip ;
  wire \oc8051_top_1.int_ack ;
  wire [7:0] \oc8051_top_1.int_src ;
  wire \oc8051_top_1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.mem_act ;
  wire [16:0] \oc8051_top_1.oc8051_alu1.ABINPUT ;
  wire [16:0] \oc8051_top_1.oc8051_alu1.ABINPUT000 ;
  wire \oc8051_top_1.oc8051_alu1.clk ;
  wire \oc8051_top_1.oc8051_alu1.divOv ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.divsrc1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.divsrc2 ;
  wire \oc8051_top_1.oc8051_alu1.mulOv ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.mulsrc1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.mulsrc2 ;
  wire \oc8051_top_1.oc8051_alu1.rst ;
  wire \oc8051_top_1.oc8051_alu1.srcAc ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.acc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.clk ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.dptr ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op1_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op2_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op3_r ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.pc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_alu_src_sel1.sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_alu_src_sel1.sel2 ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.sel3 ;
  wire [7:0] \oc8051_top_1.oc8051_comp1.acc ;
  wire \oc8051_top_1.oc8051_comp1.cy ;
  wire \oc8051_top_1.oc8051_cy_select1.cy_in ;
  wire [1:0] \oc8051_top_1.oc8051_cy_select1.cy_sel ;
  wire [3:0] \oc8051_top_1.oc8051_decoder1.alu_op ;
  wire \oc8051_top_1.oc8051_decoder1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.cy_sel ;
  wire \oc8051_top_1.oc8051_decoder1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_decoder1.op ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.psw_set ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_wr_sel ;
  wire \oc8051_top_1.oc8051_decoder1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.src_sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.src_sel2 ;
  wire \oc8051_top_1.oc8051_decoder1.src_sel3 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.state ;
  wire \oc8051_top_1.oc8051_decoder1.wait_data ;
  wire \oc8051_top_1.oc8051_decoder1.wr ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.wr_sfr ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[7] ;
  wire \oc8051_top_1.oc8051_indi_addr1.clk ;
  wire \oc8051_top_1.oc8051_indi_addr1.rst ;
  wire \oc8051_top_1.oc8051_indi_addr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.acc ;
  wire \oc8051_top_1.oc8051_memory_interface1.bit_in ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.cdata ;
  wire \oc8051_top_1.oc8051_memory_interface1.cdone ;
  wire \oc8051_top_1.oc8051_memory_interface1.clk ;
  wire \oc8051_top_1.oc8051_memory_interface1.dmem_wait ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dptr ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.iadr_t ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_cur ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_old ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_onchip ;
  wire \oc8051_top_1.oc8051_memory_interface1.imem_wait ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm2_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.in_ram ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_t ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_v ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_vec_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.istb_t ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op2_buff ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op3_buff ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.op_pos ;
  wire \oc8051_top_1.oc8051_memory_interface1.out_of_rst ;
  wire [3:0] \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_buf ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_for_ajmp ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log_prev ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_out ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_addr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_ind ;
  wire \oc8051_top_1.oc8051_memory_interface1.reti ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ri_r ;
  wire [4:0] \oc8051_top_1.oc8051_memory_interface1.rn_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.sfr ;
  wire \oc8051_top_1.oc8051_memory_interface1.sfr_bit ;
  wire \oc8051_top_1.oc8051_rom1.clk ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.cxrom_data_out ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.data_o ;
  wire \oc8051_top_1.oc8051_rom1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.b_reg ;
  wire \oc8051_top_1.oc8051_sfr1.bit_out ;
  wire \oc8051_top_1.oc8051_sfr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.cy ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_lo ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.int_ack ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ip ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ack ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.t2_int ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.uart_int ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.p ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.set ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd ;
  wire [11:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp ;
  wire [10:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.pres_ow ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.prescaler ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.psw_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.rxd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.srcAc ;
  wire \oc8051_top_1.oc8051_sfr1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.t2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.tc2_int ;
  wire \oc8051_top_1.oc8051_sfr1.tclk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.tf0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.uart_int ;
  wire \oc8051_top_1.oc8051_sfr1.wait_data ;
  wire \oc8051_top_1.oc8051_sfr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.p0_i ;
  wire [7:0] \oc8051_top_1.p0_o ;
  wire [7:0] \oc8051_top_1.p1_i ;
  wire [7:0] \oc8051_top_1.p1_o ;
  wire [7:0] \oc8051_top_1.p2_i ;
  wire [7:0] \oc8051_top_1.p2_o ;
  wire [7:0] \oc8051_top_1.p3_i ;
  wire [7:0] \oc8051_top_1.p3_o ;
  wire [15:0] \oc8051_top_1.pc ;
  wire [15:0] \oc8051_top_1.pc_log ;
  wire [15:0] \oc8051_top_1.pc_log_prev ;
  wire [1:0] \oc8051_top_1.psw_set ;
  wire [7:0] \oc8051_top_1.ram_data ;
  wire \oc8051_top_1.rd_ind ;
  wire \oc8051_top_1.reti ;
  wire \oc8051_top_1.rxd_i ;
  wire \oc8051_top_1.sfr_bit ;
  wire [7:0] \oc8051_top_1.sfr_out ;
  wire \oc8051_top_1.srcAc ;
  wire [2:0] \oc8051_top_1.src_sel1 ;
  wire [1:0] \oc8051_top_1.src_sel2 ;
  wire \oc8051_top_1.src_sel3 ;
  wire \oc8051_top_1.t0_i ;
  wire \oc8051_top_1.t1_i ;
  wire \oc8051_top_1.t2_i ;
  wire \oc8051_top_1.t2ex_i ;
  wire \oc8051_top_1.wait_data ;
  wire \oc8051_top_1.wb_clk_i ;
  wire \oc8051_top_1.wb_rst_i ;
  input [7:0] p0_in;
  wire [7:0] p0_out;
  input [7:0] p1_in;
  wire [7:0] p1_out;
  input [7:0] p2_in;
  wire [7:0] p2_out;
  input [7:0] p3_in;
  wire [7:0] p3_out;
  wire [15:0] pc1;
  wire [15:0] pc1_plus_2;
  wire [15:0] pc2;
  output property_invalid_ajmp;
  input rst;
  input rxd_i;
  input t0_i;
  input t1_i;
  input t2_i;
  input t2ex_i;
  input [31:0] word_in;
  not _13266_ (_04856_, rst);
  not _13267_ (_04857_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  not _13268_ (_04858_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  not _13269_ (_04859_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and _13270_ (_04860_, \oc8051_top_1.oc8051_decoder1.wr , _04859_);
  and _13271_ (_04861_, _04860_, _04858_);
  and _13272_ (_04862_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  and _13273_ (_04863_, _04862_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  and _13274_ (_04864_, _04863_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  and _13275_ (_04865_, _04864_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  and _13276_ (_04866_, _04865_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  and _13277_ (_04867_, _04866_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  not _13278_ (_04868_, _04867_);
  not _13279_ (_04869_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and _13280_ (_04870_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _04859_);
  and _13281_ (_04871_, _04870_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  and _13282_ (_04872_, _04871_, _04869_);
  or _13283_ (_04873_, _04866_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  and _13284_ (_04874_, _04873_, _04872_);
  nand _13285_ (_04875_, _04874_, _04868_);
  and _13286_ (_04876_, _04871_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  not _13287_ (_04877_, _04876_);
  not _13288_ (_04878_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  and _13289_ (_04879_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _04859_);
  and _13290_ (_04880_, _04879_, _04878_);
  and _13291_ (_04881_, _04880_, _04869_);
  nand _13292_ (_04882_, _04881_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  and _13293_ (_04883_, _04882_, _04877_);
  and _13294_ (_04884_, _04870_, _04869_);
  not _13295_ (_04885_, _04884_);
  nor _13296_ (_04886_, _04885_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  nand _13297_ (_04887_, _04886_, \oc8051_top_1.oc8051_memory_interface1.ri_r [6]);
  and _13298_ (_04888_, _04880_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  nand _13299_ (_04889_, _04888_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  and _13300_ (_04890_, _04889_, _04887_);
  and _13301_ (_04892_, _04890_, _04883_);
  and _13302_ (_04893_, _04892_, _04875_);
  nand _13303_ (_04894_, _04867_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  or _13304_ (_04895_, _04867_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  and _13305_ (_04896_, _04895_, _04894_);
  nand _13306_ (_04897_, _04896_, _04872_);
  nand _13307_ (_04898_, _04881_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  and _13308_ (_04899_, _04898_, _04877_);
  nand _13309_ (_04900_, _04886_, \oc8051_top_1.oc8051_memory_interface1.ri_r [7]);
  nand _13310_ (_04901_, _04888_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  and _13311_ (_04902_, _04901_, _04900_);
  and _13312_ (_04903_, _04902_, _04899_);
  and _13313_ (_04904_, _04903_, _04897_);
  and _13314_ (_04905_, _04904_, _04893_);
  not _13315_ (_04906_, _04865_);
  or _13316_ (_04907_, _04864_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  and _13317_ (_04908_, _04907_, _04872_);
  and _13318_ (_04909_, _04908_, _04906_);
  not _13319_ (_04910_, _04909_);
  nand _13320_ (_04911_, _04888_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  and _13321_ (_04912_, _04911_, _04877_);
  nor _13322_ (_04913_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  nor _13323_ (_04914_, _04913_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _13324_ (_04915_, _04914_, _04879_);
  nand _13325_ (_04916_, _04915_, \oc8051_top_1.oc8051_memory_interface1.rn_r [4]);
  nand _13326_ (_04917_, _04886_, \oc8051_top_1.oc8051_memory_interface1.ri_r [4]);
  and _13327_ (_04918_, _04917_, _04916_);
  nand _13328_ (_04919_, _04881_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  and _13329_ (_04920_, _04919_, _04918_);
  and _13330_ (_04921_, _04920_, _04912_);
  and _13331_ (_04922_, _04921_, _04910_);
  or _13332_ (_04923_, _04865_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nand _13333_ (_04924_, _04923_, _04872_);
  or _13334_ (_04925_, _04924_, _04866_);
  nand _13335_ (_04926_, _04888_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  nand _13336_ (_04927_, _04881_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  and _13337_ (_04928_, _04927_, _04926_);
  nand _13338_ (_04929_, _04886_, \oc8051_top_1.oc8051_memory_interface1.ri_r [5]);
  and _13339_ (_04930_, _04929_, _04877_);
  and _13340_ (_04931_, _04930_, _04928_);
  and _13341_ (_04932_, _04931_, _04925_);
  not _13342_ (_04933_, _04932_);
  nor _13343_ (_04934_, _04933_, _04922_);
  and _13344_ (_04935_, _04934_, _04905_);
  and _13345_ (_04936_, _04888_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  and _13346_ (_04937_, _04881_, \oc8051_top_1.oc8051_memory_interface1.imm_r [3]);
  nor _13347_ (_04938_, _04937_, _04936_);
  nor _13348_ (_04939_, _04863_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor _13349_ (_04940_, _04939_, _04864_);
  and _13350_ (_04941_, _04940_, _04872_);
  not _13351_ (_04942_, _04941_);
  nand _13352_ (_04943_, _04915_, \oc8051_top_1.oc8051_memory_interface1.rn_r [3]);
  nand _13353_ (_04944_, _04886_, \oc8051_top_1.oc8051_memory_interface1.ri_r [3]);
  and _13354_ (_04945_, _04944_, _04943_);
  and _13355_ (_04946_, _04945_, _04942_);
  and _13356_ (_04947_, _04946_, _04938_);
  not _13357_ (_04948_, _04947_);
  nand _13358_ (_04949_, _04888_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  nand _13359_ (_04950_, _04915_, \oc8051_top_1.oc8051_memory_interface1.rn_r [0]);
  and _13360_ (_04951_, _04950_, _04949_);
  not _13361_ (_04952_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  nand _13362_ (_04953_, _04872_, _04952_);
  nand _13363_ (_04954_, _04881_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  nand _13364_ (_04955_, _04886_, \oc8051_top_1.oc8051_memory_interface1.ri_r [0]);
  and _13365_ (_04956_, _04955_, _04954_);
  and _13366_ (_04957_, _04956_, _04953_);
  and _13367_ (_04958_, _04957_, _04951_);
  not _13368_ (_04959_, _04958_);
  nor _13369_ (_04960_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  nor _13370_ (_04961_, _04960_, _04862_);
  nand _13371_ (_04962_, _04961_, _04872_);
  nand _13372_ (_04963_, _04886_, \oc8051_top_1.oc8051_memory_interface1.ri_r [1]);
  and _13373_ (_04964_, _04963_, _04962_);
  nand _13374_ (_04965_, _04881_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  nand _13375_ (_04966_, _04888_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [1]);
  nand _13376_ (_04967_, _04915_, \oc8051_top_1.oc8051_memory_interface1.rn_r [1]);
  and _13377_ (_04968_, _04967_, _04966_);
  and _13378_ (_04969_, _04968_, _04965_);
  and _13379_ (_04971_, _04969_, _04964_);
  not _13380_ (_04972_, _04872_);
  nor _13381_ (_04973_, _04862_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  or _13382_ (_04974_, _04973_, _04863_);
  or _13383_ (_04975_, _04974_, _04972_);
  nand _13384_ (_04976_, _04886_, \oc8051_top_1.oc8051_memory_interface1.ri_r [2]);
  and _13385_ (_04977_, _04976_, _04975_);
  nand _13386_ (_04978_, _04881_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  nand _13387_ (_04979_, _04888_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [2]);
  nand _13388_ (_04980_, _04915_, \oc8051_top_1.oc8051_memory_interface1.rn_r [2]);
  and _13389_ (_04981_, _04980_, _04979_);
  and _13390_ (_04982_, _04981_, _04978_);
  and _13391_ (_04984_, _04982_, _04977_);
  and _13392_ (_04985_, _04984_, _04971_);
  and _13393_ (_04986_, _04985_, _04959_);
  and _13394_ (_04987_, _04986_, _04948_);
  and _13395_ (_04988_, _04987_, _04935_);
  and _13396_ (_04989_, _04971_, _04958_);
  and _13397_ (_04990_, _04989_, _04984_);
  and _13398_ (_04991_, _04990_, _04948_);
  and _13399_ (_04992_, _04991_, _04935_);
  and _13400_ (_04993_, _04932_, _04922_);
  and _13401_ (_04994_, _04993_, _04905_);
  and _13402_ (_04995_, _04994_, _04985_);
  not _13403_ (_04996_, _04971_);
  nor _13404_ (_04997_, _04996_, _04958_);
  and _13405_ (_04998_, _04984_, _04947_);
  and _13406_ (_04999_, _04998_, _04997_);
  and _13407_ (_05000_, _04999_, _04935_);
  and _13408_ (_05001_, _04998_, _04989_);
  and _13409_ (_05002_, _05001_, _04935_);
  or _13410_ (_05003_, _05002_, _05000_);
  or _13411_ (_05004_, _05003_, _04995_);
  or _13412_ (_05005_, _05004_, _04992_);
  or _13413_ (_05006_, _05005_, _04988_);
  nand _13414_ (_05007_, _05006_, _04861_);
  and _13415_ (_05008_, _05005_, _04861_);
  nor _13416_ (_05009_, _05008_, _05007_);
  nor _13417_ (_05010_, _05009_, _04857_);
  not _13418_ (_05011_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  not _13419_ (_05012_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  not _13420_ (_05013_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and _13421_ (_05014_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], _05013_);
  nand _13422_ (_05015_, _05014_, _05012_);
  nor _13423_ (_05016_, _05015_, _05011_);
  not _13424_ (_05017_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  or _13425_ (_05018_, _05012_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  or _13426_ (_05019_, _05018_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  nor _13427_ (_05020_, _05019_, _05017_);
  nor _13428_ (_05021_, _05020_, _05016_);
  not _13429_ (_05022_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  or _13430_ (_05023_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  or _13431_ (_05024_, _05023_, _05013_);
  nor _13432_ (_05025_, _05024_, _05022_);
  not _13433_ (_05026_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  or _13434_ (_05027_, _05018_, _05013_);
  nor _13435_ (_05028_, _05027_, _05026_);
  nor _13436_ (_05029_, _05028_, _05025_);
  and _13437_ (_05030_, _05029_, _05021_);
  not _13438_ (_05031_, \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  and _13439_ (_05032_, _05031_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r );
  nor _13440_ (_05033_, _05032_, ABINPUT[7]);
  nand _13441_ (_05034_, _05031_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r );
  nor _13442_ (_05035_, _05034_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  nor _13443_ (_05036_, _05035_, _05033_);
  nor _13444_ (_05037_, _05023_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and _13445_ (_05038_, _05037_, _05036_);
  and _13446_ (_05039_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  and _13447_ (_05040_, _05039_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and _13448_ (_05041_, _05040_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [6]);
  not _13449_ (_05042_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nand _13450_ (_05043_, _05039_, _05013_);
  nor _13451_ (_05044_, _05043_, _05042_);
  nor _13452_ (_05045_, _05044_, _05041_);
  not _13453_ (_05046_, _05045_);
  nor _13454_ (_05047_, _05046_, _05038_);
  and _13455_ (_05048_, _05047_, _05030_);
  not _13456_ (_05049_, _05048_);
  or _13457_ (_05050_, _05032_, ABINPUT[0]);
  or _13458_ (_05051_, _05034_, \oc8051_top_1.oc8051_sfr1.bit_out );
  nand _13459_ (_05052_, _05051_, _05050_);
  not _13460_ (_05053_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  nand _13461_ (_05054_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  and _13462_ (_05055_, _05054_, _05053_);
  or _13463_ (_05056_, _05055_, _05052_);
  not _13464_ (_05057_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  or _13465_ (_05058_, _05055_, _05057_);
  nand _13466_ (_05059_, _05058_, _05056_);
  not _13467_ (_05060_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  nor _13468_ (_05061_, _05015_, _05060_);
  not _13469_ (_05062_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  nor _13470_ (_05063_, _05019_, _05062_);
  nor _13471_ (_05064_, _05063_, _05061_);
  not _13472_ (_05065_, _05027_);
  and _13473_ (_05066_, _05065_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  not _13474_ (_05067_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor _13475_ (_05068_, _05024_, _05067_);
  nor _13476_ (_05069_, _05068_, _05066_);
  and _13477_ (_05070_, _05069_, _05064_);
  nor _13478_ (_05071_, _05032_, ABINPUT[5]);
  nor _13479_ (_05072_, _05034_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  nor _13480_ (_05073_, _05072_, _05071_);
  and _13481_ (_05074_, _05073_, _05037_);
  not _13482_ (_05075_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor _13483_ (_05076_, _05043_, _05075_);
  and _13484_ (_05077_, _05040_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [4]);
  nor _13485_ (_05078_, _05077_, _05076_);
  not _13486_ (_05079_, _05078_);
  nor _13487_ (_05080_, _05079_, _05074_);
  and _13488_ (_05081_, _05080_, _05070_);
  not _13489_ (_05082_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  or _13490_ (_05083_, _05015_, _05082_);
  not _13491_ (_05084_, \oc8051_top_1.oc8051_memory_interface1.imm_r [3]);
  or _13492_ (_05085_, _05019_, _05084_);
  and _13493_ (_05086_, _05085_, _05083_);
  not _13494_ (_05087_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nor _13495_ (_05088_, _05027_, _05087_);
  not _13496_ (_05089_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor _13497_ (_05090_, _05024_, _05089_);
  nor _13498_ (_05091_, _05090_, _05088_);
  and _13499_ (_05092_, _05091_, _05086_);
  not _13500_ (_05093_, _05037_);
  or _13501_ (_05094_, _05032_, ABINPUT[4]);
  or _13502_ (_05095_, _05034_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  nand _13503_ (_05096_, _05095_, _05094_);
  or _13504_ (_05097_, _05096_, _05093_);
  and _13505_ (_05098_, _05040_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [3]);
  not _13506_ (_05099_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor _13507_ (_05100_, _05043_, _05099_);
  nor _13508_ (_05101_, _05100_, _05098_);
  and _13509_ (_05102_, _05101_, _05097_);
  and _13510_ (_05103_, _05102_, _05092_);
  not _13511_ (_05104_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  or _13512_ (_05105_, _05019_, _05104_);
  not _13513_ (_05106_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  or _13514_ (_05107_, _05015_, _05106_);
  and _13515_ (_05108_, _05107_, _05105_);
  not _13516_ (_05109_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  or _13517_ (_05110_, _05027_, _05109_);
  not _13518_ (_05111_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  or _13519_ (_05112_, _05024_, _05111_);
  and _13520_ (_05114_, _05112_, _05110_);
  and _13521_ (_05115_, _05114_, _05108_);
  or _13522_ (_05117_, _05032_, ABINPUT[1]);
  or _13523_ (_05118_, _05034_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  nand _13524_ (_05119_, _05118_, _05117_);
  or _13525_ (_05120_, _05119_, _05093_);
  nand _13526_ (_05121_, _05040_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [0]);
  not _13527_ (_05122_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or _13528_ (_05123_, _05043_, _05122_);
  and _13529_ (_05124_, _05123_, _05121_);
  and _13530_ (_05125_, _05124_, _05120_);
  and _13531_ (_05126_, _05125_, _05115_);
  or _13532_ (_05128_, _05032_, ABINPUT[2]);
  or _13533_ (_05129_, _05034_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  nand _13534_ (_05130_, _05129_, _05128_);
  or _13535_ (_05131_, _05130_, _05093_);
  not _13536_ (_05132_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  or _13537_ (_05134_, _05019_, _05132_);
  not _13538_ (_05135_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [1]);
  or _13539_ (_05137_, _05015_, _05135_);
  and _13540_ (_05138_, _05137_, _05134_);
  and _13541_ (_05139_, _05138_, _05131_);
  not _13542_ (_05140_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  or _13543_ (_05141_, _05027_, _05140_);
  not _13544_ (_05142_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  or _13545_ (_05144_, _05024_, _05142_);
  and _13546_ (_05145_, _05144_, _05141_);
  nand _13547_ (_05146_, _05040_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [1]);
  not _13548_ (_05147_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or _13549_ (_05148_, _05043_, _05147_);
  and _13550_ (_05149_, _05148_, _05146_);
  and _13551_ (_05150_, _05149_, _05145_);
  and _13552_ (_05151_, _05150_, _05139_);
  not _13553_ (_05152_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  or _13554_ (_05153_, _05019_, _05152_);
  not _13555_ (_05154_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [2]);
  or _13556_ (_05155_, _05015_, _05154_);
  and _13557_ (_05156_, _05155_, _05153_);
  not _13558_ (_05157_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  or _13559_ (_05158_, _05024_, _05157_);
  not _13560_ (_05159_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  or _13561_ (_05160_, _05027_, _05159_);
  and _13562_ (_05161_, _05160_, _05158_);
  and _13563_ (_05162_, _05161_, _05156_);
  or _13564_ (_05163_, _05032_, ABINPUT[3]);
  or _13565_ (_05164_, _05034_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  nand _13566_ (_05165_, _05164_, _05163_);
  or _13567_ (_05166_, _05165_, _05093_);
  not _13568_ (_05167_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or _13569_ (_05168_, _05043_, _05167_);
  nand _13570_ (_05169_, _05040_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [2]);
  and _13571_ (_05170_, _05169_, _05168_);
  and _13572_ (_05171_, _05170_, _05166_);
  and _13573_ (_05172_, _05171_, _05162_);
  and _13574_ (_05173_, _05172_, _05151_);
  and _13575_ (_05174_, _05173_, _05126_);
  and _13576_ (_05175_, _05174_, _05103_);
  and _13577_ (_05176_, _05175_, _05081_);
  not _13578_ (_05177_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  nor _13579_ (_05178_, _05015_, _05177_);
  not _13580_ (_05179_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  nor _13581_ (_05180_, _05019_, _05179_);
  nor _13582_ (_05181_, _05180_, _05178_);
  not _13583_ (_05183_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nor _13584_ (_05184_, _05027_, _05183_);
  not _13585_ (_05185_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor _13586_ (_05186_, _05024_, _05185_);
  nor _13587_ (_05187_, _05186_, _05184_);
  and _13588_ (_05188_, _05187_, _05181_);
  nor _13589_ (_05189_, _05032_, ABINPUT[6]);
  nor _13590_ (_05190_, _05034_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  nor _13591_ (_05191_, _05190_, _05189_);
  and _13592_ (_05192_, _05191_, _05037_);
  and _13593_ (_05193_, _05040_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [5]);
  not _13594_ (_05194_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor _13595_ (_05195_, _05043_, _05194_);
  nor _13596_ (_05196_, _05195_, _05193_);
  not _13597_ (_05197_, _05196_);
  nor _13598_ (_05198_, _05197_, _05192_);
  and _13599_ (_05199_, _05198_, _05188_);
  nand _13600_ (_05201_, _05199_, _05176_);
  nand _13601_ (_05202_, _05201_, _05059_);
  not _13602_ (_05204_, _05103_);
  not _13603_ (_05205_, _05172_);
  nand _13604_ (_05206_, _05125_, _05115_);
  nand _13605_ (_05207_, _05150_, _05139_);
  and _13606_ (_05208_, _05207_, _05206_);
  and _13607_ (_05209_, _05208_, _05205_);
  and _13608_ (_05210_, _05209_, _05204_);
  nor _13609_ (_05211_, _05199_, _05081_);
  and _13610_ (_05212_, _05211_, _05210_);
  or _13611_ (_05213_, _05212_, _05059_);
  and _13612_ (_05214_, _05213_, _05202_);
  nand _13613_ (_05215_, _05214_, _05049_);
  not _13614_ (_05216_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and _13615_ (_05217_, \oc8051_top_1.oc8051_decoder1.alu_op [1], _04859_);
  and _13616_ (_05218_, _05217_, _05216_);
  and _13617_ (_05220_, \oc8051_top_1.oc8051_decoder1.alu_op [3], _04859_);
  and _13618_ (_05221_, _05220_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and _13619_ (_05223_, _05221_, _05218_);
  or _13620_ (_05224_, _05214_, _05049_);
  and _13621_ (_05225_, _05224_, _05223_);
  and _13622_ (_05226_, _05225_, _05215_);
  and _13623_ (_05227_, _05058_, _05056_);
  and _13624_ (_05228_, _05227_, _05048_);
  not _13625_ (_05229_, _05228_);
  and _13626_ (_05230_, _05217_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and _13627_ (_05231_, _05230_, _05221_);
  not _13628_ (_05232_, _05231_);
  nor _13629_ (_05233_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  and _13630_ (_05234_, _05233_, _05036_);
  not _13631_ (_05236_, _05234_);
  and _13632_ (_05237_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  and _13633_ (_05238_, _05237_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  not _13634_ (_05239_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and _13635_ (_05240_, _05239_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  and _13636_ (_05241_, _05240_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor _13637_ (_05242_, _05241_, _05238_);
  and _13638_ (_05243_, _05242_, _05236_);
  and _13639_ (_05244_, _05243_, _05059_);
  nor _13640_ (_05245_, _05244_, _05232_);
  and _13641_ (_05246_, _05245_, _05229_);
  nor _13642_ (_05247_, _05246_, _05226_);
  and _13643_ (_05248_, _05243_, _05048_);
  not _13644_ (_05249_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  and _13645_ (_05250_, _04859_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and _13646_ (_05252_, _05250_, _05249_);
  not _13647_ (_05253_, _05220_);
  nor _13648_ (_05254_, _05253_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and _13649_ (_05255_, _05254_, _05252_);
  not _13650_ (_05256_, _05255_);
  nor _13651_ (_05257_, _05256_, _05248_);
  nor _13652_ (_05258_, _05250_, _05217_);
  and _13653_ (_05259_, _05258_, _05254_);
  nor _13654_ (_05260_, _05243_, _05048_);
  nor _13655_ (_05261_, _05260_, _05248_);
  and _13656_ (_05262_, _05261_, _05259_);
  nor _13657_ (_05263_, _05262_, _05257_);
  not _13658_ (_05264_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and _13659_ (_05265_, \oc8051_top_1.oc8051_decoder1.alu_op [2], _04859_);
  and _13660_ (_05266_, _05265_, _05264_);
  and _13661_ (_05267_, _05266_, _05230_);
  and _13662_ (_05268_, _05267_, _05260_);
  and _13663_ (_05269_, _05266_, _05218_);
  and _13664_ (_05270_, _05269_, _05048_);
  nor _13665_ (_05271_, _05270_, _05268_);
  nor _13666_ (_05272_, _05265_, _05220_);
  and _13667_ (_05273_, _05272_, _05258_);
  not _13668_ (_05274_, _05273_);
  nand _13669_ (_05275_, _05272_, _05250_);
  nand _13670_ (_05276_, _05266_, _05249_);
  and _13671_ (_05277_, _05276_, _05275_);
  and _13672_ (_05278_, _05277_, _05274_);
  and _13673_ (_05279_, _05221_, _05249_);
  and _13674_ (_05280_, _05254_, _05217_);
  nor _13675_ (_05281_, _05280_, _05279_);
  and _13676_ (_05282_, _05281_, _05278_);
  nor _13677_ (_05283_, _05282_, _05048_);
  not _13678_ (_05284_, _05283_);
  and _13679_ (_05285_, _05284_, _05271_);
  and _13680_ (_05286_, _05285_, _05263_);
  and _13681_ (_05287_, _05286_, _05247_);
  not _13682_ (_05288_, _05287_);
  and _13683_ (_05289_, _05288_, _05009_);
  or _13684_ (_05290_, _05289_, _05010_);
  and _13685_ (_13054_, _05290_, _04856_);
  and _13686_ (_05291_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], _04859_);
  and _13687_ (_05292_, _05291_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  not _13688_ (_05293_, _05292_);
  nor _13689_ (_05294_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  not _13690_ (_05295_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and _13691_ (_05296_, _05295_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _13692_ (_05297_, _05296_, _05294_);
  not _13693_ (_05298_, _05297_);
  nor _13694_ (_05299_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and _13695_ (_05300_, _05022_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _13696_ (_05301_, _05300_, _05299_);
  not _13697_ (_05303_, _05301_);
  nor _13698_ (_05304_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and _13699_ (_05305_, _05185_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _13700_ (_05306_, _05305_, _05304_);
  not _13701_ (_05307_, _05306_);
  nor _13702_ (_05308_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and _13703_ (_05309_, _05089_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _13704_ (_05310_, _05309_, _05308_);
  nor _13705_ (_05312_, _05032_, ABINPUT[8]);
  nor _13706_ (_05313_, _05034_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  nor _13707_ (_05314_, _05313_, _05312_);
  and _13708_ (_05315_, _05314_, _05233_);
  not _13709_ (_05316_, _05315_);
  and _13710_ (_05317_, _05237_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  and _13711_ (_05318_, _05240_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor _13712_ (_05319_, _05318_, _05317_);
  and _13713_ (_05320_, _05319_, _05316_);
  not _13714_ (_05321_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  nor _13715_ (_05322_, _05019_, _05321_);
  not _13716_ (_05323_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  nor _13717_ (_05324_, _05015_, _05323_);
  nor _13718_ (_05325_, _05324_, _05322_);
  nor _13719_ (_05326_, _05024_, _05295_);
  not _13720_ (_05327_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor _13721_ (_05328_, _05027_, _05327_);
  nor _13722_ (_05329_, _05328_, _05326_);
  and _13723_ (_05330_, _05329_, _05325_);
  and _13724_ (_05331_, _05314_, _05037_);
  not _13725_ (_05332_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor _13726_ (_05333_, _05043_, _05332_);
  and _13727_ (_05334_, _05040_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [7]);
  nor _13728_ (_05335_, _05334_, _05333_);
  not _13729_ (_05336_, _05335_);
  nor _13730_ (_05337_, _05336_, _05331_);
  and _13731_ (_05338_, _05337_, _05330_);
  nor _13732_ (_05339_, _05338_, _05320_);
  not _13733_ (_05340_, _05339_);
  and _13734_ (_05341_, _05233_, _05073_);
  not _13735_ (_05342_, _05341_);
  and _13736_ (_05343_, _05237_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  and _13737_ (_05344_, _05240_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor _13738_ (_05345_, _05344_, _05343_);
  and _13739_ (_05346_, _05345_, _05342_);
  nor _13740_ (_05347_, _05346_, _05081_);
  and _13741_ (_05348_, _05346_, _05081_);
  nor _13742_ (_05349_, _05348_, _05347_);
  not _13743_ (_05350_, _05233_);
  nor _13744_ (_05351_, _05350_, _05096_);
  not _13745_ (_05352_, _05351_);
  and _13746_ (_05353_, _05237_, \oc8051_top_1.oc8051_memory_interface1.imm_r [3]);
  and _13747_ (_05354_, _05240_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor _13748_ (_05355_, _05354_, _05353_);
  and _13749_ (_05356_, _05355_, _05352_);
  nor _13750_ (_05357_, _05356_, _05103_);
  and _13751_ (_05359_, _05356_, _05103_);
  nor _13752_ (_05360_, _05359_, _05357_);
  not _13753_ (_05362_, _05360_);
  or _13754_ (_05363_, _05350_, _05165_);
  and _13755_ (_05365_, _05237_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  and _13756_ (_05366_, _05240_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor _13757_ (_05367_, _05366_, _05365_);
  and _13758_ (_05368_, _05367_, _05363_);
  nor _13759_ (_05369_, _05368_, _05172_);
  not _13760_ (_05370_, _05369_);
  and _13761_ (_05371_, _05368_, _05172_);
  nor _13762_ (_05372_, _05371_, _05369_);
  or _13763_ (_05373_, _05350_, _05130_);
  nand _13764_ (_05374_, _05237_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  nand _13765_ (_05375_, _05240_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and _13766_ (_05376_, _05375_, _05374_);
  nand _13767_ (_05377_, _05376_, _05373_);
  and _13768_ (_05378_, _05377_, _05207_);
  or _13769_ (_05379_, _05350_, _05119_);
  nand _13770_ (_05380_, _05237_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  nand _13771_ (_05381_, _05240_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and _13772_ (_05382_, _05381_, _05380_);
  and _13773_ (_05383_, _05382_, _05379_);
  not _13774_ (_05384_, _05383_);
  and _13775_ (_05385_, _05384_, _05206_);
  and _13776_ (_05386_, _05376_, _05373_);
  and _13777_ (_05387_, _05386_, _05151_);
  nor _13778_ (_05388_, _05387_, _05378_);
  and _13779_ (_05389_, _05388_, _05385_);
  or _13780_ (_05390_, _05389_, _05378_);
  nand _13781_ (_05391_, _05390_, _05372_);
  nand _13782_ (_05392_, _05391_, _05370_);
  and _13783_ (_05393_, _05392_, _05362_);
  nor _13784_ (_05394_, _05392_, _05362_);
  or _13785_ (_05395_, _05394_, _05393_);
  and _13786_ (_05396_, _05383_, _05126_);
  nor _13787_ (_05397_, _05396_, _05385_);
  and _13788_ (_05398_, _05397_, _05059_);
  and _13789_ (_05399_, _05398_, _05388_);
  or _13790_ (_05400_, _05390_, _05372_);
  and _13791_ (_05401_, _05400_, _05391_);
  and _13792_ (_05402_, _05401_, _05399_);
  and _13793_ (_05403_, _05402_, _05395_);
  not _13794_ (_05404_, _05359_);
  and _13795_ (_05405_, _05392_, _05404_);
  or _13796_ (_05406_, _05405_, _05357_);
  or _13797_ (_05407_, _05406_, _05403_);
  nand _13798_ (_05408_, _05407_, _05349_);
  and _13799_ (_05409_, _05233_, _05191_);
  not _13800_ (_05410_, _05409_);
  and _13801_ (_05411_, _05237_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  and _13802_ (_05412_, _05240_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor _13803_ (_05413_, _05412_, _05411_);
  and _13804_ (_05414_, _05413_, _05410_);
  nor _13805_ (_05415_, _05414_, _05199_);
  and _13806_ (_05416_, _05414_, _05199_);
  nor _13807_ (_05417_, _05416_, _05415_);
  and _13808_ (_05418_, _05417_, _05347_);
  nor _13809_ (_05419_, _05417_, _05347_);
  nor _13810_ (_05420_, _05419_, _05418_);
  not _13811_ (_05421_, _05420_);
  or _13812_ (_05422_, _05421_, _05408_);
  not _13813_ (_05423_, _05261_);
  nor _13814_ (_05424_, _05418_, _05415_);
  nor _13815_ (_05425_, _05424_, _05423_);
  and _13816_ (_05426_, _05424_, _05423_);
  nor _13817_ (_05427_, _05426_, _05425_);
  not _13818_ (_05428_, _05427_);
  or _13819_ (_05429_, _05428_, _05422_);
  nor _13820_ (_05430_, _05425_, _05260_);
  and _13821_ (_05431_, _05430_, _05429_);
  and _13822_ (_05432_, _05338_, _05320_);
  or _13823_ (_05433_, _05432_, _05431_);
  nand _13824_ (_05434_, _05433_, _05340_);
  nor _13825_ (_05435_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and _13826_ (_05436_, _05111_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _13827_ (_05437_, _05436_, _05435_);
  and _13828_ (_05438_, _05437_, _05434_);
  nor _13829_ (_05439_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and _13830_ (_05440_, _05142_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _13831_ (_05441_, _05440_, _05439_);
  and _13832_ (_05442_, _05441_, _05438_);
  nor _13833_ (_05443_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and _13834_ (_05444_, _05157_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _13835_ (_05445_, _05444_, _05443_);
  and _13836_ (_05446_, _05445_, _05442_);
  and _13837_ (_05447_, _05446_, _05310_);
  nor _13838_ (_05448_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and _13839_ (_05449_, _05067_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _13840_ (_05450_, _05449_, _05448_);
  nand _13841_ (_05451_, _05450_, _05447_);
  or _13842_ (_05452_, _05451_, _05307_);
  or _13843_ (_05453_, _05452_, _05303_);
  or _13844_ (_05454_, _05453_, _05298_);
  and _13845_ (_05455_, _05272_, _05252_);
  nand _13846_ (_05456_, _05453_, _05298_);
  and _13847_ (_05457_, _05456_, _05455_);
  and _13848_ (_05458_, _05457_, _05454_);
  not _13849_ (_05459_, _05320_);
  nor _13850_ (_05460_, _05243_, _05059_);
  nor _13851_ (_05461_, _05460_, _05244_);
  and _13852_ (_05462_, _05199_, _05048_);
  and _13853_ (_05463_, _05338_, _05462_);
  and _13854_ (_05464_, _05463_, _05176_);
  and _13855_ (_05465_, _05464_, _05383_);
  and _13856_ (_05466_, _05465_, _05386_);
  and _13857_ (_05467_, _05466_, _05368_);
  and _13858_ (_05468_, _05467_, _05356_);
  and _13859_ (_05469_, _05468_, _05346_);
  and _13860_ (_05470_, _05414_, _05059_);
  nand _13861_ (_05471_, _05470_, _05469_);
  not _13862_ (_05472_, _05368_);
  nor _13863_ (_05473_, _05338_, _05048_);
  and _13864_ (_05474_, _05473_, _05211_);
  and _13865_ (_05475_, _05474_, _05210_);
  and _13866_ (_05476_, _05475_, _05384_);
  and _13867_ (_05477_, _05476_, _05377_);
  and _13868_ (_05478_, _05477_, _05472_);
  nor _13869_ (_05479_, _05414_, _05059_);
  nor _13870_ (_05480_, _05356_, _05346_);
  and _13871_ (_05481_, _05480_, _05479_);
  nand _13872_ (_05482_, _05481_, _05478_);
  and _13873_ (_05483_, _05482_, _05471_);
  nor _13874_ (_05484_, _05483_, _05461_);
  nand _13875_ (_05485_, _05484_, _05459_);
  or _13876_ (_05486_, _05484_, _05459_);
  and _13877_ (_05487_, _05486_, _05485_);
  and _13878_ (_05488_, _05487_, _05223_);
  and _13879_ (_05489_, _05254_, _05230_);
  not _13880_ (_05490_, _05489_);
  nor _13881_ (_05491_, _05490_, _05103_);
  and _13882_ (_05492_, _05231_, _05227_);
  or _13883_ (_05493_, _05492_, _05273_);
  and _13884_ (_05494_, _05493_, _05459_);
  or _13885_ (_05495_, _05232_, _05227_);
  nor _13886_ (_05496_, _05495_, _05338_);
  and _13887_ (_05497_, _05266_, _05258_);
  and _13888_ (_05498_, _05497_, ABINPUT001[16]);
  and _13889_ (_05499_, _05272_, _05230_);
  and _13890_ (_05500_, _05499_, ABINPUT000[16]);
  or _13891_ (_05501_, _05500_, _05498_);
  or _13892_ (_05502_, _05501_, _05496_);
  or _13893_ (_05503_, _05502_, _05494_);
  or _13894_ (_05504_, _05503_, _05491_);
  or _13895_ (_05506_, _05504_, _05488_);
  or _13896_ (_05507_, _05506_, _05458_);
  or _13897_ (_05509_, _05507_, _05293_);
  and _13898_ (_05510_, _04861_, _04885_);
  and _13899_ (_05512_, _05510_, _04947_);
  not _13900_ (_05513_, _04893_);
  nor _13901_ (_05515_, _04904_, _05513_);
  and _13902_ (_05517_, _05515_, _04993_);
  nor _13903_ (_05519_, _04971_, _04958_);
  and _13904_ (_05520_, _05519_, _04984_);
  and _13905_ (_05522_, _05520_, _05517_);
  and _13906_ (_05524_, _05522_, _05512_);
  nor _13907_ (_05525_, _05338_, _05274_);
  nor _13908_ (_05526_, _05338_, _05059_);
  nor _13909_ (_05527_, _05320_, _05227_);
  or _13910_ (_05528_, _05527_, _05526_);
  and _13911_ (_05529_, _05528_, _05231_);
  not _13912_ (_05530_, _05338_);
  nor _13913_ (_05531_, _05227_, _05048_);
  nor _13914_ (_05532_, _05531_, _05228_);
  and _13915_ (_05533_, _05532_, _05214_);
  nor _13916_ (_05534_, _05533_, _05530_);
  and _13917_ (_05535_, _05533_, _05530_);
  nor _13918_ (_05536_, _05535_, _05534_);
  and _13919_ (_05537_, _05536_, _05223_);
  nor _13920_ (_05538_, _05537_, _05529_);
  and _13921_ (_05540_, _05252_, _05221_);
  and _13922_ (_05541_, _05540_, _05059_);
  and _13923_ (_05542_, _05258_, _05221_);
  and _13924_ (_05543_, _05542_, _05206_);
  nor _13925_ (_05544_, _05543_, _05541_);
  nand _13926_ (_05545_, _05544_, _05538_);
  and _13927_ (_05546_, _05280_, _05049_);
  not _13928_ (_05547_, _05546_);
  nor _13929_ (_05548_, _05432_, _05256_);
  nor _13930_ (_05549_, _05432_, _05339_);
  and _13931_ (_05550_, _05549_, _05259_);
  nor _13932_ (_05551_, _05550_, _05548_);
  nand _13933_ (_05552_, _05551_, _05547_);
  or _13934_ (_05553_, _05552_, _05545_);
  and _13935_ (_05554_, _05339_, _05267_);
  and _13936_ (_05555_, _05338_, _05269_);
  nor _13937_ (_05556_, _05555_, _05554_);
  and _13938_ (_05557_, _05266_, _05252_);
  not _13939_ (_05558_, _05557_);
  nor _13940_ (_05559_, _05173_, _05103_);
  and _13941_ (_05560_, _05559_, _05557_);
  not _13942_ (_05561_, _05560_);
  or _13943_ (_05562_, _05338_, _05462_);
  and _13944_ (_05563_, _05562_, _05227_);
  and _13945_ (_05564_, _05563_, _05561_);
  not _13946_ (_05565_, _05081_);
  and _13947_ (_05567_, _05560_, _05565_);
  nor _13948_ (_05568_, _05567_, _05564_);
  and _13949_ (_05569_, _05568_, _05462_);
  or _13950_ (_05570_, _05569_, _05564_);
  and _13951_ (_05571_, _05570_, _05338_);
  nor _13952_ (_05572_, _05570_, _05338_);
  or _13953_ (_05573_, _05572_, _05571_);
  nor _13954_ (_05574_, _05573_, _05558_);
  and _13955_ (_05576_, _05497_, ABINPUT001[8]);
  nor _13956_ (_05577_, _05576_, _05574_);
  nand _13957_ (_05578_, _05577_, _05556_);
  and _13958_ (_05579_, _05549_, _05431_);
  nor _13959_ (_05580_, _05549_, _05431_);
  or _13960_ (_05581_, _05580_, _05579_);
  and _13961_ (_05582_, _05581_, _05455_);
  and _13962_ (_05583_, _05272_, _05218_);
  not _13963_ (_05584_, _05583_);
  not _13964_ (_05585_, _05549_);
  and _13965_ (_05586_, _05243_, _05049_);
  not _13966_ (_05587_, _05199_);
  and _13967_ (_05588_, _05414_, _05587_);
  not _13968_ (_05589_, _05346_);
  and _13969_ (_05590_, _05589_, _05081_);
  nor _13970_ (_05591_, _05417_, _05590_);
  nor _13971_ (_05592_, _05591_, _05588_);
  nor _13972_ (_05593_, _05592_, _05261_);
  nor _13973_ (_05594_, _05593_, _05586_);
  and _13974_ (_05595_, _05592_, _05261_);
  nor _13975_ (_05596_, _05595_, _05593_);
  not _13976_ (_05597_, _05596_);
  and _13977_ (_05598_, _05417_, _05590_);
  nor _13978_ (_05599_, _05598_, _05591_);
  not _13979_ (_05600_, _05599_);
  not _13980_ (_05601_, _05349_);
  nor _13981_ (_05602_, _05472_, _05172_);
  or _13982_ (_05603_, _05377_, _05151_);
  and _13983_ (_05604_, _05384_, _05126_);
  or _13984_ (_05605_, _05604_, _05388_);
  nand _13985_ (_05606_, _05605_, _05603_);
  not _13986_ (_05607_, _05606_);
  nor _13987_ (_05608_, _05607_, _05372_);
  nor _13988_ (_05609_, _05608_, _05602_);
  nor _13989_ (_05610_, _05609_, _05360_);
  and _13990_ (_05611_, _05609_, _05360_);
  or _13991_ (_05612_, _05611_, _05610_);
  and _13992_ (_05613_, _05607_, _05372_);
  or _13993_ (_05614_, _05613_, _05608_);
  and _13994_ (_05615_, _05604_, _05388_);
  not _13995_ (_05616_, _05615_);
  nand _13996_ (_05617_, _05616_, _05605_);
  nor _13997_ (_05618_, _05397_, _05227_);
  and _13998_ (_05619_, _05618_, _05617_);
  and _13999_ (_05620_, _05619_, _05614_);
  and _14000_ (_05621_, _05620_, _05612_);
  not _14001_ (_05622_, _05356_);
  or _14002_ (_05623_, _05622_, _05103_);
  and _14003_ (_05624_, _05622_, _05103_);
  or _14004_ (_05625_, _05609_, _05624_);
  and _14005_ (_05626_, _05625_, _05623_);
  or _14006_ (_05627_, _05626_, _05621_);
  and _14007_ (_05628_, _05627_, _05601_);
  and _14008_ (_05629_, _05628_, _05600_);
  and _14009_ (_05630_, _05629_, _05597_);
  or _14010_ (_05631_, _05630_, _05594_);
  and _14011_ (_05632_, _05631_, _05585_);
  nor _14012_ (_05633_, _05631_, _05585_);
  nor _14013_ (_05634_, _05633_, _05632_);
  nor _14014_ (_05635_, _05634_, _05584_);
  and _14015_ (_05636_, _05499_, ABINPUT000[8]);
  or _14016_ (_05637_, _05636_, _05635_);
  or _14017_ (_05638_, _05637_, _05582_);
  or _14018_ (_05639_, _05638_, _05578_);
  or _14019_ (_05640_, _05639_, _05553_);
  or _14020_ (_05641_, _05640_, _05525_);
  and _14021_ (_05642_, _05641_, _05524_);
  not _14022_ (_05643_, _05524_);
  and _14023_ (_05644_, _05643_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or _14024_ (_05645_, _05644_, _05292_);
  or _14025_ (_05646_, _05645_, _05642_);
  and _14026_ (_05647_, _05646_, _04856_);
  and _14027_ (_03221_, _05647_, _05509_);
  nor _14028_ (_05648_, _05356_, _05232_);
  nand _14029_ (_05649_, _05209_, _05227_);
  nand _14030_ (_05650_, _05174_, _05059_);
  and _14031_ (_05651_, _05650_, _05649_);
  nand _14032_ (_05652_, _05651_, _05103_);
  or _14033_ (_05653_, _05651_, _05103_);
  and _14034_ (_05654_, _05653_, _05223_);
  and _14035_ (_05655_, _05654_, _05652_);
  nor _14036_ (_05656_, _05655_, _05648_);
  nor _14037_ (_05657_, _05282_, _05103_);
  not _14038_ (_05658_, _05657_);
  and _14039_ (_05659_, _05360_, _05259_);
  not _14040_ (_05660_, _05659_);
  nor _14041_ (_05661_, _05359_, _05256_);
  not _14042_ (_05662_, _05661_);
  and _14043_ (_05663_, _05357_, _05267_);
  and _14044_ (_05664_, _05269_, _05103_);
  nor _14045_ (_05665_, _05664_, _05663_);
  and _14046_ (_05666_, _05665_, _05662_);
  and _14047_ (_05667_, _05666_, _05660_);
  and _14048_ (_05668_, _05667_, _05658_);
  and _14049_ (_05669_, _05668_, _05656_);
  not _14050_ (_05670_, _05669_);
  and _14051_ (_05671_, _05002_, _04861_);
  and _14052_ (_05672_, _05671_, _05670_);
  not _14053_ (_05673_, _04861_);
  and _14054_ (_05674_, _04991_, _04994_);
  and _14055_ (_05675_, _04999_, _04994_);
  and _14056_ (_05676_, _05001_, _04994_);
  or _14057_ (_05677_, _05676_, _05675_);
  nor _14058_ (_05678_, _05677_, _05674_);
  and _14059_ (_05679_, _04994_, _04987_);
  nor _14060_ (_05680_, _05002_, _05679_);
  and _14061_ (_05681_, _05680_, _05678_);
  or _14062_ (_05682_, _05681_, _05673_);
  or _14063_ (_05683_, _05682_, _04995_);
  and _14064_ (_05684_, _05683_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  or _14065_ (_05685_, _05684_, _05672_);
  and _14066_ (_04850_, _05685_, _04856_);
  and _14067_ (_05686_, _05199_, _05227_);
  not _14068_ (_05687_, _05686_);
  nor _14069_ (_05688_, _05470_, _05232_);
  and _14070_ (_05689_, _05688_, _05687_);
  and _14071_ (_05690_, _05081_, _05227_);
  not _14072_ (_05692_, _05690_);
  and _14073_ (_05693_, _05210_, _05227_);
  or _14074_ (_05694_, _05693_, _05176_);
  and _14075_ (_05696_, _05694_, _05692_);
  or _14076_ (_05698_, _05587_, _05696_);
  nand _14077_ (_05699_, _05587_, _05696_);
  and _14078_ (_05700_, _05699_, _05223_);
  and _14079_ (_05701_, _05700_, _05698_);
  nor _14080_ (_05702_, _05701_, _05689_);
  nor _14081_ (_05703_, _05282_, _05199_);
  not _14082_ (_05704_, _05703_);
  and _14083_ (_05705_, _05417_, _05259_);
  not _14084_ (_05707_, _05705_);
  nor _14085_ (_05708_, _05416_, _05256_);
  not _14086_ (_05710_, _05708_);
  and _14087_ (_05711_, _05415_, _05267_);
  and _14088_ (_05713_, _05269_, _05199_);
  nor _14089_ (_05714_, _05713_, _05711_);
  and _14090_ (_05715_, _05714_, _05710_);
  and _14091_ (_05716_, _05715_, _05707_);
  and _14092_ (_05717_, _05716_, _05704_);
  nand _14093_ (_05718_, _05717_, _05702_);
  and _14094_ (_05719_, _05000_, _04861_);
  and _14095_ (_05720_, _05719_, _05718_);
  nand _14096_ (_05721_, _05004_, _04861_);
  not _14097_ (_05722_, _05721_);
  nand _14098_ (_05723_, _05722_, _05682_);
  and _14099_ (_05724_, _05723_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  or _14100_ (_05725_, _05724_, _05720_);
  and _14101_ (_04852_, _05725_, _04856_);
  not _14102_ (_05726_, \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  nor _14103_ (_05727_, \oc8051_top_1.oc8051_memory_interface1.imem_wait , \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  and _14104_ (_05728_, _05727_, _05726_);
  nor _14105_ (_05729_, \oc8051_top_1.oc8051_decoder1.state [0], \oc8051_top_1.oc8051_decoder1.state [1]);
  and _14106_ (_05730_, _05729_, _04859_);
  and _14107_ (_05731_, _05730_, _05728_);
  not _14108_ (_05732_, _05731_);
  not _14109_ (_05733_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  not _14110_ (_05734_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  not _14111_ (_05735_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  not _14112_ (_05736_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  not _14113_ (_05737_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  nor _14114_ (_05738_, _05737_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nand _14115_ (_05739_, _05738_, _05736_);
  or _14116_ (_05740_, _05739_, _05735_);
  and _14117_ (_05741_, _05737_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _14118_ (_05742_, _05741_, _05736_);
  nand _14119_ (_05743_, _05742_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  and _14120_ (_05744_, _05743_, _05740_);
  not _14121_ (_05745_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nand _14122_ (_05746_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  or _14123_ (_05747_, _05746_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  or _14124_ (_05748_, _05747_, _05745_);
  not _14125_ (_05749_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  or _14126_ (_05750_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  or _14127_ (_05751_, _05750_, _05736_);
  or _14128_ (_05752_, _05751_, _05749_);
  and _14129_ (_05753_, _05752_, _05748_);
  not _14130_ (_05754_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nor _14131_ (_05755_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  or _14132_ (_05756_, _05755_, _05736_);
  or _14133_ (_05757_, _05756_, _05754_);
  and _14134_ (_05758_, _05755_, _05736_);
  nand _14135_ (_05759_, _05758_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  and _14136_ (_05760_, _05759_, _05757_);
  and _14137_ (_05761_, _05760_, _05753_);
  nand _14138_ (_05762_, _05761_, _05744_);
  nand _14139_ (_05763_, _05762_, _05734_);
  nand _14140_ (_05764_, _05763_, _05733_);
  nor _14141_ (_05765_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], _05733_);
  not _14142_ (_05766_, _05765_);
  and _14143_ (_05767_, _05766_, _05764_);
  or _14144_ (_05768_, _05767_, _05732_);
  not _14145_ (_05769_, _05728_);
  nor _14146_ (_05770_, _05730_, \oc8051_top_1.oc8051_decoder1.op [0]);
  nor _14147_ (_05771_, _05770_, _05769_);
  and _14148_ (_05772_, _05771_, _05768_);
  not _14149_ (_05773_, _05772_);
  not _14150_ (_05774_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  or _14151_ (_05775_, _05747_, _05774_);
  nand _14152_ (_05776_, _05742_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  and _14153_ (_05777_, _05776_, _05775_);
  not _14154_ (_05778_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  or _14155_ (_05779_, _05756_, _05778_);
  nand _14156_ (_05780_, _05758_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  and _14157_ (_05781_, _05780_, _05779_);
  not _14158_ (_05782_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  or _14159_ (_05783_, _05751_, _05782_);
  not _14160_ (_05784_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  or _14161_ (_05785_, _05739_, _05784_);
  and _14162_ (_05786_, _05785_, _05783_);
  and _14163_ (_05787_, _05786_, _05781_);
  nand _14164_ (_05788_, _05787_, _05777_);
  nand _14165_ (_05789_, _05788_, _05734_);
  nand _14166_ (_05790_, _05789_, _05733_);
  nor _14167_ (_05791_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], _05733_);
  not _14168_ (_05792_, _05791_);
  and _14169_ (_05793_, _05792_, _05790_);
  or _14170_ (_05794_, _05793_, _05732_);
  nor _14171_ (_05795_, _05730_, \oc8051_top_1.oc8051_decoder1.op [2]);
  nor _14172_ (_05796_, _05795_, _05769_);
  nand _14173_ (_05797_, _05796_, _05794_);
  and _14174_ (_05798_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], \oc8051_top_1.oc8051_memory_interface1.cdone );
  not _14175_ (_05799_, _05798_);
  nand _14176_ (_05800_, _05758_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  nand _14177_ (_05801_, _05742_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  and _14178_ (_05802_, _05801_, _05800_);
  not _14179_ (_05803_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  or _14180_ (_05804_, _05756_, _05803_);
  not _14181_ (_05805_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  or _14182_ (_05806_, _05751_, _05805_);
  and _14183_ (_05807_, _05806_, _05804_);
  not _14184_ (_05808_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  or _14185_ (_05810_, _05747_, _05808_);
  not _14186_ (_05811_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  or _14187_ (_05812_, _05739_, _05811_);
  and _14188_ (_05813_, _05812_, _05810_);
  and _14189_ (_05814_, _05813_, _05807_);
  and _14190_ (_05815_, _05814_, _05802_);
  or _14191_ (_05816_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  or _14192_ (_05817_, _05816_, _05815_);
  nand _14193_ (_05818_, _05817_, _05799_);
  or _14194_ (_05819_, _05818_, _05732_);
  nor _14195_ (_05820_, _05730_, \oc8051_top_1.oc8051_decoder1.op [3]);
  nor _14196_ (_05821_, _05820_, _05769_);
  nand _14197_ (_05822_, _05821_, _05819_);
  and _14198_ (_05823_, _05822_, _05797_);
  not _14199_ (_05824_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  or _14200_ (_05825_, _05751_, _05824_);
  not _14201_ (_05826_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  or _14202_ (_05827_, _05747_, _05826_);
  and _14203_ (_05828_, _05827_, _05825_);
  not _14204_ (_05829_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  or _14205_ (_05830_, _05739_, _05829_);
  and _14206_ (_05831_, _05830_, _05828_);
  nand _14207_ (_05832_, _05742_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  and _14208_ (_05833_, _05832_, _05734_);
  not _14209_ (_05834_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  or _14210_ (_05835_, _05756_, _05834_);
  nand _14211_ (_05836_, _05758_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  and _14212_ (_05837_, _05836_, _05835_);
  and _14213_ (_05838_, _05837_, _05833_);
  nand _14214_ (_05839_, _05838_, _05831_);
  or _14215_ (_05840_, _05839_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor _14216_ (_05841_, _05733_, \oc8051_top_1.oc8051_memory_interface1.cdata [1]);
  not _14217_ (_05842_, _05841_);
  and _14218_ (_05843_, _05842_, _05840_);
  or _14219_ (_05844_, _05843_, _05732_);
  nor _14220_ (_05845_, _05730_, \oc8051_top_1.oc8051_decoder1.op [1]);
  nor _14221_ (_05846_, _05845_, _05769_);
  and _14222_ (_05847_, _05846_, _05844_);
  and _14223_ (_05848_, _05847_, _05823_);
  and _14224_ (_05849_, _05848_, _05773_);
  not _14225_ (_05850_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  or _14226_ (_05851_, _05751_, _05850_);
  not _14227_ (_05852_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  or _14228_ (_05853_, _05747_, _05852_);
  and _14229_ (_05854_, _05853_, _05851_);
  not _14230_ (_05855_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  or _14231_ (_05856_, _05739_, _05855_);
  and _14232_ (_05857_, _05856_, _05854_);
  nand _14233_ (_05858_, _05742_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  and _14234_ (_05860_, _05858_, _05734_);
  not _14235_ (_05861_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  or _14236_ (_05862_, _05756_, _05861_);
  nand _14237_ (_05863_, _05758_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  and _14238_ (_05864_, _05863_, _05862_);
  and _14239_ (_05865_, _05864_, _05860_);
  nand _14240_ (_05866_, _05865_, _05857_);
  or _14241_ (_05867_, _05866_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor _14242_ (_05868_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], _05733_);
  not _14243_ (_05869_, _05868_);
  and _14244_ (_05870_, _05869_, _05867_);
  or _14245_ (_05871_, _05870_, _05732_);
  nor _14246_ (_05872_, _05730_, \oc8051_top_1.oc8051_decoder1.op [4]);
  nor _14247_ (_05873_, _05872_, _05769_);
  and _14248_ (_05874_, _05873_, _05871_);
  not _14249_ (_05875_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  or _14250_ (_05876_, _05739_, _05875_);
  nand _14251_ (_05877_, _05742_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  and _14252_ (_05878_, _05877_, _05876_);
  not _14253_ (_05879_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  or _14254_ (_05880_, _05747_, _05879_);
  not _14255_ (_05881_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  or _14256_ (_05882_, _05751_, _05881_);
  and _14257_ (_05883_, _05882_, _05880_);
  not _14258_ (_05884_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  or _14259_ (_05885_, _05756_, _05884_);
  nand _14260_ (_05886_, _05758_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  and _14261_ (_05888_, _05886_, _05885_);
  and _14262_ (_05889_, _05888_, _05883_);
  nand _14263_ (_05890_, _05889_, _05878_);
  and _14264_ (_05891_, _05890_, _05734_);
  or _14265_ (_05892_, _05891_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor _14266_ (_05893_, \oc8051_top_1.oc8051_memory_interface1.cdata [5], _05733_);
  not _14267_ (_05894_, _05893_);
  and _14268_ (_05895_, _05894_, _05892_);
  or _14269_ (_05896_, _05895_, _05732_);
  nor _14270_ (_05897_, _05730_, \oc8051_top_1.oc8051_decoder1.op [5]);
  nor _14271_ (_05898_, _05897_, _05769_);
  and _14272_ (_05899_, _05898_, _05896_);
  not _14273_ (_05900_, _05899_);
  nand _14274_ (_05901_, _05758_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  nand _14275_ (_05902_, _05742_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  and _14276_ (_05903_, _05902_, _05901_);
  not _14277_ (_05904_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  or _14278_ (_05905_, _05756_, _05904_);
  not _14279_ (_05906_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  or _14280_ (_05907_, _05747_, _05906_);
  and _14281_ (_05908_, _05907_, _05905_);
  not _14282_ (_05909_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  or _14283_ (_05910_, _05751_, _05909_);
  not _14284_ (_05911_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  or _14285_ (_05912_, _05739_, _05911_);
  and _14286_ (_05913_, _05912_, _05910_);
  and _14287_ (_05914_, _05913_, _05908_);
  and _14288_ (_05915_, _05914_, _05903_);
  or _14289_ (_05916_, _05915_, _05816_);
  and _14290_ (_05917_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  not _14291_ (_05918_, _05917_);
  nand _14292_ (_05919_, _05918_, _05916_);
  or _14293_ (_05920_, _05919_, _05732_);
  nor _14294_ (_05921_, _05730_, \oc8051_top_1.oc8051_decoder1.op [7]);
  nor _14295_ (_05922_, _05921_, _05769_);
  nand _14296_ (_05923_, _05922_, _05920_);
  and _14297_ (_05924_, _05758_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  and _14298_ (_05925_, _05742_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  or _14299_ (_05926_, _05925_, _05924_);
  and _14300_ (_05927_, _05750_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and _14301_ (_05928_, _05927_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nor _14302_ (_05929_, _05746_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and _14303_ (_05930_, _05929_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  or _14304_ (_05932_, _05930_, _05928_);
  and _14305_ (_05933_, _05755_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and _14306_ (_05934_, _05933_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and _14307_ (_05935_, _05738_, _05736_);
  and _14308_ (_05936_, _05935_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  or _14309_ (_05937_, _05936_, _05934_);
  or _14310_ (_05938_, _05937_, _05932_);
  or _14311_ (_05939_, _05938_, _05926_);
  not _14312_ (_05940_, _05939_);
  nor _14313_ (_05941_, _05940_, _05816_);
  and _14314_ (_05942_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], \oc8051_top_1.oc8051_memory_interface1.cdone );
  or _14315_ (_05943_, _05942_, _05941_);
  or _14316_ (_05944_, _05943_, _05732_);
  nor _14317_ (_05945_, _05730_, \oc8051_top_1.oc8051_decoder1.op [6]);
  nor _14318_ (_05946_, _05945_, _05769_);
  nand _14319_ (_05947_, _05946_, _05944_);
  and _14320_ (_05948_, _05947_, _05923_);
  and _14321_ (_05949_, _05948_, _05900_);
  and _14322_ (_05950_, _05949_, _05874_);
  and _14323_ (_05951_, _05950_, _05849_);
  not _14324_ (_05952_, _05847_);
  and _14325_ (_05953_, _05772_, _05952_);
  and _14326_ (_05954_, _05953_, _05823_);
  and _14327_ (_05955_, _05954_, _05874_);
  or _14328_ (_05956_, _05955_, _05951_);
  not _14329_ (_05957_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and _14330_ (_05958_, \oc8051_top_1.oc8051_decoder1.state [1], _04859_);
  and _14331_ (_05959_, _05958_, _05957_);
  and _14332_ (_05960_, _05959_, _05956_);
  or _14333_ (_05961_, _05960_, \oc8051_top_1.oc8051_sfr1.wait_data );
  or _14334_ (_05962_, _05729_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and _14335_ (_05963_, _05796_, _05794_);
  and _14336_ (_05964_, _05847_, _05963_);
  and _14337_ (_05965_, _05964_, _05822_);
  and _14338_ (_05966_, _05965_, _05949_);
  and _14339_ (_05967_, _05946_, _05944_);
  and _14340_ (_05968_, _05967_, _05899_);
  and _14341_ (_05969_, _05968_, _05874_);
  and _14342_ (_05970_, _05969_, _05965_);
  or _14343_ (_05971_, _05970_, _05966_);
  not _14344_ (_05972_, _05874_);
  and _14345_ (_05973_, _05822_, _05972_);
  and _14346_ (_05974_, _05973_, _05964_);
  and _14347_ (_05976_, _05922_, _05920_);
  and _14348_ (_05977_, _05947_, _05976_);
  and _14349_ (_05978_, _05977_, _05899_);
  and _14350_ (_05979_, _05978_, _05974_);
  or _14351_ (_05980_, _05979_, _05971_);
  nor _14352_ (_05982_, _05772_, _05847_);
  and _14353_ (_05983_, _05982_, _05823_);
  and _14354_ (_05984_, _05967_, _05900_);
  and _14355_ (_05985_, _05984_, _05976_);
  and _14356_ (_05986_, _05985_, _05972_);
  and _14357_ (_05987_, _05986_, _05983_);
  and _14358_ (_05988_, _05985_, _05965_);
  or _14359_ (_05989_, _05988_, _05987_);
  or _14360_ (_05990_, _05989_, _05980_);
  or _14361_ (_05991_, _05990_, _05956_);
  and _14362_ (_05992_, _05991_, _05962_);
  not _14363_ (_05993_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and _14364_ (_05994_, \oc8051_top_1.oc8051_decoder1.state [0], _04859_);
  and _14365_ (_05995_, _05994_, _05993_);
  and _14366_ (_05996_, _05978_, _05972_);
  and _14367_ (_05997_, _05822_, _05963_);
  and _14368_ (_05998_, _05982_, _05997_);
  and _14369_ (_05999_, _05998_, _05996_);
  and _14370_ (_06000_, _05977_, _05900_);
  and _14371_ (_06001_, _06000_, _05972_);
  and _14372_ (_06002_, _06001_, _05998_);
  nor _14373_ (_06003_, _06002_, _05999_);
  not _14374_ (_06004_, _06003_);
  and _14375_ (_06005_, _06004_, _05995_);
  or _14376_ (_06006_, _06005_, _05992_);
  or _14377_ (_06007_, _06006_, _05961_);
  or _14378_ (_06008_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _04859_);
  and _14379_ (_06009_, _06008_, _04856_);
  and _14380_ (_04891_, _06009_, _06007_);
  nor _14381_ (_06010_, _05282_, _05151_);
  not _14382_ (_06011_, _06010_);
  and _14383_ (_06012_, _05151_, _05059_);
  and _14384_ (_06013_, _05207_, _05227_);
  nor _14385_ (_06014_, _06013_, _06012_);
  or _14386_ (_06015_, _06014_, _05126_);
  nand _14387_ (_06016_, _06014_, _05126_);
  and _14388_ (_06017_, _06016_, _05223_);
  nand _14389_ (_06018_, _06017_, _06015_);
  not _14390_ (_06019_, _05259_);
  or _14391_ (_06020_, _05387_, _05378_);
  or _14392_ (_06021_, _06020_, _06019_);
  or _14393_ (_06022_, _05387_, _05256_);
  nand _14394_ (_06023_, _05378_, _05267_);
  and _14395_ (_06024_, _05377_, _05231_);
  and _14396_ (_06025_, _05269_, _05151_);
  nor _14397_ (_06026_, _06025_, _06024_);
  and _14398_ (_06027_, _06026_, _06023_);
  and _14399_ (_06028_, _06027_, _06022_);
  and _14400_ (_06029_, _06028_, _06021_);
  and _14401_ (_06030_, _06029_, _06018_);
  and _14402_ (_06032_, _06030_, _06011_);
  not _14403_ (_06033_, _06032_);
  and _14404_ (_06034_, _06033_, _05009_);
  not _14405_ (_06035_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  nor _14406_ (_06036_, _05009_, _06035_);
  or _14407_ (_06037_, _06036_, _06034_);
  and _14408_ (_04983_, _06037_, _04856_);
  nand _14409_ (_06038_, _05008_, _05678_);
  or _14410_ (_06039_, _05003_, _05679_);
  and _14411_ (_06040_, _06039_, _04861_);
  or _14412_ (_06041_, _06040_, _06038_);
  and _14413_ (_06042_, _06041_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  and _14414_ (_06043_, _04992_, _04861_);
  and _14415_ (_06044_, _06043_, _06033_);
  or _14416_ (_06045_, _06044_, _06042_);
  and _14417_ (_05235_, _06045_, _04856_);
  not _14418_ (_06046_, _05675_);
  and _14419_ (_06047_, _06046_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  nor _14420_ (_06048_, _06032_, _06046_);
  or _14421_ (_06049_, _06048_, _05673_);
  or _14422_ (_06050_, _06049_, _06047_);
  or _14423_ (_06051_, _04861_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  and _14424_ (_06052_, _06051_, _04856_);
  and _14425_ (_06640_, _06052_, _06050_);
  and _14426_ (_06053_, _05338_, _05459_);
  nor _14427_ (_06054_, _05632_, _06053_);
  or _14428_ (_06055_, _06054_, _05584_);
  nand _14429_ (_06056_, _05434_, _05455_);
  nor _14430_ (_06057_, _05572_, _05059_);
  nand _14431_ (_06058_, _05572_, _05059_);
  nand _14432_ (_06059_, _06058_, _05557_);
  or _14433_ (_06060_, _06059_, _06057_);
  nor _14434_ (_06061_, _05338_, _05490_);
  not _14435_ (_06062_, _05052_);
  and _14436_ (_06063_, _05055_, _06062_);
  and _14437_ (_06064_, _05254_, _05218_);
  and _14438_ (_06065_, _05267_, _06062_);
  nor _14439_ (_06066_, _06065_, _06064_);
  nor _14440_ (_06067_, _06066_, _06063_);
  nor _14441_ (_06068_, _06067_, _06061_);
  and _14442_ (_06069_, _05058_, _05052_);
  and _14443_ (_06070_, _05259_, _05056_);
  nor _14444_ (_06071_, _06070_, _05255_);
  nor _14445_ (_06072_, _06071_, _06069_);
  not _14446_ (_06073_, _06072_);
  and _14447_ (_06074_, _05540_, _05206_);
  not _14448_ (_06075_, _05269_);
  and _14449_ (_06076_, _06075_, _05227_);
  and _14450_ (_06077_, _05542_, _05052_);
  nor _14451_ (_06078_, _06077_, _05273_);
  and _14452_ (_06079_, _06078_, _05059_);
  nor _14453_ (_06080_, _06079_, _06076_);
  nor _14454_ (_06081_, _06080_, _06074_);
  and _14455_ (_06082_, _06081_, _06073_);
  and _14456_ (_06083_, _06082_, _06068_);
  and _14457_ (_06084_, _06083_, _05561_);
  and _14458_ (_06086_, _06084_, _06060_);
  and _14459_ (_06087_, _06086_, _06056_);
  and _14460_ (_06088_, _06087_, _06055_);
  not _14461_ (_06089_, _05517_);
  not _14462_ (_06090_, _04984_);
  and _14463_ (_06091_, _04997_, _06090_);
  and _14464_ (_06092_, _04860_, _04885_);
  and _14465_ (_06093_, _06092_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  not _14466_ (_06094_, _06093_);
  nor _14467_ (_06095_, _06094_, _04947_);
  nand _14468_ (_06096_, _06095_, _06091_);
  nor _14469_ (_06097_, _06096_, _06089_);
  nand _14470_ (_06098_, _06097_, _06088_);
  not _14471_ (_06099_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  nor _14472_ (_06100_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff , _06099_);
  not _14473_ (_06101_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  not _14474_ (_06102_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  and _14475_ (_06103_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  not _14476_ (_06104_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and _14477_ (_06105_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _06104_);
  nor _14478_ (_06106_, _06105_, _06103_);
  nor _14479_ (_06107_, _06106_, _06102_);
  or _14480_ (_06108_, _06107_, _06101_);
  and _14481_ (_06109_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and _14482_ (_06110_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _06104_);
  nor _14483_ (_06112_, _06110_, _06109_);
  nor _14484_ (_06113_, _06112_, _06102_);
  and _14485_ (_06114_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and _14486_ (_06115_, _06104_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  or _14487_ (_06116_, _06115_, _06114_);
  not _14488_ (_06117_, _06116_);
  nand _14489_ (_06118_, _06117_, _06113_);
  or _14490_ (_06119_, _06118_, _06108_);
  and _14491_ (_06120_, _06119_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or _14492_ (_06121_, _06120_, _06100_);
  or _14493_ (_06122_, _06121_, _06097_);
  and _14494_ (_06123_, _06122_, _06098_);
  not _14495_ (_06124_, _05510_);
  nor _14496_ (_06125_, _06124_, _04947_);
  and _14497_ (_06126_, _06125_, _04990_);
  and _14498_ (_06127_, _06126_, _05517_);
  or _14499_ (_06128_, _06127_, _06123_);
  not _14500_ (_06129_, _06127_);
  or _14501_ (_06130_, _06129_, _05718_);
  and _14502_ (_06131_, _06130_, _04856_);
  and _14503_ (_08562_, _06131_, _06128_);
  and _14504_ (_06132_, _04932_, _04893_);
  not _14505_ (_06133_, _04904_);
  and _14506_ (_06134_, _06095_, _04922_);
  and _14507_ (_06135_, _06134_, _06133_);
  and _14508_ (_06136_, _06135_, _06132_);
  nand _14509_ (_06137_, _06136_, _04958_);
  and _14510_ (_06138_, _06137_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or _14511_ (_06139_, _06138_, _06127_);
  and _14512_ (_06140_, _04948_, _04922_);
  nor _14513_ (_06141_, _06094_, _04904_);
  and _14514_ (_06142_, _06141_, _06140_);
  and _14515_ (_06143_, _06142_, _06132_);
  nand _14516_ (_06144_, _06087_, _06055_);
  and _14517_ (_06145_, _04996_, _04958_);
  and _14518_ (_06146_, _06145_, _06090_);
  and _14519_ (_06147_, _06146_, _06144_);
  and _14520_ (_06148_, _04984_, _04958_);
  or _14521_ (_06149_, _04989_, _06148_);
  and _14522_ (_06150_, _06149_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or _14523_ (_06151_, _06150_, _06147_);
  and _14524_ (_06152_, _06151_, _06143_);
  or _14525_ (_06153_, _06152_, _06139_);
  nand _14526_ (_06154_, _06127_, _05287_);
  and _14527_ (_06155_, _06154_, _04856_);
  and _14528_ (_08584_, _06155_, _06153_);
  nand _14529_ (_06156_, _06107_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  and _14530_ (_06157_, _06116_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  or _14531_ (_06159_, _06157_, _06113_);
  or _14532_ (_06160_, _06159_, _06156_);
  nand _14533_ (_06161_, _06160_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  nand _14534_ (_06162_, _06161_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and _14535_ (_06163_, _05517_, _04987_);
  and _14536_ (_06164_, _06163_, _06093_);
  or _14537_ (_06165_, _06164_, _06162_);
  and _14538_ (_06166_, _06165_, _06129_);
  nand _14539_ (_06168_, _06164_, _06088_);
  and _14540_ (_06169_, _06168_, _06166_);
  nor _14541_ (_06170_, _06129_, _06032_);
  or _14542_ (_06171_, _06170_, _06169_);
  and _14543_ (_08683_, _06171_, _04856_);
  and _14544_ (_06172_, \oc8051_top_1.oc8051_memory_interface1.reti , \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  and _14545_ (_06173_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _06104_);
  and _14546_ (_06174_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _14547_ (_06175_, _06174_, _06173_);
  and _14548_ (_06176_, _06175_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  nor _14549_ (_06177_, _06176_, _06102_);
  and _14550_ (_06178_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and _14551_ (_06179_, _06178_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  not _14552_ (_06180_, _06179_);
  and _14553_ (_06181_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and _14554_ (_06182_, _06181_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and _14555_ (_06183_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and _14556_ (_06184_, _06183_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  nor _14557_ (_06185_, _06184_, _06182_);
  and _14558_ (_06186_, _06185_, _06180_);
  not _14559_ (_06187_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  nor _14560_ (_06188_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  nor _14561_ (_06189_, _06188_, _06187_);
  nand _14562_ (_06190_, _06189_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  not _14563_ (_06191_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  nor _14564_ (_06192_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  nor _14565_ (_06193_, _06192_, _06191_);
  and _14566_ (_06194_, _06193_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  not _14567_ (_06195_, _06194_);
  and _14568_ (_06196_, _06195_, _06190_);
  and _14569_ (_06197_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and _14570_ (_06198_, _06197_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  not _14571_ (_06199_, _06198_);
  and _14572_ (_06200_, _06199_, _06196_);
  and _14573_ (_06201_, _06200_, _06186_);
  nor _14574_ (_06202_, _06201_, _06177_);
  and _14575_ (_06203_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _06102_);
  not _14576_ (_06204_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and _14577_ (_06205_, _06178_, _06204_);
  not _14578_ (_06206_, _06205_);
  not _14579_ (_06207_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and _14580_ (_06208_, _06181_, _06207_);
  not _14581_ (_06209_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and _14582_ (_06210_, _06183_, _06209_);
  nor _14583_ (_06211_, _06210_, _06208_);
  and _14584_ (_06212_, _06211_, _06206_);
  not _14585_ (_06213_, _06212_);
  and _14586_ (_06214_, _06213_, _06203_);
  not _14587_ (_06215_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and _14588_ (_06216_, _06189_, _06215_);
  not _14589_ (_06217_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and _14590_ (_06218_, _06193_, _06217_);
  nor _14591_ (_06219_, _06218_, _06216_);
  not _14592_ (_06220_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and _14593_ (_06221_, _06197_, _06220_);
  not _14594_ (_06222_, _06221_);
  nand _14595_ (_06223_, _06222_, _06219_);
  and _14596_ (_06224_, _06223_, _06203_);
  or _14597_ (_06225_, _06224_, _06214_);
  nor _14598_ (_06226_, _06225_, _06202_);
  and _14599_ (_06227_, _06226_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  not _14600_ (_06228_, _06202_);
  nor _14601_ (_06229_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _06104_);
  and _14602_ (_06230_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _06104_);
  nor _14603_ (_06231_, _06230_, _06229_);
  nor _14604_ (_06232_, _06231_, _06228_);
  or _14605_ (_06233_, _06232_, _06227_);
  or _14606_ (_06234_, _06233_, _06172_);
  not _14607_ (_06235_, _06172_);
  or _14608_ (_06236_, _06231_, _06235_);
  and _14609_ (_06237_, _06236_, _04856_);
  and _14610_ (_09163_, _06237_, _06234_);
  and _14611_ (_06238_, _05731_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  and _14612_ (_06240_, _06238_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  not _14613_ (_06241_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _14614_ (_06242_, _06238_, _06241_);
  or _14615_ (_06243_, _06242_, _06240_);
  and _14616_ (_09192_, _06243_, _04856_);
  nand _14617_ (_06244_, _06228_, _06214_);
  or _14618_ (_06245_, _06186_, _06177_);
  and _14619_ (_06246_, _06245_, _06235_);
  and _14620_ (_06248_, _06246_, _06244_);
  nor _14621_ (_06249_, _06172_, _06104_);
  nor _14622_ (_06250_, _06235_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  nor _14623_ (_06251_, _06250_, _06249_);
  or _14624_ (_06252_, _06251_, _06248_);
  or _14625_ (_06253_, _06224_, _06202_);
  not _14626_ (_06254_, _06200_);
  or _14627_ (_06255_, _06245_, _06254_);
  and _14628_ (_06256_, _06255_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and _14629_ (_06257_, _06256_, _06253_);
  or _14630_ (_06258_, _06257_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  and _14631_ (_06259_, _06258_, _04856_);
  and _14632_ (_09318_, _06259_, _06252_);
  and _14633_ (_06260_, _06238_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  not _14634_ (_06261_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor _14635_ (_06262_, _06238_, _06261_);
  or _14636_ (_06263_, _06262_, _06260_);
  and _14637_ (_09528_, _06263_, _04856_);
  nand _14638_ (_06264_, _06201_, _06102_);
  or _14639_ (_06265_, _06264_, _06225_);
  nand _14640_ (_06266_, _06229_, _06172_);
  and _14641_ (_06267_, _06266_, _04856_);
  and _14642_ (_10162_, _06267_, _06265_);
  and _14643_ (_06268_, _05519_, _06090_);
  and _14644_ (_06269_, _04933_, _04893_);
  and _14645_ (_06270_, _06269_, _06142_);
  and _14646_ (_06271_, _06270_, _06268_);
  or _14647_ (_06272_, _06271_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and _14648_ (_06273_, _04933_, _04922_);
  and _14649_ (_06274_, _06273_, _05515_);
  and _14650_ (_06275_, _06274_, _06126_);
  not _14651_ (_06276_, _06275_);
  and _14652_ (_06277_, _06276_, _06272_);
  nand _14653_ (_06278_, _06271_, _06088_);
  and _14654_ (_06279_, _06278_, _06277_);
  nor _14655_ (_06280_, _05338_, _05282_);
  not _14656_ (_06281_, _06280_);
  and _14657_ (_06282_, _06281_, _05556_);
  and _14658_ (_06283_, _06282_, _05551_);
  and _14659_ (_06284_, _06283_, _05538_);
  nor _14660_ (_06285_, _06284_, _06276_);
  or _14661_ (_06286_, _06285_, _06279_);
  and _14662_ (_10217_, _06286_, _04856_);
  not _14663_ (_06287_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  nor _14664_ (_06288_, _06172_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _14665_ (_06289_, _06288_, _06287_);
  or _14666_ (_06290_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], _06104_);
  or _14667_ (_06291_, _06253_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  and _14668_ (_06292_, _06291_, _06290_);
  and _14669_ (_06293_, _06292_, _06248_);
  or _14670_ (_06294_, _06293_, _06289_);
  and _14671_ (_10318_, _06294_, _04856_);
  nor _14672_ (_06295_, _04947_, _04922_);
  and _14673_ (_06296_, _06295_, _06141_);
  and _14674_ (_06297_, _06296_, _06269_);
  and _14675_ (_06298_, _06297_, _06268_);
  nand _14676_ (_06299_, _06298_, _06088_);
  or _14677_ (_06300_, _06298_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and _14678_ (_06301_, _06268_, _05512_);
  nor _14679_ (_06302_, _04932_, _04922_);
  and _14680_ (_06303_, _06302_, _05515_);
  and _14681_ (_06304_, _06303_, _06301_);
  not _14682_ (_06305_, _06304_);
  and _14683_ (_06306_, _06305_, _06300_);
  and _14684_ (_06307_, _06306_, _06299_);
  nor _14685_ (_06308_, _06305_, _06284_);
  or _14686_ (_06309_, _06308_, _06307_);
  and _14687_ (_10339_, _06309_, _04856_);
  and _14688_ (_06310_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _04856_);
  and _14689_ (_10459_, _06310_, _06172_);
  and _14690_ (_06311_, _06268_, _06095_);
  and _14691_ (_06312_, _06311_, _05517_);
  nand _14692_ (_06313_, _06312_, _06088_);
  nor _14693_ (_06314_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  nor _14694_ (_06316_, _06314_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf );
  nand _14695_ (_06317_, _06157_, _06112_);
  or _14696_ (_06318_, _06317_, _06108_);
  and _14697_ (_06319_, _06318_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or _14698_ (_06320_, _06319_, _06316_);
  or _14699_ (_06321_, _06320_, _06312_);
  and _14700_ (_06322_, _06321_, _06129_);
  and _14701_ (_06323_, _06322_, _06313_);
  nor _14702_ (_06324_, _06284_, _06129_);
  or _14703_ (_06325_, _06324_, _06323_);
  and _14704_ (_10480_, _06325_, _04856_);
  and _14705_ (_10675_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _04856_);
  and _14706_ (_06326_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  or _14707_ (_06327_, _06156_, _06118_);
  and _14708_ (_06328_, _06327_, _06326_);
  and _14709_ (_06329_, _05520_, _04948_);
  and _14710_ (_06330_, _06329_, _05517_);
  and _14711_ (_06331_, _06330_, _06093_);
  or _14712_ (_06332_, _06331_, _06328_);
  and _14713_ (_06333_, _06332_, _06129_);
  nand _14714_ (_06334_, _06331_, _06088_);
  and _14715_ (_06335_, _06334_, _06333_);
  nor _14716_ (_06336_, _06129_, _05669_);
  or _14717_ (_06337_, _06336_, _06335_);
  and _14718_ (_10816_, _06337_, _04856_);
  and _14719_ (_06338_, \oc8051_top_1.oc8051_sfr1.prescaler [0], \oc8051_top_1.oc8051_sfr1.prescaler [1]);
  or _14720_ (_06339_, \oc8051_top_1.oc8051_sfr1.prescaler [0], \oc8051_top_1.oc8051_sfr1.prescaler [1]);
  nand _14721_ (_06340_, _06339_, _04856_);
  nor _14722_ (_11292_, _06340_, _06338_);
  nor _14723_ (_11844_, \oc8051_top_1.oc8051_sfr1.prescaler [0], rst);
  or _14724_ (_06341_, _06238_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  not _14725_ (_06342_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nand _14726_ (_06343_, _06238_, _06342_);
  and _14727_ (_06344_, _06343_, _04856_);
  and _14728_ (_12295_, _06344_, _06341_);
  not _14729_ (_06345_, \oc8051_top_1.oc8051_sfr1.prescaler [2]);
  and _14730_ (_06346_, _06338_, _06345_);
  and _14731_ (_06347_, _06346_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  nor _14732_ (_06348_, _06338_, _06345_);
  or _14733_ (_06349_, _06348_, _06346_);
  nand _14734_ (_06350_, _06349_, _04856_);
  nor _14735_ (_12580_, _06350_, _06347_);
  or _14736_ (_06351_, _04992_, _05003_);
  and _14737_ (_06352_, _06351_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  and _14738_ (_06353_, _06352_, _04861_);
  or _14739_ (_06354_, _05007_, _04995_);
  and _14740_ (_06355_, _06354_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  or _14741_ (_06356_, _05385_, _06019_);
  and _14742_ (_06357_, _06356_, _05256_);
  or _14743_ (_06358_, _06357_, _05396_);
  nand _14744_ (_06359_, _05385_, _05267_);
  or _14745_ (_06360_, _06075_, _05206_);
  and _14746_ (_06361_, _06360_, _06359_);
  or _14747_ (_06362_, _05383_, _05232_);
  not _14748_ (_06363_, _05223_);
  or _14749_ (_06364_, _06363_, _05206_);
  and _14750_ (_06365_, _06364_, _06362_);
  or _14751_ (_06366_, _05282_, _05126_);
  and _14752_ (_06367_, _06366_, _06365_);
  and _14753_ (_06368_, _06367_, _06361_);
  and _14754_ (_06369_, _06368_, _06358_);
  nor _14755_ (_06370_, _06369_, _05673_);
  and _14756_ (_06371_, _06370_, _04988_);
  or _14757_ (_06372_, _06371_, _06355_);
  or _14758_ (_06373_, _06372_, _06353_);
  and _14759_ (_13213_, _06373_, _04856_);
  and _14760_ (_06374_, _06354_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  and _14761_ (_06375_, _05718_, _04988_);
  and _14762_ (_06376_, _06351_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  or _14763_ (_06377_, _06376_, _06375_);
  and _14764_ (_06378_, _06377_, _04861_);
  or _14765_ (_06379_, _06378_, _06374_);
  and _14766_ (_01164_, _06379_, _04856_);
  and _14767_ (_06380_, _06038_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  and _14768_ (_06381_, _06370_, _04992_);
  and _14769_ (_06382_, _04861_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  and _14770_ (_06383_, _06382_, _06039_);
  or _14771_ (_06384_, _06383_, _06381_);
  or _14772_ (_06385_, _06384_, _06380_);
  and _14773_ (_01432_, _06385_, _04856_);
  nand _14774_ (_06386_, _05721_, _05008_);
  and _14775_ (_06387_, _06386_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  nor _14776_ (_06388_, _05282_, _05081_);
  not _14777_ (_06389_, _06388_);
  not _14778_ (_06390_, _05693_);
  nand _14779_ (_06391_, _05175_, _05059_);
  nand _14780_ (_06392_, _06391_, _06390_);
  nand _14781_ (_06393_, _06392_, _05565_);
  or _14782_ (_06395_, _06392_, _05565_);
  and _14783_ (_06396_, _06395_, _05223_);
  nand _14784_ (_06397_, _06396_, _06393_);
  nand _14785_ (_06398_, _05349_, _05259_);
  and _14786_ (_06399_, _05347_, _05267_);
  and _14787_ (_06400_, _05269_, _05081_);
  nor _14788_ (_06401_, _06400_, _06399_);
  and _14789_ (_06402_, _05346_, _05059_);
  nor _14790_ (_06403_, _06402_, _05232_);
  and _14791_ (_06404_, _06403_, _05692_);
  nor _14792_ (_06405_, _05348_, _05256_);
  nor _14793_ (_06406_, _06405_, _06404_);
  and _14794_ (_06407_, _06406_, _06401_);
  and _14795_ (_06408_, _06407_, _06398_);
  and _14796_ (_06409_, _06408_, _06397_);
  nand _14797_ (_06410_, _06409_, _06389_);
  and _14798_ (_06411_, _06410_, _06043_);
  or _14799_ (_06412_, _06411_, _06387_);
  and _14800_ (_01517_, _06412_, _04856_);
  and _14801_ (_06413_, _06354_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  and _14802_ (_06414_, _06410_, _04988_);
  and _14803_ (_06415_, _06351_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  or _14804_ (_06416_, _06415_, _06414_);
  and _14805_ (_06417_, _06416_, _04861_);
  or _14806_ (_06418_, _06417_, _06413_);
  and _14807_ (_01547_, _06418_, _04856_);
  and _14808_ (_06419_, _05719_, _05670_);
  and _14809_ (_06420_, _05723_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  or _14810_ (_06421_, _06420_, _06419_);
  and _14811_ (_01669_, _06421_, _04856_);
  and _14812_ (_06422_, _06041_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  and _14813_ (_06423_, _06043_, _05670_);
  or _14814_ (_06424_, _06423_, _06422_);
  and _14815_ (_01710_, _06424_, _04856_);
  and _14816_ (_06425_, _06041_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  and _14817_ (_06426_, _06043_, _05288_);
  or _14818_ (_06427_, _06426_, _06425_);
  and _14819_ (_01955_, _06427_, _04856_);
  nand _14820_ (_06428_, _05452_, _05303_);
  and _14821_ (_06429_, _06428_, _05453_);
  nand _14822_ (_06430_, _06429_, _05455_);
  and _14823_ (_06431_, _05483_, _05243_);
  not _14824_ (_06432_, _06431_);
  nor _14825_ (_06433_, _05483_, _05243_);
  nor _14826_ (_06434_, _06433_, _06363_);
  and _14827_ (_06435_, _06434_, _06432_);
  nor _14828_ (_06436_, _05531_, _05460_);
  nor _14829_ (_06437_, _06436_, _05232_);
  not _14830_ (_06438_, _06437_);
  nor _14831_ (_06439_, _05490_, _05172_);
  not _14832_ (_06440_, _06439_);
  nor _14833_ (_06441_, _05274_, _05243_);
  and _14834_ (_06442_, _05497_, ABINPUT001[15]);
  and _14835_ (_06443_, _05499_, ABINPUT000[15]);
  nor _14836_ (_06444_, _06443_, _06442_);
  not _14837_ (_06445_, _06444_);
  nor _14838_ (_06446_, _06445_, _06441_);
  and _14839_ (_06448_, _06446_, _06440_);
  and _14840_ (_06449_, _06448_, _06438_);
  not _14841_ (_06450_, _06449_);
  nor _14842_ (_06451_, _06450_, _06435_);
  nand _14843_ (_06452_, _06451_, _06430_);
  or _14844_ (_06453_, _06452_, _05293_);
  not _14845_ (_06454_, _05455_);
  and _14846_ (_06455_, _05428_, _05422_);
  nor _14847_ (_06456_, _06455_, _06454_);
  and _14848_ (_06457_, _06456_, _05429_);
  not _14849_ (_06458_, _06457_);
  nor _14850_ (_06459_, _05629_, _05597_);
  nor _14851_ (_06460_, _06459_, _05630_);
  nor _14852_ (_06461_, _06460_, _05584_);
  and _14853_ (_06462_, _05568_, _05199_);
  nor _14854_ (_06463_, _06462_, _05048_);
  nor _14855_ (_06464_, _06463_, _05569_);
  nor _14856_ (_06466_, _06464_, _05558_);
  not _14857_ (_06468_, _05279_);
  or _14858_ (_06469_, _05338_, _06468_);
  and _14859_ (_06470_, _05499_, ABINPUT000[7]);
  not _14860_ (_06471_, _06470_);
  and _14861_ (_06473_, _06471_, _06469_);
  and _14862_ (_06474_, _05280_, _05587_);
  nor _14863_ (_06475_, _05274_, _05048_);
  and _14864_ (_06476_, _05497_, ABINPUT001[7]);
  or _14865_ (_06477_, _06476_, _06475_);
  nor _14866_ (_06478_, _06477_, _06474_);
  and _14867_ (_06479_, _06478_, _05271_);
  and _14868_ (_06480_, _06479_, _06473_);
  and _14869_ (_06481_, _06480_, _05263_);
  not _14870_ (_06482_, _06481_);
  nor _14871_ (_06483_, _06482_, _06466_);
  and _14872_ (_06485_, _06483_, _05247_);
  not _14873_ (_06486_, _06485_);
  nor _14874_ (_06487_, _06486_, _06461_);
  and _14875_ (_06488_, _06487_, _06458_);
  nor _14876_ (_06489_, _06488_, _05643_);
  and _14877_ (_06490_, _05643_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or _14878_ (_06491_, _06490_, _05292_);
  or _14879_ (_06492_, _06491_, _06489_);
  and _14880_ (_06493_, _06492_, _04856_);
  and _14881_ (_02380_, _06493_, _06453_);
  and _14882_ (_06494_, _06145_, _04984_);
  and _14883_ (_06495_, _06494_, _05512_);
  and _14884_ (_06496_, _06495_, _05517_);
  nor _14885_ (_06497_, _06496_, _05292_);
  not _14886_ (_06498_, _06497_);
  nand _14887_ (_06499_, _06498_, _06488_);
  or _14888_ (_06500_, _06498_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and _14889_ (_06501_, _06500_, _04856_);
  and _14890_ (_02512_, _06501_, _06499_);
  nor _14891_ (_06502_, _05401_, _05399_);
  not _14892_ (_06503_, _06502_);
  nor _14893_ (_06504_, _05402_, _06454_);
  and _14894_ (_06505_, _06504_, _06503_);
  not _14895_ (_06506_, _06505_);
  nor _14896_ (_06507_, _05619_, _05614_);
  nor _14897_ (_06508_, _06507_, _05620_);
  nor _14898_ (_06509_, _06508_, _05584_);
  not _14899_ (_06510_, _06509_);
  and _14900_ (_06511_, _05173_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor _14901_ (_06512_, _05559_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor _14902_ (_06513_, _06512_, _05207_);
  nor _14903_ (_06514_, _06513_, _05172_);
  nor _14904_ (_06515_, _06514_, _06511_);
  nor _14905_ (_06516_, _06515_, _05558_);
  nor _14906_ (_06517_, _05371_, _05256_);
  and _14907_ (_06518_, _05372_, _05259_);
  or _14908_ (_06519_, _06518_, _06517_);
  not _14909_ (_06520_, _06519_);
  and _14910_ (_06521_, _05280_, _05207_);
  and _14911_ (_06522_, _05497_, ABINPUT001[3]);
  and _14912_ (_06523_, _05499_, ABINPUT000[3]);
  nor _14913_ (_06524_, _06523_, _06522_);
  not _14914_ (_06525_, _06524_);
  nor _14915_ (_06526_, _06525_, _06521_);
  or _14916_ (_06527_, _06468_, _05103_);
  nor _14917_ (_06528_, _05274_, _05172_);
  not _14918_ (_06529_, _06528_);
  and _14919_ (_06530_, _06529_, _06527_);
  and _14920_ (_06531_, _06530_, _06526_);
  and _14921_ (_06532_, _06531_, _06520_);
  not _14922_ (_06533_, _06532_);
  nor _14923_ (_06534_, _06533_, _06516_);
  not _14924_ (_06535_, _06534_);
  or _14925_ (_06536_, _06012_, _05206_);
  or _14926_ (_06537_, _06013_, _05126_);
  nand _14927_ (_06538_, _06537_, _06536_);
  or _14928_ (_06539_, _06538_, _05172_);
  nand _14929_ (_06540_, _06538_, _05172_);
  and _14930_ (_06541_, _06540_, _05223_);
  and _14931_ (_06542_, _06541_, _06539_);
  nor _14932_ (_06543_, _05368_, _05232_);
  or _14933_ (_06544_, _06543_, _06542_);
  not _14934_ (_06545_, _06544_);
  and _14935_ (_06546_, _05369_, _05267_);
  and _14936_ (_06547_, _05269_, _05172_);
  nor _14937_ (_06548_, _06547_, _06546_);
  nand _14938_ (_06549_, _06548_, _06545_);
  nor _14939_ (_06550_, _06549_, _06535_);
  and _14940_ (_06551_, _06550_, _06510_);
  and _14941_ (_06552_, _06551_, _06506_);
  nand _14942_ (_06553_, _06552_, _06498_);
  or _14943_ (_06554_, _06498_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and _14944_ (_06555_, _06554_, _04856_);
  and _14945_ (_02954_, _06555_, _06553_);
  nor _14946_ (_06556_, _05402_, _05395_);
  or _14947_ (_06557_, _06556_, _06454_);
  nor _14948_ (_06558_, _06557_, _05403_);
  not _14949_ (_06559_, _06558_);
  nor _14950_ (_06560_, _05620_, _05612_);
  nor _14951_ (_06561_, _06560_, _05621_);
  nor _14952_ (_06562_, _06561_, _05584_);
  not _14953_ (_06563_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor _14954_ (_06564_, _05173_, _06563_);
  nor _14955_ (_06565_, _06564_, _05204_);
  or _14956_ (_06566_, _06565_, _05558_);
  nor _14957_ (_06567_, _06566_, _05559_);
  and _14958_ (_06568_, _05280_, _05205_);
  and _14959_ (_06569_, _05497_, ABINPUT001[4]);
  and _14960_ (_06570_, _05499_, ABINPUT000[4]);
  nor _14961_ (_06571_, _06570_, _06569_);
  not _14962_ (_06572_, _06571_);
  nor _14963_ (_06573_, _06572_, _06568_);
  nor _14964_ (_06574_, _05274_, _05103_);
  not _14965_ (_06575_, _06574_);
  or _14966_ (_06576_, _06468_, _05081_);
  and _14967_ (_06578_, _06576_, _06575_);
  and _14968_ (_06579_, _06578_, _06573_);
  not _14969_ (_06580_, _06579_);
  nor _14970_ (_06581_, _06580_, _06567_);
  and _14971_ (_06582_, _06581_, _05667_);
  and _14972_ (_06583_, _06582_, _05656_);
  not _14973_ (_06584_, _06583_);
  nor _14974_ (_06585_, _06584_, _06562_);
  and _14975_ (_06586_, _06585_, _06559_);
  nand _14976_ (_06587_, _06586_, _06498_);
  not _14977_ (_06588_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  nand _14978_ (_06589_, _06497_, _06588_);
  and _14979_ (_06590_, _06589_, _04856_);
  and _14980_ (_03036_, _06590_, _06587_);
  and _14981_ (_06591_, _05683_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  and _14982_ (_06592_, _05671_, _05288_);
  or _14983_ (_06593_, _06592_, _06591_);
  and _14984_ (_03190_, _06593_, _04856_);
  and _14985_ (_06594_, _05985_, _05874_);
  and _14986_ (_06595_, _06594_, _05849_);
  and _14987_ (_06596_, _05968_, _05923_);
  and _14988_ (_06597_, _06596_, _05972_);
  and _14989_ (_06598_, _05848_, _05772_);
  and _14990_ (_06599_, _06598_, _06597_);
  and _14991_ (_06600_, _06597_, _05849_);
  or _14992_ (_06601_, _06600_, _06599_);
  nor _14993_ (_06602_, _06601_, _06595_);
  and _14994_ (_06603_, _05985_, _05983_);
  nor _14995_ (_06604_, _06603_, _05951_);
  nand _14996_ (_06605_, _06604_, _06602_);
  and _14997_ (_06606_, _05997_, _05953_);
  and _14998_ (_06607_, _06606_, _05969_);
  and _14999_ (_06608_, _05949_, _05972_);
  and _15000_ (_06609_, _06606_, _06608_);
  and _15001_ (_06610_, _06594_, _06606_);
  or _15002_ (_06611_, _06610_, _06609_);
  and _15003_ (_06612_, _05978_, _05874_);
  and _15004_ (_06613_, _06612_, _05849_);
  and _15005_ (_06614_, _05986_, _05849_);
  nor _15006_ (_06615_, _06614_, _06613_);
  not _15007_ (_06616_, _06615_);
  or _15008_ (_06617_, _06616_, _06611_);
  or _15009_ (_06618_, _06617_, _06607_);
  and _15010_ (_06619_, _05984_, _05923_);
  and _15011_ (_06620_, _06619_, _05972_);
  and _15012_ (_06621_, _06598_, _06620_);
  and _15013_ (_06622_, _06620_, _05849_);
  or _15014_ (_06623_, _06622_, _06621_);
  and _15015_ (_06624_, _06000_, _05874_);
  and _15016_ (_06625_, _06624_, _05849_);
  and _15017_ (_06626_, _06606_, _06001_);
  or _15018_ (_06627_, _06626_, _06625_);
  and _15019_ (_06628_, _06606_, _05986_);
  and _15020_ (_06629_, _06606_, _05950_);
  or _15021_ (_06630_, _06629_, _06628_);
  or _15022_ (_06631_, _06630_, _06627_);
  or _15023_ (_06632_, _06631_, _06623_);
  or _15024_ (_06633_, _06632_, _06618_);
  or _15025_ (_06634_, _06633_, _06605_);
  and _15026_ (_06635_, _06619_, _05874_);
  and _15027_ (_06636_, _06635_, _05848_);
  not _15028_ (_06637_, _05822_);
  or _15029_ (_06638_, _05964_, _06637_);
  and _15030_ (_06639_, _06638_, _06001_);
  or _15031_ (_06641_, _06639_, _06636_);
  or _15032_ (_06642_, _06641_, _05955_);
  or _15033_ (_06643_, _06642_, _06634_);
  and _15034_ (_06644_, _06643_, _05730_);
  and _15035_ (_06645_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _15036_ (_06646_, _06005_, _05960_);
  not _15037_ (_06647_, _05959_);
  nand _15038_ (_06648_, _05983_, _05950_);
  nor _15039_ (_06649_, _06648_, _06647_);
  or _15040_ (_06650_, _06649_, _06646_);
  or _15041_ (_06651_, _06650_, _06645_);
  or _15042_ (_06652_, _06651_, _06644_);
  and _15043_ (_03594_, _06652_, _04856_);
  not _15044_ (_06653_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and _15045_ (_06654_, _05291_, _06653_);
  and _15046_ (_06655_, _06654_, _05507_);
  not _15047_ (_06656_, _06654_);
  and _15048_ (_06657_, _06268_, _06144_);
  nor _15049_ (_06658_, _06268_, _05332_);
  or _15050_ (_06659_, _06658_, _06657_);
  nor _15051_ (_06660_, _06653_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1]);
  and _15052_ (_06661_, _06660_, _04859_);
  nor _15053_ (_06662_, _04904_, _04893_);
  and _15054_ (_06663_, _06662_, _06273_);
  and _15055_ (_06664_, _06663_, _05001_);
  and _15056_ (_06665_, _06664_, _05510_);
  nor _15057_ (_06666_, _06665_, _06661_);
  and _15058_ (_06667_, _06666_, _06656_);
  nor _15059_ (_06668_, _04948_, _04904_);
  and _15060_ (_06669_, _06668_, _04922_);
  nor _15061_ (_06670_, _04932_, _04893_);
  and _15062_ (_06671_, _06670_, _06093_);
  and _15063_ (_06672_, _06671_, _06669_);
  and _15064_ (_06673_, _06672_, _06667_);
  nand _15065_ (_06674_, _06673_, _06659_);
  not _15066_ (_06675_, _06666_);
  and _15067_ (_06676_, _06675_, _05641_);
  not _15068_ (_06677_, _06672_);
  and _15069_ (_06678_, _06677_, _06667_);
  and _15070_ (_06679_, _06678_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor _15071_ (_06680_, _06679_, _06676_);
  nand _15072_ (_06681_, _06680_, _06674_);
  and _15073_ (_06682_, _06681_, _06656_);
  or _15074_ (_06684_, _06682_, _06655_);
  and _15075_ (_04014_, _06684_, _04856_);
  not _15076_ (_06685_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  and _15077_ (_06686_, _05679_, _04861_);
  nor _15078_ (_06687_, _06686_, _06685_);
  not _15079_ (_06688_, _06686_);
  nor _15080_ (_06689_, _06688_, _05287_);
  or _15081_ (_06690_, _06689_, _06687_);
  and _15082_ (_04065_, _06690_, _04856_);
  or _15083_ (_06691_, _06497_, _05641_);
  or _15084_ (_06692_, _06498_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and _15085_ (_06693_, _06692_, _04856_);
  and _15086_ (_04848_, _06693_, _06691_);
  and _15087_ (_06694_, _06033_, _05671_);
  and _15088_ (_06695_, _04995_, _04861_);
  or _15089_ (_06696_, _06695_, _05682_);
  and _15090_ (_06697_, _06696_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  or _15091_ (_06698_, _06697_, _06694_);
  and _15092_ (_04849_, _06698_, _04856_);
  or _15093_ (_06699_, _06238_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nand _15094_ (_06700_, _06238_, _05185_);
  and _15095_ (_06701_, _06700_, _04856_);
  and _15096_ (_04851_, _06701_, _06699_);
  and _15097_ (_06702_, _06386_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  nor _15098_ (_06703_, _05282_, _05172_);
  or _15099_ (_06704_, _06703_, _06519_);
  or _15100_ (_06705_, _06704_, _06549_);
  and _15101_ (_06706_, _06705_, _06043_);
  or _15102_ (_06707_, _06706_, _06702_);
  and _15103_ (_04853_, _06707_, _04856_);
  not _15104_ (_06708_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  nor _15105_ (_06709_, _05675_, _06708_);
  and _15106_ (_06710_, _06705_, _05675_);
  or _15107_ (_06711_, _06710_, _06709_);
  or _15108_ (_06712_, _06711_, _05673_);
  or _15109_ (_06713_, _04861_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  and _15110_ (_06714_, _06713_, _04856_);
  and _15111_ (_04854_, _06714_, _06712_);
  and _15112_ (_06715_, _05723_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  and _15113_ (_06716_, _06705_, _05719_);
  or _15114_ (_06717_, _06716_, _06715_);
  and _15115_ (_04855_, _06717_, _04856_);
  and _15116_ (_06718_, _06033_, _05719_);
  and _15117_ (_06719_, _05723_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  or _15118_ (_06720_, _06719_, _06718_);
  and _15119_ (_04970_, _06720_, _04856_);
  and _15120_ (_06721_, _04856_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and _15121_ (_06722_, _06721_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and _15122_ (_06723_, _05998_, _06608_);
  or _15123_ (_06724_, _06723_, _06611_);
  and _15124_ (_06725_, _05998_, _05950_);
  or _15125_ (_06726_, _06725_, _06629_);
  or _15126_ (_06727_, _06726_, _06724_);
  nand _15127_ (_06728_, _06612_, _05983_);
  not _15128_ (_06729_, _06728_);
  or _15129_ (_06730_, _05847_, _06637_);
  nor _15130_ (_06731_, _06730_, _05797_);
  and _15131_ (_06732_, _06620_, _06731_);
  and _15132_ (_06733_, _06732_, _05772_);
  or _15133_ (_06734_, _06733_, _06729_);
  and _15134_ (_06735_, _06732_, _05773_);
  and _15135_ (_06736_, _06620_, _05848_);
  and _15136_ (_06737_, _05969_, _05923_);
  and _15137_ (_06738_, _06737_, _05849_);
  or _15138_ (_06739_, _06738_, _06736_);
  or _15139_ (_06740_, _06739_, _06735_);
  or _15140_ (_06741_, _06740_, _06734_);
  or _15141_ (_06742_, _06741_, _06727_);
  nor _15142_ (_06743_, _05822_, _05874_);
  and _15143_ (_06744_, _06743_, _05949_);
  or _15144_ (_06745_, _06594_, _05950_);
  and _15145_ (_06746_, _06745_, _06637_);
  or _15146_ (_06747_, _06746_, _06744_);
  nor _15147_ (_06748_, _06601_, _05966_);
  not _15148_ (_06749_, _06748_);
  and _15149_ (_06750_, _06743_, _06596_);
  and _15150_ (_06751_, _06598_, _05948_);
  or _15151_ (_06752_, _06751_, _06750_);
  or _15152_ (_06753_, _06752_, _06749_);
  or _15153_ (_06754_, _06753_, _06747_);
  and _15154_ (_06755_, _06597_, _05965_);
  and _15155_ (_06756_, _06620_, _05965_);
  or _15156_ (_06757_, _06756_, _06755_);
  or _15157_ (_06758_, _06757_, _05988_);
  and _15158_ (_06759_, _05998_, _05986_);
  or _15159_ (_06760_, _06759_, _06628_);
  and _15160_ (_06761_, _06597_, _06731_);
  and _15161_ (_06762_, _05983_, _05996_);
  and _15162_ (_06763_, _06743_, _05984_);
  or _15163_ (_06764_, _06763_, _06762_);
  or _15164_ (_06765_, _06764_, _06761_);
  or _15165_ (_06766_, _06765_, _06760_);
  or _15166_ (_06767_, _06766_, _06758_);
  or _15167_ (_06768_, _06767_, _06754_);
  or _15168_ (_06769_, _06768_, _06742_);
  and _15169_ (_06770_, _05730_, _04856_);
  and _15170_ (_06771_, _06770_, _06769_);
  or _15171_ (_05113_, _06771_, _06722_);
  and _15172_ (_06772_, _05968_, _05976_);
  and _15173_ (_06773_, _06772_, _05874_);
  nand _15174_ (_06774_, _06773_, _05848_);
  nand _15175_ (_06775_, _06773_, _05983_);
  and _15176_ (_06776_, _06775_, _06774_);
  and _15177_ (_06777_, _06772_, _05972_);
  and _15178_ (_06778_, _06777_, _05983_);
  and _15179_ (_06779_, _06777_, _05848_);
  nor _15180_ (_06780_, _06779_, _06778_);
  and _15181_ (_06781_, _06780_, _06776_);
  not _15182_ (_06782_, _06770_);
  and _15183_ (_06783_, _06598_, _06000_);
  or _15184_ (_06784_, _06783_, _06782_);
  or _15185_ (_05116_, _06784_, _06781_);
  and _15186_ (_06786_, _06598_, _05996_);
  and _15187_ (_06787_, _06624_, _05983_);
  or _15188_ (_06788_, _06787_, _06786_);
  and _15189_ (_06789_, _06763_, _05976_);
  or _15190_ (_06790_, _06789_, _05988_);
  or _15191_ (_06791_, _06790_, _06760_);
  or _15192_ (_06792_, _06791_, _06788_);
  and _15193_ (_06793_, _06792_, _05730_);
  and _15194_ (_06794_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _15195_ (_06795_, _06794_, _06005_);
  or _15196_ (_06796_, _06795_, _06793_);
  and _15197_ (_05127_, _06796_, _04856_);
  and _15198_ (_06797_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  not _15199_ (_06798_, _06797_);
  not _15200_ (_06799_, _05962_);
  or _15201_ (_06800_, _06737_, _06624_);
  and _15202_ (_06801_, _06800_, _06598_);
  nor _15203_ (_06802_, _06801_, _06786_);
  and _15204_ (_06803_, _06802_, _06003_);
  nor _15205_ (_06804_, _06803_, _06799_);
  not _15206_ (_06805_, _06804_);
  and _15207_ (_06806_, _05983_, _06596_);
  and _15208_ (_06807_, _06806_, _05959_);
  and _15209_ (_06808_, _06619_, _05983_);
  and _15210_ (_06809_, _06808_, _05959_);
  nor _15211_ (_06810_, _06809_, _06807_);
  not _15212_ (_06811_, _06810_);
  not _15213_ (_06812_, _05729_);
  nor _15214_ (_06813_, _06003_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and _15215_ (_06814_, _06813_, _06812_);
  nor _15216_ (_06815_, _06814_, _06811_);
  nand _15217_ (_06816_, _06815_, _06805_);
  nand _15218_ (_06817_, _06816_, _04859_);
  and _15219_ (_06818_, _06817_, _06798_);
  not _15220_ (_06819_, _06818_);
  and _15221_ (_06820_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  not _15222_ (_06821_, _06820_);
  and _15223_ (_06822_, _05948_, _05899_);
  and _15224_ (_06823_, _06822_, _05849_);
  not _15225_ (_06824_, _06823_);
  nand _15226_ (_06825_, _06001_, _05965_);
  and _15227_ (_06826_, _06825_, _06824_);
  nand _15228_ (_06827_, _06594_, _05983_);
  nand _15229_ (_06828_, _06777_, _05965_);
  and _15230_ (_06829_, _06828_, _06827_);
  and _15231_ (_06830_, _06829_, _06826_);
  and _15232_ (_06831_, _05965_, _05874_);
  and _15233_ (_06832_, _06619_, _06831_);
  and _15234_ (_06833_, _06822_, _05965_);
  or _15235_ (_06834_, _06833_, _06832_);
  and _15236_ (_06835_, _06000_, _06831_);
  and _15237_ (_06836_, _06612_, _05965_);
  nor _15238_ (_06837_, _06836_, _05966_);
  not _15239_ (_06838_, _06837_);
  or _15240_ (_06839_, _06838_, _06835_);
  nor _15241_ (_06840_, _06839_, _06834_);
  and _15242_ (_06841_, _06840_, _06830_);
  not _15243_ (_06842_, _06802_);
  nor _15244_ (_06843_, _06842_, _06758_);
  nand _15245_ (_06844_, _06843_, _06841_);
  nand _15246_ (_06845_, _06844_, _05962_);
  and _15247_ (_06846_, _05994_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and _15248_ (_06847_, _06823_, _06846_);
  nor _15249_ (_06848_, _06847_, _06807_);
  nand _15250_ (_06849_, _06848_, _06845_);
  nand _15251_ (_06850_, _06849_, _04859_);
  nand _15252_ (_06851_, _06850_, _06821_);
  and _15253_ (_06852_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  not _15254_ (_06853_, _06852_);
  and _15255_ (_06854_, _06822_, _05972_);
  nand _15256_ (_06855_, _06854_, _05983_);
  not _15257_ (_06856_, _06855_);
  and _15258_ (_06857_, _06822_, _05874_);
  nand _15259_ (_06858_, _06857_, _05983_);
  nand _15260_ (_06859_, _06858_, _06648_);
  nor _15261_ (_06860_, _06859_, _06856_);
  and _15262_ (_06861_, _06612_, _06606_);
  and _15263_ (_06862_, _06624_, _06606_);
  nor _15264_ (_06863_, _06862_, _06861_);
  and _15265_ (_06864_, _06863_, _06860_);
  and _15266_ (_06865_, _06001_, _05849_);
  or _15267_ (_06866_, _06865_, _06636_);
  nand _15268_ (_06867_, _06635_, _06606_);
  nand _15269_ (_06868_, _06822_, _06606_);
  nand _15270_ (_06869_, _06868_, _06867_);
  nor _15271_ (_06870_, _06869_, _06866_);
  and _15272_ (_06871_, _06777_, _06606_);
  and _15273_ (_06872_, _05996_, _05849_);
  nor _15274_ (_06873_, _06872_, _06871_);
  and _15275_ (_06875_, _06873_, _06870_);
  and _15276_ (_06876_, _06875_, _06864_);
  nor _15277_ (_06877_, _06609_, _05979_);
  or _15278_ (_06878_, _06762_, _06738_);
  nor _15279_ (_06879_, _06878_, _06623_);
  nand _15280_ (_06880_, _06620_, _06606_);
  and _15281_ (_06882_, _06880_, _06728_);
  nor _15282_ (_06883_, _06610_, _06629_);
  and _15283_ (_06885_, _06883_, _06615_);
  and _15284_ (_06886_, _06885_, _06882_);
  and _15285_ (_06887_, _06886_, _06879_);
  and _15286_ (_06888_, _06597_, _06606_);
  or _15287_ (_06889_, _06888_, _06628_);
  nor _15288_ (_06890_, _06889_, _06603_);
  and _15289_ (_06891_, _06890_, _06824_);
  and _15290_ (_06892_, _06743_, _05978_);
  nor _15291_ (_06893_, _06892_, _06627_);
  and _15292_ (_06894_, _06893_, _06602_);
  and _15293_ (_06895_, _06894_, _06891_);
  and _15294_ (_06897_, _06895_, _06887_);
  and _15295_ (_06898_, _06897_, _06877_);
  nand _15296_ (_06899_, _06898_, _06876_);
  nand _15297_ (_06900_, _06899_, _05962_);
  not _15298_ (_06901_, _06847_);
  and _15299_ (_06902_, _06901_, _06810_);
  nand _15300_ (_06903_, _06902_, _06900_);
  nand _15301_ (_06904_, _06903_, _04859_);
  and _15302_ (_06905_, _06904_, _06853_);
  or _15303_ (_06906_, _06905_, _06851_);
  or _15304_ (_06907_, _06906_, _06819_);
  nor _15305_ (_06908_, _05730_, _05104_);
  and _15306_ (_06910_, _05730_, _05734_);
  not _15307_ (_06911_, _06910_);
  and _15308_ (_06912_, _05929_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and _15309_ (_06913_, _05935_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor _15310_ (_06915_, _06913_, _06912_);
  and _15311_ (_06916_, _05927_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and _15312_ (_06917_, _05742_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor _15313_ (_06918_, _06917_, _06916_);
  and _15314_ (_06919_, _05758_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  and _15315_ (_06920_, _05933_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nor _15316_ (_06921_, _06920_, _06919_);
  and _15317_ (_06922_, _06921_, _06918_);
  and _15318_ (_06923_, _06922_, _06915_);
  nor _15319_ (_06924_, _06923_, _06911_);
  nor _15320_ (_06925_, _06924_, _06908_);
  or _15321_ (_06926_, _06925_, _06907_);
  and _15322_ (_06928_, _06905_, _06851_);
  and _15323_ (_06929_, _06928_, _06818_);
  not _15324_ (_06930_, _04922_);
  and _15325_ (_06931_, _05510_, _05001_);
  and _15326_ (_06932_, _06931_, _04934_);
  and _15327_ (_06934_, _06932_, _06662_);
  not _15328_ (_06935_, _06934_);
  and _15329_ (_06936_, _06935_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and _15330_ (_06937_, _06934_, _06410_);
  nor _15331_ (_06938_, _06937_, _06936_);
  nor _15332_ (_06940_, _06938_, _06930_);
  and _15333_ (_06941_, _06938_, _06930_);
  nor _15334_ (_06943_, _06941_, _06940_);
  and _15335_ (_06944_, _06935_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  nor _15336_ (_06946_, _06935_, _05669_);
  nor _15337_ (_06947_, _06946_, _06944_);
  and _15338_ (_06948_, _06947_, _04948_);
  or _15339_ (_06949_, _06947_, _04948_);
  nor _15340_ (_06950_, _05772_, _04958_);
  and _15341_ (_06951_, _05772_, _04958_);
  or _15342_ (_06952_, _06951_, _05007_);
  nor _15343_ (_06953_, _06952_, _06950_);
  nand _15344_ (_06955_, _06953_, _06949_);
  nor _15345_ (_06956_, _06955_, _06948_);
  and _15346_ (_06957_, _06956_, _06943_);
  and _15347_ (_06958_, _06957_, _06369_);
  not _15348_ (_06959_, _06938_);
  nor _15349_ (_06960_, _06947_, _05773_);
  and _15350_ (_06961_, _06960_, _06959_);
  and _15351_ (_06962_, _06961_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  and _15352_ (_06963_, _06947_, _05773_);
  and _15353_ (_06964_, _06963_, _06938_);
  and _15354_ (_06965_, _06964_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  nor _15355_ (_06966_, _06965_, _06962_);
  nor _15356_ (_06967_, _06947_, _05772_);
  and _15357_ (_06968_, _06967_, _06959_);
  and _15358_ (_06969_, _06968_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  and _15359_ (_06970_, _06960_, _06938_);
  and _15360_ (_06971_, _06970_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  nor _15361_ (_06972_, _06971_, _06969_);
  and _15362_ (_06973_, _06972_, _06966_);
  not _15363_ (_06974_, _06957_);
  and _15364_ (_06976_, _06963_, _06959_);
  nand _15365_ (_06977_, _06976_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  and _15366_ (_06978_, _06947_, _05772_);
  and _15367_ (_06979_, _06978_, _06938_);
  nand _15368_ (_06980_, _06979_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  and _15369_ (_06981_, _06980_, _06977_);
  not _15370_ (_06982_, _06978_);
  nor _15371_ (_06983_, _06982_, _06938_);
  nand _15372_ (_06984_, _06983_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  and _15373_ (_06985_, _06967_, _06938_);
  nand _15374_ (_06986_, _06985_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  and _15375_ (_06987_, _06986_, _06984_);
  and _15376_ (_06988_, _06987_, _06981_);
  and _15377_ (_06989_, _06988_, _06974_);
  and _15378_ (_06990_, _06989_, _06973_);
  nor _15379_ (_06991_, _06990_, _06958_);
  nand _15380_ (_06992_, _06991_, _06929_);
  and _15381_ (_06993_, _06992_, _06926_);
  nand _15382_ (_06994_, _06904_, _06853_);
  and _15383_ (_06995_, _06994_, _06851_);
  nand _15384_ (_06996_, _06995_, _06818_);
  not _15385_ (_06997_, _06369_);
  and _15386_ (_06998_, _05510_, _04999_);
  and _15387_ (_06999_, _06998_, _05517_);
  nand _15388_ (_07000_, _06999_, _06997_);
  or _15389_ (_07001_, _06999_, _04952_);
  and _15390_ (_07002_, _07001_, _07000_);
  and _15391_ (_07003_, _07002_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  nor _15392_ (_07004_, _07002_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  nor _15393_ (_07005_, _07004_, _07003_);
  nor _15394_ (_07006_, _07005_, _04872_);
  not _15395_ (_07007_, _07006_);
  and _15396_ (_07008_, _07007_, _04953_);
  nor _15397_ (_07009_, _07008_, _06999_);
  not _15398_ (_07010_, _07009_);
  and _15399_ (_07011_, _07010_, _07000_);
  or _15400_ (_07012_, _07011_, _06996_);
  and _15401_ (_07013_, _06850_, _06821_);
  and _15402_ (_07014_, _06905_, _07013_);
  nand _15403_ (_07015_, _07014_, _06818_);
  or _15404_ (_07016_, _07015_, _05773_);
  and _15405_ (_07017_, _07016_, _07012_);
  and _15406_ (_07018_, _07017_, _06993_);
  nor _15407_ (_07019_, _05730_, _05132_);
  and _15408_ (_07020_, _05929_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and _15409_ (_07021_, _05935_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor _15410_ (_07022_, _07021_, _07020_);
  and _15411_ (_07023_, _05927_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and _15412_ (_07024_, _05742_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor _15413_ (_07025_, _07024_, _07023_);
  and _15414_ (_07026_, _05758_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  and _15415_ (_07027_, _05933_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor _15416_ (_07028_, _07027_, _07026_);
  and _15417_ (_07029_, _07028_, _07025_);
  and _15418_ (_07030_, _07029_, _07022_);
  nor _15419_ (_07031_, _07030_, _06911_);
  nor _15420_ (_07032_, _07031_, _07019_);
  or _15421_ (_07033_, _07032_, _06907_);
  or _15422_ (_07034_, _07015_, _05952_);
  and _15423_ (_07035_, _07034_, _07033_);
  and _15424_ (_07036_, _06957_, _06032_);
  and _15425_ (_07037_, _06976_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  and _15426_ (_07038_, _06985_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  nor _15427_ (_07039_, _07038_, _07037_);
  and _15428_ (_07040_, _06961_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  and _15429_ (_07041_, _06979_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  nor _15430_ (_07042_, _07041_, _07040_);
  and _15431_ (_07043_, _07042_, _07039_);
  nand _15432_ (_07044_, _06983_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  nand _15433_ (_07045_, _06964_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  and _15434_ (_07046_, _07045_, _07044_);
  nand _15435_ (_07047_, _06968_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  nand _15436_ (_07048_, _06970_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  and _15437_ (_07049_, _07048_, _07047_);
  and _15438_ (_07050_, _07049_, _07046_);
  and _15439_ (_07051_, _07050_, _06974_);
  and _15440_ (_07052_, _07051_, _07043_);
  nor _15441_ (_07053_, _07052_, _07036_);
  nand _15442_ (_07054_, _07053_, _06929_);
  not _15443_ (_07055_, _06999_);
  or _15444_ (_07056_, _07055_, _06032_);
  not _15445_ (_07057_, _04962_);
  nand _15446_ (_07058_, _07055_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  and _15447_ (_07059_, _07058_, _07056_);
  and _15448_ (_07060_, _07059_, _07003_);
  nor _15449_ (_07061_, _07059_, _07003_);
  nor _15450_ (_07062_, _07061_, _07060_);
  nor _15451_ (_07063_, _07062_, _04872_);
  nor _15452_ (_07064_, _07063_, _07057_);
  nor _15453_ (_07065_, _07064_, _06999_);
  not _15454_ (_07066_, _07065_);
  and _15455_ (_07067_, _07066_, _07056_);
  or _15456_ (_07068_, _07067_, _06996_);
  or _15457_ (_07069_, _06994_, _07013_);
  or _15458_ (_07070_, _07069_, _06818_);
  and _15459_ (_07071_, _07070_, _07068_);
  and _15460_ (_07072_, _07071_, _07054_);
  nand _15461_ (_07073_, _07072_, _07035_);
  and _15462_ (_07074_, _07073_, _07018_);
  or _15463_ (_07075_, _07015_, _05797_);
  nor _15464_ (_07076_, _05730_, _05152_);
  and _15465_ (_07077_, _05929_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and _15466_ (_07078_, _05935_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor _15467_ (_07079_, _07078_, _07077_);
  and _15468_ (_07080_, _05927_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and _15469_ (_07081_, _05758_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  nor _15470_ (_07082_, _07081_, _07080_);
  and _15471_ (_07083_, _05933_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and _15472_ (_07084_, _05742_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor _15473_ (_07085_, _07084_, _07083_);
  and _15474_ (_07086_, _07085_, _07082_);
  and _15475_ (_07087_, _07086_, _07079_);
  nor _15476_ (_07088_, _07087_, _06911_);
  nor _15477_ (_07089_, _07088_, _07076_);
  or _15478_ (_07090_, _07089_, _06907_);
  and _15479_ (_07091_, _07090_, _07075_);
  and _15480_ (_07092_, _06995_, _06818_);
  nand _15481_ (_07093_, _06999_, _06705_);
  nand _15482_ (_07094_, _07055_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  and _15483_ (_07095_, _07094_, _07093_);
  and _15484_ (_07096_, _07095_, _07060_);
  nor _15485_ (_07097_, _07095_, _07060_);
  or _15486_ (_07098_, _07097_, _07096_);
  nand _15487_ (_07099_, _07098_, _04972_);
  nand _15488_ (_07100_, _07099_, _04975_);
  nand _15489_ (_07101_, _07100_, _07055_);
  nand _15490_ (_07102_, _07101_, _07093_);
  nand _15491_ (_07103_, _07102_, _07092_);
  or _15492_ (_07104_, _06974_, _06705_);
  nand _15493_ (_07105_, _06968_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  nand _15494_ (_07106_, _06983_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  and _15495_ (_07108_, _07106_, _07105_);
  nand _15496_ (_07109_, _06979_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  nand _15497_ (_07110_, _06985_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  and _15498_ (_07111_, _07110_, _07109_);
  and _15499_ (_07112_, _07111_, _07108_);
  not _15500_ (_07113_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  nand _15501_ (_07114_, _06960_, _06959_);
  or _15502_ (_07115_, _07114_, _07113_);
  nand _15503_ (_07116_, _06970_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  and _15504_ (_07117_, _07116_, _07115_);
  nand _15505_ (_07118_, _06976_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  nand _15506_ (_07119_, _06964_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  and _15507_ (_07120_, _07119_, _07118_);
  and _15508_ (_07121_, _07120_, _07117_);
  and _15509_ (_07122_, _07121_, _06974_);
  nand _15510_ (_07123_, _07122_, _07112_);
  and _15511_ (_07124_, _07123_, _07104_);
  nand _15512_ (_07125_, _07124_, _06929_);
  and _15513_ (_07126_, _07125_, _07103_);
  and _15514_ (_07127_, _07126_, _07091_);
  or _15515_ (_07128_, _07015_, _06947_);
  nor _15516_ (_07129_, _05730_, _05084_);
  and _15517_ (_07130_, _05929_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and _15518_ (_07131_, _05935_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor _15519_ (_07132_, _07131_, _07130_);
  and _15520_ (_07133_, _05927_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and _15521_ (_07134_, _05758_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor _15522_ (_07135_, _07134_, _07133_);
  and _15523_ (_07136_, _05933_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and _15524_ (_07137_, _05742_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor _15525_ (_07138_, _07137_, _07136_);
  and _15526_ (_07139_, _07138_, _07135_);
  and _15527_ (_07140_, _07139_, _07132_);
  nor _15528_ (_07141_, _07140_, _06911_);
  nor _15529_ (_07142_, _07141_, _07129_);
  or _15530_ (_07143_, _07142_, _06907_);
  and _15531_ (_07144_, _07143_, _07128_);
  nor _15532_ (_07145_, _07055_, _05669_);
  and _15533_ (_07146_, _07055_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor _15534_ (_07147_, _07146_, _07145_);
  and _15535_ (_07148_, _07147_, _07096_);
  nor _15536_ (_07149_, _07147_, _07096_);
  or _15537_ (_07150_, _07149_, _07148_);
  nand _15538_ (_07151_, _07150_, _04972_);
  nand _15539_ (_07152_, _07151_, _04942_);
  and _15540_ (_07153_, _07152_, _07055_);
  nor _15541_ (_07154_, _07153_, _07145_);
  or _15542_ (_07155_, _07154_, _06996_);
  and _15543_ (_07156_, _06957_, _05669_);
  and _15544_ (_07157_, _06976_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  and _15545_ (_07158_, _06985_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  nor _15546_ (_07159_, _07158_, _07157_);
  and _15547_ (_07160_, _06961_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  and _15548_ (_07161_, _06979_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  nor _15549_ (_07162_, _07161_, _07160_);
  and _15550_ (_07163_, _07162_, _07159_);
  nand _15551_ (_07164_, _06983_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  nand _15552_ (_07165_, _06964_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  and _15553_ (_07166_, _07165_, _07164_);
  nand _15554_ (_07167_, _06968_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  nand _15555_ (_07168_, _06970_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  and _15556_ (_07169_, _07168_, _07167_);
  and _15557_ (_07170_, _07169_, _07166_);
  and _15558_ (_07171_, _07170_, _06974_);
  and _15559_ (_07172_, _07171_, _07163_);
  nor _15560_ (_07173_, _07172_, _07156_);
  nand _15561_ (_07174_, _07173_, _06929_);
  and _15562_ (_07175_, _07174_, _07155_);
  and _15563_ (_07176_, _07175_, _07144_);
  and _15564_ (_07177_, _07176_, _07127_);
  nor _15565_ (_07178_, _05730_, _05062_);
  and _15566_ (_07179_, _05929_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and _15567_ (_07180_, _05935_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor _15568_ (_07181_, _07180_, _07179_);
  and _15569_ (_07182_, _05927_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and _15570_ (_07183_, _05742_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor _15571_ (_07184_, _07183_, _07182_);
  and _15572_ (_07185_, _05758_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  and _15573_ (_07186_, _05933_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nor _15574_ (_07187_, _07186_, _07185_);
  and _15575_ (_07188_, _07187_, _07184_);
  and _15576_ (_07189_, _07188_, _07181_);
  nor _15577_ (_07190_, _06911_, _07189_);
  nor _15578_ (_07191_, _07190_, _07178_);
  or _15579_ (_07192_, _07191_, _06907_);
  or _15580_ (_07193_, _07015_, _06938_);
  and _15581_ (_07194_, _07193_, _07192_);
  nor _15582_ (_07195_, _06974_, _06410_);
  and _15583_ (_07196_, _06976_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  and _15584_ (_07197_, _06985_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  nor _15585_ (_07198_, _07197_, _07196_);
  and _15586_ (_07199_, _06961_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  and _15587_ (_07200_, _06979_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  nor _15588_ (_07201_, _07200_, _07199_);
  and _15589_ (_07202_, _07201_, _07198_);
  nand _15590_ (_07203_, _06983_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  nand _15591_ (_07204_, _06964_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  and _15592_ (_07205_, _07204_, _07203_);
  nand _15593_ (_07206_, _06968_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  nand _15594_ (_07207_, _06970_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  and _15595_ (_07208_, _07207_, _07206_);
  and _15596_ (_07209_, _07208_, _07205_);
  and _15597_ (_07210_, _07209_, _06974_);
  and _15598_ (_07211_, _07210_, _07202_);
  nor _15599_ (_07212_, _07211_, _07195_);
  nand _15600_ (_07213_, _07212_, _06929_);
  and _15601_ (_07214_, _06999_, _06410_);
  and _15602_ (_07215_, _07055_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  nor _15603_ (_07216_, _07215_, _07214_);
  nand _15604_ (_07217_, _07216_, _07148_);
  or _15605_ (_07218_, _07216_, _07148_);
  nand _15606_ (_07219_, _07218_, _07217_);
  nand _15607_ (_07220_, _07219_, _04972_);
  nand _15608_ (_07221_, _07220_, _04910_);
  and _15609_ (_07222_, _07221_, _07055_);
  or _15610_ (_07223_, _07222_, _07214_);
  nand _15611_ (_07224_, _07223_, _07092_);
  or _15612_ (_07225_, _06851_, _06818_);
  and _15613_ (_07226_, _07225_, _07224_);
  and _15614_ (_07227_, _07226_, _07213_);
  and _15615_ (_07228_, _07227_, _07194_);
  or _15616_ (_07229_, _06974_, _05718_);
  nand _15617_ (_07230_, _06964_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  nand _15618_ (_07231_, _06979_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  and _15619_ (_07232_, _07231_, _07230_);
  nand _15620_ (_07233_, _06983_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  nand _15621_ (_07234_, _06985_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  and _15622_ (_07235_, _07234_, _07233_);
  and _15623_ (_07236_, _07235_, _07232_);
  nand _15624_ (_07237_, _06970_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  nand _15625_ (_07238_, _06976_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  and _15626_ (_07239_, _07238_, _07237_);
  nand _15627_ (_07240_, _06961_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  nand _15628_ (_07241_, _06968_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  and _15629_ (_07242_, _07241_, _07240_);
  and _15630_ (_07243_, _07242_, _07239_);
  and _15631_ (_07244_, _07243_, _06974_);
  nand _15632_ (_07245_, _07244_, _07236_);
  and _15633_ (_07246_, _07245_, _07229_);
  nand _15634_ (_07247_, _07246_, _06929_);
  nor _15635_ (_07248_, _05730_, _05179_);
  and _15636_ (_07249_, _05929_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and _15637_ (_07250_, _05935_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor _15638_ (_07251_, _07250_, _07249_);
  and _15639_ (_07252_, _05927_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and _15640_ (_07253_, _05758_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor _15641_ (_07254_, _07253_, _07252_);
  and _15642_ (_07255_, _05933_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and _15643_ (_07256_, _05742_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor _15644_ (_07257_, _07256_, _07255_);
  and _15645_ (_07258_, _07257_, _07254_);
  and _15646_ (_07259_, _07258_, _07251_);
  nor _15647_ (_07260_, _07259_, _06911_);
  nor _15648_ (_07261_, _07260_, _07248_);
  or _15649_ (_07262_, _07261_, _06907_);
  and _15650_ (_07263_, _07262_, _07247_);
  and _15651_ (_07264_, _06999_, _05718_);
  and _15652_ (_07265_, _07216_, _07148_);
  and _15653_ (_07266_, _07055_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor _15654_ (_07267_, _07266_, _07264_);
  nand _15655_ (_07268_, _07267_, _07265_);
  or _15656_ (_07269_, _07267_, _07265_);
  nand _15657_ (_07270_, _07269_, _07268_);
  nand _15658_ (_07271_, _07270_, _04972_);
  nand _15659_ (_07272_, _07271_, _04925_);
  and _15660_ (_07273_, _07272_, _07055_);
  nor _15661_ (_07274_, _07273_, _07264_);
  or _15662_ (_07275_, _07274_, _07013_);
  nand _15663_ (_07276_, _07275_, _06818_);
  and _15664_ (_07277_, _07069_, _06906_);
  nand _15665_ (_07278_, _07277_, _07276_);
  and _15666_ (_07279_, _07278_, _07263_);
  or _15667_ (_07280_, _06928_, _06818_);
  nor _15668_ (_07281_, _05730_, _05017_);
  and _15669_ (_07282_, _05929_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and _15670_ (_07283_, _05935_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor _15671_ (_07284_, _07283_, _07282_);
  and _15672_ (_07285_, _05927_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and _15673_ (_07286_, _05758_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor _15674_ (_07287_, _07286_, _07285_);
  and _15675_ (_07288_, _05933_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and _15676_ (_07289_, _05742_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor _15677_ (_07290_, _07289_, _07288_);
  and _15678_ (_07291_, _07290_, _07287_);
  and _15679_ (_07292_, _07291_, _07284_);
  nor _15680_ (_07293_, _07292_, _06911_);
  nor _15681_ (_07294_, _07293_, _07281_);
  or _15682_ (_07295_, _07294_, _06907_);
  and _15683_ (_07296_, _07295_, _07280_);
  nor _15684_ (_07297_, _07055_, _05287_);
  and _15685_ (_07299_, _07267_, _07265_);
  and _15686_ (_07300_, _07055_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor _15687_ (_07301_, _07300_, _07297_);
  or _15688_ (_07303_, _07301_, _07299_);
  nand _15689_ (_07304_, _07301_, _07299_);
  nand _15690_ (_07305_, _07304_, _07303_);
  nand _15691_ (_07306_, _07305_, _04972_);
  nand _15692_ (_07308_, _07306_, _04875_);
  and _15693_ (_07309_, _07308_, _07055_);
  or _15694_ (_07310_, _07309_, _07297_);
  nand _15695_ (_07311_, _07310_, _07092_);
  nand _15696_ (_07312_, _06957_, _05287_);
  or _15697_ (_07314_, _07114_, _04857_);
  nand _15698_ (_07315_, _06979_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  and _15699_ (_07316_, _07315_, _07314_);
  nand _15700_ (_07317_, _06968_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  nand _15701_ (_07319_, _06970_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  and _15702_ (_07320_, _07319_, _07317_);
  and _15703_ (_07321_, _07320_, _07316_);
  nand _15704_ (_07322_, _06983_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  nand _15705_ (_07323_, _06964_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  and _15706_ (_07325_, _07323_, _07322_);
  nand _15707_ (_07326_, _06976_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  nand _15708_ (_07327_, _06985_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  and _15709_ (_07328_, _07327_, _07326_);
  and _15710_ (_07330_, _07328_, _07325_);
  and _15711_ (_07331_, _07330_, _06974_);
  nand _15712_ (_07333_, _07331_, _07321_);
  and _15713_ (_07334_, _07333_, _07312_);
  nand _15714_ (_07335_, _07334_, _06929_);
  and _15715_ (_07336_, _07335_, _07311_);
  and _15716_ (_07337_, _07336_, _07296_);
  and _15717_ (_07338_, _06999_, _06284_);
  and _15718_ (_07339_, _07055_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  or _15719_ (_07340_, _07339_, _07304_);
  nand _15720_ (_07341_, _07339_, _07304_);
  nand _15721_ (_07342_, _07341_, _07340_);
  nand _15722_ (_07343_, _07342_, _04972_);
  and _15723_ (_07344_, _07055_, _04897_);
  and _15724_ (_07345_, _07344_, _07343_);
  nor _15725_ (_07346_, _07345_, _07338_);
  nand _15726_ (_07347_, _07346_, _06995_);
  nand _15727_ (_07348_, _06957_, _06284_);
  and _15728_ (_07349_, _06968_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  and _15729_ (_07350_, _06979_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  or _15730_ (_07351_, _07350_, _07349_);
  and _15731_ (_07352_, _06961_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  and _15732_ (_07353_, _06983_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  or _15733_ (_07354_, _07353_, _07352_);
  or _15734_ (_07355_, _07354_, _07351_);
  nand _15735_ (_07356_, _06970_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  nand _15736_ (_07357_, _06964_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  and _15737_ (_07358_, _07357_, _07356_);
  nand _15738_ (_07359_, _06976_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  nand _15739_ (_07360_, _06985_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  and _15740_ (_07361_, _07360_, _07359_);
  and _15741_ (_07362_, _07361_, _07358_);
  nand _15742_ (_07363_, _07362_, _06974_);
  or _15743_ (_07364_, _07363_, _07355_);
  and _15744_ (_07365_, _07364_, _07348_);
  nand _15745_ (_07366_, _07365_, _06929_);
  nor _15746_ (_07367_, _05730_, _05321_);
  and _15747_ (_07368_, _05929_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and _15748_ (_07369_, _05935_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor _15749_ (_07370_, _07369_, _07368_);
  and _15750_ (_07371_, _05927_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and _15751_ (_07372_, _05758_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  nor _15752_ (_07373_, _07372_, _07371_);
  and _15753_ (_07374_, _05933_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and _15754_ (_07375_, _05742_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor _15755_ (_07376_, _07375_, _07374_);
  and _15756_ (_07377_, _07376_, _07373_);
  and _15757_ (_07378_, _07377_, _07370_);
  nor _15758_ (_07379_, _07378_, _06911_);
  nor _15759_ (_07380_, _07379_, _07367_);
  or _15760_ (_07381_, _07380_, _06906_);
  and _15761_ (_07382_, _07381_, _06818_);
  and _15762_ (_07383_, _07382_, _07366_);
  nand _15763_ (_07384_, _07383_, _07347_);
  and _15764_ (_07385_, _07384_, _07337_);
  and _15765_ (_07386_, _07385_, _07279_);
  and _15766_ (_07387_, _07386_, _07228_);
  and _15767_ (_07388_, _07387_, _07177_);
  and _15768_ (_07389_, _07388_, _07074_);
  and _15769_ (_07390_, _07389_, _05292_);
  not _15770_ (_07391_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  nand _15771_ (_07392_, _07017_, _06993_);
  or _15772_ (_07393_, _07073_, _07392_);
  nand _15773_ (_07394_, _07175_, _07144_);
  and _15774_ (_07395_, _07394_, _07127_);
  not _15775_ (_07396_, _07395_);
  or _15776_ (_07397_, _07396_, _07393_);
  nand _15777_ (_07398_, _07227_, _07194_);
  nand _15778_ (_07399_, _07278_, _07263_);
  and _15779_ (_07400_, _07383_, _07347_);
  or _15780_ (_07401_, _07400_, _07337_);
  or _15781_ (_07402_, _07401_, _07399_);
  or _15782_ (_07403_, _07402_, _07398_);
  or _15783_ (_07404_, _07403_, _07397_);
  nor _15784_ (_07405_, _07404_, _07391_);
  nand _15785_ (_07406_, _07126_, _07091_);
  and _15786_ (_07407_, _07394_, _07406_);
  not _15787_ (_07408_, _07407_);
  or _15788_ (_07409_, _07408_, _07393_);
  or _15789_ (_07410_, _07409_, _07403_);
  not _15790_ (_07411_, _07410_);
  and _15791_ (_07412_, _07411_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  or _15792_ (_07414_, _07412_, _07405_);
  and _15793_ (_07415_, _07072_, _07035_);
  or _15794_ (_07417_, _07415_, _07392_);
  or _15795_ (_07418_, _07417_, _07396_);
  or _15796_ (_07420_, _07418_, _07403_);
  not _15797_ (_07422_, _07420_);
  and _15798_ (_07424_, _07422_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  or _15799_ (_07425_, _07073_, _07018_);
  or _15800_ (_07426_, _07408_, _07425_);
  or _15801_ (_07428_, _07426_, _07403_);
  not _15802_ (_07429_, _07428_);
  and _15803_ (_07430_, _07429_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  or _15804_ (_07432_, _07430_, _07424_);
  or _15805_ (_07433_, _07432_, _07414_);
  nand _15806_ (_07435_, _07386_, _07228_);
  or _15807_ (_07436_, _07397_, _07435_);
  not _15808_ (_07437_, _07436_);
  and _15809_ (_07438_, _07437_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  or _15810_ (_07439_, _07415_, _07018_);
  or _15811_ (_07440_, _07439_, _07396_);
  or _15812_ (_07441_, _07403_, _07440_);
  not _15813_ (_07442_, _07441_);
  and _15814_ (_07443_, _07442_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  or _15815_ (_07444_, _07443_, _07438_);
  and _15816_ (_07445_, _07415_, _07018_);
  and _15817_ (_07446_, _07395_, _07445_);
  and _15818_ (_07447_, _07385_, _07399_);
  and _15819_ (_07448_, _07447_, _07228_);
  and _15820_ (_07449_, _07448_, _07446_);
  and _15821_ (_07450_, _07449_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and _15822_ (_07451_, _07447_, _07398_);
  and _15823_ (_07452_, _07073_, _07392_);
  and _15824_ (_07453_, _07452_, _07406_);
  and _15825_ (_07454_, _07453_, _07176_);
  and _15826_ (_07455_, _07454_, _07451_);
  and _15827_ (_07456_, _07455_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  or _15828_ (_07457_, _07456_, _07450_);
  or _15829_ (_07458_, _07457_, _07444_);
  or _15830_ (_07459_, _07458_, _07433_);
  not _15831_ (_07460_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and _15832_ (_07461_, _07415_, _07392_);
  and _15833_ (_07462_, _07461_, _07395_);
  nand _15834_ (_07463_, _07462_, _07387_);
  nor _15835_ (_07464_, _07463_, _07460_);
  or _15836_ (_07465_, _07440_, _07435_);
  not _15837_ (_07466_, _07465_);
  and _15838_ (_07467_, _07466_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  or _15839_ (_07468_, _07467_, _07464_);
  or _15840_ (_07469_, _07418_, _07435_);
  not _15841_ (_07470_, _07469_);
  and _15842_ (_07471_, _07470_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  or _15843_ (_07472_, _07426_, _07435_);
  not _15844_ (_07473_, _07472_);
  and _15845_ (_07474_, _07473_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  or _15846_ (_07475_, _07474_, _07471_);
  or _15847_ (_07476_, _07475_, _07468_);
  nor _15848_ (_07477_, _07409_, _07435_);
  and _15849_ (_07478_, _07477_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and _15850_ (_07479_, _07454_, _07387_);
  and _15851_ (_07480_, _07479_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  or _15852_ (_07481_, _07480_, _07478_);
  and _15853_ (_07482_, _07386_, _07398_);
  nand _15854_ (_07483_, _07482_, _07462_);
  not _15855_ (_07484_, _07483_);
  and _15856_ (_07485_, _07484_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  nand _15857_ (_07486_, _07482_, _07446_);
  not _15858_ (_07487_, _07486_);
  and _15859_ (_07488_, _07487_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or _15860_ (_07489_, _07488_, _07485_);
  or _15861_ (_07490_, _07489_, _07481_);
  or _15862_ (_07491_, _07490_, _07476_);
  or _15863_ (_07492_, _07491_, _07459_);
  and _15864_ (_07493_, _07389_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and _15865_ (_07494_, _07388_, _07452_);
  and _15866_ (_07495_, _07494_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or _15867_ (_07496_, _07495_, _07493_);
  and _15868_ (_07497_, _07445_, _07177_);
  and _15869_ (_07498_, _07497_, _07398_);
  nor _15870_ (_07499_, _07401_, _07279_);
  and _15871_ (_07500_, _07499_, _07498_);
  and _15872_ (_07501_, _07500_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nand _15873_ (_07502_, _07387_, _07177_);
  or _15874_ (_07503_, _07502_, _07425_);
  nor _15875_ (_07504_, _07503_, _07011_);
  or _15876_ (_07505_, _07504_, _07501_);
  or _15877_ (_07506_, _07505_, _07496_);
  and _15878_ (_07507_, _07448_, _07497_);
  and _15879_ (_07508_, _06635_, _06731_);
  nor _15880_ (_07509_, _07508_, _06866_);
  and _15881_ (_07510_, _06637_, _05874_);
  and _15882_ (_07511_, _07510_, _05985_);
  nor _15883_ (_07512_, _07511_, _06744_);
  and _15884_ (_07513_, _06635_, _05965_);
  nor _15885_ (_07514_, _06619_, _05950_);
  nor _15886_ (_07515_, _07514_, _05822_);
  nor _15887_ (_07516_, _07515_, _07513_);
  nor _15888_ (_07518_, _06756_, _06750_);
  and _15889_ (_07519_, _07518_, _07516_);
  and _15890_ (_07521_, _07519_, _07512_);
  nor _15891_ (_07522_, _06888_, _06609_);
  nor _15892_ (_07523_, _06755_, _06595_);
  and _15893_ (_07525_, _07523_, _07522_);
  and _15894_ (_07526_, _07525_, _06748_);
  and _15895_ (_07527_, _07526_, _07521_);
  and _15896_ (_07528_, _07527_, _06887_);
  and _15897_ (_07530_, _07528_, _07509_);
  nor _15898_ (_07531_, _07530_, _06799_);
  or _15899_ (_07532_, _07531_, p2_in[0]);
  not _15900_ (_07533_, _07531_);
  or _15901_ (_07535_, _07533_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and _15902_ (_07536_, _07535_, _07532_);
  and _15903_ (_07538_, _07536_, _07507_);
  and _15904_ (_07539_, _07451_, _07497_);
  or _15905_ (_07541_, _07531_, p3_in[0]);
  or _15906_ (_07542_, _07533_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and _15907_ (_07544_, _07542_, _07541_);
  and _15908_ (_07545_, _07544_, _07539_);
  or _15909_ (_07546_, _07545_, _07538_);
  and _15910_ (_07547_, _07387_, _07497_);
  or _15911_ (_07548_, _07531_, p0_in[0]);
  or _15912_ (_07549_, _07533_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  and _15913_ (_07550_, _07549_, _07548_);
  and _15914_ (_07551_, _07550_, _07547_);
  and _15915_ (_07552_, _07482_, _07497_);
  or _15916_ (_07553_, _07531_, p1_in[0]);
  or _15917_ (_07554_, _07533_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and _15918_ (_07555_, _07554_, _07553_);
  and _15919_ (_07556_, _07555_, _07552_);
  or _15920_ (_07557_, _07556_, _07551_);
  or _15921_ (_07558_, _07557_, _07546_);
  or _15922_ (_07559_, _07558_, _07506_);
  not _15923_ (_07560_, _07402_);
  and _15924_ (_07561_, _07560_, _07498_);
  nor _15925_ (_07562_, _06666_, _06488_);
  and _15926_ (_07563_, _06678_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor _15927_ (_07564_, _07563_, _07562_);
  nor _15928_ (_07565_, _07564_, _06654_);
  not _15929_ (_07566_, _07565_);
  and _15930_ (_07567_, _06654_, _06452_);
  not _15931_ (_07568_, _06673_);
  nor _15932_ (_07569_, _06146_, _05042_);
  nor _15933_ (_07570_, _07569_, _06147_);
  nor _15934_ (_07571_, _07570_, _07568_);
  nor _15935_ (_07572_, _07571_, _07567_);
  nand _15936_ (_07573_, _07572_, _07566_);
  nand _15937_ (_07574_, _07573_, _06684_);
  or _15938_ (_07575_, _07573_, _06684_);
  and _15939_ (_07576_, _07575_, _07574_);
  or _15940_ (_07577_, _05445_, _05442_);
  nor _15941_ (_07578_, _05446_, _06454_);
  nand _15942_ (_07579_, _07578_, _07577_);
  nor _15943_ (_07580_, _05466_, _05227_);
  nor _15944_ (_07581_, _05477_, _05059_);
  nor _15945_ (_07582_, _07581_, _07580_);
  and _15946_ (_07583_, _07582_, _05368_);
  nor _15947_ (_07584_, _07582_, _05368_);
  or _15948_ (_07585_, _07584_, _07583_);
  and _15949_ (_07586_, _07585_, _05223_);
  nor _15950_ (_07587_, _05490_, _05048_);
  nor _15951_ (_07588_, _05368_, _05274_);
  and _15952_ (_07589_, _05497_, ABINPUT001[11]);
  or _15953_ (_07590_, _07589_, _07588_);
  nor _15954_ (_07591_, _07590_, _07587_);
  nor _15955_ (_07592_, _05232_, _05172_);
  and _15956_ (_07593_, _05499_, ABINPUT000[11]);
  nor _15957_ (_07594_, _07593_, _07592_);
  and _15958_ (_07595_, _07594_, _07591_);
  not _15959_ (_07596_, _07595_);
  nor _15960_ (_07597_, _07596_, _07586_);
  nand _15961_ (_07598_, _07597_, _07579_);
  nand _15962_ (_07599_, _07598_, _06654_);
  nor _15963_ (_07600_, _06672_, _05167_);
  nor _15964_ (_07601_, _07600_, _06675_);
  and _15965_ (_07602_, _06494_, _06144_);
  nor _15966_ (_07603_, _06494_, _05167_);
  or _15967_ (_07604_, _07603_, _07602_);
  nand _15968_ (_07605_, _07604_, _06672_);
  and _15969_ (_07606_, _07605_, _07601_);
  nor _15970_ (_07607_, _06654_, _06552_);
  nor _15971_ (_07609_, _07607_, _06667_);
  or _15972_ (_07610_, _07609_, _07606_);
  nand _15973_ (_07612_, _07610_, _07599_);
  or _15974_ (_07613_, _05446_, _05310_);
  nor _15975_ (_07614_, _05447_, _06454_);
  nand _15976_ (_07616_, _07614_, _07613_);
  and _15977_ (_07617_, _05478_, _05227_);
  and _15978_ (_07619_, _05467_, _05059_);
  nor _15979_ (_07620_, _07619_, _07617_);
  and _15980_ (_07621_, _07620_, _05356_);
  not _15981_ (_07622_, _07621_);
  nor _15982_ (_07624_, _07620_, _05356_);
  nor _15983_ (_07625_, _07624_, _06363_);
  and _15984_ (_07626_, _07625_, _07622_);
  nor _15985_ (_07628_, _05356_, _05274_);
  and _15986_ (_07629_, _05497_, ABINPUT001[12]);
  or _15987_ (_07631_, _07629_, _07628_);
  nor _15988_ (_07632_, _07631_, _06061_);
  nor _15989_ (_07633_, _05232_, _05103_);
  and _15990_ (_07634_, _05499_, ABINPUT000[12]);
  nor _15991_ (_07636_, _07634_, _07633_);
  and _15992_ (_07637_, _07636_, _07632_);
  not _15993_ (_07638_, _07637_);
  nor _15994_ (_07639_, _07638_, _07626_);
  nand _15995_ (_07640_, _07639_, _07616_);
  or _15996_ (_07641_, _07640_, _06656_);
  and _15997_ (_07642_, _06144_, _05520_);
  nor _15998_ (_07643_, _05520_, _05099_);
  or _15999_ (_07644_, _07643_, _07642_);
  nand _16000_ (_07645_, _07644_, _06673_);
  nor _16001_ (_07646_, _06666_, _06586_);
  and _16002_ (_07647_, _06678_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor _16003_ (_07648_, _07647_, _07646_);
  and _16004_ (_07649_, _07648_, _07645_);
  nand _16005_ (_07650_, _07649_, _06656_);
  nand _16006_ (_07651_, _07650_, _07641_);
  nand _16007_ (_07652_, _07651_, _07612_);
  or _16008_ (_07653_, _07651_, _07612_);
  and _16009_ (_07654_, _07653_, _07652_);
  or _16010_ (_07655_, _05437_, _05434_);
  nor _16011_ (_07656_, _05438_, _06454_);
  nand _16012_ (_07657_, _07656_, _07655_);
  and _16013_ (_07658_, _05464_, _05059_);
  and _16014_ (_07659_, _05475_, _05227_);
  nor _16015_ (_07660_, _07659_, _07658_);
  and _16016_ (_07661_, _07660_, _05383_);
  nor _16017_ (_07662_, _07660_, _05383_);
  nor _16018_ (_07663_, _07662_, _07661_);
  and _16019_ (_07664_, _07663_, _05223_);
  nor _16020_ (_07665_, _05490_, _05081_);
  nor _16021_ (_07666_, _05383_, _05274_);
  and _16022_ (_07667_, _05497_, ABINPUT001[9]);
  or _16023_ (_07668_, _07667_, _07666_);
  nor _16024_ (_07669_, _07668_, _07665_);
  and _16025_ (_07670_, _05231_, _05206_);
  and _16026_ (_07671_, _05499_, ABINPUT000[9]);
  nor _16027_ (_07672_, _07671_, _07670_);
  and _16028_ (_07673_, _07672_, _07669_);
  not _16029_ (_07674_, _07673_);
  nor _16030_ (_07675_, _07674_, _07664_);
  nand _16031_ (_07676_, _07675_, _07657_);
  and _16032_ (_07677_, _07676_, _06654_);
  nor _16033_ (_07678_, _05397_, _05059_);
  nor _16034_ (_07679_, _07678_, _05398_);
  not _16035_ (_07680_, _07679_);
  nor _16036_ (_07681_, _05455_, _05583_);
  nor _16037_ (_07682_, _07681_, _07680_);
  not _16038_ (_07683_, _07682_);
  and _16039_ (_07684_, _05530_, _06064_);
  and _16040_ (_07685_, _05489_, _05059_);
  and _16041_ (_07686_, _05497_, ABINPUT001[1]);
  and _16042_ (_07687_, _05499_, ABINPUT000[1]);
  nor _16043_ (_07688_, _07687_, _07686_);
  not _16044_ (_07689_, _07688_);
  nor _16045_ (_07690_, _07689_, _07685_);
  not _16046_ (_07691_, _07690_);
  nor _16047_ (_07692_, _07691_, _07684_);
  or _16048_ (_07693_, _06468_, _05151_);
  nor _16049_ (_07694_, _05557_, _05273_);
  nor _16050_ (_07695_, _07694_, _05126_);
  not _16051_ (_07696_, _07695_);
  and _16052_ (_07697_, _07696_, _07693_);
  and _16053_ (_07698_, _07697_, _07692_);
  and _16054_ (_07699_, _07698_, _06365_);
  and _16055_ (_07700_, _07699_, _06361_);
  and _16056_ (_07701_, _07700_, _06358_);
  and _16057_ (_07702_, _07701_, _07683_);
  nor _16058_ (_07703_, _07702_, _06666_);
  and _16059_ (_07704_, _06678_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor _16060_ (_07705_, _07704_, _07703_);
  nor _16061_ (_07706_, _07705_, _06654_);
  nor _16062_ (_07707_, _07706_, _07677_);
  and _16063_ (_07708_, _06144_, _04990_);
  nor _16064_ (_07709_, _04990_, _05122_);
  or _16065_ (_07710_, _07709_, _07708_);
  nand _16066_ (_07711_, _07710_, _06673_);
  and _16067_ (_07712_, _07711_, _07707_);
  and _16068_ (_07713_, _06144_, _04986_);
  nor _16069_ (_07714_, _04986_, _05147_);
  or _16070_ (_07715_, _07714_, _07713_);
  nand _16071_ (_07716_, _07715_, _06673_);
  or _16072_ (_07717_, _05441_, _05438_);
  nor _16073_ (_07718_, _05442_, _06454_);
  nand _16074_ (_07719_, _07718_, _07717_);
  and _16075_ (_07720_, _05476_, _05227_);
  and _16076_ (_07721_, _05465_, _05059_);
  nor _16077_ (_07722_, _07721_, _07720_);
  nor _16078_ (_07723_, _07722_, _05377_);
  and _16079_ (_07724_, _07722_, _05377_);
  nor _16080_ (_07725_, _07724_, _07723_);
  nor _16081_ (_07726_, _07725_, _06363_);
  nor _16082_ (_07727_, _05490_, _05199_);
  and _16083_ (_07729_, _05377_, _05273_);
  and _16084_ (_07730_, _05497_, ABINPUT001[10]);
  or _16085_ (_07732_, _07730_, _07729_);
  nor _16086_ (_07733_, _07732_, _07727_);
  and _16087_ (_07735_, _05231_, _05207_);
  and _16088_ (_07736_, _05499_, ABINPUT000[10]);
  nor _16089_ (_07737_, _07736_, _07735_);
  and _16090_ (_07739_, _07737_, _07733_);
  not _16091_ (_07740_, _07739_);
  nor _16092_ (_07741_, _07740_, _07726_);
  nand _16093_ (_07743_, _07741_, _07719_);
  and _16094_ (_07744_, _07743_, _06654_);
  nor _16095_ (_07746_, _05618_, _05617_);
  nor _16096_ (_07748_, _07746_, _05619_);
  nor _16097_ (_07749_, _07748_, _05584_);
  not _16098_ (_07751_, _07749_);
  or _16099_ (_07752_, _06468_, _05172_);
  and _16100_ (_07753_, _05497_, ABINPUT001[2]);
  and _16101_ (_07754_, _05499_, ABINPUT000[2]);
  nor _16102_ (_07755_, _07754_, _07753_);
  and _16103_ (_07756_, _07755_, _07752_);
  and _16104_ (_07757_, _05273_, _05207_);
  and _16105_ (_07758_, _05280_, _05206_);
  nor _16106_ (_07759_, _07758_, _07757_);
  and _16107_ (_07760_, _07759_, _07756_);
  and _16108_ (_07761_, _07760_, _06030_);
  and _16109_ (_07762_, _06512_, _05207_);
  nor _16110_ (_07763_, _07762_, _06513_);
  nor _16111_ (_07764_, _07763_, _05558_);
  not _16112_ (_07765_, _05385_);
  and _16113_ (_07766_, _06020_, _07765_);
  or _16114_ (_07767_, _07766_, _05389_);
  and _16115_ (_07768_, _07767_, _05398_);
  nor _16116_ (_07769_, _07767_, _05398_);
  or _16117_ (_07770_, _07769_, _07768_);
  and _16118_ (_07771_, _07770_, _05455_);
  nor _16119_ (_07772_, _07771_, _07764_);
  and _16120_ (_07773_, _07772_, _07761_);
  and _16121_ (_07774_, _07773_, _07751_);
  nor _16122_ (_07775_, _07774_, _06666_);
  and _16123_ (_07776_, _06678_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor _16124_ (_07777_, _07776_, _07775_);
  nor _16125_ (_07778_, _07777_, _06654_);
  nor _16126_ (_07779_, _07778_, _07744_);
  nand _16127_ (_07780_, _07779_, _07716_);
  nand _16128_ (_07781_, _07780_, _07712_);
  or _16129_ (_07782_, _07780_, _07712_);
  nand _16130_ (_07783_, _07782_, _07781_);
  nand _16131_ (_07784_, _07783_, _07654_);
  or _16132_ (_07785_, _07783_, _07654_);
  nand _16133_ (_07786_, _07785_, _07784_);
  nor _16134_ (_07787_, _05627_, _05349_);
  and _16135_ (_07788_, _05627_, _05349_);
  nor _16136_ (_07789_, _07788_, _07787_);
  and _16137_ (_07790_, _07789_, _05583_);
  not _16138_ (_07791_, _07790_);
  nor _16139_ (_07792_, _05407_, _05349_);
  nor _16140_ (_07793_, _07792_, _06454_);
  and _16141_ (_07794_, _07793_, _05408_);
  nor _16142_ (_07795_, _05560_, _05565_);
  not _16143_ (_07796_, _07795_);
  nor _16144_ (_07797_, _05567_, _05558_);
  and _16145_ (_07798_, _07797_, _07796_);
  and _16146_ (_07799_, _05280_, _05204_);
  and _16147_ (_07800_, _05497_, ABINPUT001[5]);
  and _16148_ (_07801_, _05499_, ABINPUT000[5]);
  nor _16149_ (_07802_, _07801_, _07800_);
  not _16150_ (_07803_, _07802_);
  nor _16151_ (_07804_, _07803_, _07799_);
  or _16152_ (_07805_, _06468_, _05199_);
  not _16153_ (_07806_, _07805_);
  nor _16154_ (_07807_, _05274_, _05081_);
  nor _16155_ (_07808_, _07807_, _07806_);
  and _16156_ (_07809_, _07808_, _07804_);
  not _16157_ (_07810_, _07809_);
  nor _16158_ (_07811_, _07810_, _07798_);
  and _16159_ (_07812_, _07811_, _06409_);
  not _16160_ (_07813_, _07812_);
  nor _16161_ (_07814_, _07813_, _07794_);
  and _16162_ (_07815_, _07814_, _07791_);
  nor _16163_ (_07816_, _07815_, _06666_);
  and _16164_ (_07817_, _06678_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor _16165_ (_07818_, _07817_, _07816_);
  nor _16166_ (_07819_, _07818_, _06654_);
  not _16167_ (_07820_, _07819_);
  or _16168_ (_07821_, _05450_, _05447_);
  and _16169_ (_07822_, _05451_, _05455_);
  and _16170_ (_07823_, _07822_, _07821_);
  and _16171_ (_07824_, _05468_, _05059_);
  and _16172_ (_07825_, _07617_, _05622_);
  nor _16173_ (_07826_, _07825_, _07824_);
  nand _16174_ (_07828_, _07826_, _05346_);
  or _16175_ (_07829_, _07826_, _05346_);
  and _16176_ (_07831_, _07829_, _07828_);
  and _16177_ (_07832_, _07831_, _05223_);
  and _16178_ (_07833_, _05489_, _05206_);
  nand _16179_ (_07835_, _05081_, _05059_);
  and _16180_ (_07836_, _05346_, _05227_);
  nor _16181_ (_07838_, _07836_, _05232_);
  and _16182_ (_07840_, _07838_, _07835_);
  nor _16183_ (_07841_, _05346_, _05274_);
  and _16184_ (_07843_, _05497_, ABINPUT001[13]);
  and _16185_ (_07845_, _05499_, ABINPUT000[13]);
  or _16186_ (_07846_, _07845_, _07843_);
  or _16187_ (_07847_, _07846_, _07841_);
  or _16188_ (_07848_, _07847_, _07840_);
  or _16189_ (_07850_, _07848_, _07833_);
  or _16190_ (_07851_, _07850_, _07832_);
  or _16191_ (_07853_, _07851_, _07823_);
  nand _16192_ (_07854_, _07853_, _06654_);
  and _16193_ (_07855_, _04989_, _06090_);
  and _16194_ (_07857_, _07855_, _06144_);
  nor _16195_ (_07858_, _07855_, _05075_);
  or _16196_ (_07859_, _07858_, _07857_);
  nand _16197_ (_07860_, _07859_, _06673_);
  and _16198_ (_07861_, _07860_, _07854_);
  nand _16199_ (_07862_, _07861_, _07820_);
  nor _16200_ (_07863_, _06672_, _05194_);
  nor _16201_ (_07864_, _07863_, _06675_);
  and _16202_ (_07865_, _06091_, _06144_);
  nor _16203_ (_07866_, _06091_, _05194_);
  or _16204_ (_07867_, _07866_, _07865_);
  nand _16205_ (_07868_, _07867_, _06673_);
  and _16206_ (_07869_, _07868_, _07864_);
  nor _16207_ (_07870_, _05628_, _05600_);
  nor _16208_ (_07871_, _07870_, _05629_);
  nor _16209_ (_07872_, _07871_, _05584_);
  not _16210_ (_07873_, _07872_);
  and _16211_ (_07874_, _05421_, _05408_);
  nor _16212_ (_07875_, _07874_, _06454_);
  and _16213_ (_07876_, _07875_, _05422_);
  nor _16214_ (_07877_, _05568_, _05199_);
  nor _16215_ (_07878_, _07877_, _06462_);
  nor _16216_ (_07879_, _07878_, _05558_);
  and _16217_ (_07880_, _05280_, _05565_);
  and _16218_ (_07881_, _05497_, ABINPUT001[6]);
  and _16219_ (_07882_, _05499_, ABINPUT000[6]);
  nor _16220_ (_07883_, _07882_, _07881_);
  not _16221_ (_07884_, _07883_);
  nor _16222_ (_07885_, _07884_, _07880_);
  or _16223_ (_07886_, _06468_, _05048_);
  nor _16224_ (_07887_, _05274_, _05199_);
  not _16225_ (_07888_, _07887_);
  and _16226_ (_07889_, _07888_, _07886_);
  and _16227_ (_07890_, _07889_, _07885_);
  and _16228_ (_07891_, _07890_, _05716_);
  not _16229_ (_07892_, _07891_);
  nor _16230_ (_07893_, _07892_, _07879_);
  and _16231_ (_07894_, _07893_, _05702_);
  not _16232_ (_07895_, _07894_);
  nor _16233_ (_07896_, _07895_, _07876_);
  and _16234_ (_07897_, _07896_, _07873_);
  and _16235_ (_07898_, _07897_, _06675_);
  or _16236_ (_07899_, _07898_, _07869_);
  nand _16237_ (_07900_, _07899_, _06656_);
  nand _16238_ (_07901_, _05451_, _05307_);
  and _16239_ (_07902_, _05452_, _05455_);
  and _16240_ (_07903_, _07902_, _07901_);
  not _16241_ (_07904_, _05414_);
  nor _16242_ (_07905_, _07825_, _05469_);
  nor _16243_ (_07906_, _07905_, _07836_);
  or _16244_ (_07907_, _07906_, _07904_);
  nand _16245_ (_07908_, _07906_, _07904_);
  and _16246_ (_07909_, _07908_, _07907_);
  and _16247_ (_07910_, _07909_, _05223_);
  and _16248_ (_07911_, _05489_, _05207_);
  nor _16249_ (_07912_, _05199_, _05227_);
  or _16250_ (_07913_, _07912_, _05479_);
  and _16251_ (_07914_, _07913_, _05231_);
  nor _16252_ (_07915_, _05414_, _05274_);
  and _16253_ (_07916_, _05497_, ABINPUT001[14]);
  and _16254_ (_07917_, _05499_, ABINPUT000[14]);
  or _16255_ (_07918_, _07917_, _07916_);
  or _16256_ (_07919_, _07918_, _07915_);
  or _16257_ (_07920_, _07919_, _07914_);
  or _16258_ (_07921_, _07920_, _07911_);
  or _16259_ (_07922_, _07921_, _07910_);
  or _16260_ (_07924_, _07922_, _07903_);
  or _16261_ (_07925_, _07924_, _06656_);
  nand _16262_ (_07927_, _07925_, _07900_);
  nand _16263_ (_07928_, _07927_, _07862_);
  or _16264_ (_07929_, _07927_, _07862_);
  nand _16265_ (_07931_, _07929_, _07928_);
  nand _16266_ (_07932_, _07931_, _07786_);
  or _16267_ (_07933_, _07931_, _07786_);
  nand _16268_ (_07935_, _07933_, _07932_);
  nor _16269_ (_07936_, _07935_, _07576_);
  and _16270_ (_07937_, _07935_, _07576_);
  or _16271_ (_07939_, _07937_, _07936_);
  and _16272_ (_07940_, _07939_, _07561_);
  and _16273_ (_07942_, _07499_, _07228_);
  and _16274_ (_07943_, _07942_, _07497_);
  and _16275_ (_07944_, _07943_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or _16276_ (_07945_, _07944_, _07940_);
  or _16277_ (_07947_, _07945_, _07559_);
  or _16278_ (_07948_, _07947_, _07492_);
  nor _16279_ (_07949_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  not _16280_ (_07951_, _07949_);
  nand _16281_ (_07952_, _07951_, _07561_);
  or _16282_ (_07953_, _07502_, _07439_);
  or _16283_ (_07954_, _07953_, _05293_);
  nand _16284_ (_07955_, _07943_, _06654_);
  and _16285_ (_07956_, _07955_, _07954_);
  nand _16286_ (_07957_, _07956_, _07952_);
  nand _16287_ (_07958_, _07957_, _04859_);
  or _16288_ (_07959_, _07228_, _06930_);
  or _16289_ (_07960_, _07398_, _04922_);
  nand _16290_ (_07961_, _07960_, _07959_);
  or _16291_ (_07962_, _07392_, _04958_);
  or _16292_ (_07963_, _07018_, _04959_);
  nand _16293_ (_07964_, _07963_, _07962_);
  nor _16294_ (_07965_, _07964_, _07961_);
  or _16295_ (_07966_, _07073_, _04971_);
  or _16296_ (_07967_, _07279_, _04932_);
  or _16297_ (_07968_, _07399_, _04933_);
  and _16298_ (_07969_, _07968_, _07967_);
  or _16299_ (_07970_, _07337_, _04893_);
  nand _16300_ (_07971_, _07336_, _07296_);
  or _16301_ (_07972_, _07971_, _05513_);
  and _16302_ (_07973_, _07972_, _07970_);
  nor _16303_ (_07974_, _07973_, _07969_);
  and _16304_ (_07975_, _07974_, _07966_);
  and _16305_ (_07976_, _07975_, _07965_);
  or _16306_ (_07977_, _07176_, _04947_);
  or _16307_ (_07978_, _07394_, _04948_);
  and _16308_ (_07979_, _07978_, _07977_);
  or _16309_ (_07980_, _07400_, _04904_);
  or _16310_ (_07981_, _07384_, _06133_);
  and _16311_ (_07982_, _07981_, _07980_);
  nor _16312_ (_07983_, _07982_, _07979_);
  or _16313_ (_07984_, _07127_, _06090_);
  or _16314_ (_07985_, _07406_, _04984_);
  nand _16315_ (_07986_, _07985_, _07984_);
  or _16316_ (_07987_, _07415_, _04996_);
  nand _16317_ (_07988_, _07987_, _06092_);
  nor _16318_ (_07989_, _07988_, _07986_);
  and _16319_ (_07990_, _07989_, _07983_);
  nand _16320_ (_07991_, _07990_, _07976_);
  or _16321_ (_07992_, _04904_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  or _16322_ (_07993_, _07992_, _07991_);
  not _16323_ (_07994_, _07961_);
  and _16324_ (_07995_, _07974_, _07994_);
  and _16325_ (_07996_, _07995_, _07983_);
  not _16326_ (_07997_, _07453_);
  and _16327_ (_07998_, _07997_, _06141_);
  nand _16328_ (_07999_, _07998_, _07996_);
  nand _16329_ (_08000_, _07943_, _06660_);
  and _16330_ (_08001_, _08000_, _07999_);
  nand _16331_ (_08002_, _08001_, _07993_);
  nand _16332_ (_08003_, _08002_, _04859_);
  and _16333_ (_08004_, _08003_, _07958_);
  and _16334_ (_08005_, _08004_, _07948_);
  and _16335_ (_08006_, _07410_, _07404_);
  and _16336_ (_08007_, _07428_, _07420_);
  and _16337_ (_08008_, _08007_, _08006_);
  and _16338_ (_08009_, _07441_, _07436_);
  nor _16339_ (_08010_, _07455_, _07449_);
  and _16340_ (_08011_, _08010_, _08009_);
  and _16341_ (_08012_, _08011_, _08008_);
  and _16342_ (_08013_, _07465_, _07463_);
  and _16343_ (_08014_, _07472_, _07469_);
  and _16344_ (_08015_, _08014_, _08013_);
  nor _16345_ (_08016_, _07479_, _07477_);
  and _16346_ (_08017_, _07486_, _07483_);
  and _16347_ (_08018_, _08017_, _08016_);
  and _16348_ (_08019_, _08018_, _08015_);
  and _16349_ (_08021_, _08019_, _08012_);
  nor _16350_ (_08022_, _07943_, _07561_);
  nand _16351_ (_08024_, _07385_, _07497_);
  or _16352_ (_08025_, _07502_, _07417_);
  and _16353_ (_08027_, _07953_, _08025_);
  and _16354_ (_08028_, _07388_, _07461_);
  nor _16355_ (_08029_, _08028_, _07500_);
  and _16356_ (_08031_, _08029_, _08027_);
  and _16357_ (_08032_, _08031_, _08024_);
  and _16358_ (_08033_, _08032_, _08022_);
  nand _16359_ (_08034_, _08033_, _08021_);
  and _16360_ (_08036_, _08034_, _07958_);
  nand _16361_ (_08037_, _08036_, _08003_);
  and _16362_ (_08038_, _08037_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  or _16363_ (_08040_, _08038_, _08005_);
  or _16364_ (_08041_, _08040_, _07390_);
  nand _16365_ (_08043_, _07390_, _07702_);
  and _16366_ (_08044_, _08043_, _04856_);
  and _16367_ (_05133_, _08044_, _08041_);
  and _16368_ (_08046_, _06721_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and _16369_ (_08047_, _06624_, _05998_);
  or _16370_ (_08048_, _08047_, _06838_);
  or _16371_ (_08049_, _08048_, _06727_);
  and _16372_ (_08050_, _07510_, _05978_);
  or _16373_ (_08051_, _08050_, _06747_);
  and _16374_ (_08052_, _06612_, _05998_);
  or _16375_ (_08053_, _08052_, _06788_);
  or _16376_ (_08054_, _08053_, _08051_);
  or _16377_ (_08055_, _08054_, _08049_);
  and _16378_ (_08056_, _08055_, _06770_);
  or _16379_ (_05136_, _08056_, _08046_);
  nor _16380_ (_08057_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , rst);
  and _16381_ (_08058_, _08057_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  not _16382_ (_08059_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  nor _16383_ (_08060_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  nor _16384_ (_08061_, _08060_, _08059_);
  and _16385_ (_08062_, _08061_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re );
  not _16386_ (_08063_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  nor _16387_ (_08064_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _08063_);
  not _16388_ (_08065_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  nor _16389_ (_08066_, _08065_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  and _16390_ (_08067_, _08066_, _08064_);
  not _16391_ (_08068_, _08067_);
  and _16392_ (_08069_, _08068_, _08062_);
  not _16393_ (_08070_, _08060_);
  and _16394_ (_08071_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and _16395_ (_08072_, _08071_, _08070_);
  not _16396_ (_08073_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  nor _16397_ (_08074_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0], _08073_);
  and _16398_ (_08075_, _08074_, _08059_);
  and _16399_ (_08076_, _08075_, _08060_);
  nor _16400_ (_08077_, _08076_, _08062_);
  not _16401_ (_08078_, _08077_);
  nor _16402_ (_08079_, _08078_, _08072_);
  nor _16403_ (_08080_, _08079_, _08069_);
  and _16404_ (_08081_, _08060_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  and _16405_ (_08082_, _08081_, \oc8051_top_1.oc8051_sfr1.pres_ow );
  or _16406_ (_08083_, _08082_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  or _16407_ (_08084_, _08083_, _08080_);
  and _16408_ (_08085_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _04856_);
  and _16409_ (_08086_, _08067_, _08062_);
  nor _16410_ (_08087_, _08086_, _08082_);
  or _16411_ (_08088_, _08087_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  and _16412_ (_08089_, _08088_, _08085_);
  and _16413_ (_08090_, _08089_, _08084_);
  or _16414_ (_05143_, _08090_, _08058_);
  not _16415_ (_08091_, _05843_);
  not _16416_ (_08092_, _05818_);
  and _16417_ (_08093_, _08092_, _05793_);
  and _16418_ (_08094_, _08093_, _08091_);
  and _16419_ (_08095_, _08094_, _05767_);
  not _16420_ (_08096_, _05895_);
  and _16421_ (_08097_, _08096_, _05870_);
  and _16422_ (_08098_, _05943_, _05919_);
  and _16423_ (_08099_, _08098_, _08097_);
  and _16424_ (_08100_, _08099_, _08095_);
  not _16425_ (_08101_, _05919_);
  nor _16426_ (_08102_, _05943_, _08101_);
  and _16427_ (_08103_, _05895_, _05870_);
  and _16428_ (_08104_, _08103_, _08102_);
  and _16429_ (_08105_, _08104_, _08094_);
  nor _16430_ (_08106_, _08105_, _08100_);
  nor _16431_ (_08107_, _05818_, _05793_);
  nor _16432_ (_08108_, _05767_, _05843_);
  and _16433_ (_08109_, _08108_, _08107_);
  nor _16434_ (_08110_, _05943_, _05919_);
  and _16435_ (_08111_, _08110_, _08097_);
  not _16436_ (_08112_, _05870_);
  and _16437_ (_08113_, _05895_, _08112_);
  and _16438_ (_08114_, _08113_, _08110_);
  or _16439_ (_08115_, _08114_, _08111_);
  and _16440_ (_08116_, _08115_, _08109_);
  not _16441_ (_08117_, _05767_);
  and _16442_ (_08119_, _08107_, _05843_);
  and _16443_ (_08120_, _08119_, _08117_);
  and _16444_ (_08121_, _08110_, _08096_);
  and _16445_ (_08122_, _08121_, _08120_);
  nor _16446_ (_08123_, _08122_, _08116_);
  nand _16447_ (_08124_, _08123_, _08106_);
  and _16448_ (_08125_, _05943_, _08101_);
  and _16449_ (_08126_, _08125_, _08103_);
  and _16450_ (_08127_, _08126_, _08109_);
  and _16451_ (_08128_, _08107_, _08091_);
  not _16452_ (_08130_, _08128_);
  and _16453_ (_08131_, _08125_, _08113_);
  nor _16454_ (_08132_, _08131_, _05767_);
  nor _16455_ (_08133_, _08132_, _08130_);
  nor _16456_ (_08134_, _08133_, _08127_);
  nor _16457_ (_08135_, _05895_, _05870_);
  and _16458_ (_08136_, _08135_, _08102_);
  and _16459_ (_08137_, _08136_, _08109_);
  and _16460_ (_08138_, _08098_, _08096_);
  and _16461_ (_08139_, _05818_, _05870_);
  and _16462_ (_08140_, _08139_, _08138_);
  nor _16463_ (_08142_, _08140_, _08137_);
  nand _16464_ (_08143_, _08142_, _08134_);
  or _16465_ (_08144_, _08143_, _08124_);
  or _16466_ (_08145_, _08119_, _08109_);
  and _16467_ (_08146_, _08125_, _08097_);
  and _16468_ (_08147_, _08146_, _08109_);
  and _16469_ (_08149_, _08098_, _05895_);
  or _16470_ (_08150_, _08149_, _08147_);
  and _16471_ (_08151_, _08150_, _08145_);
  not _16472_ (_08152_, _08109_);
  and _16473_ (_08153_, _08110_, _08103_);
  and _16474_ (_08154_, _08125_, _08135_);
  nor _16475_ (_08155_, _08154_, _08153_);
  nor _16476_ (_08156_, _08155_, _08152_);
  and _16477_ (_08157_, _08108_, _08093_);
  and _16478_ (_08158_, _08102_, _08112_);
  and _16479_ (_08159_, _08158_, _08157_);
  and _16480_ (_08160_, _08119_, _05767_);
  and _16481_ (_08161_, _08160_, _08126_);
  or _16482_ (_08162_, _08161_, _08159_);
  or _16483_ (_08163_, _08162_, _08156_);
  and _16484_ (_08164_, _08153_, _08120_);
  and _16485_ (_08165_, _08102_, _08096_);
  and _16486_ (_08166_, _08160_, _08165_);
  or _16487_ (_08167_, _08166_, _08164_);
  and _16488_ (_08168_, _08120_, _08114_);
  and _16489_ (_08169_, _08102_, _05895_);
  and _16490_ (_08170_, _05843_, _05870_);
  and _16491_ (_08171_, _08170_, _08093_);
  or _16492_ (_08172_, _08171_, _08139_);
  and _16493_ (_08173_, _08172_, _08169_);
  or _16494_ (_08174_, _08173_, _08168_);
  or _16495_ (_08175_, _08174_, _08167_);
  or _16496_ (_08176_, _08175_, _08163_);
  or _16497_ (_08177_, _08176_, _08151_);
  or _16498_ (_08178_, _08177_, _08144_);
  and _16499_ (_08179_, _08178_, _05731_);
  and _16500_ (_08180_, _05728_, _04859_);
  and _16501_ (_08181_, _08180_, _05957_);
  nor _16502_ (_08182_, _08181_, _05993_);
  or _16503_ (_08183_, _08182_, rst);
  or _16504_ (_05182_, _08183_, _08179_);
  and _16505_ (_08184_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and _16506_ (_08185_, _06626_, _05730_);
  or _16507_ (_08186_, _08185_, _08184_);
  or _16508_ (_08187_, _08186_, _06005_);
  and _16509_ (_05200_, _08187_, _04856_);
  and _16510_ (_08188_, _06410_, _05719_);
  and _16511_ (_08189_, _05723_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  or _16512_ (_08190_, _08189_, _08188_);
  and _16513_ (_05203_, _08190_, _04856_);
  and _16514_ (_08191_, _06721_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  or _16515_ (_08192_, _05986_, _05950_);
  and _16516_ (_08193_, _08192_, _05965_);
  or _16517_ (_08194_, _06789_, _06628_);
  or _16518_ (_08195_, _08194_, _06872_);
  or _16519_ (_08196_, _08195_, _08193_);
  or _16520_ (_08197_, _06786_, _06610_);
  and _16521_ (_08198_, _06594_, _05848_);
  or _16522_ (_08199_, _06613_, _08198_);
  or _16523_ (_08200_, _06746_, _06726_);
  or _16524_ (_08201_, _08200_, _08199_);
  or _16525_ (_08202_, _08201_, _08197_);
  or _16526_ (_08203_, _08202_, _08196_);
  and _16527_ (_08204_, _08203_, _06770_);
  or _16528_ (_05219_, _08204_, _08191_);
  and _16529_ (_08205_, _06721_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _16530_ (_08206_, _06808_, _06806_);
  not _16531_ (_08207_, _08206_);
  and _16532_ (_08208_, _06777_, _05998_);
  and _16533_ (_08209_, _06598_, _05986_);
  or _16534_ (_08210_, _08209_, _08208_);
  or _16535_ (_08211_, _08210_, _08207_);
  and _16536_ (_08212_, _06783_, _05972_);
  and _16537_ (_08213_, _06001_, _05983_);
  not _16538_ (_08214_, _06858_);
  or _16539_ (_08215_, _08214_, _08198_);
  or _16540_ (_08216_, _08215_, _08213_);
  and _16541_ (_08217_, _06855_, _06648_);
  not _16542_ (_08218_, _08217_);
  or _16543_ (_08219_, _08218_, _06614_);
  or _16544_ (_08220_, _08219_, _08216_);
  or _16545_ (_08221_, _08220_, _08212_);
  or _16546_ (_08222_, _08221_, _08211_);
  and _16547_ (_08223_, _08222_, _06770_);
  or _16548_ (_05222_, _08223_, _08205_);
  and _16549_ (_08224_, _06688_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  and _16550_ (_08225_, _06686_, _06410_);
  or _16551_ (_08226_, _08225_, _08224_);
  and _16552_ (_05251_, _08226_, _04856_);
  and _16553_ (_08228_, _05969_, _06637_);
  or _16554_ (_08229_, _08228_, _05955_);
  or _16555_ (_08231_, _06892_, _06790_);
  or _16556_ (_08232_, _08231_, _08229_);
  or _16557_ (_08233_, _06641_, _05980_);
  or _16558_ (_08235_, _08233_, _06747_);
  or _16559_ (_08236_, _08235_, _08232_);
  or _16560_ (_08237_, _08236_, _06634_);
  and _16561_ (_08238_, _08237_, _05730_);
  and _16562_ (_08239_, \oc8051_top_1.oc8051_decoder1.wr , \oc8051_top_1.oc8051_sfr1.wait_data );
  or _16563_ (_08240_, _08239_, _06650_);
  or _16564_ (_08241_, _08240_, _08238_);
  and _16565_ (_05302_, _08241_, _04856_);
  and _16566_ (_08242_, _06822_, _06731_);
  and _16567_ (_08243_, _06822_, _06637_);
  or _16568_ (_08244_, _08243_, _08242_);
  and _16569_ (_08245_, _06624_, _05965_);
  and _16570_ (_08246_, _07510_, _06000_);
  or _16571_ (_08247_, _08246_, _06833_);
  or _16572_ (_08248_, _08247_, _08245_);
  or _16573_ (_08249_, _08248_, _08244_);
  or _16574_ (_08250_, _08047_, _06862_);
  or _16575_ (_08251_, _08250_, _08249_);
  and _16576_ (_08252_, _08251_, _05730_);
  and _16577_ (_08253_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _16578_ (_08254_, _08253_, _06813_);
  or _16579_ (_08255_, _08254_, _08252_);
  and _16580_ (_05311_, _08255_, _04856_);
  and _16581_ (_05358_, _05919_, _04856_);
  nor _16582_ (_05361_, _07380_, rst);
  nor _16583_ (_08256_, _05730_, _05323_);
  not _16584_ (_08257_, _05730_);
  and _16585_ (_08258_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and _16586_ (_08259_, _05933_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and _16587_ (_08260_, _05742_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor _16588_ (_08261_, _08260_, _08259_);
  and _16589_ (_08262_, _05927_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and _16590_ (_08263_, _05935_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor _16591_ (_08264_, _08263_, _08262_);
  and _16592_ (_08265_, _05758_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  and _16593_ (_08266_, _05929_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nor _16594_ (_08267_, _08266_, _08265_);
  and _16595_ (_08268_, _08267_, _08264_);
  and _16596_ (_08269_, _08268_, _08261_);
  nor _16597_ (_08270_, _08269_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _16598_ (_08271_, _08270_, _08258_);
  nor _16599_ (_08272_, _08271_, _08257_);
  nor _16600_ (_08273_, _08272_, _08256_);
  nor _16601_ (_05364_, _08273_, rst);
  nor _16602_ (_08274_, _04948_, _04922_);
  and _16603_ (_08275_, _04932_, _05513_);
  and _16604_ (_08276_, _08275_, _08274_);
  and _16605_ (_08277_, _08276_, _06141_);
  and _16606_ (_08278_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  or _16607_ (_08280_, _08278_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and _16608_ (_08281_, _05627_, _05583_);
  and _16609_ (_08282_, _05407_, _05455_);
  nand _16610_ (_08284_, _05273_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nand _16611_ (_08285_, _08284_, _08278_);
  or _16612_ (_08286_, _08285_, _08282_);
  or _16613_ (_08287_, _08286_, _08281_);
  and _16614_ (_08288_, _08287_, _08280_);
  or _16615_ (_08289_, _08288_, _08277_);
  or _16616_ (_08290_, _06146_, _06563_);
  nand _16617_ (_08291_, _08290_, _08277_);
  or _16618_ (_08292_, _08291_, _06147_);
  and _16619_ (_08294_, _08292_, _08289_);
  or _16620_ (_08295_, _08294_, _06934_);
  nand _16621_ (_08296_, _06934_, _05287_);
  and _16622_ (_08298_, _08296_, _04856_);
  and _16623_ (_05505_, _08298_, _08295_);
  and _16624_ (_05508_, _05767_, _04856_);
  and _16625_ (_05511_, _05843_, _04856_);
  and _16626_ (_05514_, _05793_, _04856_);
  and _16627_ (_05516_, _05818_, _04856_);
  and _16628_ (_05518_, _05870_, _04856_);
  and _16629_ (_05521_, _05895_, _04856_);
  and _16630_ (_05523_, _05943_, _04856_);
  and _16631_ (_08304_, _08277_, _06091_);
  nand _16632_ (_08305_, _08304_, _06088_);
  or _16633_ (_08306_, _08304_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and _16634_ (_08308_, _08306_, _06935_);
  and _16635_ (_08309_, _08308_, _08305_);
  and _16636_ (_08310_, _06934_, _05718_);
  or _16637_ (_08311_, _08310_, _08309_);
  and _16638_ (_05539_, _08311_, _04856_);
  nand _16639_ (_08312_, _07897_, _06498_);
  not _16640_ (_08313_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  nand _16641_ (_08314_, _06497_, _08313_);
  and _16642_ (_08315_, _08314_, _04856_);
  and _16643_ (_05566_, _08315_, _08312_);
  nand _16644_ (_08316_, _07815_, _06498_);
  or _16645_ (_08317_, _06498_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and _16646_ (_08318_, _08317_, _04856_);
  and _16647_ (_05575_, _08318_, _08316_);
  or _16648_ (_08319_, _07676_, _05293_);
  or _16649_ (_08320_, _05524_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  nand _16650_ (_08321_, _07702_, _05524_);
  and _16651_ (_08322_, _08321_, _08320_);
  or _16652_ (_08323_, _08322_, _05292_);
  and _16653_ (_08324_, _08323_, _04856_);
  and _16654_ (_05691_, _08324_, _08319_);
  or _16655_ (_08325_, _07924_, _05293_);
  nor _16656_ (_08326_, _07897_, _05643_);
  not _16657_ (_08327_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  nor _16658_ (_08328_, _05524_, _08327_);
  or _16659_ (_08329_, _08328_, _05292_);
  or _16660_ (_08330_, _08329_, _08326_);
  and _16661_ (_08331_, _08330_, _04856_);
  and _16662_ (_05695_, _08331_, _08325_);
  or _16663_ (_08332_, _07853_, _05293_);
  nor _16664_ (_08333_, _07815_, _05643_);
  and _16665_ (_08334_, _05643_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or _16666_ (_08335_, _08334_, _05292_);
  or _16667_ (_08336_, _08335_, _08333_);
  and _16668_ (_08337_, _08336_, _04856_);
  and _16669_ (_05697_, _08337_, _08332_);
  or _16670_ (_08338_, _07743_, _05293_);
  nor _16671_ (_08339_, _07774_, _05643_);
  not _16672_ (_08340_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  nor _16673_ (_08341_, _05524_, _08340_);
  or _16674_ (_08342_, _08341_, _05292_);
  or _16675_ (_08343_, _08342_, _08339_);
  and _16676_ (_08344_, _08343_, _04856_);
  and _16677_ (_05706_, _08344_, _08338_);
  or _16678_ (_08345_, _07640_, _05293_);
  nor _16679_ (_08346_, _06586_, _05643_);
  not _16680_ (_08347_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  nor _16681_ (_08348_, _05524_, _08347_);
  or _16682_ (_08349_, _08348_, _05292_);
  or _16683_ (_08350_, _08349_, _08346_);
  and _16684_ (_08351_, _08350_, _04856_);
  and _16685_ (_05709_, _08351_, _08345_);
  or _16686_ (_08352_, _07598_, _05293_);
  nor _16687_ (_08353_, _06552_, _05643_);
  and _16688_ (_08354_, _05643_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or _16689_ (_08355_, _08354_, _05292_);
  or _16690_ (_08356_, _08355_, _08353_);
  and _16691_ (_08357_, _08356_, _04856_);
  and _16692_ (_05712_, _08357_, _08352_);
  nor _16693_ (_08358_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  not _16694_ (_08359_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor _16695_ (_08360_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _08359_);
  nor _16696_ (_08361_, _08360_, _08358_);
  not _16697_ (_08363_, \oc8051_symbolic_cxrom1.regvalid [13]);
  not _16698_ (_08364_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and _16699_ (_08365_, _05746_, _05736_);
  nor _16700_ (_08366_, _08365_, _08257_);
  nor _16701_ (_08367_, _08366_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  nor _16702_ (_08368_, _08367_, _08364_);
  and _16703_ (_08369_, _08368_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor _16704_ (_08370_, _08368_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor _16705_ (_08371_, _08370_, _08369_);
  nor _16706_ (_08372_, _08371_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor _16707_ (_08373_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _08359_);
  nor _16708_ (_08375_, _08373_, _08372_);
  and _16709_ (_08376_, _08375_, _08363_);
  nor _16710_ (_08377_, _08375_, \oc8051_symbolic_cxrom1.regvalid [5]);
  or _16711_ (_08378_, _08377_, _08376_);
  not _16712_ (_08380_, _08378_);
  nor _16713_ (_08381_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor _16714_ (_08382_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _08359_);
  nor _16715_ (_08383_, _08382_, _08381_);
  not _16716_ (_08385_, _08383_);
  and _16717_ (_08386_, _08367_, _08364_);
  nor _16718_ (_08387_, _08386_, _08368_);
  nor _16719_ (_08389_, _08387_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor _16720_ (_08390_, _08359_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2]);
  nor _16721_ (_08392_, _08390_, _08389_);
  and _16722_ (_08393_, _08392_, _08385_);
  nand _16723_ (_08394_, _08393_, _08380_);
  and _16724_ (_08396_, _08394_, _08361_);
  nor _16725_ (_08397_, _08392_, _08385_);
  not _16726_ (_08398_, _08397_);
  not _16727_ (_08399_, \oc8051_symbolic_cxrom1.regvalid [3]);
  nor _16728_ (_08401_, _08375_, _08399_);
  and _16729_ (_08403_, _08375_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor _16730_ (_08404_, _08403_, _08401_);
  nor _16731_ (_08405_, _08404_, _08398_);
  and _16732_ (_08406_, _08392_, _08383_);
  not _16733_ (_08407_, _08406_);
  not _16734_ (_08408_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and _16735_ (_08409_, _08375_, _08408_);
  nor _16736_ (_08410_, _08375_, \oc8051_symbolic_cxrom1.regvalid [7]);
  or _16737_ (_08411_, _08410_, _08409_);
  nor _16738_ (_08412_, _08411_, _08407_);
  nor _16739_ (_08413_, _08412_, _08405_);
  not _16740_ (_08414_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and _16741_ (_08415_, _08375_, _08414_);
  nor _16742_ (_08416_, _08392_, _08383_);
  not _16743_ (_08417_, _08416_);
  nor _16744_ (_08418_, _08375_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or _16745_ (_08419_, _08418_, _08417_);
  or _16746_ (_08420_, _08419_, _08415_);
  and _16747_ (_08421_, _08420_, _08413_);
  and _16748_ (_08422_, _08421_, _08396_);
  not _16749_ (_08423_, _08392_);
  and _16750_ (_08424_, _08375_, \oc8051_symbolic_cxrom1.regvalid [12]);
  not _16751_ (_08425_, _08375_);
  and _16752_ (_08426_, _08425_, \oc8051_symbolic_cxrom1.regvalid [4]);
  nor _16753_ (_08427_, _08426_, _08424_);
  nor _16754_ (_08428_, _08427_, _08423_);
  nor _16755_ (_08429_, _08392_, _08375_);
  and _16756_ (_08430_, _08429_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and _16757_ (_08431_, _08423_, _08375_);
  and _16758_ (_08432_, _08431_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor _16759_ (_08433_, _08432_, _08430_);
  not _16760_ (_08434_, _08433_);
  nor _16761_ (_08435_, _08434_, _08428_);
  nor _16762_ (_08436_, _08435_, _08383_);
  and _16763_ (_08437_, _08429_, _08383_);
  and _16764_ (_08438_, _08437_, \oc8051_symbolic_cxrom1.regvalid [2]);
  not _16765_ (_08439_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and _16766_ (_08440_, _08375_, _08439_);
  nor _16767_ (_08441_, _08375_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or _16768_ (_08442_, _08441_, _08440_);
  nor _16769_ (_08443_, _08442_, _08407_);
  and _16770_ (_08444_, _08375_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and _16771_ (_08445_, _08444_, _08397_);
  or _16772_ (_08446_, _08445_, _08361_);
  or _16773_ (_08447_, _08446_, _08443_);
  or _16774_ (_08448_, _08447_, _08438_);
  nor _16775_ (_08449_, _08448_, _08436_);
  nor _16776_ (_08450_, _08449_, _08422_);
  not _16777_ (_08451_, _08450_);
  and _16778_ (_08452_, _08451_, word_in[7]);
  not _16779_ (_08453_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  nand _16780_ (_08454_, _08361_, _08453_);
  or _16781_ (_08455_, _08361_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  and _16782_ (_08456_, _08455_, _08454_);
  and _16783_ (_08457_, _08456_, _08406_);
  not _16784_ (_08458_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  nand _16785_ (_08459_, _08361_, _08458_);
  or _16786_ (_08460_, _08361_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  and _16787_ (_08461_, _08460_, _08459_);
  and _16788_ (_08462_, _08461_, _08397_);
  or _16789_ (_08463_, _08462_, _08457_);
  not _16790_ (_08464_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  nand _16791_ (_08465_, _08361_, _08464_);
  or _16792_ (_08466_, _08361_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  and _16793_ (_08467_, _08466_, _08465_);
  and _16794_ (_08468_, _08467_, _08393_);
  not _16795_ (_08469_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  nand _16796_ (_08470_, _08361_, _08469_);
  or _16797_ (_08471_, _08361_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  and _16798_ (_08472_, _08471_, _08470_);
  and _16799_ (_08473_, _08472_, _08416_);
  or _16800_ (_08474_, _08473_, _08468_);
  or _16801_ (_08475_, _08474_, _08463_);
  and _16802_ (_08476_, _08475_, _08375_);
  not _16803_ (_08477_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  nand _16804_ (_08478_, _08361_, _08477_);
  or _16805_ (_08479_, _08361_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  and _16806_ (_08480_, _08479_, _08478_);
  and _16807_ (_08481_, _08480_, _08437_);
  and _16808_ (_08482_, _08406_, _08425_);
  not _16809_ (_08483_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  nand _16810_ (_08484_, _08361_, _08483_);
  or _16811_ (_08485_, _08361_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  and _16812_ (_08486_, _08485_, _08484_);
  and _16813_ (_08487_, _08486_, _08482_);
  not _16814_ (_08488_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  nand _16815_ (_08489_, _08361_, _08488_);
  or _16816_ (_08490_, _08361_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  and _16817_ (_08491_, _08490_, _08489_);
  and _16818_ (_08493_, _08491_, _08393_);
  not _16819_ (_08494_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  nand _16820_ (_08495_, _08361_, _08494_);
  or _16821_ (_08496_, _08361_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  and _16822_ (_08498_, _08496_, _08495_);
  and _16823_ (_08500_, _08498_, _08416_);
  or _16824_ (_08502_, _08500_, _08493_);
  and _16825_ (_08503_, _08502_, _08425_);
  or _16826_ (_08505_, _08503_, _08487_);
  or _16827_ (_08506_, _08505_, _08481_);
  or _16828_ (_08507_, _08506_, _08476_);
  and _16829_ (_08509_, _08507_, _08450_);
  or _16830_ (\oc8051_symbolic_cxrom1.cxrom_data_out [7], _08509_, _08452_);
  and _16831_ (_08511_, _08385_, _08361_);
  not _16832_ (_08512_, _08511_);
  and _16833_ (_08514_, _08383_, _08361_);
  nor _16834_ (_08515_, _08514_, _08392_);
  and _16835_ (_08516_, _08514_, _08392_);
  nor _16836_ (_08517_, _08516_, _08515_);
  not _16837_ (_08518_, _08517_);
  nor _16838_ (_08519_, _08518_, _08442_);
  nor _16839_ (_08520_, _08516_, _08425_);
  and _16840_ (_08521_, _08516_, _08425_);
  nor _16841_ (_08522_, _08521_, _08520_);
  nor _16842_ (_08523_, _08522_, _08517_);
  and _16843_ (_08524_, _08523_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and _16844_ (_08525_, _08522_, _08518_);
  and _16845_ (_08526_, _08525_, \oc8051_symbolic_cxrom1.regvalid [2]);
  or _16846_ (_08527_, _08526_, _08524_);
  nor _16847_ (_08528_, _08527_, _08519_);
  nor _16848_ (_08529_, _08528_, _08512_);
  not _16849_ (_08530_, _08529_);
  not _16850_ (_08531_, _08514_);
  nor _16851_ (_08532_, _08518_, _08427_);
  and _16852_ (_08533_, _08525_, \oc8051_symbolic_cxrom1.regvalid [0]);
  nor _16853_ (_08534_, _08533_, _08532_);
  or _16854_ (_08535_, _08534_, _08531_);
  nand _16855_ (_08536_, _08521_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and _16856_ (_08537_, _08536_, _08535_);
  and _16857_ (_08538_, _08537_, _08530_);
  not _16858_ (_08539_, _08361_);
  and _16859_ (_08540_, _08383_, _08539_);
  not _16860_ (_08541_, _08540_);
  nor _16861_ (_08542_, _08518_, _08411_);
  and _16862_ (_08543_, _08523_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and _16863_ (_08544_, _08525_, \oc8051_symbolic_cxrom1.regvalid [3]);
  or _16864_ (_08545_, _08544_, _08543_);
  nor _16865_ (_08546_, _08545_, _08542_);
  nor _16866_ (_08547_, _08546_, _08541_);
  nor _16867_ (_08548_, _08383_, _08361_);
  not _16868_ (_08549_, _08548_);
  nor _16869_ (_08550_, _08518_, _08378_);
  and _16870_ (_08551_, _08523_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and _16871_ (_08552_, _08525_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or _16872_ (_08553_, _08552_, _08551_);
  nor _16873_ (_08554_, _08553_, _08550_);
  nor _16874_ (_08555_, _08554_, _08549_);
  nor _16875_ (_08556_, _08555_, _08547_);
  and _16876_ (_08557_, _08556_, _08538_);
  or _16877_ (_08558_, _08514_, _08548_);
  not _16878_ (_08559_, _08558_);
  not _16879_ (_08560_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  nand _16880_ (_08561_, _08361_, _08560_);
  or _16881_ (_08563_, _08361_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  and _16882_ (_08564_, _08563_, _08561_);
  and _16883_ (_08565_, _08564_, _08559_);
  not _16884_ (_08566_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  nand _16885_ (_08567_, _08361_, _08566_);
  or _16886_ (_08568_, _08361_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  and _16887_ (_08569_, _08568_, _08567_);
  and _16888_ (_08570_, _08569_, _08558_);
  or _16889_ (_08571_, _08570_, _08565_);
  and _16890_ (_08572_, _08571_, _08523_);
  and _16891_ (_08573_, _08517_, _08375_);
  not _16892_ (_08574_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  nand _16893_ (_08575_, _08361_, _08574_);
  or _16894_ (_08576_, _08361_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  and _16895_ (_08577_, _08576_, _08575_);
  and _16896_ (_08578_, _08577_, _08559_);
  not _16897_ (_08579_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  nand _16898_ (_08580_, _08361_, _08579_);
  or _16899_ (_08581_, _08361_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  and _16900_ (_08583_, _08581_, _08580_);
  and _16901_ (_08585_, _08583_, _08558_);
  or _16902_ (_08586_, _08585_, _08578_);
  and _16903_ (_08587_, _08586_, _08573_);
  or _16904_ (_08588_, _08587_, _08572_);
  and _16905_ (_08589_, _08361_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  nor _16906_ (_08590_, _08361_, _08494_);
  or _16907_ (_08591_, _08590_, _08589_);
  and _16908_ (_08592_, _08591_, _08558_);
  not _16909_ (_08593_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  nand _16910_ (_08594_, _08361_, _08593_);
  or _16911_ (_08595_, _08361_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  and _16912_ (_08596_, _08595_, _08594_);
  and _16913_ (_08597_, _08596_, _08559_);
  or _16914_ (_08598_, _08597_, _08592_);
  and _16915_ (_08599_, _08598_, _08525_);
  and _16916_ (_08600_, _08517_, _08425_);
  not _16917_ (_08601_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  nand _16918_ (_08602_, _08361_, _08601_);
  or _16919_ (_08603_, _08361_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  and _16920_ (_08604_, _08603_, _08602_);
  and _16921_ (_08605_, _08604_, _08558_);
  not _16922_ (_08606_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  nand _16923_ (_08607_, _08361_, _08606_);
  or _16924_ (_08608_, _08361_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  and _16925_ (_08609_, _08608_, _08607_);
  and _16926_ (_08610_, _08609_, _08559_);
  or _16927_ (_08611_, _08610_, _08605_);
  and _16928_ (_08612_, _08611_, _08600_);
  or _16929_ (_08613_, _08612_, _08599_);
  nor _16930_ (_08614_, _08613_, _08588_);
  nor _16931_ (_08615_, _08614_, _08557_);
  and _16932_ (_08616_, _08557_, word_in[15]);
  or _16933_ (\oc8051_symbolic_cxrom1.cxrom_data_out [15], _08616_, _08615_);
  nor _16934_ (_08617_, _08406_, _08416_);
  and _16935_ (_08618_, _08407_, _08375_);
  or _16936_ (_08619_, _08618_, _08482_);
  nor _16937_ (_08620_, _08619_, _08617_);
  and _16938_ (_08621_, _08620_, \oc8051_symbolic_cxrom1.regvalid [2]);
  not _16939_ (_08622_, _08621_);
  not _16940_ (_08623_, _08617_);
  nor _16941_ (_08624_, _08623_, _08442_);
  and _16942_ (_08625_, _08619_, _08623_);
  and _16943_ (_08626_, _08625_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor _16944_ (_08627_, _08626_, _08624_);
  and _16945_ (_08628_, _08627_, _08622_);
  nor _16946_ (_08629_, _08628_, _08549_);
  not _16947_ (_08630_, _08629_);
  nor _16948_ (_08631_, _08623_, _08427_);
  and _16949_ (_08632_, _08620_, \oc8051_symbolic_cxrom1.regvalid [0]);
  nor _16950_ (_08633_, _08632_, _08631_);
  or _16951_ (_08634_, _08633_, _08541_);
  or _16952_ (_08635_, _08375_, _08361_);
  nor _16953_ (_08636_, _08635_, _08407_);
  nand _16954_ (_08637_, _08636_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and _16955_ (_08638_, _08637_, _08634_);
  and _16956_ (_08639_, _08638_, _08630_);
  nor _16957_ (_08640_, _08623_, _08378_);
  and _16958_ (_08641_, _08620_, \oc8051_symbolic_cxrom1.regvalid [1]);
  and _16959_ (_08642_, _08625_, \oc8051_symbolic_cxrom1.regvalid [9]);
  or _16960_ (_08643_, _08642_, _08641_);
  nor _16961_ (_08644_, _08643_, _08640_);
  nor _16962_ (_08645_, _08644_, _08531_);
  and _16963_ (_08646_, _08620_, \oc8051_symbolic_cxrom1.regvalid [3]);
  not _16964_ (_08647_, _08646_);
  nor _16965_ (_08648_, _08623_, _08411_);
  and _16966_ (_08649_, _08625_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor _16967_ (_08650_, _08649_, _08648_);
  and _16968_ (_08651_, _08650_, _08647_);
  nor _16969_ (_08652_, _08651_, _08512_);
  nor _16970_ (_08653_, _08652_, _08645_);
  and _16971_ (_08654_, _08653_, _08639_);
  and _16972_ (_08655_, _08486_, _08393_);
  and _16973_ (_08656_, _08498_, _08375_);
  or _16974_ (_08657_, _08656_, _08655_);
  and _16975_ (_08658_, _08491_, _08397_);
  and _16976_ (_08659_, _08480_, _08416_);
  or _16977_ (_08660_, _08659_, _08658_);
  nor _16978_ (_08661_, _08660_, _08657_);
  nor _16979_ (_08662_, _08661_, _08619_);
  and _16980_ (_08663_, _08467_, _08397_);
  and _16981_ (_08664_, _08461_, _08416_);
  or _16982_ (_08665_, _08664_, _08663_);
  and _16983_ (_08666_, _08456_, _08393_);
  and _16984_ (_08667_, _08472_, _08406_);
  or _16985_ (_08668_, _08667_, _08666_);
  or _16986_ (_08669_, _08668_, _08665_);
  and _16987_ (_08670_, _08669_, _08619_);
  nor _16988_ (_08671_, _08670_, _08662_);
  nor _16989_ (_08672_, _08671_, _08654_);
  and _16990_ (_08673_, _08654_, word_in[23]);
  or _16991_ (\oc8051_symbolic_cxrom1.cxrom_data_out [23], _08673_, _08672_);
  and _16992_ (_08674_, _08516_, _08375_);
  and _16993_ (_08675_, _08674_, \oc8051_symbolic_cxrom1.regvalid [2]);
  and _16994_ (_08676_, _08549_, _08392_);
  nor _16995_ (_08677_, _08549_, _08392_);
  nor _16996_ (_08678_, _08677_, _08676_);
  not _16997_ (_08679_, _08678_);
  nor _16998_ (_08680_, _08442_, _08679_);
  and _16999_ (_08681_, _08676_, _08375_);
  nor _17000_ (_08682_, _08676_, _08375_);
  nor _17001_ (_08684_, _08682_, _08681_);
  and _17002_ (_08685_, _08684_, _08679_);
  and _17003_ (_08686_, _08685_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor _17004_ (_08687_, _08686_, _08680_);
  nor _17005_ (_08688_, _08687_, _08531_);
  nor _17006_ (_08689_, _08679_, _08427_);
  nor _17007_ (_08690_, _08684_, _08678_);
  and _17008_ (_08692_, _08690_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and _17009_ (_08693_, _08685_, \oc8051_symbolic_cxrom1.regvalid [8]);
  or _17010_ (_08695_, _08693_, _08692_);
  nor _17011_ (_08696_, _08695_, _08689_);
  nor _17012_ (_08698_, _08696_, _08512_);
  or _17013_ (_08699_, _08698_, _08688_);
  nor _17014_ (_08700_, _08699_, _08675_);
  nor _17015_ (_08701_, _08679_, _08378_);
  and _17016_ (_08703_, _08685_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and _17017_ (_08704_, _08690_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or _17018_ (_08706_, _08704_, _08703_);
  nor _17019_ (_08707_, _08706_, _08701_);
  nor _17020_ (_08708_, _08707_, _08541_);
  nor _17021_ (_08710_, _08679_, _08411_);
  and _17022_ (_08711_, _08685_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor _17023_ (_08712_, _08711_, _08710_);
  nor _17024_ (_08713_, _08712_, _08549_);
  and _17025_ (_08714_, _08677_, _08401_);
  or _17026_ (_08715_, _08714_, _08713_);
  nor _17027_ (_08716_, _08715_, _08708_);
  and _17028_ (_08717_, _08716_, _08700_);
  and _17029_ (_08718_, _08569_, _08559_);
  and _17030_ (_08719_, _08564_, _08558_);
  or _17031_ (_08720_, _08719_, _08718_);
  and _17032_ (_08721_, _08720_, _08685_);
  and _17033_ (_08722_, _08591_, _08559_);
  and _17034_ (_08723_, _08596_, _08558_);
  or _17035_ (_08724_, _08723_, _08722_);
  and _17036_ (_08725_, _08724_, _08690_);
  and _17037_ (_08726_, _08678_, _08425_);
  and _17038_ (_08727_, _08604_, _08559_);
  and _17039_ (_08728_, _08609_, _08558_);
  or _17040_ (_08729_, _08728_, _08727_);
  and _17041_ (_08730_, _08729_, _08726_);
  and _17042_ (_08731_, _08678_, _08375_);
  and _17043_ (_08732_, _08583_, _08559_);
  and _17044_ (_08733_, _08577_, _08558_);
  or _17045_ (_08734_, _08733_, _08732_);
  and _17046_ (_08735_, _08734_, _08731_);
  or _17047_ (_08736_, _08735_, _08730_);
  or _17048_ (_08737_, _08736_, _08725_);
  nor _17049_ (_08738_, _08737_, _08721_);
  nor _17050_ (_08739_, _08738_, _08717_);
  and _17051_ (_08740_, _08717_, word_in[31]);
  or _17052_ (\oc8051_symbolic_cxrom1.cxrom_data_out [31], _08740_, _08739_);
  and _17053_ (_08741_, _08392_, _08375_);
  or _17054_ (_08742_, _08741_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and _17055_ (_05809_, _08742_, _04856_);
  and _17056_ (_08743_, _08717_, _04856_);
  and _17057_ (_08744_, _08743_, _08678_);
  and _17058_ (_08745_, _08744_, _08684_);
  and _17059_ (_08746_, _08745_, _08548_);
  and _17060_ (_08747_, _08654_, _04856_);
  and _17061_ (_08748_, _08747_, _08617_);
  and _17062_ (_08749_, _08748_, _08619_);
  and _17063_ (_08750_, _08749_, _08511_);
  and _17064_ (_08751_, _08557_, _04856_);
  and _17065_ (_08752_, _08751_, _08540_);
  and _17066_ (_08753_, _08752_, _08573_);
  and _17067_ (_08754_, _08422_, _04856_);
  and _17068_ (_08755_, _08754_, _08383_);
  nor _17069_ (_08756_, _08450_, rst);
  and _17070_ (_08757_, _08756_, _08741_);
  and _17071_ (_08758_, _08757_, _08755_);
  nor _17072_ (_08759_, _08758_, _08453_);
  and _17073_ (_08760_, _08756_, word_in[7]);
  and _17074_ (_08761_, _08760_, _08758_);
  or _17075_ (_08762_, _08761_, _08759_);
  or _17076_ (_08763_, _08762_, _08753_);
  not _17077_ (_08764_, word_in[15]);
  nand _17078_ (_08765_, _08753_, _08764_);
  and _17079_ (_08766_, _08765_, _08763_);
  or _17080_ (_08767_, _08766_, _08750_);
  not _17081_ (_08768_, _08750_);
  and _17082_ (_08769_, _08747_, word_in[23]);
  or _17083_ (_08770_, _08769_, _08768_);
  and _17084_ (_08771_, _08770_, _08767_);
  or _17085_ (_08772_, _08771_, _08746_);
  not _17086_ (_08773_, _08746_);
  and _17087_ (_08774_, _08743_, word_in[31]);
  or _17088_ (_08775_, _08774_, _08773_);
  and _17089_ (_13255_, _08775_, _08772_);
  or _17090_ (_08776_, _08690_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and _17091_ (_05859_, _08776_, _04856_);
  and _17092_ (_08777_, _08690_, _08540_);
  and _17093_ (_08778_, _08416_, _08425_);
  or _17094_ (_08779_, _08778_, _08674_);
  or _17095_ (_08780_, _08779_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or _17096_ (_08781_, _08780_, _08777_);
  and _17097_ (_05887_, _08781_, _04856_);
  and _17098_ (_08782_, _08726_, _08540_);
  or _17099_ (_08783_, _08782_, \oc8051_symbolic_cxrom1.regvalid [2]);
  or _17100_ (_08784_, _08779_, _08783_);
  and _17101_ (_05931_, _08784_, _04856_);
  and _17102_ (_08785_, _08037_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  not _17103_ (_08786_, _07390_);
  nand _17104_ (_08787_, _08003_, _07958_);
  not _17105_ (_08788_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or _17106_ (_08789_, _07410_, _08788_);
  not _17107_ (_08790_, _07404_);
  nand _17108_ (_08791_, _08790_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and _17109_ (_08792_, _08791_, _08789_);
  nand _17110_ (_08793_, _07422_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  not _17111_ (_08794_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or _17112_ (_08795_, _07428_, _08794_);
  and _17113_ (_08796_, _08795_, _08793_);
  and _17114_ (_08797_, _08796_, _08792_);
  nand _17115_ (_08798_, _07437_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  nand _17116_ (_08799_, _07442_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and _17117_ (_08800_, _08799_, _08798_);
  nand _17118_ (_08801_, _07449_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  nand _17119_ (_08802_, _07455_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and _17120_ (_08803_, _08802_, _08801_);
  and _17121_ (_08804_, _08803_, _08800_);
  and _17122_ (_08805_, _08804_, _08797_);
  not _17123_ (_08806_, _07463_);
  nand _17124_ (_08807_, _08806_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  not _17125_ (_08808_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  or _17126_ (_08809_, _07465_, _08808_);
  and _17127_ (_08810_, _08809_, _08807_);
  nand _17128_ (_08811_, _07470_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  not _17129_ (_08812_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or _17130_ (_08813_, _07472_, _08812_);
  and _17131_ (_08814_, _08813_, _08811_);
  and _17132_ (_08815_, _08814_, _08810_);
  not _17133_ (_08816_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  or _17134_ (_08817_, _07486_, _08816_);
  nand _17135_ (_08818_, _07484_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  and _17136_ (_08819_, _08818_, _08817_);
  nand _17137_ (_08820_, _07477_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  nand _17138_ (_08821_, _07479_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  and _17139_ (_08822_, _08821_, _08820_);
  and _17140_ (_08823_, _08822_, _08819_);
  and _17141_ (_08824_, _08823_, _08815_);
  and _17142_ (_08825_, _08824_, _08805_);
  or _17143_ (_08826_, _07503_, _07154_);
  nand _17144_ (_08827_, _07500_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and _17145_ (_08828_, _08827_, _08826_);
  or _17146_ (_08829_, _08025_, _06588_);
  or _17147_ (_08830_, _07953_, _08347_);
  and _17148_ (_08831_, _08830_, _08829_);
  and _17149_ (_08832_, _08831_, _08828_);
  nor _17150_ (_08833_, _07531_, p0_in[3]);
  not _17151_ (_08834_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and _17152_ (_08835_, _07531_, _08834_);
  nor _17153_ (_08836_, _08835_, _08833_);
  nand _17154_ (_08837_, _08836_, _07547_);
  nor _17155_ (_08838_, _07531_, p1_in[3]);
  not _17156_ (_08839_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and _17157_ (_08840_, _07531_, _08839_);
  nor _17158_ (_08841_, _08840_, _08838_);
  nand _17159_ (_08842_, _08841_, _07552_);
  and _17160_ (_08843_, _08842_, _08837_);
  nor _17161_ (_08844_, _07531_, p2_in[3]);
  not _17162_ (_08845_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and _17163_ (_08846_, _07531_, _08845_);
  nor _17164_ (_08847_, _08846_, _08844_);
  nand _17165_ (_08848_, _08847_, _07507_);
  nor _17166_ (_08849_, _07531_, p3_in[3]);
  not _17167_ (_08850_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and _17168_ (_08851_, _07531_, _08850_);
  nor _17169_ (_08852_, _08851_, _08849_);
  nand _17170_ (_08853_, _08852_, _07539_);
  and _17171_ (_08854_, _08853_, _08848_);
  and _17172_ (_08855_, _08854_, _08843_);
  and _17173_ (_08856_, _08855_, _08832_);
  nand _17174_ (_08857_, _07943_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nand _17175_ (_08858_, _07561_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and _17176_ (_08859_, _08858_, _08857_);
  and _17177_ (_08860_, _08859_, _08856_);
  and _17178_ (_08861_, _08860_, _08825_);
  or _17179_ (_08862_, _08861_, _08787_);
  nand _17180_ (_08863_, _08862_, _08786_);
  or _17181_ (_08864_, _08863_, _08785_);
  nand _17182_ (_08865_, _07390_, _06586_);
  and _17183_ (_08866_, _08865_, _04856_);
  and _17184_ (_05975_, _08866_, _08864_);
  or _17185_ (_08867_, _08429_, \oc8051_symbolic_cxrom1.regvalid [3]);
  and _17186_ (_05981_, _08867_, _04856_);
  not _17187_ (_08868_, _08429_);
  nor _17188_ (_08869_, _08423_, _08375_);
  and _17189_ (_08870_, _08869_, _08548_);
  or _17190_ (_08871_, _08870_, \oc8051_symbolic_cxrom1.regvalid [4]);
  and _17191_ (_08872_, _08871_, _08868_);
  or _17192_ (_08873_, _08512_, _08392_);
  nor _17193_ (_08874_, _08873_, _08375_);
  and _17194_ (_08875_, _08677_, _08426_);
  or _17195_ (_08876_, _08875_, _08437_);
  or _17196_ (_08877_, _08876_, _08874_);
  or _17197_ (_08878_, _08877_, _08872_);
  and _17198_ (_06031_, _08878_, _04856_);
  and _17199_ (_08880_, _08514_, _08429_);
  or _17200_ (_08882_, _08870_, _08880_);
  or _17201_ (_08883_, _08406_, _08375_);
  or _17202_ (_08884_, _08883_, _08882_);
  and _17203_ (_08885_, _08884_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and _17204_ (_08886_, _08869_, _08511_);
  and _17205_ (_08887_, _08782_, \oc8051_symbolic_cxrom1.regvalid [5]);
  or _17206_ (_08888_, _08887_, _08886_);
  nor _17207_ (_08889_, _08888_, _08885_);
  nor _17208_ (_08890_, _08889_, _08682_);
  and _17209_ (_08891_, _08778_, \oc8051_symbolic_cxrom1.regvalid [5]);
  or _17210_ (_08892_, _08891_, _08782_);
  or _17211_ (_08893_, _08892_, _08870_);
  or _17212_ (_08894_, _08893_, _08880_);
  or _17213_ (_08895_, _08894_, _08890_);
  and _17214_ (_06085_, _08895_, _04856_);
  and _17215_ (_08896_, _08037_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  and _17216_ (_08897_, _08790_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  not _17217_ (_08898_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  nor _17218_ (_08899_, _07410_, _08898_);
  or _17219_ (_08900_, _08899_, _08897_);
  not _17220_ (_08901_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  nor _17221_ (_08902_, _07428_, _08901_);
  and _17222_ (_08903_, _07422_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  or _17223_ (_08904_, _08903_, _08902_);
  or _17224_ (_08905_, _08904_, _08900_);
  and _17225_ (_08906_, _07437_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and _17226_ (_08907_, _07442_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  or _17227_ (_08908_, _08907_, _08906_);
  and _17228_ (_08909_, _07449_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and _17229_ (_08910_, _07455_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or _17230_ (_08911_, _08910_, _08909_);
  or _17231_ (_08912_, _08911_, _08908_);
  or _17232_ (_08913_, _08912_, _08905_);
  and _17233_ (_08914_, _08806_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and _17234_ (_08915_, _07466_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  or _17235_ (_08916_, _08915_, _08914_);
  and _17236_ (_08917_, _07470_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  and _17237_ (_08918_, _07473_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  or _17238_ (_08919_, _08918_, _08917_);
  or _17239_ (_08920_, _08919_, _08916_);
  and _17240_ (_08921_, _07484_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  not _17241_ (_08922_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  nor _17242_ (_08923_, _07486_, _08922_);
  or _17243_ (_08924_, _08923_, _08921_);
  and _17244_ (_08925_, _07477_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _17245_ (_08926_, _07479_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  or _17246_ (_08927_, _08926_, _08925_);
  or _17247_ (_08928_, _08927_, _08924_);
  or _17248_ (_08929_, _08928_, _08920_);
  or _17249_ (_08930_, _08929_, _08913_);
  and _17250_ (_08931_, _07500_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and _17251_ (_08932_, _08028_, _07102_);
  or _17252_ (_08933_, _08932_, _08931_);
  and _17253_ (_08934_, _07494_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  and _17254_ (_08935_, _07389_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  or _17255_ (_08936_, _08935_, _08934_);
  or _17256_ (_08937_, _08936_, _08933_);
  or _17257_ (_08938_, _07531_, p1_in[2]);
  or _17258_ (_08939_, _07533_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and _17259_ (_08940_, _08939_, _08938_);
  and _17260_ (_08941_, _08940_, _07552_);
  or _17261_ (_08942_, _07531_, p0_in[2]);
  or _17262_ (_08943_, _07533_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and _17263_ (_08944_, _08943_, _08942_);
  and _17264_ (_08945_, _08944_, _07547_);
  or _17265_ (_08946_, _08945_, _08941_);
  or _17266_ (_08947_, _07531_, p3_in[2]);
  or _17267_ (_08948_, _07533_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and _17268_ (_08949_, _08948_, _08947_);
  and _17269_ (_08950_, _08949_, _07539_);
  or _17270_ (_08951_, _07531_, p2_in[2]);
  or _17271_ (_08952_, _07533_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and _17272_ (_08953_, _08952_, _08951_);
  and _17273_ (_08954_, _08953_, _07507_);
  or _17274_ (_08955_, _08954_, _08950_);
  or _17275_ (_08956_, _08955_, _08946_);
  or _17276_ (_08957_, _08956_, _08937_);
  and _17277_ (_08958_, _07943_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and _17278_ (_08959_, _07561_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or _17279_ (_08960_, _08959_, _08958_);
  or _17280_ (_08961_, _08960_, _08957_);
  or _17281_ (_08962_, _08961_, _08930_);
  and _17282_ (_08963_, _08962_, _08004_);
  or _17283_ (_08964_, _08963_, _07390_);
  or _17284_ (_08965_, _08964_, _08896_);
  nand _17285_ (_08966_, _07390_, _06552_);
  and _17286_ (_08967_, _08966_, _04856_);
  and _17287_ (_06111_, _08967_, _08965_);
  and _17288_ (_08968_, _08676_, _08425_);
  or _17289_ (_08969_, _08520_, _08968_);
  and _17290_ (_08970_, _08868_, \oc8051_symbolic_cxrom1.regvalid [6]);
  and _17291_ (_08971_, _08970_, _08635_);
  or _17292_ (_08972_, _08971_, _08636_);
  and _17293_ (_08973_, _08972_, _08883_);
  and _17294_ (_08974_, _08882_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or _17295_ (_08975_, _08974_, _08886_);
  or _17296_ (_08976_, _08975_, _08973_);
  and _17297_ (_08977_, _08976_, _08969_);
  or _17298_ (_08978_, _08974_, _08972_);
  and _17299_ (_08979_, _08978_, _08674_);
  and _17300_ (_08980_, _08782_, \oc8051_symbolic_cxrom1.regvalid [6]);
  and _17301_ (_08981_, _08778_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or _17302_ (_08982_, _08981_, _08880_);
  or _17303_ (_08983_, _08982_, _08980_);
  or _17304_ (_08984_, _08983_, _08870_);
  or _17305_ (_08985_, _08984_, _08979_);
  or _17306_ (_08986_, _08985_, _08977_);
  and _17307_ (_06158_, _08986_, _04856_);
  and _17308_ (_08987_, _06668_, _06132_);
  and _17309_ (_08988_, _08987_, _04922_);
  and _17310_ (_08989_, _08988_, _06268_);
  nand _17311_ (_08990_, _08989_, _06088_);
  or _17312_ (_08991_, _08989_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and _17313_ (_08992_, _08991_, _06093_);
  and _17314_ (_08993_, _08992_, _08990_);
  and _17315_ (_08994_, _05517_, _05001_);
  nand _17316_ (_08995_, _08994_, _06284_);
  or _17317_ (_08996_, _08994_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and _17318_ (_08997_, _08996_, _05510_);
  and _17319_ (_08998_, _08997_, _08995_);
  not _17320_ (_08999_, _06092_);
  and _17321_ (_09000_, _08999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  or _17322_ (_09001_, _09000_, rst);
  or _17323_ (_09002_, _09001_, _08998_);
  or _17324_ (_06167_, _09002_, _08993_);
  or _17325_ (_09003_, _08516_, _08375_);
  and _17326_ (_09004_, _08429_, \oc8051_symbolic_cxrom1.regvalid [7]);
  or _17327_ (_09005_, _08636_, _08375_);
  and _17328_ (_09006_, _09005_, \oc8051_symbolic_cxrom1.regvalid [7]);
  and _17329_ (_09007_, _08385_, \oc8051_symbolic_cxrom1.regvalid [7]);
  and _17330_ (_09008_, _09007_, _08869_);
  or _17331_ (_09009_, _09008_, _08521_);
  or _17332_ (_09010_, _09009_, _09006_);
  or _17333_ (_09011_, _09010_, _09004_);
  and _17334_ (_09012_, _09011_, _09003_);
  or _17335_ (_09013_, _09004_, _08870_);
  or _17336_ (_09014_, _09013_, _08886_);
  or _17337_ (_09015_, _09014_, _08636_);
  or _17338_ (_09016_, _09015_, _09012_);
  and _17339_ (_06239_, _09016_, _04856_);
  and _17340_ (_09017_, _08987_, _06930_);
  and _17341_ (_09018_, _09017_, _06268_);
  nand _17342_ (_09019_, _09018_, _06088_);
  or _17343_ (_09020_, _09018_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and _17344_ (_09021_, _09020_, _06093_);
  and _17345_ (_09022_, _09021_, _09019_);
  and _17346_ (_09023_, _05515_, _04934_);
  and _17347_ (_09024_, _09023_, _05001_);
  nand _17348_ (_09025_, _09024_, _06284_);
  or _17349_ (_09026_, _09024_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and _17350_ (_09027_, _09026_, _05510_);
  and _17351_ (_09028_, _09027_, _09025_);
  and _17352_ (_09029_, _08999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  or _17353_ (_09030_, _09029_, rst);
  or _17354_ (_09031_, _09030_, _09028_);
  or _17355_ (_06247_, _09031_, _09022_);
  nor _17356_ (_09032_, _08726_, _08685_);
  and _17357_ (_09033_, _09032_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and _17358_ (_09034_, _08559_, _08869_);
  and _17359_ (_09035_, _09034_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and _17360_ (_09037_, _08677_, _08375_);
  and _17361_ (_09038_, _08726_, \oc8051_symbolic_cxrom1.regvalid [8]);
  or _17362_ (_09039_, _09038_, _09037_);
  or _17363_ (_09040_, _09039_, _09035_);
  or _17364_ (_09041_, _09040_, _09033_);
  and _17365_ (_09042_, _09041_, _08375_);
  and _17366_ (_09043_, _08429_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and _17367_ (_09044_, _08870_, \oc8051_symbolic_cxrom1.regvalid [8]);
  or _17368_ (_09045_, _08886_, _08521_);
  or _17369_ (_09046_, _09045_, _09044_);
  or _17370_ (_09047_, _09046_, _09043_);
  or _17371_ (_09048_, _09047_, _08636_);
  or _17372_ (_09049_, _09048_, _09042_);
  and _17373_ (_06315_, _09049_, _04856_);
  not _17374_ (_09050_, _08677_);
  and _17375_ (_09051_, _08520_, _09050_);
  or _17376_ (_09052_, _09051_, _08674_);
  nor _17377_ (_09053_, _08873_, _08425_);
  and _17378_ (_09054_, _08883_, \oc8051_symbolic_cxrom1.regvalid [9]);
  or _17379_ (_09055_, _09054_, _09053_);
  and _17380_ (_09056_, _09055_, _09052_);
  or _17381_ (_09057_, _08886_, _08726_);
  and _17382_ (_09058_, _09057_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor _17383_ (_09059_, _08635_, _08417_);
  and _17384_ (_09060_, _09059_, \oc8051_symbolic_cxrom1.regvalid [9]);
  or _17385_ (_09061_, _09060_, _08636_);
  or _17386_ (_09062_, _09061_, _09058_);
  or _17387_ (_09063_, _09062_, _08521_);
  or _17388_ (_09064_, _09063_, _09037_);
  or _17389_ (_09065_, _09064_, _09056_);
  and _17390_ (_06394_, _09065_, _04856_);
  and _17391_ (_09066_, _06612_, _06731_);
  or _17392_ (_09067_, _08208_, _09066_);
  and _17393_ (_09068_, _06773_, _05998_);
  or _17394_ (_09069_, _09068_, _06002_);
  or _17395_ (_09070_, _06594_, _05949_);
  and _17396_ (_09071_, _09070_, _05998_);
  or _17397_ (_09072_, _09071_, _09069_);
  or _17398_ (_09074_, _09072_, _09067_);
  and _17399_ (_09075_, _06857_, _06731_);
  or _17400_ (_09076_, _09075_, _05999_);
  or _17401_ (_09077_, _09076_, _06783_);
  and _17402_ (_09078_, _07510_, _06619_);
  or _17403_ (_09079_, _09078_, _08243_);
  or _17404_ (_09080_, _09079_, _07508_);
  or _17405_ (_09081_, _09080_, _09077_);
  and _17406_ (_09082_, _06635_, _05849_);
  and _17407_ (_09083_, _06597_, _05998_);
  or _17408_ (_09084_, _09083_, _09082_);
  or _17409_ (_09085_, _09084_, _08245_);
  or _17410_ (_09086_, _06759_, _06751_);
  or _17411_ (_09087_, _09086_, _08250_);
  and _17412_ (_09088_, _06737_, _06598_);
  and _17413_ (_09089_, _06737_, _05998_);
  or _17414_ (_09090_, _09089_, _09088_);
  and _17415_ (_09091_, _06773_, _06606_);
  and _17416_ (_09092_, _06620_, _05998_);
  or _17417_ (_09093_, _09092_, _09091_);
  or _17418_ (_09094_, _09093_, _09090_);
  or _17419_ (_09095_, _09094_, _09087_);
  or _17420_ (_09096_, _09095_, _09085_);
  and _17421_ (_09097_, _08242_, _05972_);
  or _17422_ (_09098_, _09097_, _05970_);
  or _17423_ (_09099_, _08247_, _07513_);
  or _17424_ (_09100_, _09099_, _09098_);
  or _17425_ (_09101_, _09100_, _08229_);
  or _17426_ (_09102_, _09101_, _05951_);
  or _17427_ (_09103_, _09102_, _09096_);
  or _17428_ (_09104_, _09103_, _09081_);
  or _17429_ (_09105_, _09104_, _09074_);
  and _17430_ (_09106_, _09105_, _05730_);
  and _17431_ (_09107_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _17432_ (_09108_, _06003_, _05962_);
  not _17433_ (_09109_, _06783_);
  nand _17434_ (_09110_, _09109_, _06780_);
  and _17435_ (_09111_, _09110_, _05995_);
  or _17436_ (_09112_, _09111_, _09108_);
  or _17437_ (_09113_, _09112_, _09107_);
  or _17438_ (_09114_, _09113_, _09106_);
  and _17439_ (_06447_, _09114_, _04856_);
  and _17440_ (_06465_, _07612_, _04856_);
  and _17441_ (_09115_, _05515_, _04947_);
  and _17442_ (_09116_, _09115_, _06302_);
  and _17443_ (_09117_, _09116_, _06268_);
  or _17444_ (_09118_, _09117_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and _17445_ (_09119_, _09118_, _06093_);
  nand _17446_ (_09120_, _09117_, _06088_);
  and _17447_ (_09121_, _09120_, _09119_);
  and _17448_ (_09122_, _06302_, _05001_);
  and _17449_ (_09123_, _09122_, _05515_);
  not _17450_ (_09124_, _09123_);
  nor _17451_ (_09125_, _09124_, _06284_);
  and _17452_ (_09126_, _09124_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or _17453_ (_09127_, _09126_, _09125_);
  and _17454_ (_09128_, _09127_, _05510_);
  and _17455_ (_09129_, _08999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or _17456_ (_09130_, _09129_, rst);
  or _17457_ (_09131_, _09130_, _09128_);
  or _17458_ (_06467_, _09131_, _09121_);
  and _17459_ (_09132_, _09115_, _06273_);
  and _17460_ (_09133_, _09132_, _06268_);
  nand _17461_ (_09134_, _09133_, _06088_);
  or _17462_ (_09135_, _09133_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and _17463_ (_09136_, _09135_, _06093_);
  and _17464_ (_09137_, _09136_, _09134_);
  and _17465_ (_09138_, _06274_, _05001_);
  not _17466_ (_09139_, _09138_);
  nor _17467_ (_09140_, _09139_, _06284_);
  and _17468_ (_09141_, _09139_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or _17469_ (_09142_, _09141_, _09140_);
  and _17470_ (_09143_, _09142_, _05510_);
  and _17471_ (_09144_, _08999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or _17472_ (_09145_, _09144_, rst);
  or _17473_ (_09146_, _09145_, _09143_);
  or _17474_ (_06472_, _09146_, _09137_);
  and _17475_ (_09147_, _08540_, _08731_);
  not _17476_ (_09148_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor _17477_ (_09149_, _08558_, _09148_);
  and _17478_ (_09150_, _09149_, _08726_);
  or _17479_ (_09151_, _09150_, _09147_);
  and _17480_ (_09152_, _08600_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nand _17481_ (_09153_, _08515_, _08873_);
  and _17482_ (_09154_, _09153_, _08444_);
  or _17483_ (_09155_, _09154_, _09152_);
  or _17484_ (_09156_, _09155_, _09151_);
  or _17485_ (_09157_, _08521_, _09037_);
  and _17486_ (_09158_, _09157_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and _17487_ (_09159_, _09059_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or _17488_ (_09160_, _09159_, _09158_);
  or _17489_ (_09161_, _09160_, _09156_);
  and _17490_ (_09162_, _08520_, _08417_);
  and _17491_ (_09164_, _09162_, _09161_);
  or _17492_ (_09165_, _09158_, _09053_);
  or _17493_ (_09166_, _09165_, _09164_);
  and _17494_ (_09167_, _09166_, _09051_);
  and _17495_ (_09168_, _09161_, _08674_);
  and _17496_ (_09169_, _08617_, _08425_);
  and _17497_ (_09170_, _09169_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and _17498_ (_09171_, _08636_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and _17499_ (_09172_, _08778_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or _17500_ (_09173_, _09172_, _08521_);
  or _17501_ (_09174_, _09173_, _09171_);
  or _17502_ (_09175_, _09174_, _09037_);
  or _17503_ (_09176_, _09175_, _09170_);
  or _17504_ (_09177_, _09176_, _09168_);
  or _17505_ (_09178_, _09177_, _09167_);
  and _17506_ (_06484_, _09178_, _04856_);
  and _17507_ (_09179_, _08514_, _08731_);
  and _17508_ (_09180_, _08741_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or _17509_ (_09181_, _09180_, _09179_);
  and _17510_ (_09182_, _08559_, _08429_);
  or _17511_ (_09183_, _09059_, _08521_);
  or _17512_ (_09184_, _09183_, _09182_);
  and _17513_ (_09185_, _09184_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and _17514_ (_09186_, _08600_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or _17515_ (_09187_, _09186_, _09037_);
  or _17516_ (_09188_, _09187_, _09147_);
  or _17517_ (_09189_, _09188_, _09185_);
  or _17518_ (_09190_, _09189_, _09181_);
  or _17519_ (_09191_, _09190_, _09053_);
  and _17520_ (_06577_, _09191_, _04856_);
  not _17521_ (_09193_, \oc8051_symbolic_cxrom1.regvalid [12]);
  nor _17522_ (_09194_, _09052_, _09193_);
  and _17523_ (_09195_, _08681_, \oc8051_symbolic_cxrom1.regvalid [12]);
  or _17524_ (_09196_, _09195_, _08731_);
  or _17525_ (_09197_, _09196_, _09194_);
  and _17526_ (_06683_, _09197_, _04856_);
  and _17527_ (_09198_, _08619_, _08617_);
  or _17528_ (_09199_, _09198_, \oc8051_symbolic_cxrom1.regvalid [13]);
  and _17529_ (_06785_, _09199_, _04856_);
  and _17530_ (_09200_, _06301_, _05517_);
  or _17531_ (_09201_, _09200_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  and _17532_ (_09202_, _09201_, _04856_);
  not _17533_ (_09203_, _09200_);
  or _17534_ (_09204_, _09203_, _06705_);
  and _17535_ (_06874_, _09204_, _09202_);
  and _17536_ (_09205_, _05510_, _04987_);
  and _17537_ (_09206_, _09205_, _09023_);
  and _17538_ (_09207_, _09206_, _08060_);
  and _17539_ (_09208_, _09207_, _06410_);
  and _17540_ (_09209_, \oc8051_top_1.oc8051_sfr1.pres_ow , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  and _17541_ (_09210_, _09209_, _08060_);
  and _17542_ (_09211_, _08070_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr );
  and _17543_ (_09212_, _09211_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  nor _17544_ (_09213_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  nor _17545_ (_09214_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  and _17546_ (_09215_, _09214_, _09213_);
  and _17547_ (_09216_, _09215_, _09212_);
  nor _17548_ (_09217_, _09216_, _09210_);
  not _17549_ (_09218_, _09217_);
  and _17550_ (_09219_, _09218_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  and _17551_ (_09220_, _09217_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  nor _17552_ (_09221_, _09220_, _09219_);
  nor _17553_ (_09222_, _09221_, _09206_);
  and _17554_ (_09223_, _09206_, _08070_);
  and _17555_ (_09224_, _09223_, _05670_);
  or _17556_ (_09225_, _09224_, _09222_);
  or _17557_ (_09226_, _09225_, _09208_);
  and _17558_ (_06881_, _09226_, _04856_);
  and _17559_ (_09227_, _09218_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  nor _17560_ (_09228_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  nor _17561_ (_09229_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  and _17562_ (_09230_, _09229_, _09228_);
  nor _17563_ (_09231_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  nor _17564_ (_09232_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  nor _17565_ (_09233_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  and _17566_ (_09234_, _09233_, _09232_);
  and _17567_ (_09235_, _09234_, _09231_);
  and _17568_ (_09236_, _09235_, _09230_);
  and _17569_ (_09237_, _09236_, _09210_);
  or _17570_ (_09238_, _09237_, _09217_);
  and _17571_ (_09239_, _09238_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  nor _17572_ (_09240_, _09239_, _09227_);
  nor _17573_ (_09241_, _09240_, _09206_);
  nor _17574_ (_09242_, _08070_, _06369_);
  and _17575_ (_09243_, _09242_, _09206_);
  or _17576_ (_09244_, _09243_, _09241_);
  and _17577_ (_06884_, _09244_, _04856_);
  or _17578_ (_09245_, _08573_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and _17579_ (_06896_, _09245_, _04856_);
  and _17580_ (_09246_, _05719_, _05288_);
  and _17581_ (_09247_, _05723_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  or _17582_ (_09248_, _09247_, _09246_);
  and _17583_ (_06909_, _09248_, _04856_);
  not _17584_ (_09249_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor _17585_ (_09250_, _08072_, _08062_);
  or _17586_ (_09251_, _09250_, _09249_);
  and _17587_ (_09252_, _09251_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  and _17588_ (_09253_, _08062_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and _17589_ (_09254_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  nor _17590_ (_09255_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  nor _17591_ (_09256_, _09255_, _09254_);
  and _17592_ (_09257_, _09256_, _09253_);
  or _17593_ (_09258_, _09257_, _09252_);
  and _17594_ (_06914_, _09258_, _04856_);
  and _17595_ (_09259_, _06296_, _06132_);
  and _17596_ (_09260_, _09259_, _06146_);
  nand _17597_ (_09261_, _09260_, _06088_);
  or _17598_ (_09262_, _09260_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  and _17599_ (_09263_, _09023_, _06126_);
  not _17600_ (_09264_, _09263_);
  and _17601_ (_09265_, _09264_, _09262_);
  and _17602_ (_09266_, _09265_, _09261_);
  nor _17603_ (_09267_, _09264_, _05287_);
  or _17604_ (_09268_, _09267_, _09266_);
  and _17605_ (_06927_, _09268_, _04856_);
  or _17606_ (_09269_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  or _17607_ (_09270_, _09269_, _09259_);
  not _17608_ (_09271_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  or _17609_ (_09272_, _04986_, _09271_);
  nand _17610_ (_09273_, _09272_, _09259_);
  or _17611_ (_09274_, _09273_, _07713_);
  and _17612_ (_09275_, _09274_, _09270_);
  or _17613_ (_09276_, _09275_, _09263_);
  nand _17614_ (_09277_, _09263_, _06032_);
  and _17615_ (_09278_, _09277_, _04856_);
  and _17616_ (_06933_, _09278_, _09276_);
  or _17617_ (_09279_, _09200_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  and _17618_ (_09280_, _09279_, _04856_);
  nand _17619_ (_09281_, _09200_, _05669_);
  and _17620_ (_06939_, _09281_, _09280_);
  not _17621_ (_09282_, _06284_);
  and _17622_ (_09283_, _09207_, _09282_);
  and _17623_ (_09284_, _09218_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  and _17624_ (_09285_, _09217_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  nor _17625_ (_09286_, _09285_, _09284_);
  nor _17626_ (_09287_, _09286_, _09206_);
  and _17627_ (_09288_, _09223_, _05288_);
  or _17628_ (_09289_, _09288_, _09287_);
  or _17629_ (_09290_, _09289_, _09283_);
  and _17630_ (_06942_, _09290_, _04856_);
  nand _17631_ (_09291_, _09223_, _06369_);
  nand _17632_ (_09292_, _09207_, _06032_);
  and _17633_ (_09293_, _09218_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  and _17634_ (_09294_, _09217_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  or _17635_ (_09295_, _09294_, _09293_);
  or _17636_ (_09296_, _09295_, _09206_);
  and _17637_ (_09297_, _09296_, _04856_);
  and _17638_ (_09298_, _09297_, _09292_);
  and _17639_ (_06945_, _09298_, _09291_);
  and _17640_ (_09299_, _08057_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  and _17641_ (_09300_, _08085_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  or _17642_ (_06954_, _09300_, _09299_);
  or _17643_ (_09301_, _09218_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  or _17644_ (_09302_, _09217_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  and _17645_ (_09303_, _09302_, _09301_);
  or _17646_ (_09304_, _09303_, _09206_);
  and _17647_ (_09305_, _09304_, _04856_);
  nand _17648_ (_09306_, _09223_, _06284_);
  and _17649_ (_06975_, _09306_, _09305_);
  or _17650_ (_09307_, _06607_, _05999_);
  or _17651_ (_09308_, _06636_, _06599_);
  or _17652_ (_09309_, _09308_, _09307_);
  and _17653_ (_09310_, _08228_, _05976_);
  or _17654_ (_09311_, _09310_, _08245_);
  or _17655_ (_09312_, _09088_, _06621_);
  or _17656_ (_09313_, _09312_, _09311_);
  or _17657_ (_09314_, _09313_, _09309_);
  and _17658_ (_09315_, _06772_, _06831_);
  and _17659_ (_09316_, _06598_, _06624_);
  or _17660_ (_09317_, _06787_, _09316_);
  or _17661_ (_09319_, _09317_, _09315_);
  or _17662_ (_09320_, _09319_, _09099_);
  or _17663_ (_09321_, _09079_, _06869_);
  or _17664_ (_09322_, _09321_, _09087_);
  or _17665_ (_09323_, _09322_, _09320_);
  or _17666_ (_09324_, _09323_, _09314_);
  or _17667_ (_09325_, _09324_, _09074_);
  and _17668_ (_09326_, _09325_, _05730_);
  and _17669_ (_09327_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _17670_ (_09328_, _09327_, _09112_);
  or _17671_ (_09329_, _09328_, _09326_);
  and _17672_ (_07107_, _09329_, _04856_);
  and _17673_ (_09330_, _08751_, _08674_);
  not _17674_ (_09331_, _09330_);
  not _17675_ (_09332_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  and _17676_ (_09333_, _08756_, _08383_);
  not _17677_ (_09334_, _09333_);
  not _17678_ (_09335_, _08754_);
  and _17679_ (_09336_, _08756_, _09335_);
  and _17680_ (_09337_, _09336_, _09334_);
  and _17681_ (_09338_, _09337_, _08429_);
  nor _17682_ (_09339_, _09338_, _09332_);
  and _17683_ (_09340_, _09338_, word_in[0]);
  or _17684_ (_09341_, _09340_, _09339_);
  and _17685_ (_09342_, _09341_, _09331_);
  and _17686_ (_09343_, _09330_, word_in[8]);
  or _17687_ (_09344_, _09343_, _09342_);
  nand _17688_ (_09345_, _08747_, _08777_);
  and _17689_ (_09346_, _09345_, _09344_);
  and _17690_ (_09347_, _08511_, _08741_);
  and _17691_ (_09348_, _09347_, _08743_);
  and _17692_ (_09349_, _08747_, word_in[16]);
  and _17693_ (_09350_, _09349_, _08777_);
  or _17694_ (_09351_, _09350_, _09348_);
  or _17695_ (_09352_, _09351_, _09346_);
  not _17696_ (_09353_, _09348_);
  or _17697_ (_09354_, _09353_, word_in[24]);
  and _17698_ (_07298_, _09354_, _09352_);
  not _17699_ (_09355_, _09338_);
  or _17700_ (_09356_, _09355_, word_in[1]);
  or _17701_ (_09357_, _09338_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  and _17702_ (_09358_, _09357_, _09331_);
  and _17703_ (_09359_, _09358_, _09356_);
  and _17704_ (_09360_, _09330_, word_in[9]);
  nor _17705_ (_09361_, _09360_, _09359_);
  nand _17706_ (_09362_, _09361_, _09345_);
  or _17707_ (_09363_, _09345_, word_in[17]);
  and _17708_ (_09364_, _09363_, _09353_);
  and _17709_ (_09365_, _09364_, _09362_);
  and _17710_ (_09366_, _08743_, word_in[25]);
  and _17711_ (_09367_, _09366_, _09348_);
  or _17712_ (_07302_, _09367_, _09365_);
  and _17713_ (_09368_, _08743_, word_in[26]);
  and _17714_ (_09369_, _09368_, _09348_);
  or _17715_ (_09370_, _09355_, word_in[2]);
  or _17716_ (_09371_, _09338_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  and _17717_ (_09372_, _09371_, _09331_);
  and _17718_ (_09373_, _09372_, _09370_);
  and _17719_ (_09374_, _09330_, word_in[10]);
  nor _17720_ (_09375_, _09374_, _09373_);
  nand _17721_ (_09376_, _09375_, _09345_);
  or _17722_ (_09377_, _09345_, word_in[18]);
  and _17723_ (_09378_, _09377_, _09353_);
  and _17724_ (_09379_, _09378_, _09376_);
  or _17725_ (_07307_, _09379_, _09369_);
  and _17726_ (_09380_, _08743_, word_in[27]);
  and _17727_ (_09381_, _09380_, _09348_);
  or _17728_ (_09382_, _09355_, word_in[3]);
  or _17729_ (_09383_, _09338_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  and _17730_ (_09384_, _09383_, _09331_);
  and _17731_ (_09385_, _09384_, _09382_);
  and _17732_ (_09386_, _09330_, word_in[11]);
  nor _17733_ (_09387_, _09386_, _09385_);
  nand _17734_ (_09388_, _09387_, _09345_);
  or _17735_ (_09389_, _09345_, word_in[19]);
  and _17736_ (_09390_, _09389_, _09353_);
  and _17737_ (_09391_, _09390_, _09388_);
  or _17738_ (_07313_, _09391_, _09381_);
  or _17739_ (_09392_, _09355_, word_in[4]);
  or _17740_ (_09393_, _09338_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  and _17741_ (_09394_, _09393_, _09331_);
  and _17742_ (_09395_, _09394_, _09392_);
  and _17743_ (_09396_, _09330_, word_in[12]);
  nor _17744_ (_09397_, _09396_, _09395_);
  nand _17745_ (_09398_, _09397_, _09345_);
  or _17746_ (_09399_, _09345_, word_in[20]);
  and _17747_ (_09400_, _09399_, _09353_);
  and _17748_ (_09401_, _09400_, _09398_);
  and _17749_ (_09402_, _08743_, word_in[28]);
  and _17750_ (_09403_, _09402_, _09348_);
  or _17751_ (_07318_, _09403_, _09401_);
  or _17752_ (_09404_, _09355_, word_in[5]);
  or _17753_ (_09405_, _09338_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  and _17754_ (_09406_, _09405_, _09331_);
  and _17755_ (_09407_, _09406_, _09404_);
  and _17756_ (_09408_, _09330_, word_in[13]);
  nor _17757_ (_09409_, _09408_, _09407_);
  nand _17758_ (_09410_, _09409_, _09345_);
  or _17759_ (_09411_, _09345_, word_in[21]);
  and _17760_ (_09412_, _09411_, _09353_);
  and _17761_ (_09413_, _09412_, _09410_);
  and _17762_ (_09414_, _08743_, word_in[29]);
  and _17763_ (_09415_, _09414_, _09348_);
  or _17764_ (_07324_, _09415_, _09413_);
  or _17765_ (_09416_, _09355_, word_in[6]);
  or _17766_ (_09417_, _09338_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  and _17767_ (_09418_, _09417_, _09331_);
  and _17768_ (_09419_, _09418_, _09416_);
  and _17769_ (_09420_, _09330_, word_in[14]);
  nor _17770_ (_09421_, _09420_, _09419_);
  nand _17771_ (_09422_, _09421_, _09345_);
  or _17772_ (_09423_, _09345_, word_in[22]);
  and _17773_ (_09424_, _09423_, _09353_);
  and _17774_ (_09425_, _09424_, _09422_);
  and _17775_ (_09426_, _08743_, word_in[30]);
  and _17776_ (_09427_, _09426_, _09348_);
  or _17777_ (_07329_, _09427_, _09425_);
  and _17778_ (_09428_, _09348_, word_in[31]);
  or _17779_ (_09429_, _09355_, word_in[7]);
  or _17780_ (_09430_, _09338_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  and _17781_ (_09431_, _09430_, _09331_);
  and _17782_ (_09432_, _09431_, _09429_);
  and _17783_ (_09433_, _09330_, word_in[15]);
  nor _17784_ (_09434_, _09433_, _09432_);
  nand _17785_ (_09435_, _09434_, _09345_);
  or _17786_ (_09436_, _09345_, word_in[23]);
  and _17787_ (_09437_, _09436_, _09353_);
  and _17788_ (_09438_, _09437_, _09435_);
  or _17789_ (_07332_, _09438_, _09428_);
  and _17790_ (_09439_, _08747_, _08514_);
  and _17791_ (_09440_, _09439_, _08620_);
  and _17792_ (_09441_, _08751_, _08548_);
  and _17793_ (_09442_, _09441_, _08525_);
  not _17794_ (_09443_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  and _17795_ (_09444_, _08756_, _08868_);
  and _17796_ (_09445_, _08754_, _08385_);
  not _17797_ (_09446_, _09445_);
  nor _17798_ (_09447_, _09446_, _09444_);
  nor _17799_ (_09448_, _09447_, _09443_);
  and _17800_ (_09449_, _08756_, word_in[0]);
  and _17801_ (_09450_, _09447_, _09449_);
  or _17802_ (_09451_, _09450_, _09448_);
  or _17803_ (_09452_, _09451_, _09442_);
  not _17804_ (_09453_, _09442_);
  or _17805_ (_09454_, _09453_, word_in[8]);
  and _17806_ (_09455_, _09454_, _09452_);
  or _17807_ (_09456_, _09455_, _09440_);
  and _17808_ (_09457_, _08743_, _08777_);
  not _17809_ (_09458_, _09457_);
  not _17810_ (_09459_, _09440_);
  or _17811_ (_09460_, _09459_, _09349_);
  and _17812_ (_09461_, _09460_, _09458_);
  and _17813_ (_09462_, _09461_, _09456_);
  and _17814_ (_09463_, _09457_, word_in[24]);
  or _17815_ (_07413_, _09463_, _09462_);
  and _17816_ (_09464_, _08747_, word_in[17]);
  and _17817_ (_09465_, _09440_, _09464_);
  and _17818_ (_09466_, _08756_, word_in[1]);
  and _17819_ (_09467_, _09447_, _09466_);
  not _17820_ (_09468_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  nor _17821_ (_09469_, _09447_, _09468_);
  nor _17822_ (_09470_, _09469_, _09467_);
  nor _17823_ (_09471_, _09470_, _09442_);
  and _17824_ (_09472_, _09442_, word_in[9]);
  or _17825_ (_09473_, _09472_, _09471_);
  and _17826_ (_09474_, _09473_, _09459_);
  or _17827_ (_09475_, _09474_, _09465_);
  and _17828_ (_09476_, _09475_, _09458_);
  and _17829_ (_09477_, _09457_, word_in[25]);
  or _17830_ (_07416_, _09477_, _09476_);
  and _17831_ (_09478_, _08747_, word_in[18]);
  and _17832_ (_09479_, _09440_, _09478_);
  and _17833_ (_09480_, _08756_, word_in[2]);
  and _17834_ (_09481_, _09447_, _09480_);
  not _17835_ (_09482_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  nor _17836_ (_09483_, _09447_, _09482_);
  nor _17837_ (_09484_, _09483_, _09481_);
  nor _17838_ (_09485_, _09484_, _09442_);
  and _17839_ (_09486_, _09442_, word_in[10]);
  or _17840_ (_09487_, _09486_, _09485_);
  and _17841_ (_09488_, _09487_, _09459_);
  or _17842_ (_09489_, _09488_, _09479_);
  and _17843_ (_09490_, _09489_, _09458_);
  and _17844_ (_09491_, _09457_, word_in[26]);
  or _17845_ (_07419_, _09491_, _09490_);
  and _17846_ (_09493_, _08747_, word_in[19]);
  and _17847_ (_09494_, _09440_, _09493_);
  and _17848_ (_09495_, _08756_, word_in[3]);
  and _17849_ (_09496_, _09447_, _09495_);
  not _17850_ (_09497_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  nor _17851_ (_09498_, _09447_, _09497_);
  nor _17852_ (_09499_, _09498_, _09496_);
  nor _17853_ (_09500_, _09499_, _09442_);
  and _17854_ (_09501_, _09442_, word_in[11]);
  or _17855_ (_09502_, _09501_, _09500_);
  and _17856_ (_09503_, _09502_, _09459_);
  or _17857_ (_09504_, _09503_, _09494_);
  and _17858_ (_09505_, _09504_, _09458_);
  and _17859_ (_09506_, _09457_, word_in[27]);
  or _17860_ (_07421_, _09506_, _09505_);
  and _17861_ (_09507_, _09457_, word_in[28]);
  not _17862_ (_09508_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  nor _17863_ (_09509_, _09447_, _09508_);
  and _17864_ (_09510_, _08756_, word_in[4]);
  and _17865_ (_09511_, _09447_, _09510_);
  or _17866_ (_09512_, _09511_, _09509_);
  or _17867_ (_09514_, _09512_, _09442_);
  or _17868_ (_09515_, _09453_, word_in[12]);
  and _17869_ (_09516_, _09515_, _09514_);
  or _17870_ (_09517_, _09516_, _09440_);
  and _17871_ (_09518_, _08747_, word_in[20]);
  or _17872_ (_09519_, _09459_, _09518_);
  and _17873_ (_09520_, _09519_, _09458_);
  and _17874_ (_09522_, _09520_, _09517_);
  or _17875_ (_07423_, _09522_, _09507_);
  and _17876_ (_09523_, _08747_, word_in[21]);
  and _17877_ (_09524_, _09440_, _09523_);
  and _17878_ (_09525_, _08756_, word_in[5]);
  and _17879_ (_09526_, _09447_, _09525_);
  not _17880_ (_09527_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  nor _17881_ (_09530_, _09447_, _09527_);
  nor _17882_ (_09531_, _09530_, _09526_);
  nor _17883_ (_09532_, _09531_, _09442_);
  and _17884_ (_09533_, _09442_, word_in[13]);
  or _17885_ (_09534_, _09533_, _09532_);
  and _17886_ (_09535_, _09534_, _09459_);
  or _17887_ (_09536_, _09535_, _09524_);
  and _17888_ (_09537_, _09536_, _09458_);
  and _17889_ (_09538_, _09457_, word_in[29]);
  or _17890_ (_07427_, _09538_, _09537_);
  not _17891_ (_09539_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  nor _17892_ (_09540_, _09447_, _09539_);
  and _17893_ (_09541_, _08756_, word_in[6]);
  and _17894_ (_09542_, _09447_, _09541_);
  or _17895_ (_09543_, _09542_, _09540_);
  or _17896_ (_09544_, _09543_, _09442_);
  or _17897_ (_09545_, _09453_, word_in[14]);
  and _17898_ (_09546_, _09545_, _09544_);
  or _17899_ (_09547_, _09546_, _09440_);
  and _17900_ (_09548_, _08747_, word_in[22]);
  or _17901_ (_09549_, _09459_, _09548_);
  and _17902_ (_09550_, _09549_, _09458_);
  and _17903_ (_09551_, _09550_, _09547_);
  and _17904_ (_09552_, _09457_, word_in[30]);
  or _17905_ (_07431_, _09552_, _09551_);
  and _17906_ (_09553_, _09440_, _08769_);
  and _17907_ (_09554_, _09447_, _08760_);
  nor _17908_ (_09555_, _09447_, _08494_);
  or _17909_ (_09556_, _09555_, _09554_);
  or _17910_ (_09557_, _09556_, _09442_);
  nand _17911_ (_09558_, _09442_, _08764_);
  and _17912_ (_09559_, _09558_, _09459_);
  and _17913_ (_09560_, _09559_, _09557_);
  or _17914_ (_09561_, _09560_, _09553_);
  and _17915_ (_09562_, _09561_, _09458_);
  and _17916_ (_09563_, _09457_, word_in[31]);
  or _17917_ (_07434_, _09563_, _09562_);
  and _17918_ (_09564_, _08743_, _08674_);
  and _17919_ (_09565_, _08747_, _08548_);
  and _17920_ (_09566_, _09565_, _08620_);
  not _17921_ (_09567_, _09566_);
  or _17922_ (_09568_, _09567_, _09349_);
  and _17923_ (_09569_, _08751_, _08511_);
  and _17924_ (_09570_, _09569_, _08525_);
  not _17925_ (_09571_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  and _17926_ (_09572_, _09333_, _09335_);
  and _17927_ (_09573_, _09572_, _08429_);
  nor _17928_ (_09574_, _09573_, _09571_);
  and _17929_ (_09575_, _09573_, _09449_);
  or _17930_ (_09576_, _09575_, _09574_);
  or _17931_ (_09577_, _09576_, _09570_);
  not _17932_ (_09578_, _09570_);
  or _17933_ (_09579_, _09578_, word_in[8]);
  and _17934_ (_09580_, _09579_, _09577_);
  or _17935_ (_09581_, _09580_, _09566_);
  and _17936_ (_09582_, _09581_, _09568_);
  or _17937_ (_09583_, _09582_, _09564_);
  not _17938_ (_09584_, _09564_);
  or _17939_ (_09585_, _09584_, word_in[24]);
  and _17940_ (_07517_, _09585_, _09583_);
  not _17941_ (_09586_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  nor _17942_ (_09587_, _09573_, _09586_);
  and _17943_ (_09588_, _09573_, _09466_);
  or _17944_ (_09589_, _09588_, _09587_);
  or _17945_ (_09590_, _09589_, _09570_);
  or _17946_ (_09591_, _09578_, word_in[9]);
  and _17947_ (_09592_, _09591_, _09590_);
  or _17948_ (_09593_, _09592_, _09566_);
  or _17949_ (_09594_, _09567_, _09464_);
  and _17950_ (_09595_, _09594_, _09584_);
  and _17951_ (_09596_, _09595_, _09593_);
  and _17952_ (_09597_, _09564_, word_in[25]);
  or _17953_ (_07520_, _09597_, _09596_);
  or _17954_ (_09598_, _09567_, _09478_);
  not _17955_ (_09599_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  nor _17956_ (_09600_, _09573_, _09599_);
  and _17957_ (_09601_, _09573_, _09480_);
  or _17958_ (_09602_, _09601_, _09600_);
  or _17959_ (_09603_, _09602_, _09570_);
  or _17960_ (_09604_, _09578_, word_in[10]);
  and _17961_ (_09605_, _09604_, _09603_);
  or _17962_ (_09606_, _09605_, _09566_);
  and _17963_ (_09607_, _09606_, _09598_);
  or _17964_ (_09608_, _09607_, _09564_);
  or _17965_ (_09609_, _09584_, word_in[26]);
  and _17966_ (_07524_, _09609_, _09608_);
  not _17967_ (_09610_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  nor _17968_ (_09611_, _09573_, _09610_);
  and _17969_ (_09612_, _09573_, _09495_);
  or _17970_ (_09613_, _09612_, _09611_);
  or _17971_ (_09614_, _09613_, _09570_);
  or _17972_ (_09615_, _09578_, word_in[11]);
  and _17973_ (_09616_, _09615_, _09614_);
  or _17974_ (_09617_, _09616_, _09566_);
  or _17975_ (_09618_, _09567_, _09493_);
  and _17976_ (_09619_, _09618_, _09584_);
  and _17977_ (_09620_, _09619_, _09617_);
  and _17978_ (_09621_, _09564_, word_in[27]);
  or _17979_ (_07529_, _09621_, _09620_);
  not _17980_ (_09622_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  nor _17981_ (_09623_, _09573_, _09622_);
  and _17982_ (_09624_, _09573_, _09510_);
  or _17983_ (_09625_, _09624_, _09623_);
  or _17984_ (_09626_, _09625_, _09570_);
  or _17985_ (_09627_, _09578_, word_in[12]);
  and _17986_ (_09628_, _09627_, _09626_);
  or _17987_ (_09629_, _09628_, _09566_);
  or _17988_ (_09630_, _09567_, _09518_);
  and _17989_ (_09631_, _09630_, _09584_);
  and _17990_ (_09632_, _09631_, _09629_);
  and _17991_ (_09633_, _09564_, word_in[28]);
  or _17992_ (_07534_, _09633_, _09632_);
  or _17993_ (_09634_, _09567_, _09523_);
  not _17994_ (_09635_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  nor _17995_ (_09636_, _09573_, _09635_);
  and _17996_ (_09637_, _09573_, _09525_);
  or _17997_ (_09638_, _09637_, _09636_);
  or _17998_ (_09639_, _09638_, _09570_);
  or _17999_ (_09640_, _09578_, word_in[13]);
  and _18000_ (_09641_, _09640_, _09639_);
  or _18001_ (_09642_, _09641_, _09566_);
  and _18002_ (_09643_, _09642_, _09634_);
  or _18003_ (_09644_, _09643_, _09564_);
  or _18004_ (_09645_, _09584_, word_in[29]);
  and _18005_ (_07537_, _09645_, _09644_);
  or _18006_ (_09646_, _09567_, _09548_);
  not _18007_ (_09647_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  nor _18008_ (_09648_, _09573_, _09647_);
  and _18009_ (_09649_, _09573_, _09541_);
  or _18010_ (_09650_, _09649_, _09648_);
  or _18011_ (_09651_, _09650_, _09570_);
  or _18012_ (_09652_, _09578_, word_in[14]);
  and _18013_ (_09653_, _09652_, _09651_);
  or _18014_ (_09654_, _09653_, _09566_);
  and _18015_ (_09655_, _09654_, _09646_);
  or _18016_ (_09656_, _09655_, _09564_);
  or _18017_ (_09657_, _09584_, word_in[30]);
  and _18018_ (_07540_, _09657_, _09656_);
  nor _18019_ (_09658_, _09573_, _08593_);
  and _18020_ (_09659_, _09573_, _08760_);
  or _18021_ (_09660_, _09659_, _09658_);
  or _18022_ (_09661_, _09660_, _09570_);
  nand _18023_ (_09662_, _09570_, _08764_);
  and _18024_ (_09663_, _09662_, _09661_);
  or _18025_ (_09664_, _09663_, _09566_);
  or _18026_ (_09665_, _09567_, _08769_);
  and _18027_ (_09666_, _09665_, _09584_);
  and _18028_ (_09667_, _09666_, _09664_);
  and _18029_ (_09668_, _09564_, word_in[31]);
  or _18030_ (_07543_, _09668_, _09667_);
  and _18031_ (_09669_, _08747_, _08511_);
  and _18032_ (_09670_, _09669_, _08620_);
  not _18033_ (_09671_, _09670_);
  and _18034_ (_09672_, _08752_, _08525_);
  not _18035_ (_09673_, _08755_);
  nor _18036_ (_09674_, _09444_, _09673_);
  and _18037_ (_09675_, _09674_, _09449_);
  not _18038_ (_09676_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  nor _18039_ (_09677_, _09674_, _09676_);
  nor _18040_ (_09678_, _09677_, _09675_);
  nor _18041_ (_09679_, _09678_, _09672_);
  and _18042_ (_09680_, _09672_, word_in[8]);
  or _18043_ (_09681_, _09680_, _09679_);
  and _18044_ (_09682_, _09681_, _09671_);
  and _18045_ (_09683_, _08743_, _09059_);
  and _18046_ (_09684_, _09670_, _09349_);
  or _18047_ (_09685_, _09684_, _09683_);
  or _18048_ (_09686_, _09685_, _09682_);
  not _18049_ (_09687_, _09683_);
  or _18050_ (_09688_, _09687_, word_in[24]);
  and _18051_ (_07608_, _09688_, _09686_);
  and _18052_ (_09689_, _09670_, _09464_);
  and _18053_ (_09690_, _09674_, _09466_);
  not _18054_ (_09691_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  nor _18055_ (_09692_, _09674_, _09691_);
  nor _18056_ (_09693_, _09692_, _09690_);
  nor _18057_ (_09694_, _09693_, _09672_);
  and _18058_ (_09695_, _09672_, word_in[9]);
  or _18059_ (_09696_, _09695_, _09694_);
  and _18060_ (_09697_, _09696_, _09671_);
  or _18061_ (_09698_, _09697_, _09689_);
  and _18062_ (_09699_, _09698_, _09687_);
  and _18063_ (_09700_, _09683_, word_in[25]);
  or _18064_ (_07611_, _09700_, _09699_);
  and _18065_ (_09701_, _09683_, word_in[26]);
  not _18066_ (_09702_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  nor _18067_ (_09703_, _09674_, _09702_);
  and _18068_ (_09704_, _09674_, _09480_);
  or _18069_ (_09705_, _09704_, _09703_);
  or _18070_ (_09706_, _09705_, _09672_);
  not _18071_ (_09707_, _09672_);
  or _18072_ (_09708_, _09707_, word_in[10]);
  and _18073_ (_09709_, _09708_, _09706_);
  or _18074_ (_09710_, _09709_, _09670_);
  or _18075_ (_09711_, _09671_, _09478_);
  and _18076_ (_09712_, _09711_, _09687_);
  and _18077_ (_09713_, _09712_, _09710_);
  or _18078_ (_07615_, _09713_, _09701_);
  and _18079_ (_09714_, _09683_, word_in[27]);
  not _18080_ (_09715_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  nor _18081_ (_09716_, _09674_, _09715_);
  and _18082_ (_09717_, _09674_, _09495_);
  or _18083_ (_09718_, _09717_, _09716_);
  or _18084_ (_09719_, _09718_, _09672_);
  or _18085_ (_09720_, _09707_, word_in[11]);
  and _18086_ (_09721_, _09720_, _09719_);
  or _18087_ (_09722_, _09721_, _09670_);
  or _18088_ (_09723_, _09671_, _09493_);
  and _18089_ (_09724_, _09723_, _09687_);
  and _18090_ (_09725_, _09724_, _09722_);
  or _18091_ (_07618_, _09725_, _09714_);
  and _18092_ (_09726_, _09670_, _09518_);
  and _18093_ (_09727_, _09674_, _09510_);
  not _18094_ (_09728_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  nor _18095_ (_09729_, _09674_, _09728_);
  nor _18096_ (_09730_, _09729_, _09727_);
  nor _18097_ (_09731_, _09730_, _09672_);
  and _18098_ (_09732_, _09672_, word_in[12]);
  or _18099_ (_09733_, _09732_, _09731_);
  and _18100_ (_09734_, _09733_, _09671_);
  or _18101_ (_09735_, _09734_, _09726_);
  and _18102_ (_09736_, _09735_, _09687_);
  and _18103_ (_09737_, _09683_, word_in[28]);
  or _18104_ (_07623_, _09737_, _09736_);
  and _18105_ (_09738_, _09683_, word_in[29]);
  and _18106_ (_09739_, _09674_, _09525_);
  not _18107_ (_09740_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  nor _18108_ (_09741_, _09674_, _09740_);
  nor _18109_ (_09742_, _09741_, _09739_);
  nor _18110_ (_09743_, _09742_, _09672_);
  and _18111_ (_09744_, _09672_, word_in[13]);
  or _18112_ (_09745_, _09744_, _09743_);
  or _18113_ (_09746_, _09745_, _09670_);
  or _18114_ (_09747_, _09671_, _09523_);
  and _18115_ (_09748_, _09747_, _09687_);
  and _18116_ (_09749_, _09748_, _09746_);
  or _18117_ (_07627_, _09749_, _09738_);
  and _18118_ (_09750_, _09683_, word_in[30]);
  and _18119_ (_09751_, _09674_, _09541_);
  not _18120_ (_09752_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  nor _18121_ (_09753_, _09674_, _09752_);
  nor _18122_ (_09754_, _09753_, _09751_);
  nor _18123_ (_09755_, _09754_, _09672_);
  and _18124_ (_09756_, _09672_, word_in[14]);
  or _18125_ (_09757_, _09756_, _09755_);
  and _18126_ (_09758_, _09757_, _09671_);
  and _18127_ (_09759_, _09670_, _09548_);
  or _18128_ (_09760_, _09759_, _09758_);
  and _18129_ (_09761_, _09760_, _09687_);
  or _18130_ (_07630_, _09761_, _09750_);
  and _18131_ (_09762_, _09670_, _08769_);
  and _18132_ (_09763_, _09674_, _08760_);
  nor _18133_ (_09764_, _09674_, _08477_);
  or _18134_ (_09765_, _09764_, _09763_);
  or _18135_ (_09766_, _09765_, _09672_);
  nand _18136_ (_09767_, _09672_, _08764_);
  and _18137_ (_09768_, _09767_, _09671_);
  and _18138_ (_09769_, _09768_, _09766_);
  or _18139_ (_09770_, _09769_, _09762_);
  and _18140_ (_09771_, _09770_, _09687_);
  and _18141_ (_09772_, _09683_, word_in[31]);
  or _18142_ (_07635_, _09772_, _09771_);
  not _18143_ (_09773_, _08684_);
  and _18144_ (_09774_, _08744_, _09773_);
  and _18145_ (_09775_, _09774_, _08511_);
  not _18146_ (_09776_, _09775_);
  not _18147_ (_09777_, _08619_);
  and _18148_ (_09778_, _08748_, _09777_);
  and _18149_ (_09779_, _09778_, _08540_);
  and _18150_ (_09780_, _09779_, _09349_);
  not _18151_ (_09781_, _09779_);
  and _18152_ (_09783_, _08751_, _08880_);
  not _18153_ (_09784_, _09783_);
  nor _18154_ (_09785_, _09333_, _08754_);
  and _18155_ (_09786_, _08756_, _08869_);
  and _18156_ (_09787_, _09786_, _09785_);
  and _18157_ (_09789_, _09787_, word_in[0]);
  not _18158_ (_09790_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  nor _18159_ (_09792_, _09787_, _09790_);
  or _18160_ (_09793_, _09792_, _09789_);
  and _18161_ (_09795_, _09793_, _09784_);
  and _18162_ (_09796_, _09783_, word_in[8]);
  or _18163_ (_09797_, _09796_, _09795_);
  and _18164_ (_09798_, _09797_, _09781_);
  or _18165_ (_09799_, _09798_, _09780_);
  and _18166_ (_09800_, _09799_, _09776_);
  and _18167_ (_09801_, _08743_, word_in[24]);
  and _18168_ (_09802_, _09775_, _09801_);
  or _18169_ (_07728_, _09802_, _09800_);
  or _18170_ (_09803_, _09784_, word_in[9]);
  not _18171_ (_09804_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  nor _18172_ (_09805_, _09787_, _09804_);
  and _18173_ (_09807_, _09787_, word_in[1]);
  or _18174_ (_09808_, _09807_, _09805_);
  or _18175_ (_09809_, _09808_, _09783_);
  and _18176_ (_09811_, _09809_, _09803_);
  or _18177_ (_09812_, _09811_, _09779_);
  or _18178_ (_09814_, _09781_, _09464_);
  and _18179_ (_09815_, _09814_, _09812_);
  or _18180_ (_09816_, _09815_, _09775_);
  or _18181_ (_09817_, _09776_, _09366_);
  and _18182_ (_07731_, _09817_, _09816_);
  not _18183_ (_09818_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  nor _18184_ (_09819_, _09787_, _09818_);
  and _18185_ (_09821_, _09787_, word_in[2]);
  or _18186_ (_09823_, _09821_, _09819_);
  and _18187_ (_09824_, _09823_, _09784_);
  and _18188_ (_09825_, _09783_, word_in[10]);
  or _18189_ (_09826_, _09825_, _09824_);
  and _18190_ (_09827_, _09826_, _09781_);
  and _18191_ (_09828_, _09779_, _09478_);
  or _18192_ (_09829_, _09828_, _09775_);
  or _18193_ (_09830_, _09829_, _09827_);
  or _18194_ (_09832_, _09776_, _09368_);
  and _18195_ (_07734_, _09832_, _09830_);
  and _18196_ (_09833_, _09779_, _09493_);
  not _18197_ (_09834_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  nor _18198_ (_09835_, _09787_, _09834_);
  and _18199_ (_09836_, _09787_, word_in[3]);
  or _18200_ (_09837_, _09836_, _09835_);
  and _18201_ (_09838_, _09837_, _09784_);
  and _18202_ (_09839_, _09783_, word_in[11]);
  or _18203_ (_09840_, _09839_, _09838_);
  and _18204_ (_09841_, _09840_, _09781_);
  or _18205_ (_09842_, _09841_, _09833_);
  and _18206_ (_09843_, _09842_, _09776_);
  and _18207_ (_09844_, _09775_, _09380_);
  or _18208_ (_07738_, _09844_, _09843_);
  and _18209_ (_09845_, _09779_, _09518_);
  not _18210_ (_09846_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  nor _18211_ (_09847_, _09787_, _09846_);
  and _18212_ (_09848_, _09787_, word_in[4]);
  or _18213_ (_09849_, _09848_, _09847_);
  and _18214_ (_09850_, _09849_, _09784_);
  and _18215_ (_09851_, _09783_, word_in[12]);
  or _18216_ (_09852_, _09851_, _09850_);
  and _18217_ (_09853_, _09852_, _09781_);
  or _18218_ (_09854_, _09853_, _09845_);
  and _18219_ (_09855_, _09854_, _09776_);
  and _18220_ (_09856_, _09775_, _09402_);
  or _18221_ (_07742_, _09856_, _09855_);
  and _18222_ (_09857_, _09779_, _09523_);
  not _18223_ (_09858_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  nor _18224_ (_09859_, _09787_, _09858_);
  and _18225_ (_09860_, _09787_, word_in[5]);
  or _18226_ (_09861_, _09860_, _09859_);
  and _18227_ (_09862_, _09861_, _09784_);
  and _18228_ (_09863_, _09783_, word_in[13]);
  or _18229_ (_09864_, _09863_, _09862_);
  and _18230_ (_09865_, _09864_, _09781_);
  or _18231_ (_09866_, _09865_, _09857_);
  and _18232_ (_09867_, _09866_, _09776_);
  and _18233_ (_09868_, _09775_, _09414_);
  or _18234_ (_07745_, _09868_, _09867_);
  and _18235_ (_09869_, _09779_, _09548_);
  not _18236_ (_09870_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  nor _18237_ (_09871_, _09787_, _09870_);
  and _18238_ (_09872_, _09787_, word_in[6]);
  or _18239_ (_09873_, _09872_, _09871_);
  and _18240_ (_09874_, _09873_, _09784_);
  and _18241_ (_09875_, _09783_, word_in[14]);
  or _18242_ (_09876_, _09875_, _09874_);
  and _18243_ (_09877_, _09876_, _09781_);
  or _18244_ (_09878_, _09877_, _09869_);
  and _18245_ (_09879_, _09878_, _09776_);
  and _18246_ (_09880_, _09775_, _09426_);
  or _18247_ (_07747_, _09880_, _09879_);
  and _18248_ (_09881_, _09779_, _08769_);
  nor _18249_ (_09882_, _09787_, _08601_);
  and _18250_ (_09883_, _09787_, word_in[7]);
  or _18251_ (_09884_, _09883_, _09882_);
  and _18252_ (_09885_, _09884_, _09784_);
  and _18253_ (_09886_, _09783_, word_in[15]);
  or _18254_ (_09887_, _09886_, _09885_);
  and _18255_ (_09888_, _09887_, _09781_);
  or _18256_ (_09889_, _09888_, _09881_);
  and _18257_ (_09890_, _09889_, _09776_);
  and _18258_ (_09891_, _09775_, _08774_);
  or _18259_ (_07750_, _09891_, _09890_);
  and _18260_ (_09892_, _09774_, _08540_);
  not _18261_ (_09893_, _09892_);
  and _18262_ (_09894_, _09778_, _08514_);
  and _18263_ (_09895_, _09894_, _09349_);
  not _18264_ (_09896_, _09894_);
  and _18265_ (_09897_, _09441_, _08600_);
  and _18266_ (_09898_, _09786_, _09445_);
  and _18267_ (_09899_, _09898_, _09449_);
  not _18268_ (_09900_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  nor _18269_ (_09901_, _09898_, _09900_);
  nor _18270_ (_09902_, _09901_, _09899_);
  nor _18271_ (_09903_, _09902_, _09897_);
  and _18272_ (_09904_, _09897_, word_in[8]);
  or _18273_ (_09905_, _09904_, _09903_);
  and _18274_ (_09906_, _09905_, _09896_);
  or _18275_ (_09907_, _09906_, _09895_);
  and _18276_ (_09908_, _09907_, _09893_);
  and _18277_ (_09909_, _09892_, _09801_);
  or _18278_ (_07827_, _09909_, _09908_);
  or _18279_ (_09910_, _09896_, _09464_);
  not _18280_ (_09911_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  nor _18281_ (_09912_, _09898_, _09911_);
  and _18282_ (_09913_, _09898_, _09466_);
  or _18283_ (_09914_, _09913_, _09912_);
  or _18284_ (_09915_, _09914_, _09897_);
  not _18285_ (_09916_, _09897_);
  or _18286_ (_09917_, _09916_, word_in[9]);
  and _18287_ (_09918_, _09917_, _09915_);
  or _18288_ (_09919_, _09918_, _09894_);
  and _18289_ (_09920_, _09919_, _09910_);
  or _18290_ (_09921_, _09920_, _09892_);
  or _18291_ (_09922_, _09893_, _09366_);
  and _18292_ (_07830_, _09922_, _09921_);
  and _18293_ (_09923_, _09898_, _09480_);
  not _18294_ (_09924_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  nor _18295_ (_09925_, _09898_, _09924_);
  nor _18296_ (_09926_, _09925_, _09923_);
  nor _18297_ (_09927_, _09926_, _09897_);
  and _18298_ (_09928_, _09897_, word_in[10]);
  or _18299_ (_09929_, _09928_, _09927_);
  and _18300_ (_09930_, _09929_, _09896_);
  and _18301_ (_09931_, _09894_, _09478_);
  or _18302_ (_09932_, _09931_, _09892_);
  or _18303_ (_09933_, _09932_, _09930_);
  or _18304_ (_09934_, _09893_, _09368_);
  and _18305_ (_07834_, _09934_, _09933_);
  and _18306_ (_09935_, _06688_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  nor _18307_ (_09936_, _06688_, _05669_);
  or _18308_ (_09937_, _09936_, _09935_);
  and _18309_ (_07837_, _09937_, _04856_);
  and _18310_ (_09938_, _09898_, _09495_);
  not _18311_ (_09939_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  nor _18312_ (_09940_, _09898_, _09939_);
  nor _18313_ (_09941_, _09940_, _09938_);
  nor _18314_ (_09942_, _09941_, _09897_);
  and _18315_ (_09943_, _09897_, word_in[11]);
  or _18316_ (_09944_, _09943_, _09942_);
  and _18317_ (_09945_, _09944_, _09896_);
  and _18318_ (_09946_, _09894_, _09493_);
  or _18319_ (_09947_, _09946_, _09945_);
  and _18320_ (_09948_, _09947_, _09893_);
  and _18321_ (_09949_, _09892_, _09380_);
  or _18322_ (_07839_, _09949_, _09948_);
  or _18323_ (_09950_, _05682_, _05676_);
  and _18324_ (_09951_, _09950_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  and _18325_ (_09952_, _06997_, _05671_);
  or _18326_ (_09953_, _05674_, _05679_);
  or _18327_ (_09954_, _05675_, _09953_);
  and _18328_ (_09955_, _04861_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  and _18329_ (_09956_, _09955_, _09954_);
  or _18330_ (_09957_, _09956_, _09952_);
  or _18331_ (_09958_, _09957_, _09951_);
  and _18332_ (_07842_, _09958_, _04856_);
  and _18333_ (_09959_, _09894_, _09518_);
  and _18334_ (_09960_, _09898_, _09510_);
  not _18335_ (_09961_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  nor _18336_ (_09962_, _09898_, _09961_);
  nor _18337_ (_09963_, _09962_, _09960_);
  nor _18338_ (_09964_, _09963_, _09897_);
  and _18339_ (_09965_, _09897_, word_in[12]);
  or _18340_ (_09966_, _09965_, _09964_);
  and _18341_ (_09967_, _09966_, _09896_);
  or _18342_ (_09968_, _09967_, _09959_);
  and _18343_ (_09969_, _09968_, _09893_);
  and _18344_ (_09970_, _09892_, _09402_);
  or _18345_ (_07844_, _09970_, _09969_);
  not _18346_ (_09971_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  nor _18347_ (_09972_, _09898_, _09971_);
  and _18348_ (_09973_, _09898_, _09525_);
  or _18349_ (_09974_, _09973_, _09972_);
  or _18350_ (_09975_, _09974_, _09897_);
  or _18351_ (_09976_, _09916_, word_in[13]);
  and _18352_ (_09977_, _09976_, _09975_);
  or _18353_ (_09978_, _09977_, _09894_);
  or _18354_ (_09979_, _09896_, _09523_);
  and _18355_ (_09980_, _09979_, _09978_);
  or _18356_ (_09981_, _09980_, _09892_);
  or _18357_ (_09982_, _09893_, _09414_);
  and _18358_ (_07849_, _09982_, _09981_);
  not _18359_ (_09983_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  nor _18360_ (_09985_, _09898_, _09983_);
  and _18361_ (_09986_, _09898_, _09541_);
  or _18362_ (_09987_, _09986_, _09985_);
  or _18363_ (_09988_, _09987_, _09897_);
  or _18364_ (_09989_, _09916_, word_in[14]);
  and _18365_ (_09990_, _09989_, _09988_);
  and _18366_ (_09991_, _09990_, _09896_);
  and _18367_ (_09992_, _09894_, _09548_);
  or _18368_ (_09993_, _09992_, _09892_);
  or _18369_ (_09994_, _09993_, _09991_);
  or _18370_ (_09995_, _09893_, _09426_);
  and _18371_ (_07852_, _09995_, _09994_);
  and _18372_ (_09997_, _09894_, _08769_);
  and _18373_ (_09998_, _09898_, _08760_);
  nor _18374_ (_09999_, _09898_, _08488_);
  nor _18375_ (_10000_, _09999_, _09998_);
  nor _18376_ (_10001_, _10000_, _09897_);
  and _18377_ (_10002_, _09897_, word_in[15]);
  or _18378_ (_10003_, _10002_, _10001_);
  and _18379_ (_10004_, _10003_, _09896_);
  or _18380_ (_10005_, _10004_, _09997_);
  and _18381_ (_10006_, _10005_, _09893_);
  and _18382_ (_10007_, _09892_, _08774_);
  or _18383_ (_07856_, _10007_, _10006_);
  and _18384_ (_10008_, _09774_, _08514_);
  not _18385_ (_10009_, _10008_);
  and _18386_ (_10010_, _09778_, _08548_);
  and _18387_ (_10011_, _10010_, _09349_);
  not _18388_ (_10012_, _10010_);
  and _18389_ (_10013_, _09569_, _08600_);
  and _18390_ (_10014_, _09572_, _08869_);
  and _18391_ (_10015_, _10014_, word_in[0]);
  not _18392_ (_10016_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  nor _18393_ (_10017_, _10014_, _10016_);
  nor _18394_ (_10018_, _10017_, _10015_);
  nor _18395_ (_10019_, _10018_, _10013_);
  and _18396_ (_10020_, _10013_, word_in[8]);
  or _18397_ (_10021_, _10020_, _10019_);
  and _18398_ (_10022_, _10021_, _10012_);
  or _18399_ (_10023_, _10022_, _10011_);
  and _18400_ (_10024_, _10023_, _10009_);
  and _18401_ (_10025_, _10008_, _09801_);
  or _18402_ (_07923_, _10025_, _10024_);
  not _18403_ (_10026_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  nor _18404_ (_10027_, _10014_, _10026_);
  and _18405_ (_10028_, _10014_, word_in[1]);
  or _18406_ (_10029_, _10028_, _10027_);
  or _18407_ (_10030_, _10029_, _10013_);
  not _18408_ (_10031_, _10013_);
  or _18409_ (_10032_, _10031_, word_in[9]);
  and _18410_ (_10033_, _10032_, _10030_);
  or _18411_ (_10034_, _10033_, _10010_);
  or _18412_ (_10035_, _10012_, _09464_);
  and _18413_ (_10036_, _10035_, _10009_);
  and _18414_ (_10037_, _10036_, _10034_);
  and _18415_ (_10038_, _10008_, _09366_);
  or _18416_ (_07926_, _10038_, _10037_);
  and _18417_ (_10039_, _10010_, _09478_);
  not _18418_ (_10040_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  nor _18419_ (_10041_, _10014_, _10040_);
  and _18420_ (_10042_, _10014_, word_in[2]);
  nor _18421_ (_10043_, _10042_, _10041_);
  nor _18422_ (_10044_, _10043_, _10013_);
  and _18423_ (_10045_, _10013_, word_in[10]);
  or _18424_ (_10046_, _10045_, _10044_);
  and _18425_ (_10048_, _10046_, _10012_);
  or _18426_ (_10049_, _10048_, _10039_);
  and _18427_ (_10050_, _10049_, _10009_);
  and _18428_ (_10051_, _10008_, _09368_);
  or _18429_ (_07930_, _10051_, _10050_);
  or _18430_ (_10052_, _10031_, word_in[11]);
  not _18431_ (_10053_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  nor _18432_ (_10054_, _10014_, _10053_);
  and _18433_ (_10055_, _10014_, word_in[3]);
  or _18434_ (_10056_, _10055_, _10054_);
  or _18435_ (_10057_, _10056_, _10013_);
  and _18436_ (_10058_, _10057_, _10052_);
  or _18437_ (_10059_, _10058_, _10010_);
  or _18438_ (_10061_, _10012_, _09493_);
  and _18439_ (_10062_, _10061_, _10059_);
  or _18440_ (_10063_, _10062_, _10008_);
  or _18441_ (_10064_, _10009_, _09380_);
  and _18442_ (_07934_, _10064_, _10063_);
  and _18443_ (_10065_, _10010_, _09518_);
  not _18444_ (_10066_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  nor _18445_ (_10068_, _10014_, _10066_);
  and _18446_ (_10069_, _10014_, word_in[4]);
  nor _18447_ (_10070_, _10069_, _10068_);
  nor _18448_ (_10071_, _10070_, _10013_);
  and _18449_ (_10073_, _10013_, word_in[12]);
  or _18450_ (_10074_, _10073_, _10071_);
  and _18451_ (_10075_, _10074_, _10012_);
  or _18452_ (_10076_, _10075_, _10065_);
  and _18453_ (_10077_, _10076_, _10009_);
  and _18454_ (_10078_, _10008_, _09402_);
  or _18455_ (_07938_, _10078_, _10077_);
  and _18456_ (_10079_, _10010_, _09523_);
  not _18457_ (_10080_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  nor _18458_ (_10081_, _10014_, _10080_);
  and _18459_ (_10082_, _10014_, word_in[5]);
  nor _18460_ (_10083_, _10082_, _10081_);
  nor _18461_ (_10084_, _10083_, _10013_);
  and _18462_ (_10085_, _10013_, word_in[13]);
  or _18463_ (_10086_, _10085_, _10084_);
  and _18464_ (_10087_, _10086_, _10012_);
  or _18465_ (_10088_, _10087_, _10079_);
  and _18466_ (_10089_, _10088_, _10009_);
  and _18467_ (_10090_, _10008_, _09414_);
  or _18468_ (_07941_, _10090_, _10089_);
  and _18469_ (_10091_, _10010_, _09548_);
  not _18470_ (_10092_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  nor _18471_ (_10093_, _10014_, _10092_);
  and _18472_ (_10094_, _10014_, word_in[6]);
  nor _18473_ (_10095_, _10094_, _10093_);
  nor _18474_ (_10096_, _10095_, _10013_);
  and _18475_ (_10097_, _10013_, word_in[14]);
  or _18476_ (_10098_, _10097_, _10096_);
  and _18477_ (_10099_, _10098_, _10012_);
  or _18478_ (_10100_, _10099_, _10091_);
  and _18479_ (_10101_, _10100_, _10009_);
  and _18480_ (_10102_, _10008_, _09426_);
  or _18481_ (_07946_, _10102_, _10101_);
  and _18482_ (_10103_, _10010_, _08769_);
  nor _18483_ (_10104_, _10014_, _08606_);
  and _18484_ (_10105_, _10014_, word_in[7]);
  nor _18485_ (_10106_, _10105_, _10104_);
  nor _18486_ (_10107_, _10106_, _10013_);
  and _18487_ (_10108_, _10013_, word_in[15]);
  or _18488_ (_10109_, _10108_, _10107_);
  and _18489_ (_10110_, _10109_, _10012_);
  or _18490_ (_10111_, _10110_, _10103_);
  and _18491_ (_10112_, _10111_, _10009_);
  and _18492_ (_10113_, _10008_, _08774_);
  or _18493_ (_07950_, _10113_, _10112_);
  and _18494_ (_10115_, _09774_, _08548_);
  not _18495_ (_10116_, _10115_);
  and _18496_ (_10117_, _09778_, _08511_);
  and _18497_ (_10118_, _10117_, _09349_);
  not _18498_ (_10119_, _10117_);
  and _18499_ (_10120_, _08752_, _08600_);
  and _18500_ (_10121_, _09786_, _08755_);
  and _18501_ (_10122_, _10121_, word_in[0]);
  not _18502_ (_10123_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  nor _18503_ (_10124_, _10121_, _10123_);
  nor _18504_ (_10125_, _10124_, _10122_);
  nor _18505_ (_10126_, _10125_, _10120_);
  and _18506_ (_10127_, _10120_, word_in[8]);
  or _18507_ (_10128_, _10127_, _10126_);
  and _18508_ (_10129_, _10128_, _10119_);
  or _18509_ (_10130_, _10129_, _10118_);
  and _18510_ (_10131_, _10130_, _10116_);
  and _18511_ (_10132_, _10115_, _09801_);
  or _18512_ (_08020_, _10132_, _10131_);
  and _18513_ (_10133_, _10121_, word_in[1]);
  not _18514_ (_10134_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  nor _18515_ (_10136_, _10121_, _10134_);
  nor _18516_ (_10137_, _10136_, _10133_);
  nor _18517_ (_10138_, _10137_, _10120_);
  and _18518_ (_10139_, _10120_, word_in[9]);
  or _18519_ (_10140_, _10139_, _10138_);
  and _18520_ (_10141_, _10140_, _10119_);
  and _18521_ (_10142_, _10117_, _09464_);
  or _18522_ (_10144_, _10142_, _10141_);
  and _18523_ (_10145_, _10144_, _10116_);
  and _18524_ (_10147_, _10115_, _09366_);
  or _18525_ (_08023_, _10147_, _10145_);
  and _18526_ (_10148_, _10121_, word_in[2]);
  not _18527_ (_10149_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  nor _18528_ (_10150_, _10121_, _10149_);
  nor _18529_ (_10151_, _10150_, _10148_);
  nor _18530_ (_10152_, _10151_, _10120_);
  and _18531_ (_10153_, _10120_, word_in[10]);
  or _18532_ (_10154_, _10153_, _10152_);
  and _18533_ (_10155_, _10154_, _10119_);
  and _18534_ (_10156_, _10117_, _09478_);
  or _18535_ (_10157_, _10156_, _10155_);
  and _18536_ (_10158_, _10157_, _10116_);
  and _18537_ (_10159_, _10115_, _09368_);
  or _18538_ (_08026_, _10159_, _10158_);
  not _18539_ (_10160_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  nor _18540_ (_10161_, _10121_, _10160_);
  and _18541_ (_10163_, _10121_, _09495_);
  or _18542_ (_10164_, _10163_, _10161_);
  or _18543_ (_10165_, _10164_, _10120_);
  not _18544_ (_10166_, _10120_);
  or _18545_ (_10167_, _10166_, word_in[11]);
  and _18546_ (_10168_, _10167_, _10165_);
  or _18547_ (_10169_, _10168_, _10117_);
  or _18548_ (_10170_, _10119_, _09493_);
  and _18549_ (_10171_, _10170_, _10169_);
  or _18550_ (_10172_, _10171_, _10115_);
  or _18551_ (_10173_, _10116_, _09380_);
  and _18552_ (_08030_, _10173_, _10172_);
  not _18553_ (_10175_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  nor _18554_ (_10176_, _10121_, _10175_);
  and _18555_ (_10177_, _10121_, _09510_);
  or _18556_ (_10178_, _10177_, _10176_);
  or _18557_ (_10179_, _10178_, _10120_);
  or _18558_ (_10180_, _10166_, word_in[12]);
  and _18559_ (_10181_, _10180_, _10179_);
  or _18560_ (_10182_, _10181_, _10117_);
  or _18561_ (_10183_, _10119_, _09518_);
  and _18562_ (_10184_, _10183_, _10182_);
  or _18563_ (_10185_, _10184_, _10115_);
  or _18564_ (_10186_, _10116_, _09402_);
  and _18565_ (_08035_, _10186_, _10185_);
  not _18566_ (_10187_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  nor _18567_ (_10188_, _10121_, _10187_);
  and _18568_ (_10189_, _10121_, _09525_);
  or _18569_ (_10191_, _10189_, _10188_);
  or _18570_ (_10192_, _10191_, _10120_);
  or _18571_ (_10194_, _10166_, word_in[13]);
  and _18572_ (_10195_, _10194_, _10192_);
  or _18573_ (_10196_, _10195_, _10117_);
  or _18574_ (_10197_, _10119_, _09523_);
  and _18575_ (_10198_, _10197_, _10196_);
  or _18576_ (_10200_, _10198_, _10115_);
  or _18577_ (_10201_, _10116_, _09414_);
  and _18578_ (_08039_, _10201_, _10200_);
  not _18579_ (_10203_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  nor _18580_ (_10204_, _10121_, _10203_);
  and _18581_ (_10205_, _10121_, _09541_);
  or _18582_ (_10206_, _10205_, _10204_);
  or _18583_ (_10207_, _10206_, _10120_);
  or _18584_ (_10209_, _10166_, word_in[14]);
  and _18585_ (_10210_, _10209_, _10207_);
  or _18586_ (_10211_, _10210_, _10117_);
  or _18587_ (_10212_, _10119_, _09548_);
  and _18588_ (_10213_, _10212_, _10211_);
  or _18589_ (_10215_, _10213_, _10115_);
  or _18590_ (_10216_, _10116_, _09426_);
  and _18591_ (_08042_, _10216_, _10215_);
  nor _18592_ (_10218_, _10121_, _08483_);
  and _18593_ (_10219_, _10121_, _08760_);
  or _18594_ (_10220_, _10219_, _10218_);
  or _18595_ (_10222_, _10220_, _10120_);
  nand _18596_ (_10223_, _10120_, _08764_);
  and _18597_ (_10224_, _10223_, _10222_);
  or _18598_ (_10225_, _10224_, _10117_);
  or _18599_ (_10226_, _10119_, _08769_);
  and _18600_ (_10227_, _10226_, _10225_);
  or _18601_ (_10228_, _10227_, _10115_);
  or _18602_ (_10229_, _10116_, _08774_);
  and _18603_ (_08045_, _10229_, _10228_);
  nor _18604_ (_10230_, _08076_, _08072_);
  nor _18605_ (_10231_, _10230_, _08062_);
  not _18606_ (_10232_, _08087_);
  or _18607_ (_10233_, _10232_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  or _18608_ (_10234_, _10233_, _10231_);
  or _18609_ (_10235_, _08087_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  and _18610_ (_10236_, _10235_, _08085_);
  and _18611_ (_10237_, _10236_, _10234_);
  or _18612_ (_08118_, _10237_, _09299_);
  and _18613_ (_10238_, _08743_, _08685_);
  and _18614_ (_10239_, _10238_, _08511_);
  not _18615_ (_10240_, _10239_);
  and _18616_ (_10241_, _08747_, _08636_);
  and _18617_ (_10242_, _10241_, word_in[16]);
  not _18618_ (_10243_, _10241_);
  and _18619_ (_10244_, _08751_, _08521_);
  not _18620_ (_10245_, _10244_);
  not _18621_ (_10246_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  and _18622_ (_10248_, _08756_, _08431_);
  and _18623_ (_10249_, _10248_, _09785_);
  nor _18624_ (_10251_, _10249_, _10246_);
  and _18625_ (_10252_, _10249_, word_in[0]);
  or _18626_ (_10253_, _10252_, _10251_);
  and _18627_ (_10254_, _10253_, _10245_);
  and _18628_ (_10255_, _10244_, word_in[8]);
  or _18629_ (_10256_, _10255_, _10254_);
  and _18630_ (_10258_, _10256_, _10243_);
  or _18631_ (_10259_, _10258_, _10242_);
  and _18632_ (_10260_, _10259_, _10240_);
  and _18633_ (_10261_, _10239_, word_in[24]);
  or _18634_ (_08129_, _10261_, _10260_);
  and _18635_ (_10262_, _10241_, word_in[17]);
  not _18636_ (_10263_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  nor _18637_ (_10264_, _10249_, _10263_);
  and _18638_ (_10266_, _10249_, word_in[1]);
  or _18639_ (_10267_, _10266_, _10264_);
  and _18640_ (_10268_, _10267_, _10245_);
  and _18641_ (_10269_, _10244_, word_in[9]);
  or _18642_ (_10270_, _10269_, _10268_);
  and _18643_ (_10271_, _10270_, _10243_);
  or _18644_ (_10272_, _10271_, _10262_);
  and _18645_ (_10273_, _10272_, _10240_);
  and _18646_ (_10274_, _10239_, word_in[25]);
  or _18647_ (_13256_, _10274_, _10273_);
  and _18648_ (_10275_, _10241_, word_in[18]);
  not _18649_ (_10276_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  nor _18650_ (_10277_, _10249_, _10276_);
  and _18651_ (_10278_, _10249_, word_in[2]);
  or _18652_ (_10279_, _10278_, _10277_);
  and _18653_ (_10280_, _10279_, _10245_);
  and _18654_ (_10281_, _10244_, word_in[10]);
  or _18655_ (_10282_, _10281_, _10280_);
  and _18656_ (_10283_, _10282_, _10243_);
  or _18657_ (_10284_, _10283_, _10275_);
  and _18658_ (_10285_, _10284_, _10240_);
  and _18659_ (_10286_, _10239_, word_in[26]);
  or _18660_ (_13257_, _10286_, _10285_);
  and _18661_ (_10287_, _10241_, word_in[19]);
  not _18662_ (_10288_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  nor _18663_ (_10289_, _10249_, _10288_);
  and _18664_ (_10290_, _10249_, word_in[3]);
  or _18665_ (_10291_, _10290_, _10289_);
  and _18666_ (_10292_, _10291_, _10245_);
  and _18667_ (_10293_, _10244_, word_in[11]);
  or _18668_ (_10294_, _10293_, _10292_);
  and _18669_ (_10295_, _10294_, _10243_);
  or _18670_ (_10296_, _10295_, _10287_);
  and _18671_ (_10298_, _10296_, _10240_);
  and _18672_ (_10299_, _10239_, word_in[27]);
  or _18673_ (_08141_, _10299_, _10298_);
  and _18674_ (_10300_, _10241_, word_in[20]);
  not _18675_ (_10302_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  nor _18676_ (_10303_, _10249_, _10302_);
  and _18677_ (_10304_, _10249_, word_in[4]);
  or _18678_ (_10305_, _10304_, _10303_);
  and _18679_ (_10306_, _10305_, _10245_);
  and _18680_ (_10307_, _10244_, word_in[12]);
  or _18681_ (_10308_, _10307_, _10306_);
  and _18682_ (_10309_, _10308_, _10243_);
  or _18683_ (_10311_, _10309_, _10300_);
  and _18684_ (_10312_, _10311_, _10240_);
  and _18685_ (_10313_, _10239_, word_in[28]);
  or _18686_ (_13258_, _10313_, _10312_);
  and _18687_ (_10314_, _10241_, word_in[21]);
  not _18688_ (_10315_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  nor _18689_ (_10316_, _10249_, _10315_);
  and _18690_ (_10317_, _10249_, word_in[5]);
  or _18691_ (_10319_, _10317_, _10316_);
  and _18692_ (_10320_, _10319_, _10245_);
  and _18693_ (_10321_, _10244_, word_in[13]);
  or _18694_ (_10322_, _10321_, _10320_);
  and _18695_ (_10323_, _10322_, _10243_);
  or _18696_ (_10324_, _10323_, _10314_);
  and _18697_ (_10325_, _10324_, _10240_);
  and _18698_ (_10326_, _10239_, word_in[29]);
  or _18699_ (_13259_, _10326_, _10325_);
  and _18700_ (_10327_, _10241_, word_in[22]);
  not _18701_ (_10328_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  nor _18702_ (_10329_, _10249_, _10328_);
  and _18703_ (_10330_, _10249_, word_in[6]);
  or _18704_ (_10331_, _10330_, _10329_);
  and _18705_ (_10332_, _10331_, _10245_);
  and _18706_ (_10333_, _10244_, word_in[14]);
  or _18707_ (_10334_, _10333_, _10332_);
  and _18708_ (_10335_, _10334_, _10243_);
  or _18709_ (_10336_, _10335_, _10327_);
  and _18710_ (_10338_, _10336_, _10240_);
  and _18711_ (_10340_, _10239_, word_in[30]);
  or _18712_ (_08148_, _10340_, _10338_);
  and _18713_ (_10341_, _10241_, word_in[23]);
  nor _18714_ (_10342_, _10249_, _08566_);
  and _18715_ (_10343_, _10249_, word_in[7]);
  or _18716_ (_10345_, _10343_, _10342_);
  and _18717_ (_10346_, _10345_, _10245_);
  and _18718_ (_10347_, _10244_, word_in[15]);
  or _18719_ (_10348_, _10347_, _10346_);
  and _18720_ (_10349_, _10348_, _10243_);
  or _18721_ (_10350_, _10349_, _10341_);
  and _18722_ (_10351_, _10350_, _10240_);
  and _18723_ (_10352_, _10239_, word_in[31]);
  or _18724_ (_13260_, _10352_, _10351_);
  and _18725_ (_10353_, _08743_, _08636_);
  and _18726_ (_10354_, _10353_, word_in[24]);
  and _18727_ (_10355_, _09439_, _08625_);
  and _18728_ (_10356_, _09441_, _08523_);
  not _18729_ (_10357_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  and _18730_ (_10358_, _10248_, _09445_);
  nor _18731_ (_10359_, _10358_, _10357_);
  and _18732_ (_10360_, _10358_, _09449_);
  or _18733_ (_10361_, _10360_, _10359_);
  or _18734_ (_10362_, _10361_, _10356_);
  not _18735_ (_10363_, _10356_);
  or _18736_ (_10364_, _10363_, word_in[8]);
  and _18737_ (_10365_, _10364_, _10362_);
  or _18738_ (_10366_, _10365_, _10355_);
  not _18739_ (_10367_, _10353_);
  not _18740_ (_10368_, _10355_);
  or _18741_ (_10369_, _10368_, _09349_);
  and _18742_ (_10370_, _10369_, _10367_);
  and _18743_ (_10371_, _10370_, _10366_);
  or _18744_ (_13261_, _10371_, _10354_);
  or _18745_ (_10372_, _10368_, _09464_);
  not _18746_ (_10373_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  nor _18747_ (_10375_, _10358_, _10373_);
  and _18748_ (_10376_, _10358_, _09466_);
  or _18749_ (_10377_, _10376_, _10375_);
  or _18750_ (_10378_, _10377_, _10356_);
  or _18751_ (_10379_, _10363_, word_in[9]);
  and _18752_ (_10380_, _10379_, _10378_);
  or _18753_ (_10381_, _10380_, _10355_);
  and _18754_ (_10382_, _10381_, _10372_);
  or _18755_ (_10383_, _10382_, _10353_);
  or _18756_ (_10384_, _10367_, word_in[25]);
  and _18757_ (_13262_, _10384_, _10383_);
  and _18758_ (_10385_, _10358_, _09480_);
  not _18759_ (_10386_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  nor _18760_ (_10387_, _10358_, _10386_);
  nor _18761_ (_10388_, _10387_, _10385_);
  nor _18762_ (_10389_, _10388_, _10356_);
  and _18763_ (_10390_, _10356_, word_in[10]);
  or _18764_ (_10391_, _10390_, _10389_);
  and _18765_ (_10392_, _10391_, _10368_);
  and _18766_ (_10393_, _10355_, _09478_);
  or _18767_ (_10394_, _10393_, _10353_);
  or _18768_ (_10395_, _10394_, _10392_);
  or _18769_ (_10396_, _10367_, word_in[26]);
  and _18770_ (_13263_, _10396_, _10395_);
  and _18771_ (_10397_, _10358_, _09495_);
  not _18772_ (_10398_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  nor _18773_ (_10399_, _10358_, _10398_);
  nor _18774_ (_10400_, _10399_, _10397_);
  nor _18775_ (_10401_, _10400_, _10356_);
  and _18776_ (_10402_, _10356_, word_in[11]);
  or _18777_ (_10403_, _10402_, _10401_);
  and _18778_ (_10404_, _10403_, _10368_);
  and _18779_ (_10405_, _10355_, _09493_);
  or _18780_ (_10406_, _10405_, _10353_);
  or _18781_ (_10407_, _10406_, _10404_);
  or _18782_ (_10408_, _10367_, word_in[27]);
  and _18783_ (_13264_, _10408_, _10407_);
  not _18784_ (_10409_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  nor _18785_ (_10410_, _10358_, _10409_);
  and _18786_ (_10411_, _10358_, _09510_);
  or _18787_ (_10412_, _10411_, _10410_);
  or _18788_ (_10413_, _10412_, _10356_);
  or _18789_ (_10414_, _10363_, word_in[12]);
  and _18790_ (_10415_, _10414_, _10413_);
  or _18791_ (_10417_, _10415_, _10355_);
  or _18792_ (_10418_, _10368_, _09518_);
  and _18793_ (_10420_, _10418_, _10367_);
  and _18794_ (_10421_, _10420_, _10417_);
  and _18795_ (_10422_, _10353_, word_in[28]);
  or _18796_ (_13265_, _10422_, _10421_);
  and _18797_ (_10423_, _10358_, _09525_);
  not _18798_ (_10425_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  nor _18799_ (_10426_, _10358_, _10425_);
  nor _18800_ (_10428_, _10426_, _10423_);
  nor _18801_ (_10429_, _10428_, _10356_);
  and _18802_ (_10430_, _10356_, word_in[13]);
  or _18803_ (_10431_, _10430_, _10429_);
  and _18804_ (_10432_, _10431_, _10368_);
  and _18805_ (_10433_, _10355_, _09523_);
  or _18806_ (_10435_, _10433_, _10353_);
  or _18807_ (_10436_, _10435_, _10432_);
  or _18808_ (_10437_, _10367_, word_in[29]);
  and _18809_ (_08227_, _10437_, _10436_);
  or _18810_ (_10438_, _10368_, _09548_);
  not _18811_ (_10439_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  nor _18812_ (_10440_, _10358_, _10439_);
  and _18813_ (_10441_, _10358_, _09541_);
  or _18814_ (_10442_, _10441_, _10440_);
  or _18815_ (_10444_, _10442_, _10356_);
  or _18816_ (_10445_, _10363_, word_in[14]);
  and _18817_ (_10446_, _10445_, _10444_);
  or _18818_ (_10447_, _10446_, _10355_);
  and _18819_ (_10448_, _10447_, _10438_);
  or _18820_ (_10449_, _10448_, _10353_);
  or _18821_ (_10450_, _10367_, word_in[30]);
  and _18822_ (_08230_, _10450_, _10449_);
  nor _18823_ (_10451_, _10358_, _08469_);
  and _18824_ (_10452_, _10358_, _08760_);
  or _18825_ (_10453_, _10452_, _10451_);
  or _18826_ (_10454_, _10453_, _10356_);
  nand _18827_ (_10455_, _10356_, _08764_);
  and _18828_ (_10456_, _10455_, _10454_);
  or _18829_ (_10457_, _10456_, _10355_);
  or _18830_ (_10458_, _10368_, _08769_);
  and _18831_ (_10460_, _10458_, _10367_);
  and _18832_ (_10461_, _10460_, _10457_);
  and _18833_ (_10462_, _10353_, word_in[31]);
  or _18834_ (_08234_, _10462_, _10461_);
  and _18835_ (_10463_, _05007_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  and _18836_ (_10464_, _05670_, _04988_);
  and _18837_ (_10465_, _05005_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  or _18838_ (_10466_, _10465_, _10464_);
  and _18839_ (_10467_, _10466_, _04861_);
  or _18840_ (_10468_, _10467_, _10463_);
  and _18841_ (_08279_, _10468_, _04856_);
  and _18842_ (_10469_, _06688_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  and _18843_ (_10470_, _06686_, _06033_);
  or _18844_ (_10472_, _10470_, _10469_);
  and _18845_ (_08283_, _10472_, _04856_);
  and _18846_ (_10474_, _10238_, _08514_);
  and _18847_ (_10475_, _09565_, _08625_);
  not _18848_ (_10476_, _10475_);
  or _18849_ (_10477_, _10476_, _09349_);
  and _18850_ (_10479_, _09569_, _08523_);
  not _18851_ (_10481_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and _18852_ (_10482_, _09572_, _08431_);
  nor _18853_ (_10483_, _10482_, _10481_);
  and _18854_ (_10484_, _10482_, word_in[0]);
  or _18855_ (_10485_, _10484_, _10483_);
  or _18856_ (_10486_, _10485_, _10479_);
  not _18857_ (_10487_, _10479_);
  or _18858_ (_10488_, _10487_, word_in[8]);
  and _18859_ (_10489_, _10488_, _10486_);
  or _18860_ (_10490_, _10489_, _10475_);
  and _18861_ (_10491_, _10490_, _10477_);
  or _18862_ (_10492_, _10491_, _10474_);
  not _18863_ (_10493_, _10474_);
  or _18864_ (_10494_, _10493_, word_in[24]);
  and _18865_ (_08293_, _10494_, _10492_);
  not _18866_ (_10495_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  nor _18867_ (_10496_, _10482_, _10495_);
  and _18868_ (_10497_, _10482_, word_in[1]);
  or _18869_ (_10498_, _10497_, _10496_);
  or _18870_ (_10500_, _10498_, _10479_);
  or _18871_ (_10501_, _10487_, word_in[9]);
  and _18872_ (_10502_, _10501_, _10500_);
  or _18873_ (_10503_, _10502_, _10475_);
  or _18874_ (_10504_, _10476_, _09464_);
  and _18875_ (_10505_, _10504_, _10493_);
  and _18876_ (_10506_, _10505_, _10503_);
  and _18877_ (_10508_, _10474_, word_in[25]);
  or _18878_ (_08297_, _10508_, _10506_);
  or _18879_ (_10509_, _10476_, _09478_);
  not _18880_ (_10510_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  nor _18881_ (_10511_, _10482_, _10510_);
  and _18882_ (_10512_, _10482_, word_in[2]);
  or _18883_ (_10513_, _10512_, _10511_);
  or _18884_ (_10515_, _10513_, _10479_);
  or _18885_ (_10516_, _10487_, word_in[10]);
  and _18886_ (_10517_, _10516_, _10515_);
  or _18887_ (_10518_, _10517_, _10475_);
  and _18888_ (_10519_, _10518_, _10509_);
  or _18889_ (_10520_, _10519_, _10474_);
  or _18890_ (_10521_, _10493_, word_in[26]);
  and _18891_ (_08299_, _10521_, _10520_);
  not _18892_ (_10522_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  nor _18893_ (_10523_, _10482_, _10522_);
  and _18894_ (_10524_, _10482_, word_in[3]);
  or _18895_ (_10525_, _10524_, _10523_);
  or _18896_ (_10526_, _10525_, _10479_);
  or _18897_ (_10527_, _10487_, word_in[11]);
  and _18898_ (_10528_, _10527_, _10526_);
  or _18899_ (_10529_, _10528_, _10475_);
  or _18900_ (_10530_, _10476_, _09493_);
  and _18901_ (_10532_, _10530_, _10493_);
  and _18902_ (_10533_, _10532_, _10529_);
  and _18903_ (_10534_, _10474_, word_in[27]);
  or _18904_ (_08300_, _10534_, _10533_);
  not _18905_ (_10535_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  nor _18906_ (_10536_, _10482_, _10535_);
  and _18907_ (_10537_, _10482_, word_in[4]);
  or _18908_ (_10538_, _10537_, _10536_);
  or _18909_ (_10539_, _10538_, _10479_);
  or _18910_ (_10540_, _10487_, word_in[12]);
  and _18911_ (_10541_, _10540_, _10539_);
  or _18912_ (_10542_, _10541_, _10475_);
  or _18913_ (_10543_, _10476_, _09518_);
  and _18914_ (_10544_, _10543_, _10493_);
  and _18915_ (_10545_, _10544_, _10542_);
  and _18916_ (_10546_, _10474_, word_in[28]);
  or _18917_ (_08301_, _10546_, _10545_);
  not _18918_ (_10548_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  nor _18919_ (_10550_, _10482_, _10548_);
  and _18920_ (_10551_, _10482_, word_in[5]);
  or _18921_ (_10552_, _10551_, _10550_);
  or _18922_ (_10554_, _10552_, _10479_);
  or _18923_ (_10555_, _10487_, word_in[13]);
  and _18924_ (_10556_, _10555_, _10554_);
  or _18925_ (_10558_, _10556_, _10475_);
  or _18926_ (_10559_, _10476_, _09523_);
  and _18927_ (_10560_, _10559_, _10493_);
  and _18928_ (_10561_, _10560_, _10558_);
  and _18929_ (_10562_, _10474_, word_in[29]);
  or _18930_ (_08302_, _10562_, _10561_);
  or _18931_ (_10563_, _10476_, _09548_);
  not _18932_ (_10564_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  nor _18933_ (_10565_, _10482_, _10564_);
  and _18934_ (_10567_, _10482_, word_in[6]);
  or _18935_ (_10568_, _10567_, _10565_);
  or _18936_ (_10569_, _10568_, _10479_);
  or _18937_ (_10570_, _10487_, word_in[14]);
  and _18938_ (_10571_, _10570_, _10569_);
  or _18939_ (_10572_, _10571_, _10475_);
  and _18940_ (_10573_, _10572_, _10563_);
  or _18941_ (_10574_, _10573_, _10474_);
  or _18942_ (_10575_, _10493_, word_in[30]);
  and _18943_ (_08303_, _10575_, _10574_);
  nor _18944_ (_10576_, _10482_, _08560_);
  and _18945_ (_10577_, _10482_, word_in[7]);
  or _18946_ (_10578_, _10577_, _10576_);
  or _18947_ (_10579_, _10578_, _10479_);
  nand _18948_ (_10580_, _10479_, _08764_);
  and _18949_ (_10581_, _10580_, _10579_);
  or _18950_ (_10582_, _10581_, _10475_);
  or _18951_ (_10583_, _10476_, _08769_);
  and _18952_ (_10584_, _10583_, _10493_);
  and _18953_ (_10585_, _10584_, _10582_);
  and _18954_ (_10586_, _10474_, word_in[31]);
  or _18955_ (_08307_, _10586_, _10585_);
  and _18956_ (_10587_, _05676_, _04861_);
  nand _18957_ (_10588_, _10587_, _06369_);
  or _18958_ (_10589_, _10587_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  and _18959_ (_10590_, _10589_, _10588_);
  and _18960_ (_08362_, _10590_, _04856_);
  and _18961_ (_10591_, _09669_, _08625_);
  and _18962_ (_10592_, _08752_, _08523_);
  not _18963_ (_10593_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and _18964_ (_10594_, _10248_, _08755_);
  nor _18965_ (_10595_, _10594_, _10593_);
  and _18966_ (_10596_, _10594_, _09449_);
  or _18967_ (_10597_, _10596_, _10595_);
  or _18968_ (_10598_, _10597_, _10592_);
  not _18969_ (_10599_, _10592_);
  or _18970_ (_10600_, _10599_, word_in[8]);
  and _18971_ (_10601_, _10600_, _10598_);
  or _18972_ (_10602_, _10601_, _10591_);
  and _18973_ (_10603_, _10238_, _08548_);
  not _18974_ (_10604_, _10603_);
  not _18975_ (_10605_, _10591_);
  or _18976_ (_10606_, _10605_, _09349_);
  and _18977_ (_10607_, _10606_, _10604_);
  and _18978_ (_10608_, _10607_, _10602_);
  and _18979_ (_10609_, _10603_, word_in[24]);
  or _18980_ (_08374_, _10609_, _10608_);
  and _18981_ (_10610_, _10591_, _09464_);
  and _18982_ (_10611_, _10594_, _09466_);
  not _18983_ (_10612_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  nor _18984_ (_10613_, _10594_, _10612_);
  nor _18985_ (_10614_, _10613_, _10611_);
  nor _18986_ (_10615_, _10614_, _10592_);
  and _18987_ (_10616_, _10592_, word_in[9]);
  or _18988_ (_10617_, _10616_, _10615_);
  and _18989_ (_10618_, _10617_, _10605_);
  or _18990_ (_10619_, _10618_, _10610_);
  and _18991_ (_10620_, _10619_, _10604_);
  and _18992_ (_10621_, _10603_, word_in[25]);
  or _18993_ (_08379_, _10621_, _10620_);
  and _18994_ (_10622_, _10591_, _09478_);
  and _18995_ (_10623_, _10594_, _09480_);
  not _18996_ (_10624_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  nor _18997_ (_10625_, _10594_, _10624_);
  nor _18998_ (_10626_, _10625_, _10623_);
  nor _18999_ (_10627_, _10626_, _10592_);
  and _19000_ (_10628_, _10592_, word_in[10]);
  or _19001_ (_10629_, _10628_, _10627_);
  and _19002_ (_10630_, _10629_, _10605_);
  or _19003_ (_10631_, _10630_, _10622_);
  and _19004_ (_10632_, _10631_, _10604_);
  and _19005_ (_10633_, _10603_, word_in[26]);
  or _19006_ (_08384_, _10633_, _10632_);
  and _19007_ (_10634_, _10591_, _09493_);
  and _19008_ (_10635_, _10594_, _09495_);
  not _19009_ (_10636_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  nor _19010_ (_10637_, _10594_, _10636_);
  nor _19011_ (_10638_, _10637_, _10635_);
  nor _19012_ (_10639_, _10638_, _10592_);
  and _19013_ (_10640_, _10592_, word_in[11]);
  or _19014_ (_10641_, _10640_, _10639_);
  and _19015_ (_10642_, _10641_, _10605_);
  or _19016_ (_10643_, _10642_, _10634_);
  and _19017_ (_10644_, _10643_, _10604_);
  and _19018_ (_10645_, _10603_, word_in[27]);
  or _19019_ (_08388_, _10645_, _10644_);
  not _19020_ (_10646_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  nor _19021_ (_10647_, _10594_, _10646_);
  and _19022_ (_10648_, _10594_, _09510_);
  or _19023_ (_10649_, _10648_, _10647_);
  or _19024_ (_10650_, _10649_, _10592_);
  or _19025_ (_10651_, _10599_, word_in[12]);
  and _19026_ (_10652_, _10651_, _10650_);
  or _19027_ (_10653_, _10652_, _10591_);
  or _19028_ (_10654_, _10605_, _09518_);
  and _19029_ (_10655_, _10654_, _10604_);
  and _19030_ (_10656_, _10655_, _10653_);
  and _19031_ (_10657_, _10603_, word_in[28]);
  or _19032_ (_08391_, _10657_, _10656_);
  and _19033_ (_10658_, _10591_, _09523_);
  and _19034_ (_10659_, _10594_, _09525_);
  not _19035_ (_10660_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  nor _19036_ (_10661_, _10594_, _10660_);
  nor _19037_ (_10662_, _10661_, _10659_);
  nor _19038_ (_10663_, _10662_, _10592_);
  and _19039_ (_10664_, _10592_, word_in[13]);
  or _19040_ (_10665_, _10664_, _10663_);
  and _19041_ (_10666_, _10665_, _10605_);
  or _19042_ (_10667_, _10666_, _10658_);
  and _19043_ (_10668_, _10667_, _10604_);
  and _19044_ (_10669_, _10603_, word_in[29]);
  or _19045_ (_08395_, _10669_, _10668_);
  or _19046_ (_10670_, _10605_, _09548_);
  not _19047_ (_10671_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  nor _19048_ (_10672_, _10594_, _10671_);
  and _19049_ (_10673_, _10594_, _09541_);
  or _19050_ (_10674_, _10673_, _10672_);
  or _19051_ (_10676_, _10674_, _10592_);
  or _19052_ (_10677_, _10599_, word_in[14]);
  and _19053_ (_10678_, _10677_, _10676_);
  or _19054_ (_10679_, _10678_, _10591_);
  and _19055_ (_10680_, _10679_, _10670_);
  or _19056_ (_10681_, _10680_, _10603_);
  or _19057_ (_10682_, _10604_, word_in[30]);
  and _19058_ (_08400_, _10682_, _10681_);
  nor _19059_ (_10683_, _10594_, _08458_);
  and _19060_ (_10684_, _10594_, _08760_);
  or _19061_ (_10685_, _10684_, _10683_);
  or _19062_ (_10686_, _10685_, _10592_);
  nand _19063_ (_10687_, _10592_, _08764_);
  and _19064_ (_10688_, _10687_, _10686_);
  or _19065_ (_10689_, _10688_, _10591_);
  or _19066_ (_10690_, _10605_, _08769_);
  and _19067_ (_10691_, _10690_, _10604_);
  and _19068_ (_10692_, _10691_, _10689_);
  and _19069_ (_10693_, _10603_, word_in[31]);
  or _19070_ (_08402_, _10693_, _10692_);
  and _19071_ (_10694_, _08745_, _08511_);
  not _19072_ (_10695_, _10694_);
  and _19073_ (_10696_, _08749_, _08540_);
  and _19074_ (_10697_, _10696_, _09349_);
  not _19075_ (_10698_, _10696_);
  and _19076_ (_10699_, _08751_, _09179_);
  not _19077_ (_10700_, _10699_);
  and _19078_ (_10701_, _09785_, _08757_);
  and _19079_ (_10702_, _10701_, word_in[0]);
  not _19080_ (_10703_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  nor _19081_ (_10704_, _10701_, _10703_);
  or _19082_ (_10705_, _10704_, _10702_);
  and _19083_ (_10706_, _10705_, _10700_);
  and _19084_ (_10707_, _10699_, word_in[8]);
  or _19085_ (_10708_, _10707_, _10706_);
  and _19086_ (_10709_, _10708_, _10698_);
  or _19087_ (_10710_, _10709_, _10697_);
  and _19088_ (_10711_, _10710_, _10695_);
  and _19089_ (_10712_, _10694_, _09801_);
  or _19090_ (_08492_, _10712_, _10711_);
  and _19091_ (_10713_, _10696_, _09464_);
  not _19092_ (_10714_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  nor _19093_ (_10715_, _10701_, _10714_);
  and _19094_ (_10716_, _10701_, word_in[1]);
  or _19095_ (_10717_, _10716_, _10715_);
  and _19096_ (_10718_, _10717_, _10700_);
  and _19097_ (_10719_, _10699_, word_in[9]);
  or _19098_ (_10720_, _10719_, _10718_);
  and _19099_ (_10721_, _10720_, _10698_);
  or _19100_ (_10722_, _10721_, _10713_);
  and _19101_ (_10723_, _10722_, _10695_);
  and _19102_ (_10724_, _10694_, _09366_);
  or _19103_ (_08497_, _10724_, _10723_);
  and _19104_ (_10725_, _10696_, _09478_);
  not _19105_ (_10726_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  nor _19106_ (_10727_, _10701_, _10726_);
  and _19107_ (_10728_, _10701_, word_in[2]);
  or _19108_ (_10729_, _10728_, _10727_);
  and _19109_ (_10730_, _10729_, _10700_);
  and _19110_ (_10731_, _10699_, word_in[10]);
  or _19111_ (_10732_, _10731_, _10730_);
  and _19112_ (_10733_, _10732_, _10698_);
  or _19113_ (_10734_, _10733_, _10725_);
  and _19114_ (_10735_, _10734_, _10695_);
  and _19115_ (_10736_, _10694_, _09368_);
  or _19116_ (_08499_, _10736_, _10735_);
  not _19117_ (_10737_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  nor _19118_ (_10738_, _10701_, _10737_);
  and _19119_ (_10739_, _10701_, word_in[3]);
  or _19120_ (_10740_, _10739_, _10738_);
  and _19121_ (_10741_, _10740_, _10700_);
  and _19122_ (_10742_, _10699_, word_in[11]);
  or _19123_ (_10743_, _10742_, _10741_);
  and _19124_ (_10744_, _10743_, _10698_);
  and _19125_ (_10745_, _10696_, _09493_);
  or _19126_ (_10746_, _10745_, _10694_);
  or _19127_ (_10747_, _10746_, _10744_);
  or _19128_ (_10748_, _10695_, _09380_);
  and _19129_ (_08501_, _10748_, _10747_);
  not _19130_ (_10749_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  nor _19131_ (_10750_, _10701_, _10749_);
  and _19132_ (_10751_, _10701_, word_in[4]);
  or _19133_ (_10752_, _10751_, _10750_);
  and _19134_ (_10753_, _10752_, _10700_);
  and _19135_ (_10754_, _10699_, word_in[12]);
  or _19136_ (_10755_, _10754_, _10753_);
  and _19137_ (_10756_, _10755_, _10698_);
  and _19138_ (_10757_, _10696_, _09518_);
  or _19139_ (_10758_, _10757_, _10694_);
  or _19140_ (_10759_, _10758_, _10756_);
  or _19141_ (_10760_, _10695_, _09402_);
  and _19142_ (_08504_, _10760_, _10759_);
  and _19143_ (_10762_, _10696_, _09523_);
  not _19144_ (_10763_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  nor _19145_ (_10764_, _10701_, _10763_);
  and _19146_ (_10765_, _10701_, word_in[5]);
  or _19147_ (_10766_, _10765_, _10764_);
  and _19148_ (_10767_, _10766_, _10700_);
  and _19149_ (_10768_, _10699_, word_in[13]);
  or _19150_ (_10769_, _10768_, _10767_);
  and _19151_ (_10770_, _10769_, _10698_);
  or _19152_ (_10771_, _10770_, _10762_);
  and _19153_ (_10772_, _10771_, _10695_);
  and _19154_ (_10773_, _10694_, _09414_);
  or _19155_ (_08508_, _10773_, _10772_);
  and _19156_ (_10774_, _10696_, _09548_);
  not _19157_ (_10775_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  nor _19158_ (_10776_, _10701_, _10775_);
  and _19159_ (_10777_, _10701_, word_in[6]);
  or _19160_ (_10778_, _10777_, _10776_);
  and _19161_ (_10779_, _10778_, _10700_);
  and _19162_ (_10780_, _10699_, word_in[14]);
  or _19163_ (_10781_, _10780_, _10779_);
  and _19164_ (_10782_, _10781_, _10698_);
  or _19165_ (_10783_, _10782_, _10774_);
  and _19166_ (_10784_, _10783_, _10695_);
  and _19167_ (_10785_, _10694_, _09426_);
  or _19168_ (_08510_, _10785_, _10784_);
  and _19169_ (_10786_, _10696_, _08769_);
  nor _19170_ (_10787_, _10701_, _08579_);
  and _19171_ (_10788_, _10701_, word_in[7]);
  or _19172_ (_10789_, _10788_, _10787_);
  and _19173_ (_10790_, _10789_, _10700_);
  and _19174_ (_10791_, _10699_, word_in[15]);
  or _19175_ (_10792_, _10791_, _10790_);
  and _19176_ (_10793_, _10792_, _10698_);
  or _19177_ (_10794_, _10793_, _10786_);
  and _19178_ (_10795_, _10794_, _10695_);
  and _19179_ (_10796_, _10694_, _08774_);
  or _19180_ (_08513_, _10796_, _10795_);
  nand _19181_ (_10797_, _10587_, _06032_);
  or _19182_ (_10798_, _10587_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  and _19183_ (_10799_, _10798_, _04856_);
  and _19184_ (_08582_, _10799_, _10797_);
  and _19185_ (_10800_, _08745_, _08540_);
  not _19186_ (_10801_, _10800_);
  and _19187_ (_10802_, _08749_, _08514_);
  and _19188_ (_10803_, _10802_, _09349_);
  not _19189_ (_10804_, _10802_);
  and _19190_ (_10805_, _09441_, _08573_);
  and _19191_ (_10806_, _09445_, _08757_);
  and _19192_ (_10807_, _10806_, word_in[0]);
  not _19193_ (_10808_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  nor _19194_ (_10809_, _10806_, _10808_);
  nor _19195_ (_10810_, _10809_, _10807_);
  nor _19196_ (_10811_, _10810_, _10805_);
  and _19197_ (_10812_, _10805_, word_in[8]);
  or _19198_ (_10813_, _10812_, _10811_);
  and _19199_ (_10814_, _10813_, _10804_);
  or _19200_ (_10815_, _10814_, _10803_);
  and _19201_ (_10817_, _10815_, _10801_);
  and _19202_ (_10818_, _10800_, _09801_);
  or _19203_ (_13238_, _10818_, _10817_);
  not _19204_ (_10819_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  nor _19205_ (_10820_, _10806_, _10819_);
  and _19206_ (_10821_, _10806_, _09466_);
  or _19207_ (_10822_, _10821_, _10820_);
  or _19208_ (_10823_, _10822_, _10805_);
  not _19209_ (_10824_, _10805_);
  or _19210_ (_10825_, _10824_, word_in[9]);
  and _19211_ (_10826_, _10825_, _10823_);
  and _19212_ (_10827_, _10826_, _10804_);
  and _19213_ (_10828_, _10802_, _09464_);
  or _19214_ (_10829_, _10828_, _10800_);
  or _19215_ (_10830_, _10829_, _10827_);
  or _19216_ (_10831_, _10801_, _09366_);
  and _19217_ (_13239_, _10831_, _10830_);
  and _19218_ (_10832_, _10806_, word_in[2]);
  not _19219_ (_10833_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  nor _19220_ (_10834_, _10806_, _10833_);
  nor _19221_ (_10835_, _10834_, _10832_);
  nor _19222_ (_10836_, _10835_, _10805_);
  and _19223_ (_10837_, _10805_, word_in[10]);
  or _19224_ (_10838_, _10837_, _10836_);
  and _19225_ (_10839_, _10838_, _10804_);
  and _19226_ (_10840_, _10802_, _09478_);
  or _19227_ (_10841_, _10840_, _10800_);
  or _19228_ (_10842_, _10841_, _10839_);
  or _19229_ (_10843_, _10801_, _09368_);
  and _19230_ (_13240_, _10843_, _10842_);
  not _19231_ (_10844_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  nor _19232_ (_10845_, _10806_, _10844_);
  and _19233_ (_10846_, _10806_, _09495_);
  or _19234_ (_10847_, _10846_, _10845_);
  or _19235_ (_10848_, _10847_, _10805_);
  or _19236_ (_10849_, _10824_, word_in[11]);
  and _19237_ (_10851_, _10849_, _10848_);
  or _19238_ (_10852_, _10851_, _10802_);
  or _19239_ (_10853_, _10804_, _09493_);
  and _19240_ (_10854_, _10853_, _10852_);
  or _19241_ (_10855_, _10854_, _10800_);
  or _19242_ (_10856_, _10801_, _09380_);
  and _19243_ (_13241_, _10856_, _10855_);
  not _19244_ (_10857_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  nor _19245_ (_10858_, _10806_, _10857_);
  and _19246_ (_10859_, _10806_, _09510_);
  or _19247_ (_10860_, _10859_, _10858_);
  or _19248_ (_10861_, _10860_, _10805_);
  or _19249_ (_10862_, _10824_, word_in[12]);
  and _19250_ (_10863_, _10862_, _10861_);
  or _19251_ (_10864_, _10863_, _10802_);
  or _19252_ (_10865_, _10804_, _09518_);
  and _19253_ (_10867_, _10865_, _10864_);
  or _19254_ (_10868_, _10867_, _10800_);
  or _19255_ (_10870_, _10801_, _09402_);
  and _19256_ (_13242_, _10870_, _10868_);
  not _19257_ (_10871_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  nor _19258_ (_10872_, _10806_, _10871_);
  and _19259_ (_10873_, _10806_, _09525_);
  or _19260_ (_10874_, _10873_, _10872_);
  or _19261_ (_10875_, _10874_, _10805_);
  or _19262_ (_10876_, _10824_, word_in[13]);
  and _19263_ (_10877_, _10876_, _10875_);
  or _19264_ (_10878_, _10877_, _10802_);
  or _19265_ (_10879_, _10804_, _09523_);
  and _19266_ (_10880_, _10879_, _10878_);
  or _19267_ (_10881_, _10880_, _10800_);
  or _19268_ (_10882_, _10801_, _09414_);
  and _19269_ (_13243_, _10882_, _10881_);
  not _19270_ (_10884_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  nor _19271_ (_10885_, _10806_, _10884_);
  and _19272_ (_10886_, _10806_, _09541_);
  or _19273_ (_10887_, _10886_, _10885_);
  or _19274_ (_10888_, _10887_, _10805_);
  or _19275_ (_10890_, _10824_, word_in[14]);
  and _19276_ (_10891_, _10890_, _10888_);
  or _19277_ (_10892_, _10891_, _10802_);
  or _19278_ (_10894_, _10804_, _09548_);
  and _19279_ (_10895_, _10894_, _10892_);
  or _19280_ (_10896_, _10895_, _10800_);
  or _19281_ (_10897_, _10801_, _09426_);
  and _19282_ (_13244_, _10897_, _10896_);
  nor _19283_ (_10898_, _10806_, _08464_);
  and _19284_ (_10899_, _10806_, _08760_);
  or _19285_ (_10900_, _10899_, _10898_);
  or _19286_ (_10901_, _10900_, _10805_);
  nand _19287_ (_10903_, _10805_, _08764_);
  and _19288_ (_10904_, _10903_, _10901_);
  or _19289_ (_10905_, _10904_, _10802_);
  or _19290_ (_10906_, _10804_, _08769_);
  and _19291_ (_10907_, _10906_, _10905_);
  or _19292_ (_10909_, _10907_, _10800_);
  or _19293_ (_10910_, _10801_, _08774_);
  and _19294_ (_13245_, _10910_, _10909_);
  and _19295_ (_10912_, _08745_, _08514_);
  not _19296_ (_10913_, _10912_);
  and _19297_ (_10914_, _08749_, _08548_);
  and _19298_ (_10915_, _10914_, _09349_);
  not _19299_ (_10916_, _10914_);
  and _19300_ (_10917_, _09569_, _08573_);
  and _19301_ (_10918_, _09572_, _08741_);
  and _19302_ (_10920_, _10918_, word_in[0]);
  not _19303_ (_10921_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  nor _19304_ (_10922_, _10918_, _10921_);
  nor _19305_ (_10923_, _10922_, _10920_);
  nor _19306_ (_10924_, _10923_, _10917_);
  and _19307_ (_10925_, _10917_, word_in[8]);
  or _19308_ (_10926_, _10925_, _10924_);
  and _19309_ (_10927_, _10926_, _10916_);
  or _19310_ (_10928_, _10927_, _10915_);
  and _19311_ (_10929_, _10928_, _10913_);
  and _19312_ (_10930_, _10912_, _09801_);
  or _19313_ (_13246_, _10930_, _10929_);
  not _19314_ (_10931_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  nor _19315_ (_10932_, _10918_, _10931_);
  and _19316_ (_10933_, _10918_, word_in[1]);
  nor _19317_ (_10934_, _10933_, _10932_);
  nor _19318_ (_10935_, _10934_, _10917_);
  and _19319_ (_10936_, _10917_, word_in[9]);
  or _19320_ (_10937_, _10936_, _10935_);
  and _19321_ (_10938_, _10937_, _10916_);
  and _19322_ (_10939_, _10914_, _09464_);
  or _19323_ (_10940_, _10939_, _10912_);
  or _19324_ (_10941_, _10940_, _10938_);
  or _19325_ (_10942_, _10913_, _09366_);
  and _19326_ (_08691_, _10942_, _10941_);
  not _19327_ (_10943_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  nor _19328_ (_10944_, _10918_, _10943_);
  and _19329_ (_10945_, _10918_, word_in[2]);
  or _19330_ (_10946_, _10945_, _10944_);
  or _19331_ (_10947_, _10946_, _10917_);
  not _19332_ (_10948_, _10917_);
  or _19333_ (_10949_, _10948_, word_in[10]);
  and _19334_ (_10950_, _10949_, _10947_);
  or _19335_ (_10951_, _10950_, _10914_);
  or _19336_ (_10952_, _10916_, _09478_);
  and _19337_ (_10953_, _10952_, _10951_);
  or _19338_ (_10954_, _10953_, _10912_);
  or _19339_ (_10955_, _10913_, _09368_);
  and _19340_ (_08694_, _10955_, _10954_);
  or _19341_ (_10956_, _10948_, word_in[11]);
  not _19342_ (_10957_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  nor _19343_ (_10958_, _10918_, _10957_);
  and _19344_ (_10959_, _10918_, word_in[3]);
  or _19345_ (_10960_, _10959_, _10958_);
  or _19346_ (_10961_, _10960_, _10917_);
  and _19347_ (_10962_, _10961_, _10956_);
  or _19348_ (_10963_, _10962_, _10914_);
  or _19349_ (_10964_, _10916_, _09493_);
  and _19350_ (_10965_, _10964_, _10963_);
  or _19351_ (_10966_, _10965_, _10912_);
  or _19352_ (_10967_, _10913_, _09380_);
  and _19353_ (_08697_, _10967_, _10966_);
  not _19354_ (_10968_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  nor _19355_ (_10969_, _10918_, _10968_);
  and _19356_ (_10970_, _10918_, word_in[4]);
  nor _19357_ (_10971_, _10970_, _10969_);
  nor _19358_ (_10972_, _10971_, _10917_);
  and _19359_ (_10973_, _10917_, word_in[12]);
  or _19360_ (_10974_, _10973_, _10972_);
  and _19361_ (_10975_, _10974_, _10916_);
  and _19362_ (_10976_, _10914_, _09518_);
  or _19363_ (_10977_, _10976_, _10912_);
  or _19364_ (_10978_, _10977_, _10975_);
  or _19365_ (_10979_, _10913_, _09402_);
  and _19366_ (_13247_, _10979_, _10978_);
  or _19367_ (_10980_, _10916_, _09523_);
  not _19368_ (_10981_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  nor _19369_ (_10982_, _10918_, _10981_);
  and _19370_ (_10983_, _10918_, word_in[5]);
  or _19371_ (_10984_, _10983_, _10982_);
  or _19372_ (_10985_, _10984_, _10917_);
  or _19373_ (_10986_, _10948_, word_in[13]);
  and _19374_ (_10987_, _10986_, _10985_);
  or _19375_ (_10988_, _10987_, _10914_);
  and _19376_ (_10989_, _10988_, _10980_);
  or _19377_ (_10990_, _10989_, _10912_);
  or _19378_ (_10991_, _10913_, _09414_);
  and _19379_ (_08702_, _10991_, _10990_);
  and _19380_ (_10993_, _10914_, _09548_);
  not _19381_ (_10994_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  nor _19382_ (_10995_, _10918_, _10994_);
  and _19383_ (_10996_, _10918_, word_in[6]);
  nor _19384_ (_10997_, _10996_, _10995_);
  nor _19385_ (_10998_, _10997_, _10917_);
  and _19386_ (_10999_, _10917_, word_in[14]);
  or _19387_ (_11000_, _10999_, _10998_);
  and _19388_ (_11001_, _11000_, _10916_);
  or _19389_ (_11002_, _11001_, _10993_);
  and _19390_ (_11003_, _11002_, _10913_);
  and _19391_ (_11004_, _10912_, _09426_);
  or _19392_ (_08705_, _11004_, _11003_);
  nand _19393_ (_11005_, _10917_, _08764_);
  nor _19394_ (_11006_, _10918_, _08574_);
  and _19395_ (_11007_, _10918_, word_in[7]);
  or _19396_ (_11008_, _11007_, _11006_);
  or _19397_ (_11009_, _11008_, _10917_);
  and _19398_ (_11010_, _11009_, _11005_);
  or _19399_ (_11011_, _11010_, _10914_);
  or _19400_ (_11012_, _10916_, _08769_);
  and _19401_ (_11013_, _11012_, _11011_);
  or _19402_ (_11014_, _11013_, _10912_);
  or _19403_ (_11015_, _10913_, _08774_);
  and _19404_ (_08709_, _11015_, _11014_);
  and _19405_ (_11016_, _08758_, word_in[0]);
  not _19406_ (_11017_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  nor _19407_ (_11018_, _08758_, _11017_);
  nor _19408_ (_11019_, _11018_, _11016_);
  nor _19409_ (_11020_, _11019_, _08753_);
  and _19410_ (_11021_, _08753_, word_in[8]);
  or _19411_ (_11022_, _11021_, _11020_);
  and _19412_ (_11023_, _11022_, _08768_);
  and _19413_ (_11024_, _09349_, _08750_);
  or _19414_ (_11025_, _11024_, _11023_);
  and _19415_ (_11026_, _11025_, _08773_);
  and _19416_ (_11027_, _09801_, _08746_);
  or _19417_ (_13248_, _11027_, _11026_);
  not _19418_ (_11028_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  nor _19419_ (_11029_, _08758_, _11028_);
  and _19420_ (_11030_, _09466_, _08758_);
  or _19421_ (_11031_, _11030_, _11029_);
  or _19422_ (_11032_, _11031_, _08753_);
  not _19423_ (_11033_, _08753_);
  or _19424_ (_11034_, _11033_, word_in[9]);
  and _19425_ (_11035_, _11034_, _11032_);
  or _19426_ (_11036_, _11035_, _08750_);
  or _19427_ (_11037_, _09464_, _08768_);
  and _19428_ (_11038_, _11037_, _11036_);
  or _19429_ (_11039_, _11038_, _08746_);
  or _19430_ (_11040_, _09366_, _08773_);
  and _19431_ (_13249_, _11040_, _11039_);
  and _19432_ (_11041_, _08758_, word_in[2]);
  not _19433_ (_11043_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  nor _19434_ (_11044_, _08758_, _11043_);
  nor _19435_ (_11045_, _11044_, _11041_);
  nor _19436_ (_11046_, _11045_, _08753_);
  and _19437_ (_11047_, _08753_, word_in[10]);
  or _19438_ (_11048_, _11047_, _11046_);
  and _19439_ (_11049_, _11048_, _08768_);
  and _19440_ (_11050_, _09478_, _08750_);
  or _19441_ (_11051_, _11050_, _11049_);
  and _19442_ (_11052_, _11051_, _08773_);
  and _19443_ (_11053_, _09368_, _08746_);
  or _19444_ (_13250_, _11053_, _11052_);
  and _19445_ (_11054_, _08758_, word_in[3]);
  not _19446_ (_11056_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  nor _19447_ (_11057_, _08758_, _11056_);
  nor _19448_ (_11059_, _11057_, _11054_);
  nor _19449_ (_11060_, _11059_, _08753_);
  and _19450_ (_11061_, _08753_, word_in[11]);
  or _19451_ (_11062_, _11061_, _11060_);
  and _19452_ (_11063_, _11062_, _08768_);
  and _19453_ (_11064_, _09493_, _08750_);
  or _19454_ (_11065_, _11064_, _11063_);
  and _19455_ (_11066_, _11065_, _08773_);
  and _19456_ (_11067_, _09380_, _08746_);
  or _19457_ (_13251_, _11067_, _11066_);
  not _19458_ (_11068_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  nor _19459_ (_11069_, _08758_, _11068_);
  and _19460_ (_11070_, _09510_, _08758_);
  or _19461_ (_11071_, _11070_, _11069_);
  or _19462_ (_11072_, _11071_, _08753_);
  or _19463_ (_11073_, _11033_, word_in[12]);
  and _19464_ (_11074_, _11073_, _11072_);
  or _19465_ (_11075_, _11074_, _08750_);
  or _19466_ (_11076_, _09518_, _08768_);
  and _19467_ (_11077_, _11076_, _11075_);
  or _19468_ (_11078_, _11077_, _08746_);
  or _19469_ (_11079_, _09402_, _08773_);
  and _19470_ (_13252_, _11079_, _11078_);
  not _19471_ (_11080_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  nor _19472_ (_11081_, _08758_, _11080_);
  and _19473_ (_11082_, _09525_, _08758_);
  or _19474_ (_11083_, _11082_, _11081_);
  or _19475_ (_11084_, _11083_, _08753_);
  or _19476_ (_11085_, _11033_, word_in[13]);
  and _19477_ (_11086_, _11085_, _11084_);
  or _19478_ (_11087_, _11086_, _08750_);
  or _19479_ (_11088_, _09523_, _08768_);
  and _19480_ (_11090_, _11088_, _11087_);
  or _19481_ (_11091_, _11090_, _08746_);
  or _19482_ (_11092_, _09414_, _08773_);
  and _19483_ (_13253_, _11092_, _11091_);
  not _19484_ (_11093_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  nor _19485_ (_11094_, _08758_, _11093_);
  and _19486_ (_11095_, _09541_, _08758_);
  or _19487_ (_11096_, _11095_, _11094_);
  or _19488_ (_11097_, _11096_, _08753_);
  or _19489_ (_11098_, _11033_, word_in[14]);
  and _19490_ (_11099_, _11098_, _11097_);
  or _19491_ (_11100_, _11099_, _08750_);
  or _19492_ (_11101_, _09548_, _08768_);
  and _19493_ (_11102_, _11101_, _11100_);
  or _19494_ (_11103_, _11102_, _08746_);
  or _19495_ (_11104_, _09426_, _08773_);
  and _19496_ (_13254_, _11104_, _11103_);
  and _19497_ (_11105_, _06410_, _05671_);
  and _19498_ (_11106_, _06696_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  or _19499_ (_11107_, _11106_, _11105_);
  and _19500_ (_08879_, _11107_, _04856_);
  nor _19501_ (_08881_, _07651_, rst);
  and _19502_ (_11108_, _08277_, _04986_);
  nand _19503_ (_11109_, _11108_, _06088_);
  or _19504_ (_11110_, _11108_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and _19505_ (_11111_, _11110_, _06935_);
  and _19506_ (_11112_, _11111_, _11109_);
  and _19507_ (_11113_, _06934_, _06033_);
  or _19508_ (_11114_, _11113_, _11112_);
  and _19509_ (_09036_, _11114_, _04856_);
  and _19510_ (_11115_, _06688_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  and _19511_ (_11116_, _06686_, _05718_);
  or _19512_ (_11117_, _11116_, _11115_);
  and _19513_ (_09073_, _11117_, _04856_);
  and _19514_ (_11118_, _06705_, _05671_);
  and _19515_ (_11119_, _06696_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  or _19516_ (_11120_, _11119_, _11118_);
  and _19517_ (_09492_, _11120_, _04856_);
  or _19518_ (_11121_, _05793_, _06812_);
  or _19519_ (_11122_, _05729_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and _19520_ (_11123_, _11122_, _04856_);
  and _19521_ (_09513_, _11123_, _11121_);
  or _19522_ (_11124_, _05818_, _06812_);
  or _19523_ (_11125_, _05729_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and _19524_ (_11126_, _11125_, _04856_);
  and _19525_ (_09521_, _11126_, _11124_);
  or _19526_ (_11127_, _05870_, _06812_);
  or _19527_ (_11128_, _05729_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and _19528_ (_11129_, _11128_, _04856_);
  and _19529_ (_09529_, _11129_, _11127_);
  and _19530_ (_11130_, _08451_, word_in[0]);
  nand _19531_ (_11131_, _08361_, _10357_);
  or _19532_ (_11132_, _08361_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  and _19533_ (_11133_, _11132_, _11131_);
  and _19534_ (_11134_, _11133_, _08416_);
  or _19535_ (_11135_, _11134_, _08425_);
  nand _19536_ (_11136_, _08361_, _10808_);
  or _19537_ (_11137_, _08361_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  and _19538_ (_11138_, _11137_, _11136_);
  and _19539_ (_11139_, _11138_, _08393_);
  nand _19540_ (_11140_, _08361_, _11017_);
  or _19541_ (_11141_, _08361_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and _19542_ (_11142_, _11141_, _11140_);
  and _19543_ (_11143_, _11142_, _08406_);
  nand _19544_ (_11144_, _08361_, _10593_);
  or _19545_ (_11145_, _08361_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and _19546_ (_11146_, _11145_, _11144_);
  and _19547_ (_11147_, _11146_, _08397_);
  or _19548_ (_11148_, _11147_, _11143_);
  or _19549_ (_11149_, _11148_, _11139_);
  or _19550_ (_11151_, _11149_, _11135_);
  nand _19551_ (_11152_, _08361_, _09443_);
  or _19552_ (_11153_, _08361_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  and _19553_ (_11154_, _11153_, _11152_);
  and _19554_ (_11155_, _11154_, _08416_);
  or _19555_ (_11156_, _11155_, _08375_);
  nand _19556_ (_11157_, _08361_, _09900_);
  or _19557_ (_11158_, _08361_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  and _19558_ (_11159_, _11158_, _11157_);
  and _19559_ (_11160_, _11159_, _08393_);
  nand _19560_ (_11161_, _08361_, _10123_);
  or _19561_ (_11162_, _08361_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  and _19562_ (_11163_, _11162_, _11161_);
  and _19563_ (_11164_, _11163_, _08406_);
  nand _19564_ (_11165_, _08361_, _09676_);
  or _19565_ (_11166_, _08361_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  and _19566_ (_11167_, _11166_, _11165_);
  and _19567_ (_11168_, _11167_, _08397_);
  or _19568_ (_11169_, _11168_, _11164_);
  or _19569_ (_11170_, _11169_, _11160_);
  or _19570_ (_11171_, _11170_, _11156_);
  and _19571_ (_11172_, _11171_, _11151_);
  and _19572_ (_11173_, _11172_, _08450_);
  or _19573_ (\oc8051_symbolic_cxrom1.cxrom_data_out [0], _11173_, _11130_);
  and _19574_ (_11175_, _08451_, word_in[1]);
  nand _19575_ (_11176_, _08361_, _10373_);
  or _19576_ (_11177_, _08361_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  and _19577_ (_11178_, _11177_, _11176_);
  and _19578_ (_11179_, _11178_, _08416_);
  nand _19579_ (_11180_, _08361_, _10612_);
  or _19580_ (_11181_, _08361_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  and _19581_ (_11182_, _11181_, _11180_);
  and _19582_ (_11183_, _11182_, _08397_);
  nand _19583_ (_11184_, _08361_, _10819_);
  or _19584_ (_11185_, _08361_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  and _19585_ (_11186_, _11185_, _11184_);
  and _19586_ (_11187_, _11186_, _08393_);
  or _19587_ (_11188_, _11187_, _11183_);
  or _19588_ (_11189_, _11188_, _11179_);
  nand _19589_ (_11190_, _08361_, _11028_);
  or _19590_ (_11191_, _08361_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  and _19591_ (_11192_, _11191_, _11190_);
  and _19592_ (_11193_, _11192_, _08406_);
  or _19593_ (_11194_, _11193_, _08425_);
  or _19594_ (_11195_, _11194_, _11189_);
  nand _19595_ (_11196_, _08361_, _09468_);
  or _19596_ (_11197_, _08361_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  and _19597_ (_11198_, _11197_, _11196_);
  and _19598_ (_11199_, _11198_, _08416_);
  nand _19599_ (_11200_, _08361_, _09691_);
  or _19600_ (_11201_, _08361_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  and _19601_ (_11202_, _11201_, _11200_);
  and _19602_ (_11203_, _11202_, _08397_);
  nand _19603_ (_11204_, _08361_, _09911_);
  or _19604_ (_11205_, _08361_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  and _19605_ (_11206_, _11205_, _11204_);
  and _19606_ (_11207_, _11206_, _08393_);
  or _19607_ (_11208_, _11207_, _11203_);
  or _19608_ (_11209_, _11208_, _11199_);
  nand _19609_ (_11210_, _08361_, _10134_);
  or _19610_ (_11211_, _08361_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  and _19611_ (_11212_, _11211_, _11210_);
  and _19612_ (_11213_, _11212_, _08406_);
  or _19613_ (_11214_, _11213_, _08375_);
  or _19614_ (_11215_, _11214_, _11209_);
  and _19615_ (_11216_, _11215_, _11195_);
  and _19616_ (_11217_, _11216_, _08450_);
  or _19617_ (\oc8051_symbolic_cxrom1.cxrom_data_out [1], _11217_, _11175_);
  and _19618_ (_11218_, _08451_, word_in[2]);
  nand _19619_ (_11219_, _08361_, _10386_);
  or _19620_ (_11220_, _08361_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  and _19621_ (_11221_, _11220_, _11219_);
  and _19622_ (_11222_, _11221_, _08416_);
  or _19623_ (_11223_, _11222_, _08425_);
  nand _19624_ (_11224_, _08361_, _10833_);
  or _19625_ (_11225_, _08361_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  and _19626_ (_11226_, _11225_, _11224_);
  and _19627_ (_11227_, _11226_, _08393_);
  nand _19628_ (_11228_, _08361_, _11043_);
  or _19629_ (_11229_, _08361_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  and _19630_ (_11230_, _11229_, _11228_);
  and _19631_ (_11231_, _11230_, _08406_);
  nand _19632_ (_11232_, _08361_, _10624_);
  or _19633_ (_11233_, _08361_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  and _19634_ (_11234_, _11233_, _11232_);
  and _19635_ (_11235_, _11234_, _08397_);
  or _19636_ (_11237_, _11235_, _11231_);
  or _19637_ (_11238_, _11237_, _11227_);
  or _19638_ (_11239_, _11238_, _11223_);
  nand _19639_ (_11240_, _08361_, _09482_);
  or _19640_ (_11241_, _08361_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  and _19641_ (_11242_, _11241_, _11240_);
  and _19642_ (_11243_, _11242_, _08416_);
  or _19643_ (_11244_, _11243_, _08375_);
  nand _19644_ (_11245_, _08361_, _09924_);
  or _19645_ (_11246_, _08361_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  and _19646_ (_11248_, _11246_, _11245_);
  and _19647_ (_11249_, _11248_, _08393_);
  nand _19648_ (_11250_, _08361_, _10149_);
  or _19649_ (_11251_, _08361_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  and _19650_ (_11252_, _11251_, _11250_);
  and _19651_ (_11253_, _11252_, _08406_);
  nand _19652_ (_11254_, _08361_, _09702_);
  or _19653_ (_11255_, _08361_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  and _19654_ (_11256_, _11255_, _11254_);
  and _19655_ (_11257_, _11256_, _08397_);
  or _19656_ (_11258_, _11257_, _11253_);
  or _19657_ (_11259_, _11258_, _11249_);
  or _19658_ (_11260_, _11259_, _11244_);
  and _19659_ (_11261_, _11260_, _11239_);
  and _19660_ (_11262_, _11261_, _08450_);
  or _19661_ (\oc8051_symbolic_cxrom1.cxrom_data_out [2], _11262_, _11218_);
  and _19662_ (_11263_, _08451_, word_in[3]);
  nand _19663_ (_11264_, _08361_, _10398_);
  or _19664_ (_11265_, _08361_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  and _19665_ (_11266_, _11265_, _11264_);
  and _19666_ (_11267_, _11266_, _08416_);
  nand _19667_ (_11268_, _08361_, _10636_);
  or _19668_ (_11269_, _08361_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  and _19669_ (_11270_, _11269_, _11268_);
  and _19670_ (_11271_, _11270_, _08397_);
  nand _19671_ (_11272_, _08361_, _10844_);
  or _19672_ (_11273_, _08361_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  and _19673_ (_11274_, _11273_, _11272_);
  and _19674_ (_11275_, _11274_, _08393_);
  or _19675_ (_11276_, _11275_, _11271_);
  or _19676_ (_11277_, _11276_, _11267_);
  nand _19677_ (_11278_, _08361_, _11056_);
  or _19678_ (_11279_, _08361_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  and _19679_ (_11280_, _11279_, _11278_);
  and _19680_ (_11281_, _11280_, _08406_);
  or _19681_ (_11282_, _11281_, _08425_);
  or _19682_ (_11283_, _11282_, _11277_);
  nand _19683_ (_11284_, _08361_, _09497_);
  or _19684_ (_11285_, _08361_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  and _19685_ (_11286_, _11285_, _11284_);
  and _19686_ (_11287_, _11286_, _08416_);
  nand _19687_ (_11288_, _08361_, _09715_);
  or _19688_ (_11289_, _08361_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  and _19689_ (_11290_, _11289_, _11288_);
  and _19690_ (_11291_, _11290_, _08397_);
  nand _19691_ (_11293_, _08361_, _09939_);
  or _19692_ (_11294_, _08361_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  and _19693_ (_11295_, _11294_, _11293_);
  and _19694_ (_11296_, _11295_, _08393_);
  or _19695_ (_11297_, _11296_, _11291_);
  or _19696_ (_11298_, _11297_, _11287_);
  nand _19697_ (_11299_, _08361_, _10160_);
  or _19698_ (_11300_, _08361_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  and _19699_ (_11301_, _11300_, _11299_);
  and _19700_ (_11302_, _11301_, _08406_);
  or _19701_ (_11303_, _11302_, _08375_);
  or _19702_ (_11304_, _11303_, _11298_);
  and _19703_ (_11305_, _11304_, _11283_);
  and _19704_ (_11306_, _11305_, _08450_);
  or _19705_ (\oc8051_symbolic_cxrom1.cxrom_data_out [3], _11306_, _11263_);
  and _19706_ (_11307_, _08451_, word_in[4]);
  nand _19707_ (_11308_, _08361_, _10409_);
  or _19708_ (_11309_, _08361_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  and _19709_ (_11310_, _11309_, _11308_);
  and _19710_ (_11311_, _11310_, _08416_);
  nand _19711_ (_11313_, _08361_, _10646_);
  or _19712_ (_11314_, _08361_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  and _19713_ (_11315_, _11314_, _11313_);
  and _19714_ (_11316_, _11315_, _08397_);
  nand _19715_ (_11317_, _08361_, _10857_);
  or _19716_ (_11318_, _08361_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  and _19717_ (_11319_, _11318_, _11317_);
  and _19718_ (_11320_, _11319_, _08393_);
  or _19719_ (_11321_, _11320_, _11316_);
  or _19720_ (_11322_, _11321_, _11311_);
  nand _19721_ (_11323_, _08361_, _11068_);
  or _19722_ (_11324_, _08361_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  and _19723_ (_11325_, _11324_, _11323_);
  and _19724_ (_11326_, _11325_, _08406_);
  or _19725_ (_11328_, _11326_, _08425_);
  or _19726_ (_11329_, _11328_, _11322_);
  nand _19727_ (_11330_, _08361_, _09508_);
  or _19728_ (_11331_, _08361_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  and _19729_ (_11332_, _11331_, _11330_);
  and _19730_ (_11333_, _11332_, _08416_);
  nand _19731_ (_11334_, _08361_, _09728_);
  or _19732_ (_11335_, _08361_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  and _19733_ (_11336_, _11335_, _11334_);
  and _19734_ (_11337_, _11336_, _08397_);
  nand _19735_ (_11338_, _08361_, _09961_);
  or _19736_ (_11339_, _08361_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  and _19737_ (_11340_, _11339_, _11338_);
  and _19738_ (_11341_, _11340_, _08393_);
  or _19739_ (_11342_, _11341_, _11337_);
  or _19740_ (_11344_, _11342_, _11333_);
  nand _19741_ (_11345_, _08361_, _10175_);
  or _19742_ (_11346_, _08361_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  and _19743_ (_11348_, _11346_, _11345_);
  and _19744_ (_11349_, _11348_, _08406_);
  or _19745_ (_11351_, _11349_, _08375_);
  or _19746_ (_11352_, _11351_, _11344_);
  and _19747_ (_11353_, _11352_, _11329_);
  and _19748_ (_11354_, _11353_, _08450_);
  or _19749_ (\oc8051_symbolic_cxrom1.cxrom_data_out [4], _11354_, _11307_);
  and _19750_ (_11356_, _08451_, word_in[5]);
  nand _19751_ (_11358_, _08361_, _10425_);
  or _19752_ (_11359_, _08361_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  and _19753_ (_11360_, _11359_, _11358_);
  and _19754_ (_11361_, _11360_, _08416_);
  nand _19755_ (_11362_, _08361_, _10660_);
  or _19756_ (_11363_, _08361_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  and _19757_ (_11364_, _11363_, _11362_);
  and _19758_ (_11365_, _11364_, _08397_);
  nand _19759_ (_11366_, _08361_, _10871_);
  or _19760_ (_11367_, _08361_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  and _19761_ (_11368_, _11367_, _11366_);
  and _19762_ (_11369_, _11368_, _08393_);
  or _19763_ (_11371_, _11369_, _11365_);
  or _19764_ (_11372_, _11371_, _11361_);
  nand _19765_ (_11373_, _08361_, _11080_);
  or _19766_ (_11374_, _08361_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  and _19767_ (_11375_, _11374_, _11373_);
  and _19768_ (_11376_, _11375_, _08406_);
  or _19769_ (_11377_, _11376_, _08425_);
  or _19770_ (_11378_, _11377_, _11372_);
  nand _19771_ (_11379_, _08361_, _09527_);
  or _19772_ (_11380_, _08361_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  and _19773_ (_11381_, _11380_, _11379_);
  and _19774_ (_11382_, _11381_, _08416_);
  nand _19775_ (_11383_, _08361_, _09740_);
  or _19776_ (_11384_, _08361_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  and _19777_ (_11385_, _11384_, _11383_);
  and _19778_ (_11386_, _11385_, _08397_);
  nand _19779_ (_11387_, _08361_, _09971_);
  or _19780_ (_11388_, _08361_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  and _19781_ (_11389_, _11388_, _11387_);
  and _19782_ (_11390_, _11389_, _08393_);
  or _19783_ (_11391_, _11390_, _11386_);
  or _19784_ (_11392_, _11391_, _11382_);
  nand _19785_ (_11393_, _08361_, _10187_);
  or _19786_ (_11394_, _08361_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  and _19787_ (_11395_, _11394_, _11393_);
  and _19788_ (_11396_, _11395_, _08406_);
  or _19789_ (_11397_, _11396_, _08375_);
  or _19790_ (_11398_, _11397_, _11392_);
  and _19791_ (_11399_, _11398_, _11378_);
  and _19792_ (_11400_, _11399_, _08450_);
  or _19793_ (\oc8051_symbolic_cxrom1.cxrom_data_out [5], _11400_, _11356_);
  and _19794_ (_11401_, _08451_, word_in[6]);
  nand _19795_ (_11402_, _08361_, _10439_);
  or _19796_ (_11403_, _08361_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  and _19797_ (_11404_, _11403_, _11402_);
  and _19798_ (_11405_, _11404_, _08416_);
  nand _19799_ (_11407_, _08361_, _10671_);
  or _19800_ (_11408_, _08361_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  and _19801_ (_11409_, _11408_, _11407_);
  and _19802_ (_11410_, _11409_, _08397_);
  nand _19803_ (_11411_, _08361_, _10884_);
  or _19804_ (_11413_, _08361_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  and _19805_ (_11414_, _11413_, _11411_);
  and _19806_ (_11415_, _11414_, _08393_);
  or _19807_ (_11416_, _11415_, _11410_);
  or _19808_ (_11417_, _11416_, _11405_);
  nand _19809_ (_11418_, _08361_, _11093_);
  or _19810_ (_11419_, _08361_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  and _19811_ (_11420_, _11419_, _11418_);
  and _19812_ (_11421_, _11420_, _08406_);
  or _19813_ (_11422_, _11421_, _08425_);
  or _19814_ (_11423_, _11422_, _11417_);
  nand _19815_ (_11424_, _08361_, _09539_);
  or _19816_ (_11425_, _08361_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  and _19817_ (_11427_, _11425_, _11424_);
  and _19818_ (_11429_, _11427_, _08416_);
  nand _19819_ (_11430_, _08361_, _09752_);
  or _19820_ (_11431_, _08361_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  and _19821_ (_11432_, _11431_, _11430_);
  and _19822_ (_11433_, _11432_, _08397_);
  nand _19823_ (_11434_, _08361_, _09983_);
  or _19824_ (_11436_, _08361_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  and _19825_ (_11437_, _11436_, _11434_);
  and _19826_ (_11438_, _11437_, _08393_);
  or _19827_ (_11440_, _11438_, _11433_);
  or _19828_ (_11441_, _11440_, _11429_);
  nand _19829_ (_11442_, _08361_, _10203_);
  or _19830_ (_11444_, _08361_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  and _19831_ (_11445_, _11444_, _11442_);
  and _19832_ (_11446_, _11445_, _08406_);
  or _19833_ (_11447_, _11446_, _08375_);
  or _19834_ (_11448_, _11447_, _11441_);
  and _19835_ (_11449_, _11448_, _11423_);
  and _19836_ (_11450_, _11449_, _08450_);
  or _19837_ (\oc8051_symbolic_cxrom1.cxrom_data_out [6], _11450_, _11401_);
  and _19838_ (_11452_, _08557_, word_in[8]);
  nand _19839_ (_11453_, _08361_, _10481_);
  or _19840_ (_11454_, _08361_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and _19841_ (_11455_, _11454_, _11453_);
  and _19842_ (_11456_, _11455_, _08559_);
  nand _19843_ (_11457_, _08361_, _10246_);
  or _19844_ (_11458_, _08361_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  and _19845_ (_11459_, _11458_, _11457_);
  and _19846_ (_11460_, _11459_, _08558_);
  or _19847_ (_11461_, _11460_, _11456_);
  and _19848_ (_11462_, _11461_, _08523_);
  nand _19849_ (_11463_, _08361_, _09571_);
  or _19850_ (_11465_, _08361_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  and _19851_ (_11466_, _11465_, _11463_);
  and _19852_ (_11468_, _11466_, _08559_);
  nand _19853_ (_11469_, _08361_, _09332_);
  or _19854_ (_11470_, _08361_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  and _19855_ (_11471_, _11470_, _11469_);
  and _19856_ (_11472_, _11471_, _08558_);
  or _19857_ (_11473_, _11472_, _11468_);
  and _19858_ (_11474_, _11473_, _08525_);
  nand _19859_ (_11475_, _08361_, _10016_);
  or _19860_ (_11477_, _08361_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  and _19861_ (_11478_, _11477_, _11475_);
  and _19862_ (_11479_, _11478_, _08559_);
  nand _19863_ (_11480_, _08361_, _09790_);
  or _19864_ (_11481_, _08361_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  and _19865_ (_11482_, _11481_, _11480_);
  and _19866_ (_11483_, _11482_, _08558_);
  or _19867_ (_11484_, _11483_, _11479_);
  and _19868_ (_11485_, _11484_, _08600_);
  or _19869_ (_11486_, _11485_, _11474_);
  nand _19870_ (_11487_, _08361_, _10921_);
  or _19871_ (_11488_, _08361_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  and _19872_ (_11489_, _11488_, _11487_);
  and _19873_ (_11490_, _11489_, _08559_);
  nand _19874_ (_11491_, _08361_, _10703_);
  or _19875_ (_11492_, _08361_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  and _19876_ (_11493_, _11492_, _11491_);
  and _19877_ (_11494_, _11493_, _08558_);
  or _19878_ (_11495_, _11494_, _11490_);
  and _19879_ (_11496_, _11495_, _08573_);
  or _19880_ (_11497_, _11496_, _11486_);
  nor _19881_ (_11498_, _11497_, _11462_);
  nor _19882_ (_11499_, _11498_, _08557_);
  or _19883_ (\oc8051_symbolic_cxrom1.cxrom_data_out [8], _11499_, _11452_);
  and _19884_ (_11500_, _08557_, word_in[9]);
  nand _19885_ (_11501_, _08361_, _10495_);
  or _19886_ (_11502_, _08361_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  and _19887_ (_11503_, _11502_, _11501_);
  and _19888_ (_11504_, _11503_, _08559_);
  nand _19889_ (_11505_, _08361_, _10263_);
  or _19890_ (_11506_, _08361_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  and _19891_ (_11507_, _11506_, _11505_);
  and _19892_ (_11508_, _11507_, _08558_);
  or _19893_ (_11509_, _11508_, _11504_);
  and _19894_ (_11510_, _11509_, _08523_);
  nand _19895_ (_11511_, _08361_, _09586_);
  or _19896_ (_11512_, _08361_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  and _19897_ (_11513_, _11512_, _11511_);
  and _19898_ (_11514_, _11513_, _08559_);
  and _19899_ (_11515_, _08361_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  nor _19900_ (_11516_, _08361_, _09468_);
  or _19901_ (_11517_, _11516_, _11515_);
  and _19902_ (_11518_, _11517_, _08558_);
  or _19903_ (_11519_, _11518_, _11514_);
  and _19904_ (_11520_, _11519_, _08525_);
  nand _19905_ (_11521_, _08361_, _10026_);
  or _19906_ (_11523_, _08361_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  and _19907_ (_11524_, _11523_, _11521_);
  and _19908_ (_11525_, _11524_, _08559_);
  nand _19909_ (_11526_, _08361_, _09804_);
  or _19910_ (_11527_, _08361_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  and _19911_ (_11528_, _11527_, _11526_);
  and _19912_ (_11529_, _11528_, _08558_);
  or _19913_ (_11530_, _11529_, _11525_);
  and _19914_ (_11531_, _11530_, _08600_);
  or _19915_ (_11532_, _11531_, _11520_);
  nand _19916_ (_11533_, _08361_, _10931_);
  or _19917_ (_11534_, _08361_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  and _19918_ (_11535_, _11534_, _11533_);
  and _19919_ (_11536_, _11535_, _08559_);
  nand _19920_ (_11537_, _08361_, _10714_);
  or _19921_ (_11538_, _08361_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  and _19922_ (_11539_, _11538_, _11537_);
  and _19923_ (_11540_, _11539_, _08558_);
  or _19924_ (_11541_, _11540_, _11536_);
  and _19925_ (_11542_, _11541_, _08573_);
  or _19926_ (_11544_, _11542_, _11532_);
  nor _19927_ (_11545_, _11544_, _11510_);
  nor _19928_ (_11546_, _11545_, _08557_);
  or _19929_ (\oc8051_symbolic_cxrom1.cxrom_data_out [9], _11546_, _11500_);
  and _19930_ (_11547_, _08557_, word_in[10]);
  nand _19931_ (_11548_, _08361_, _10510_);
  or _19932_ (_11549_, _08361_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  and _19933_ (_11550_, _11549_, _11548_);
  and _19934_ (_11551_, _11550_, _08559_);
  nand _19935_ (_11552_, _08361_, _10276_);
  or _19936_ (_11553_, _08361_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  and _19937_ (_11554_, _11553_, _11552_);
  and _19938_ (_11555_, _11554_, _08558_);
  or _19939_ (_11556_, _11555_, _11551_);
  and _19940_ (_11557_, _11556_, _08523_);
  nand _19941_ (_11558_, _08361_, _09599_);
  or _19942_ (_11559_, _08361_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  and _19943_ (_11560_, _11559_, _11558_);
  and _19944_ (_11561_, _11560_, _08559_);
  and _19945_ (_11562_, _08361_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  nor _19946_ (_11563_, _08361_, _09482_);
  or _19947_ (_11564_, _11563_, _11562_);
  and _19948_ (_11566_, _11564_, _08558_);
  or _19949_ (_11567_, _11566_, _11561_);
  and _19950_ (_11568_, _11567_, _08525_);
  nand _19951_ (_11569_, _08361_, _10040_);
  or _19952_ (_11570_, _08361_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  and _19953_ (_11571_, _11570_, _11569_);
  and _19954_ (_11572_, _11571_, _08559_);
  nand _19955_ (_11573_, _08361_, _09818_);
  or _19956_ (_11574_, _08361_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  and _19957_ (_11575_, _11574_, _11573_);
  and _19958_ (_11576_, _11575_, _08558_);
  or _19959_ (_11577_, _11576_, _11572_);
  and _19960_ (_11578_, _11577_, _08600_);
  or _19961_ (_11580_, _11578_, _11568_);
  nand _19962_ (_11581_, _08361_, _10943_);
  or _19963_ (_11582_, _08361_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  and _19964_ (_11583_, _11582_, _11581_);
  and _19965_ (_11584_, _11583_, _08559_);
  nand _19966_ (_11585_, _08361_, _10726_);
  or _19967_ (_11586_, _08361_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  and _19968_ (_11587_, _11586_, _11585_);
  and _19969_ (_11588_, _11587_, _08558_);
  or _19970_ (_11589_, _11588_, _11584_);
  and _19971_ (_11590_, _11589_, _08573_);
  or _19972_ (_11591_, _11590_, _11580_);
  nor _19973_ (_11592_, _11591_, _11557_);
  nor _19974_ (_11593_, _11592_, _08557_);
  or _19975_ (\oc8051_symbolic_cxrom1.cxrom_data_out [10], _11593_, _11547_);
  and _19976_ (_11594_, _08557_, word_in[11]);
  nand _19977_ (_11596_, _08361_, _10522_);
  or _19978_ (_11597_, _08361_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  and _19979_ (_11599_, _11597_, _11596_);
  and _19980_ (_11600_, _11599_, _08559_);
  nand _19981_ (_11601_, _08361_, _10288_);
  or _19982_ (_11603_, _08361_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  and _19983_ (_11604_, _11603_, _11601_);
  and _19984_ (_11606_, _11604_, _08558_);
  or _19985_ (_11607_, _11606_, _11600_);
  and _19986_ (_11608_, _11607_, _08523_);
  nand _19987_ (_11609_, _08361_, _10957_);
  or _19988_ (_11611_, _08361_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  and _19989_ (_11612_, _11611_, _11609_);
  and _19990_ (_11613_, _11612_, _08559_);
  nand _19991_ (_11614_, _08361_, _10737_);
  or _19992_ (_11615_, _08361_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  and _19993_ (_11617_, _11615_, _11614_);
  and _19994_ (_11619_, _11617_, _08558_);
  or _19995_ (_11621_, _11619_, _11613_);
  and _19996_ (_11622_, _11621_, _08573_);
  nand _19997_ (_11623_, _08361_, _10053_);
  or _19998_ (_11625_, _08361_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  and _19999_ (_11626_, _11625_, _11623_);
  and _20000_ (_11627_, _11626_, _08559_);
  nand _20001_ (_11628_, _08361_, _09834_);
  or _20002_ (_11629_, _08361_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  and _20003_ (_11631_, _11629_, _11628_);
  and _20004_ (_11632_, _11631_, _08558_);
  or _20005_ (_11633_, _11632_, _11627_);
  and _20006_ (_11634_, _11633_, _08600_);
  nand _20007_ (_11635_, _08361_, _09610_);
  or _20008_ (_11636_, _08361_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  and _20009_ (_11637_, _11636_, _11635_);
  and _20010_ (_11639_, _11637_, _08559_);
  and _20011_ (_11640_, _08361_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  nor _20012_ (_11642_, _08361_, _09497_);
  or _20013_ (_11643_, _11642_, _11640_);
  and _20014_ (_11644_, _11643_, _08558_);
  or _20015_ (_11645_, _11644_, _11639_);
  and _20016_ (_11647_, _11645_, _08525_);
  or _20017_ (_11648_, _11647_, _11634_);
  or _20018_ (_11649_, _11648_, _11622_);
  nor _20019_ (_11650_, _11649_, _11608_);
  nor _20020_ (_11651_, _11650_, _08557_);
  or _20021_ (\oc8051_symbolic_cxrom1.cxrom_data_out [11], _11651_, _11594_);
  and _20022_ (_11652_, _08557_, word_in[12]);
  nand _20023_ (_11653_, _08361_, _10535_);
  or _20024_ (_11654_, _08361_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  and _20025_ (_11655_, _11654_, _11653_);
  and _20026_ (_11656_, _11655_, _08559_);
  nand _20027_ (_11657_, _08361_, _10302_);
  or _20028_ (_11659_, _08361_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  and _20029_ (_11660_, _11659_, _11657_);
  and _20030_ (_11661_, _11660_, _08558_);
  or _20031_ (_11662_, _11661_, _11656_);
  and _20032_ (_11663_, _11662_, _08523_);
  nand _20033_ (_11664_, _08361_, _09622_);
  or _20034_ (_11665_, _08361_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  and _20035_ (_11666_, _11665_, _11664_);
  and _20036_ (_11667_, _11666_, _08559_);
  and _20037_ (_11668_, _08361_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  nor _20038_ (_11669_, _08361_, _09508_);
  or _20039_ (_11670_, _11669_, _11668_);
  and _20040_ (_11671_, _11670_, _08558_);
  or _20041_ (_11672_, _11671_, _11667_);
  and _20042_ (_11673_, _11672_, _08525_);
  nand _20043_ (_11674_, _08361_, _10066_);
  or _20044_ (_11675_, _08361_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  and _20045_ (_11676_, _11675_, _11674_);
  and _20046_ (_11677_, _11676_, _08559_);
  nand _20047_ (_11678_, _08361_, _09846_);
  or _20048_ (_11679_, _08361_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  and _20049_ (_11680_, _11679_, _11678_);
  and _20050_ (_11681_, _11680_, _08558_);
  or _20051_ (_11682_, _11681_, _11677_);
  and _20052_ (_11683_, _11682_, _08600_);
  or _20053_ (_11684_, _11683_, _11673_);
  nand _20054_ (_11685_, _08361_, _10968_);
  or _20055_ (_11686_, _08361_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  and _20056_ (_11687_, _11686_, _11685_);
  and _20057_ (_11688_, _11687_, _08559_);
  nand _20058_ (_11689_, _08361_, _10749_);
  or _20059_ (_11690_, _08361_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  and _20060_ (_11691_, _11690_, _11689_);
  and _20061_ (_11692_, _11691_, _08558_);
  or _20062_ (_11693_, _11692_, _11688_);
  and _20063_ (_11694_, _11693_, _08573_);
  or _20064_ (_11695_, _11694_, _11684_);
  nor _20065_ (_11696_, _11695_, _11663_);
  nor _20066_ (_11697_, _11696_, _08557_);
  or _20067_ (\oc8051_symbolic_cxrom1.cxrom_data_out [12], _11697_, _11652_);
  and _20068_ (_11699_, _08557_, word_in[13]);
  nand _20069_ (_11700_, _08361_, _10548_);
  or _20070_ (_11701_, _08361_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  and _20071_ (_11702_, _11701_, _11700_);
  and _20072_ (_11703_, _11702_, _08559_);
  nand _20073_ (_11705_, _08361_, _10315_);
  or _20074_ (_11706_, _08361_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  and _20075_ (_11707_, _11706_, _11705_);
  and _20076_ (_11708_, _11707_, _08558_);
  or _20077_ (_11709_, _11708_, _11703_);
  and _20078_ (_11711_, _11709_, _08523_);
  nand _20079_ (_11712_, _08361_, _09635_);
  or _20080_ (_11713_, _08361_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  and _20081_ (_11714_, _11713_, _11712_);
  and _20082_ (_11716_, _11714_, _08559_);
  and _20083_ (_11717_, _08361_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  nor _20084_ (_11719_, _08361_, _09527_);
  or _20085_ (_11721_, _11719_, _11717_);
  and _20086_ (_11722_, _11721_, _08558_);
  or _20087_ (_11724_, _11722_, _11716_);
  and _20088_ (_11725_, _11724_, _08525_);
  nand _20089_ (_11727_, _08361_, _10080_);
  or _20090_ (_11728_, _08361_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  and _20091_ (_11730_, _11728_, _11727_);
  and _20092_ (_11731_, _11730_, _08559_);
  nand _20093_ (_11732_, _08361_, _09858_);
  or _20094_ (_11733_, _08361_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  and _20095_ (_11734_, _11733_, _11732_);
  and _20096_ (_11735_, _11734_, _08558_);
  or _20097_ (_11737_, _11735_, _11731_);
  and _20098_ (_11738_, _11737_, _08600_);
  or _20099_ (_11739_, _11738_, _11725_);
  nand _20100_ (_11740_, _08361_, _10981_);
  or _20101_ (_11741_, _08361_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  and _20102_ (_11742_, _11741_, _11740_);
  and _20103_ (_11743_, _11742_, _08559_);
  nand _20104_ (_11744_, _08361_, _10763_);
  or _20105_ (_11745_, _08361_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  and _20106_ (_11746_, _11745_, _11744_);
  and _20107_ (_11747_, _11746_, _08558_);
  or _20108_ (_11748_, _11747_, _11743_);
  and _20109_ (_11749_, _11748_, _08573_);
  or _20110_ (_11750_, _11749_, _11739_);
  nor _20111_ (_11752_, _11750_, _11711_);
  nor _20112_ (_11753_, _11752_, _08557_);
  or _20113_ (\oc8051_symbolic_cxrom1.cxrom_data_out [13], _11753_, _11699_);
  and _20114_ (_11755_, _08557_, word_in[14]);
  nand _20115_ (_11756_, _08361_, _10564_);
  or _20116_ (_11757_, _08361_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  and _20117_ (_11758_, _11757_, _11756_);
  and _20118_ (_11759_, _11758_, _08559_);
  nand _20119_ (_11760_, _08361_, _10328_);
  or _20120_ (_11761_, _08361_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  and _20121_ (_11762_, _11761_, _11760_);
  and _20122_ (_11763_, _11762_, _08558_);
  or _20123_ (_11764_, _11763_, _11759_);
  and _20124_ (_11765_, _11764_, _08523_);
  nand _20125_ (_11766_, _08361_, _10994_);
  or _20126_ (_11767_, _08361_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  and _20127_ (_11768_, _11767_, _11766_);
  and _20128_ (_11769_, _11768_, _08559_);
  nand _20129_ (_11770_, _08361_, _10775_);
  or _20130_ (_11771_, _08361_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  and _20131_ (_11772_, _11771_, _11770_);
  and _20132_ (_11773_, _11772_, _08558_);
  or _20133_ (_11774_, _11773_, _11769_);
  and _20134_ (_11775_, _11774_, _08573_);
  nand _20135_ (_11776_, _08361_, _10092_);
  or _20136_ (_11777_, _08361_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  and _20137_ (_11778_, _11777_, _11776_);
  and _20138_ (_11779_, _11778_, _08559_);
  nand _20139_ (_11780_, _08361_, _09870_);
  or _20140_ (_11781_, _08361_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  and _20141_ (_11782_, _11781_, _11780_);
  and _20142_ (_11783_, _11782_, _08558_);
  or _20143_ (_11784_, _11783_, _11779_);
  and _20144_ (_11785_, _11784_, _08600_);
  nand _20145_ (_11786_, _08361_, _09647_);
  or _20146_ (_11787_, _08361_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  and _20147_ (_11788_, _11787_, _11786_);
  and _20148_ (_11789_, _11788_, _08559_);
  and _20149_ (_11790_, _08361_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  nor _20150_ (_11791_, _08361_, _09539_);
  or _20151_ (_11793_, _11791_, _11790_);
  and _20152_ (_11794_, _11793_, _08558_);
  or _20153_ (_11795_, _11794_, _11789_);
  and _20154_ (_11796_, _11795_, _08525_);
  or _20155_ (_11797_, _11796_, _11785_);
  or _20156_ (_11798_, _11797_, _11775_);
  nor _20157_ (_11799_, _11798_, _11765_);
  nor _20158_ (_11800_, _11799_, _08557_);
  or _20159_ (\oc8051_symbolic_cxrom1.cxrom_data_out [14], _11800_, _11755_);
  and _20160_ (_11802_, _08654_, word_in[16]);
  and _20161_ (_11803_, _11154_, _08406_);
  and _20162_ (_11804_, _11163_, _08393_);
  or _20163_ (_11806_, _11804_, _11803_);
  and _20164_ (_11807_, _11159_, _08397_);
  and _20165_ (_11808_, _11167_, _08416_);
  or _20166_ (_11809_, _11808_, _11807_);
  or _20167_ (_11810_, _11809_, _11806_);
  or _20168_ (_11811_, _11810_, _08619_);
  and _20169_ (_11812_, _11138_, _08397_);
  and _20170_ (_11813_, _11133_, _08406_);
  or _20171_ (_11814_, _11813_, _11812_);
  and _20172_ (_11815_, _11142_, _08393_);
  and _20173_ (_11816_, _11146_, _08416_);
  or _20174_ (_11817_, _11816_, _11815_);
  nor _20175_ (_11818_, _11817_, _11814_);
  nand _20176_ (_11819_, _11818_, _08619_);
  nand _20177_ (_11820_, _11819_, _11811_);
  nor _20178_ (_11821_, _11820_, _08654_);
  or _20179_ (\oc8051_symbolic_cxrom1.cxrom_data_out [16], _11821_, _11802_);
  and _20180_ (_11822_, _08654_, word_in[17]);
  and _20181_ (_11823_, _11206_, _08397_);
  and _20182_ (_11824_, _11198_, _08406_);
  or _20183_ (_11826_, _11824_, _11823_);
  and _20184_ (_11827_, _11212_, _08393_);
  and _20185_ (_11828_, _11202_, _08416_);
  or _20186_ (_11829_, _11828_, _11827_);
  or _20187_ (_11831_, _11829_, _11826_);
  or _20188_ (_11832_, _11831_, _08619_);
  and _20189_ (_11833_, _11186_, _08397_);
  and _20190_ (_11834_, _11178_, _08406_);
  or _20191_ (_11835_, _11834_, _11833_);
  and _20192_ (_11836_, _11192_, _08393_);
  and _20193_ (_11837_, _11182_, _08416_);
  or _20194_ (_11838_, _11837_, _11836_);
  nor _20195_ (_11839_, _11838_, _11835_);
  nand _20196_ (_11840_, _11839_, _08619_);
  nand _20197_ (_11841_, _11840_, _11832_);
  nor _20198_ (_11842_, _11841_, _08654_);
  or _20199_ (\oc8051_symbolic_cxrom1.cxrom_data_out [17], _11842_, _11822_);
  and _20200_ (_11843_, _08654_, word_in[18]);
  and _20201_ (_11845_, _11248_, _08397_);
  and _20202_ (_11846_, _11242_, _08406_);
  or _20203_ (_11847_, _11846_, _11845_);
  and _20204_ (_11849_, _11252_, _08393_);
  and _20205_ (_11850_, _11256_, _08416_);
  or _20206_ (_11851_, _11850_, _11849_);
  or _20207_ (_11852_, _11851_, _11847_);
  or _20208_ (_11853_, _11852_, _08619_);
  and _20209_ (_11854_, _11226_, _08397_);
  and _20210_ (_11855_, _11221_, _08406_);
  or _20211_ (_11857_, _11855_, _11854_);
  and _20212_ (_11858_, _11230_, _08393_);
  and _20213_ (_11859_, _11234_, _08416_);
  or _20214_ (_11860_, _11859_, _11858_);
  nor _20215_ (_11861_, _11860_, _11857_);
  nand _20216_ (_11862_, _11861_, _08619_);
  nand _20217_ (_11863_, _11862_, _11853_);
  nor _20218_ (_11864_, _11863_, _08654_);
  or _20219_ (\oc8051_symbolic_cxrom1.cxrom_data_out [18], _11864_, _11843_);
  and _20220_ (_11865_, _08654_, word_in[19]);
  and _20221_ (_11866_, _11295_, _08397_);
  and _20222_ (_11867_, _11286_, _08406_);
  or _20223_ (_11868_, _11867_, _11866_);
  and _20224_ (_11869_, _11301_, _08393_);
  and _20225_ (_11870_, _11290_, _08416_);
  or _20226_ (_11871_, _11870_, _11869_);
  or _20227_ (_11872_, _11871_, _11868_);
  or _20228_ (_11873_, _11872_, _08619_);
  and _20229_ (_11874_, _11266_, _08406_);
  and _20230_ (_11875_, _11280_, _08393_);
  or _20231_ (_11876_, _11875_, _11874_);
  and _20232_ (_11878_, _11274_, _08397_);
  and _20233_ (_11879_, _11270_, _08416_);
  or _20234_ (_11880_, _11879_, _11878_);
  nor _20235_ (_11881_, _11880_, _11876_);
  nand _20236_ (_11882_, _11881_, _08619_);
  nand _20237_ (_11884_, _11882_, _11873_);
  nor _20238_ (_11885_, _11884_, _08654_);
  or _20239_ (\oc8051_symbolic_cxrom1.cxrom_data_out [19], _11885_, _11865_);
  and _20240_ (_11886_, _08654_, word_in[20]);
  and _20241_ (_11887_, _11332_, _08406_);
  and _20242_ (_11889_, _11348_, _08393_);
  or _20243_ (_11890_, _11889_, _11887_);
  and _20244_ (_11892_, _11340_, _08397_);
  and _20245_ (_11893_, _11336_, _08416_);
  or _20246_ (_11894_, _11893_, _11892_);
  or _20247_ (_11895_, _11894_, _11890_);
  or _20248_ (_11896_, _11895_, _08619_);
  and _20249_ (_11898_, _11319_, _08397_);
  and _20250_ (_11899_, _11310_, _08406_);
  or _20251_ (_11901_, _11899_, _11898_);
  and _20252_ (_11902_, _11325_, _08393_);
  and _20253_ (_11903_, _11315_, _08416_);
  or _20254_ (_11905_, _11903_, _11902_);
  nor _20255_ (_11906_, _11905_, _11901_);
  nand _20256_ (_11908_, _11906_, _08619_);
  nand _20257_ (_11909_, _11908_, _11896_);
  nor _20258_ (_11911_, _11909_, _08654_);
  or _20259_ (\oc8051_symbolic_cxrom1.cxrom_data_out [20], _11911_, _11886_);
  and _20260_ (_11912_, _08654_, word_in[21]);
  and _20261_ (_11913_, _11389_, _08397_);
  and _20262_ (_11915_, _11381_, _08406_);
  or _20263_ (_11916_, _11915_, _11913_);
  and _20264_ (_11917_, _11395_, _08393_);
  and _20265_ (_11918_, _11385_, _08416_);
  or _20266_ (_11919_, _11918_, _11917_);
  or _20267_ (_11920_, _11919_, _11916_);
  or _20268_ (_11921_, _11920_, _08619_);
  and _20269_ (_11922_, _11360_, _08406_);
  and _20270_ (_11923_, _11375_, _08393_);
  or _20271_ (_11925_, _11923_, _11922_);
  and _20272_ (_11926_, _11368_, _08397_);
  and _20273_ (_11928_, _11364_, _08416_);
  or _20274_ (_11929_, _11928_, _11926_);
  nor _20275_ (_11931_, _11929_, _11925_);
  nand _20276_ (_11932_, _11931_, _08619_);
  nand _20277_ (_11933_, _11932_, _11921_);
  nor _20278_ (_11934_, _11933_, _08654_);
  or _20279_ (\oc8051_symbolic_cxrom1.cxrom_data_out [21], _11934_, _11912_);
  and _20280_ (_11935_, _08654_, word_in[22]);
  and _20281_ (_11936_, _11427_, _08406_);
  and _20282_ (_11937_, _11445_, _08393_);
  or _20283_ (_11938_, _11937_, _11936_);
  and _20284_ (_11939_, _11437_, _08397_);
  and _20285_ (_11940_, _11432_, _08416_);
  or _20286_ (_11941_, _11940_, _11939_);
  or _20287_ (_11942_, _11941_, _11938_);
  or _20288_ (_11943_, _11942_, _08619_);
  and _20289_ (_11944_, _11404_, _08406_);
  and _20290_ (_11946_, _11420_, _08393_);
  or _20291_ (_11947_, _11946_, _11944_);
  and _20292_ (_11948_, _11414_, _08397_);
  and _20293_ (_11949_, _11409_, _08416_);
  or _20294_ (_11950_, _11949_, _11948_);
  nor _20295_ (_11951_, _11950_, _11947_);
  nand _20296_ (_11952_, _11951_, _08619_);
  nand _20297_ (_11953_, _11952_, _11943_);
  nor _20298_ (_11954_, _11953_, _08654_);
  or _20299_ (\oc8051_symbolic_cxrom1.cxrom_data_out [22], _11954_, _11935_);
  and _20300_ (_11955_, _08717_, word_in[24]);
  and _20301_ (_11956_, _11459_, _08559_);
  and _20302_ (_11957_, _11455_, _08558_);
  or _20303_ (_11958_, _11957_, _11956_);
  and _20304_ (_11959_, _11958_, _08685_);
  and _20305_ (_11960_, _11471_, _08559_);
  and _20306_ (_11961_, _11466_, _08558_);
  or _20307_ (_11962_, _11961_, _11960_);
  and _20308_ (_11963_, _11962_, _08690_);
  and _20309_ (_11964_, _11482_, _08559_);
  and _20310_ (_11965_, _11478_, _08558_);
  or _20311_ (_11966_, _11965_, _11964_);
  and _20312_ (_11967_, _11966_, _08726_);
  and _20313_ (_11968_, _11493_, _08559_);
  and _20314_ (_11969_, _11489_, _08558_);
  or _20315_ (_11970_, _11969_, _11968_);
  and _20316_ (_11971_, _11970_, _08731_);
  or _20317_ (_11972_, _11971_, _11967_);
  or _20318_ (_11973_, _11972_, _11963_);
  nor _20319_ (_11974_, _11973_, _11959_);
  nor _20320_ (_11975_, _11974_, _08717_);
  or _20321_ (\oc8051_symbolic_cxrom1.cxrom_data_out [24], _11975_, _11955_);
  and _20322_ (_11976_, _08717_, word_in[25]);
  and _20323_ (_11977_, _11507_, _08559_);
  and _20324_ (_11978_, _11503_, _08558_);
  or _20325_ (_11980_, _11978_, _11977_);
  and _20326_ (_11981_, _11980_, _08685_);
  and _20327_ (_11982_, _11517_, _08559_);
  and _20328_ (_11983_, _11513_, _08558_);
  or _20329_ (_11985_, _11983_, _11982_);
  and _20330_ (_11986_, _11985_, _08690_);
  and _20331_ (_11987_, _11528_, _08559_);
  and _20332_ (_11988_, _11524_, _08558_);
  or _20333_ (_11989_, _11988_, _11987_);
  and _20334_ (_11990_, _11989_, _08726_);
  and _20335_ (_11991_, _11539_, _08559_);
  and _20336_ (_11992_, _11535_, _08558_);
  or _20337_ (_11994_, _11992_, _11991_);
  and _20338_ (_11996_, _11994_, _08731_);
  or _20339_ (_11997_, _11996_, _11990_);
  or _20340_ (_11998_, _11997_, _11986_);
  nor _20341_ (_11999_, _11998_, _11981_);
  nor _20342_ (_12000_, _11999_, _08717_);
  or _20343_ (\oc8051_symbolic_cxrom1.cxrom_data_out [25], _12000_, _11976_);
  and _20344_ (_12002_, _08717_, word_in[26]);
  and _20345_ (_12003_, _11564_, _08559_);
  and _20346_ (_12004_, _11560_, _08558_);
  or _20347_ (_12005_, _12004_, _12003_);
  and _20348_ (_12007_, _12005_, _08690_);
  and _20349_ (_12008_, _11554_, _08559_);
  and _20350_ (_12009_, _11550_, _08558_);
  or _20351_ (_12010_, _12009_, _12008_);
  and _20352_ (_12012_, _12010_, _08685_);
  and _20353_ (_12013_, _11575_, _08559_);
  and _20354_ (_12015_, _11571_, _08558_);
  or _20355_ (_12016_, _12015_, _12013_);
  and _20356_ (_12018_, _12016_, _08726_);
  and _20357_ (_12019_, _11587_, _08559_);
  and _20358_ (_12020_, _11583_, _08558_);
  or _20359_ (_12021_, _12020_, _12019_);
  and _20360_ (_12022_, _12021_, _08731_);
  or _20361_ (_12023_, _12022_, _12018_);
  or _20362_ (_12024_, _12023_, _12012_);
  nor _20363_ (_12025_, _12024_, _12007_);
  nor _20364_ (_12026_, _12025_, _08717_);
  or _20365_ (\oc8051_symbolic_cxrom1.cxrom_data_out [26], _12026_, _12002_);
  and _20366_ (_12027_, _08717_, word_in[27]);
  and _20367_ (_12028_, _11643_, _08559_);
  and _20368_ (_12029_, _11637_, _08558_);
  or _20369_ (_12030_, _12029_, _12028_);
  and _20370_ (_12031_, _12030_, _08690_);
  and _20371_ (_12033_, _11604_, _08559_);
  and _20372_ (_12034_, _11599_, _08558_);
  or _20373_ (_12036_, _12034_, _12033_);
  and _20374_ (_12037_, _12036_, _08685_);
  and _20375_ (_12039_, _11631_, _08559_);
  and _20376_ (_12041_, _11626_, _08558_);
  or _20377_ (_12043_, _12041_, _12039_);
  and _20378_ (_12044_, _12043_, _08726_);
  and _20379_ (_12045_, _11617_, _08559_);
  and _20380_ (_12046_, _11612_, _08558_);
  or _20381_ (_12047_, _12046_, _12045_);
  and _20382_ (_12048_, _12047_, _08731_);
  or _20383_ (_12050_, _12048_, _12044_);
  or _20384_ (_12051_, _12050_, _12037_);
  nor _20385_ (_12052_, _12051_, _12031_);
  nor _20386_ (_12053_, _12052_, _08717_);
  or _20387_ (\oc8051_symbolic_cxrom1.cxrom_data_out [27], _12053_, _12027_);
  and _20388_ (_12054_, _08717_, word_in[28]);
  and _20389_ (_12055_, _11660_, _08559_);
  and _20390_ (_12056_, _11655_, _08558_);
  or _20391_ (_12057_, _12056_, _12055_);
  and _20392_ (_12058_, _12057_, _08685_);
  and _20393_ (_12059_, _11670_, _08559_);
  and _20394_ (_12060_, _11666_, _08558_);
  or _20395_ (_12061_, _12060_, _12059_);
  and _20396_ (_12062_, _12061_, _08690_);
  and _20397_ (_12063_, _11680_, _08559_);
  and _20398_ (_12064_, _11676_, _08558_);
  or _20399_ (_12065_, _12064_, _12063_);
  and _20400_ (_12066_, _12065_, _08726_);
  and _20401_ (_12067_, _11691_, _08559_);
  and _20402_ (_12068_, _11687_, _08558_);
  or _20403_ (_12069_, _12068_, _12067_);
  and _20404_ (_12070_, _12069_, _08731_);
  or _20405_ (_12071_, _12070_, _12066_);
  or _20406_ (_12072_, _12071_, _12062_);
  nor _20407_ (_12073_, _12072_, _12058_);
  nor _20408_ (_12074_, _12073_, _08717_);
  or _20409_ (\oc8051_symbolic_cxrom1.cxrom_data_out [28], _12074_, _12054_);
  and _20410_ (_12075_, _08717_, word_in[29]);
  and _20411_ (_12076_, _11707_, _08559_);
  and _20412_ (_12078_, _11702_, _08558_);
  or _20413_ (_12079_, _12078_, _12076_);
  and _20414_ (_12080_, _12079_, _08685_);
  and _20415_ (_12081_, _11721_, _08559_);
  and _20416_ (_12083_, _11714_, _08558_);
  or _20417_ (_12084_, _12083_, _12081_);
  and _20418_ (_12085_, _12084_, _08690_);
  and _20419_ (_12086_, _11734_, _08559_);
  and _20420_ (_12087_, _11730_, _08558_);
  or _20421_ (_12088_, _12087_, _12086_);
  and _20422_ (_12089_, _12088_, _08726_);
  and _20423_ (_12090_, _11746_, _08559_);
  and _20424_ (_12091_, _11742_, _08558_);
  or _20425_ (_12092_, _12091_, _12090_);
  and _20426_ (_12094_, _12092_, _08731_);
  or _20427_ (_12095_, _12094_, _12089_);
  or _20428_ (_12096_, _12095_, _12085_);
  nor _20429_ (_12097_, _12096_, _12080_);
  nor _20430_ (_12098_, _12097_, _08717_);
  or _20431_ (\oc8051_symbolic_cxrom1.cxrom_data_out [29], _12098_, _12075_);
  and _20432_ (_12099_, _08717_, word_in[30]);
  and _20433_ (_12100_, _11793_, _08559_);
  and _20434_ (_12101_, _11788_, _08558_);
  or _20435_ (_12102_, _12101_, _12100_);
  and _20436_ (_12103_, _12102_, _08690_);
  and _20437_ (_12104_, _11762_, _08559_);
  and _20438_ (_12105_, _11758_, _08558_);
  or _20439_ (_12106_, _12105_, _12104_);
  and _20440_ (_12107_, _12106_, _08685_);
  and _20441_ (_12108_, _11782_, _08559_);
  and _20442_ (_12109_, _11778_, _08558_);
  or _20443_ (_12110_, _12109_, _12108_);
  and _20444_ (_12111_, _12110_, _08726_);
  and _20445_ (_12112_, _11772_, _08559_);
  and _20446_ (_12113_, _11768_, _08558_);
  or _20447_ (_12114_, _12113_, _12112_);
  and _20448_ (_12115_, _12114_, _08731_);
  or _20449_ (_12116_, _12115_, _12111_);
  or _20450_ (_12117_, _12116_, _12107_);
  nor _20451_ (_12118_, _12117_, _12103_);
  nor _20452_ (_12120_, _12118_, _08717_);
  or _20453_ (\oc8051_symbolic_cxrom1.cxrom_data_out [30], _12120_, _12099_);
  or _20454_ (_12121_, _05843_, _06812_);
  or _20455_ (_12122_, _05729_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and _20456_ (_12123_, _12122_, _04856_);
  and _20457_ (_09782_, _12123_, _12121_);
  and _20458_ (_09788_, _06849_, _04856_);
  or _20459_ (_12124_, _05943_, _06812_);
  or _20460_ (_12125_, _05729_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and _20461_ (_12126_, _12125_, _04856_);
  and _20462_ (_09791_, _12126_, _12124_);
  or _20463_ (_12127_, _05983_, _05848_);
  and _20464_ (_12129_, _12127_, _06777_);
  nor _20465_ (_12131_, _06783_, _12129_);
  or _20466_ (_09794_, _12131_, _06782_);
  or _20467_ (_12132_, _05895_, _06812_);
  or _20468_ (_12133_, _05729_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and _20469_ (_12134_, _12133_, _04856_);
  and _20470_ (_09806_, _12134_, _12132_);
  or _20471_ (_12136_, _08164_, \oc8051_top_1.oc8051_decoder1.state [1]);
  or _20472_ (_12138_, _08168_, _08166_);
  or _20473_ (_12139_, _12138_, _08159_);
  or _20474_ (_12140_, _12139_, _12136_);
  and _20475_ (_12142_, _12140_, _08181_);
  nor _20476_ (_12143_, _08180_, _05957_);
  or _20477_ (_12144_, _12143_, rst);
  or _20478_ (_09810_, _12144_, _12142_);
  or _20479_ (_12145_, _05767_, _06812_);
  or _20480_ (_12146_, _05729_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and _20481_ (_12148_, _12146_, _04856_);
  and _20482_ (_09813_, _12148_, _12145_);
  and _20483_ (_12149_, _05983_, _06772_);
  nor _20484_ (_12150_, _06783_, _12149_);
  or _20485_ (_09820_, _12150_, _06782_);
  and _20486_ (_09822_, _06903_, _04856_);
  and _20487_ (_12152_, _09950_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  and _20488_ (_12153_, _04861_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  and _20489_ (_12155_, _12153_, _09954_);
  and _20490_ (_12157_, _05718_, _05671_);
  or _20491_ (_12158_, _12157_, _12155_);
  or _20492_ (_12159_, _12158_, _12152_);
  and _20493_ (_09831_, _12159_, _04856_);
  or _20494_ (_12160_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  nand _20495_ (_12161_, _08367_, _05906_);
  and _20496_ (_12162_, _12161_, _04856_);
  and _20497_ (_09984_, _12162_, _12160_);
  and _20498_ (_12164_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  not _20499_ (_12165_, _08367_);
  and _20500_ (_12166_, _12165_, \oc8051_top_1.oc8051_rom1.data_o [31]);
  or _20501_ (_12167_, _12166_, _12164_);
  and _20502_ (_09996_, _12167_, _04856_);
  and _20503_ (_12168_, _06818_, _04856_);
  and _20504_ (_10047_, _12168_, _06851_);
  nor _20505_ (_12170_, \oc8051_top_1.oc8051_decoder1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  and _20506_ (_12171_, _12170_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _20507_ (_10060_, _12171_, _04856_);
  and _20508_ (_02999_, \oc8051_top_1.oc8051_memory_interface1.istb_t , _04856_);
  and _20509_ (_12174_, _02999_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or _20510_ (_10067_, _12174_, _10060_);
  nand _20511_ (_12175_, _05726_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _20512_ (_10072_, _12175_, _04856_);
  and _20513_ (_10114_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , _04856_);
  nor _20514_ (_12176_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , rst);
  and _20515_ (_10135_, _12176_, \oc8051_top_1.oc8051_memory_interface1.int_ack_buff );
  and _20516_ (_12177_, _08275_, _06142_);
  and _20517_ (_12179_, _12177_, _04986_);
  or _20518_ (_12180_, _12179_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  and _20519_ (_12182_, _06662_, _04993_);
  and _20520_ (_12183_, _12182_, _06126_);
  not _20521_ (_12185_, _12183_);
  and _20522_ (_12186_, _12185_, _12180_);
  nand _20523_ (_12187_, _12179_, _06088_);
  and _20524_ (_12188_, _12187_, _12186_);
  nor _20525_ (_12189_, _12185_, _06032_);
  or _20526_ (_12190_, _12189_, _12188_);
  and _20527_ (_10143_, _12190_, _04856_);
  and _20528_ (_12191_, _12177_, _04990_);
  or _20529_ (_12192_, _12191_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and _20530_ (_12193_, _12192_, _12185_);
  nand _20531_ (_12194_, _12191_, _06088_);
  and _20532_ (_12195_, _12194_, _12193_);
  and _20533_ (_12196_, _12183_, _06997_);
  or _20534_ (_12197_, _12196_, _12195_);
  and _20535_ (_10146_, _12197_, _04856_);
  not _20536_ (_12198_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  not _20537_ (_12199_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nor _20538_ (_12200_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and _20539_ (_12201_, _12200_, _12199_);
  nor _20540_ (_12202_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  nor _20541_ (_12203_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and _20542_ (_12204_, _12203_, _12202_);
  and _20543_ (_12205_, _12204_, _12201_);
  and _20544_ (_12206_, _12205_, _12198_);
  and _20545_ (_12207_, _12206_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  or _20546_ (_12208_, _12207_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  and _20547_ (_10174_, _12208_, _04856_);
  and _20548_ (_12209_, _05940_, _05839_);
  and _20549_ (_12210_, _05815_, _05866_);
  and _20550_ (_12212_, _12210_, _12209_);
  and _20551_ (_12213_, _05731_, _04856_);
  and _20552_ (_12214_, _12213_, _05915_);
  and _20553_ (_12215_, _12214_, _05891_);
  and _20554_ (_12216_, _05763_, _05789_);
  and _20555_ (_12217_, _12216_, _12215_);
  and _20556_ (_10190_, _12217_, _12212_);
  and _20557_ (_12218_, _06134_, _04932_);
  and _20558_ (_12219_, _12218_, _06662_);
  not _20559_ (_12220_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and _20560_ (_12221_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and _20561_ (_12222_, _12221_, _12220_);
  or _20562_ (_12223_, _12222_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or _20563_ (_12224_, _12223_, _12219_);
  not _20564_ (_12225_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or _20565_ (_12226_, _06146_, _12225_);
  nand _20566_ (_12227_, _12226_, _12177_);
  or _20567_ (_12228_, _12227_, _06147_);
  and _20568_ (_12230_, _12228_, _12224_);
  or _20569_ (_12231_, _12230_, _12183_);
  nand _20570_ (_12232_, _12183_, _05287_);
  and _20571_ (_12233_, _12232_, _04856_);
  and _20572_ (_10193_, _12233_, _12231_);
  and _20573_ (_12235_, _12177_, _06091_);
  or _20574_ (_12236_, _12235_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and _20575_ (_12237_, _12236_, _12185_);
  nand _20576_ (_12238_, _12235_, _06088_);
  and _20577_ (_12240_, _12238_, _12237_);
  and _20578_ (_12241_, _12183_, _05718_);
  or _20579_ (_12242_, _12241_, _12240_);
  and _20580_ (_10199_, _12242_, _04856_);
  and _20581_ (_12243_, _12219_, _07857_);
  and _20582_ (_12244_, _12219_, _04984_);
  not _20583_ (_12245_, _12219_);
  nor _20584_ (_12246_, _04989_, _04984_);
  or _20585_ (_12247_, _12246_, _12245_);
  or _20586_ (_12248_, _12247_, _12244_);
  and _20587_ (_12249_, _12248_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  or _20588_ (_12250_, _12249_, _12183_);
  or _20589_ (_12252_, _12250_, _12243_);
  or _20590_ (_12253_, _12185_, _06410_);
  and _20591_ (_12254_, _12253_, _04856_);
  and _20592_ (_10202_, _12254_, _12252_);
  and _20593_ (_12256_, _12219_, _07642_);
  or _20594_ (_12257_, _05519_, _06090_);
  not _20595_ (_12258_, _12257_);
  and _20596_ (_12259_, _12219_, _12258_);
  not _20597_ (_12260_, _12259_);
  nand _20598_ (_12261_, _12260_, _12244_);
  and _20599_ (_12262_, _12261_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  or _20600_ (_12263_, _12262_, _12183_);
  or _20601_ (_12264_, _12263_, _12256_);
  nand _20602_ (_12265_, _12183_, _05669_);
  and _20603_ (_12266_, _12265_, _04856_);
  and _20604_ (_10208_, _12266_, _12264_);
  and _20605_ (_12268_, _06705_, _05009_);
  nor _20606_ (_12269_, _05009_, _07113_);
  or _20607_ (_12270_, _12269_, _12268_);
  and _20608_ (_10214_, _12270_, _04856_);
  nor _20609_ (_12271_, _08367_, _08257_);
  and _20610_ (_12272_, _08160_, _08154_);
  nor _20611_ (_12273_, _12272_, _08095_);
  and _20612_ (_12275_, _08103_, _08098_);
  nor _20613_ (_12276_, _12275_, _08154_);
  nor _20614_ (_12277_, _12276_, _12273_);
  not _20615_ (_12278_, _12277_);
  and _20616_ (_12279_, _08160_, _08146_);
  nor _20617_ (_12281_, _12279_, _08116_);
  and _20618_ (_12282_, _12281_, _08106_);
  and _20619_ (_12283_, _08113_, _08102_);
  nor _20620_ (_12284_, _12283_, _08138_);
  nor _20621_ (_12285_, _12284_, _08152_);
  not _20622_ (_12286_, _12285_);
  and _20623_ (_12287_, _08109_, _08104_);
  not _20624_ (_12288_, _08095_);
  and _20625_ (_12289_, _08113_, _08098_);
  nor _20626_ (_12290_, _12289_, _08110_);
  nor _20627_ (_12291_, _12290_, _12288_);
  nor _20628_ (_12292_, _12291_, _12287_);
  and _20629_ (_12293_, _12292_, _12286_);
  and _20630_ (_12294_, _12293_, _12282_);
  and _20631_ (_12296_, _12294_, _12278_);
  not _20632_ (_12297_, _12283_);
  nor _20633_ (_12298_, _08136_, _08126_);
  and _20634_ (_12299_, _12298_, _12297_);
  nor _20635_ (_12301_, _12299_, _08092_);
  not _20636_ (_12302_, _12301_);
  nor _20637_ (_12304_, _08173_, _08122_);
  and _20638_ (_12305_, _12304_, _12302_);
  and _20639_ (_12306_, _08102_, _08097_);
  not _20640_ (_12307_, _12306_);
  nor _20641_ (_12308_, _08157_, _08109_);
  nor _20642_ (_12309_, _12308_, _12307_);
  not _20643_ (_12310_, _08120_);
  or _20644_ (_12311_, _12306_, _12283_);
  not _20645_ (_12312_, _12311_);
  and _20646_ (_12313_, _08135_, _08098_);
  nor _20647_ (_12314_, _12313_, _08104_);
  and _20648_ (_12315_, _12314_, _12312_);
  nor _20649_ (_12316_, _12315_, _12310_);
  nor _20650_ (_12318_, _12316_, _12309_);
  and _20651_ (_12319_, _12318_, _12305_);
  not _20652_ (_12320_, _08147_);
  and _20653_ (_12321_, _08125_, _05895_);
  and _20654_ (_12322_, _08171_, _12321_);
  and _20655_ (_12323_, _08158_, _05843_);
  and _20656_ (_12324_, _12323_, _08093_);
  nor _20657_ (_12325_, _12324_, _12322_);
  and _20658_ (_12326_, _12325_, _12320_);
  and _20659_ (_12327_, _12326_, _08142_);
  and _20660_ (_12328_, _08146_, _08094_);
  nor _20661_ (_12329_, _12328_, _08120_);
  not _20662_ (_12330_, _08126_);
  nor _20663_ (_12331_, _08146_, _08099_);
  and _20664_ (_12332_, _12331_, _12330_);
  nor _20665_ (_12333_, _12332_, _12329_);
  not _20666_ (_12334_, _12333_);
  and _20667_ (_12335_, _12334_, _08134_);
  and _20668_ (_12336_, _12335_, _12327_);
  and _20669_ (_12337_, _08136_, _08120_);
  and _20670_ (_12339_, _08157_, _08153_);
  nor _20671_ (_12340_, _12339_, _12337_);
  nor _20672_ (_12341_, _08119_, _08094_);
  not _20673_ (_12342_, _12341_);
  and _20674_ (_12344_, _12342_, _08131_);
  not _20675_ (_12345_, _08157_);
  nor _20676_ (_12346_, _08126_, _08114_);
  nor _20677_ (_12347_, _12346_, _12345_);
  nor _20678_ (_12348_, _12347_, _12344_);
  and _20679_ (_12349_, _12348_, _12340_);
  nor _20680_ (_12350_, _12298_, _12288_);
  nor _20681_ (_12351_, _12350_, _08156_);
  and _20682_ (_12352_, _08154_, _08117_);
  and _20683_ (_12353_, _12352_, _12342_);
  nor _20684_ (_12354_, _12313_, _12306_);
  nor _20685_ (_12355_, _12354_, _12288_);
  nor _20686_ (_12356_, _12355_, _12353_);
  and _20687_ (_12357_, _12356_, _12351_);
  and _20688_ (_12358_, _12357_, _12349_);
  and _20689_ (_12359_, _12358_, _12336_);
  and _20690_ (_12360_, _12359_, _12319_);
  and _20691_ (_12361_, _12360_, _12296_);
  or _20692_ (_12362_, _12361_, _05737_);
  and _20693_ (_12363_, _08125_, _08112_);
  and _20694_ (_12364_, _12363_, _08160_);
  or _20695_ (_12365_, _12306_, _08153_);
  and _20696_ (_12366_, _12365_, _08109_);
  or _20697_ (_12367_, _12366_, _12350_);
  nor _20698_ (_12368_, _12367_, _12364_);
  and _20699_ (_12369_, _12368_, _12304_);
  nand _20700_ (_12370_, _12369_, _12282_);
  or _20701_ (_12371_, _12370_, _12361_);
  and _20702_ (_12373_, _12371_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nand _20703_ (_12374_, _12361_, _05737_);
  and _20704_ (_12375_, _12374_, _12362_);
  nand _20705_ (_12376_, _12375_, _12373_);
  nand _20706_ (_12377_, _12376_, _12362_);
  and _20707_ (_12378_, _12377_, _05730_);
  and _20708_ (_12379_, _12378_, _05736_);
  nor _20709_ (_12380_, _12378_, _05736_);
  nor _20710_ (_12381_, _12380_, _12379_);
  nor _20711_ (_12382_, _12381_, _12271_);
  and _20712_ (_12383_, _05741_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and _20713_ (_12384_, _12383_, _12271_);
  and _20714_ (_12385_, _12384_, _12370_);
  or _20715_ (_12386_, _12385_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _20716_ (_12387_, _12386_, _12382_);
  and _20717_ (_10221_, _12387_, _04856_);
  and _20718_ (_12388_, _06125_, _06091_);
  and _20719_ (_12389_, _12388_, _12182_);
  not _20720_ (_12390_, _12389_);
  nor _20721_ (_12391_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and _20722_ (_12392_, _12391_, _12221_);
  and _20723_ (_12393_, _12392_, _07391_);
  and _20724_ (_12394_, _12393_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  not _20725_ (_12395_, _12393_);
  and _20726_ (_12396_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  not _20727_ (_12397_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  and _20728_ (_12398_, \oc8051_top_1.oc8051_sfr1.pres_ow , _12397_);
  nor _20729_ (_12399_, _12398_, _12396_);
  not _20730_ (_12400_, _12399_);
  and _20731_ (_12401_, _12400_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and _20732_ (_12402_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and _20733_ (_12403_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and _20734_ (_12404_, _12403_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and _20735_ (_12405_, _12404_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and _20736_ (_12406_, _12405_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and _20737_ (_12407_, _12406_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and _20738_ (_12408_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and _20739_ (_12409_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and _20740_ (_12410_, _12409_, _12408_);
  and _20741_ (_12411_, _12410_, _12407_);
  and _20742_ (_12412_, _12411_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and _20743_ (_12413_, _12412_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and _20744_ (_12414_, _12413_, _12402_);
  and _20745_ (_12415_, _12414_, _12401_);
  nand _20746_ (_12416_, _12415_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or _20747_ (_12417_, _12415_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  and _20748_ (_12418_, _12417_, _12416_);
  and _20749_ (_12419_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  and _20750_ (_12420_, _12419_, _12414_);
  and _20751_ (_12421_, _12391_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  not _20752_ (_12422_, _12421_);
  and _20753_ (_12423_, _12422_, _12401_);
  and _20754_ (_12424_, _12423_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and _20755_ (_12425_, _12424_, _12420_);
  or _20756_ (_12426_, _12425_, _12418_);
  and _20757_ (_12427_, _12426_, _12395_);
  or _20758_ (_12428_, _12427_, _12394_);
  and _20759_ (_12429_, _07855_, _06125_);
  and _20760_ (_12430_, _12429_, _12182_);
  not _20761_ (_12431_, _12430_);
  and _20762_ (_12432_, _12431_, _12428_);
  and _20763_ (_12433_, _12430_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or _20764_ (_12434_, _12433_, _12432_);
  and _20765_ (_12435_, _12434_, _12390_);
  nor _20766_ (_12436_, _12390_, _05287_);
  or _20767_ (_12437_, _12436_, _12435_);
  and _20768_ (_10247_, _12437_, _04856_);
  and _20769_ (_12438_, _12430_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  not _20770_ (_12439_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  and _20771_ (_12440_, _12413_, _12401_);
  and _20772_ (_12441_, _12440_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  nor _20773_ (_12442_, _12441_, _12439_);
  and _20774_ (_12443_, _12441_, _12439_);
  or _20775_ (_12444_, _12443_, _12442_);
  and _20776_ (_12446_, _12423_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and _20777_ (_12447_, _12446_, _12420_);
  or _20778_ (_12448_, _12447_, _12393_);
  or _20779_ (_12449_, _12448_, _12444_);
  not _20780_ (_12450_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  nand _20781_ (_12451_, _12393_, _12450_);
  and _20782_ (_12452_, _12451_, _12449_);
  nor _20783_ (_12453_, _12430_, _12389_);
  and _20784_ (_12454_, _12453_, _12452_);
  and _20785_ (_12455_, _12389_, _05718_);
  or _20786_ (_12456_, _12455_, _12454_);
  or _20787_ (_12457_, _12456_, _12438_);
  and _20788_ (_10250_, _12457_, _04856_);
  or _20789_ (_12458_, _12395_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  nor _20790_ (_12459_, _12440_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  nor _20791_ (_12460_, _12459_, _12441_);
  or _20792_ (_12461_, _12460_, _12393_);
  and _20793_ (_12462_, _12423_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and _20794_ (_12463_, _12462_, _12420_);
  or _20795_ (_12464_, _12463_, _12461_);
  and _20796_ (_12465_, _12464_, _12458_);
  and _20797_ (_12466_, _12465_, _12453_);
  and _20798_ (_12467_, _12389_, _06410_);
  and _20799_ (_12468_, _12430_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or _20800_ (_12469_, _12468_, _12467_);
  or _20801_ (_12470_, _12469_, _12466_);
  and _20802_ (_10257_, _12470_, _04856_);
  and _20803_ (_10265_, _07384_, _04856_);
  and _20804_ (_10297_, _07365_, _04856_);
  and _20805_ (_10301_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _04856_);
  not _20806_ (_12471_, _06809_);
  and _20807_ (_12472_, _08217_, _06858_);
  and _20808_ (_12473_, _12472_, _12471_);
  nor _20809_ (_12474_, _12473_, _05994_);
  and _20810_ (_12475_, _12474_, _06810_);
  nor _20811_ (_12476_, _06268_, _06124_);
  and _20812_ (_12477_, _12476_, _07996_);
  and _20813_ (_12478_, _12477_, _12475_);
  not _20814_ (_12479_, _12478_);
  nor _20815_ (_12480_, _08206_, _05874_);
  not _20816_ (_12481_, _12474_);
  not _20817_ (_12483_, _07789_);
  and _20818_ (_12484_, _07680_, _05617_);
  and _20819_ (_12486_, _12484_, _05597_);
  and _20820_ (_12487_, _12486_, _06508_);
  and _20821_ (_12488_, _12487_, _06561_);
  and _20822_ (_12490_, _12488_, _06810_);
  and _20823_ (_12492_, _12490_, _12483_);
  and _20824_ (_12494_, _12492_, _12481_);
  and _20825_ (_12495_, _12494_, _07871_);
  and _20826_ (_12497_, _12495_, _05634_);
  not _20827_ (_12498_, _12497_);
  and _20828_ (_12499_, _12475_, _06062_);
  nor _20829_ (_12500_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor _20830_ (_12501_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and _20831_ (_12502_, _12501_, _12500_);
  nor _20832_ (_12503_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor _20833_ (_12504_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and _20834_ (_12505_, _12504_, _12503_);
  and _20835_ (_12506_, _12505_, _12502_);
  and _20836_ (_12507_, _12506_, _06807_);
  and _20837_ (_12508_, _06809_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor _20838_ (_12509_, _12508_, _12507_);
  not _20839_ (_12510_, _12509_);
  nor _20840_ (_12511_, _12510_, _12499_);
  and _20841_ (_12512_, _12511_, _12498_);
  or _20842_ (_12513_, _12512_, _08218_);
  nor _20843_ (_12514_, _12513_, _12480_);
  or _20844_ (_12515_, _06635_, _06737_);
  and _20845_ (_12516_, _12515_, _05983_);
  not _20846_ (_12517_, _12516_);
  not _20847_ (_12518_, _07511_);
  nor _20848_ (_12519_, _09066_, _06610_);
  and _20849_ (_12520_, _12519_, _12518_);
  and _20850_ (_12521_, _06638_, _06612_);
  nor _20851_ (_12522_, _12521_, _08214_);
  and _20852_ (_12523_, _12522_, _12520_);
  and _20853_ (_12524_, _12523_, _12517_);
  and _20854_ (_12525_, _12524_, _12512_);
  nor _20855_ (_12526_, _12525_, _12514_);
  nor _20856_ (_12527_, _08213_, _09088_);
  and _20857_ (_12528_, _12527_, _06824_);
  not _20858_ (_12529_, _12528_);
  nor _20859_ (_12530_, _12529_, _12526_);
  nor _20860_ (_12531_, _12530_, _06647_);
  and _20861_ (_12532_, _05949_, _05849_);
  nor _20862_ (_12533_, _12532_, _05954_);
  nor _20863_ (_12534_, _06799_, _12533_);
  nor _20864_ (_12535_, _12534_, _06847_);
  not _20865_ (_12536_, _12535_);
  nor _20866_ (_12537_, _12536_, _12531_);
  not _20867_ (_12538_, _06807_);
  nor _20868_ (_12539_, _12538_, _06678_);
  nor _20869_ (_12540_, _08277_, _07951_);
  and _20870_ (_12541_, _12540_, _06935_);
  nor _20871_ (_12542_, _12541_, _12471_);
  nor _20872_ (_12543_, _12542_, _12539_);
  not _20873_ (_12544_, _12543_);
  nor _20874_ (_12545_, _12544_, _12537_);
  and _20875_ (_12546_, _12545_, _07993_);
  and _20876_ (_12547_, _12546_, _12479_);
  nand _20877_ (_12548_, _12547_, _06901_);
  nor _20878_ (_10310_, _12548_, rst);
  not _20879_ (_12549_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  nand _20880_ (_12550_, _12393_, _12549_);
  and _20881_ (_12551_, _12407_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and _20882_ (_12552_, _12551_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and _20883_ (_12553_, _12552_, _12401_);
  and _20884_ (_12554_, _12553_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nand _20885_ (_12555_, _12554_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  or _20886_ (_12556_, _12554_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and _20887_ (_12557_, _12556_, _12555_);
  or _20888_ (_12558_, _12557_, _12393_);
  and _20889_ (_12559_, _12423_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  and _20890_ (_12560_, _12559_, _12420_);
  or _20891_ (_12561_, _12560_, _12558_);
  and _20892_ (_12562_, _12561_, _12550_);
  and _20893_ (_12563_, _12562_, _12453_);
  nor _20894_ (_12564_, _12390_, _06032_);
  and _20895_ (_12565_, _12430_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  or _20896_ (_12566_, _12565_, _12564_);
  or _20897_ (_12567_, _12566_, _12563_);
  and _20898_ (_10337_, _12567_, _04856_);
  or _20899_ (_12568_, _12395_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  nor _20900_ (_12569_, _12553_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nor _20901_ (_12570_, _12569_, _12554_);
  or _20902_ (_12571_, _12570_, _12393_);
  and _20903_ (_12572_, _12423_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  and _20904_ (_12573_, _12572_, _12420_);
  or _20905_ (_12574_, _12573_, _12571_);
  and _20906_ (_12575_, _12574_, _12568_);
  and _20907_ (_12576_, _12575_, _12453_);
  and _20908_ (_12577_, _12389_, _06997_);
  and _20909_ (_12578_, _12430_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  or _20910_ (_12579_, _12578_, _12577_);
  or _20911_ (_12581_, _12579_, _12576_);
  and _20912_ (_10344_, _12581_, _04856_);
  or _20913_ (_12582_, _12401_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and _20914_ (_12583_, _12401_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and _20915_ (_12584_, _12422_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  nand _20916_ (_12585_, _12584_, _12420_);
  nand _20917_ (_12586_, _12585_, _12583_);
  and _20918_ (_12587_, _12586_, _12582_);
  or _20919_ (_12588_, _12587_, _12393_);
  nor _20920_ (_12589_, _12395_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  nor _20921_ (_12590_, _12589_, _12430_);
  and _20922_ (_12591_, _12590_, _12588_);
  and _20923_ (_12592_, _12430_, _06997_);
  or _20924_ (_12593_, _12592_, _12389_);
  or _20925_ (_12594_, _12593_, _12591_);
  or _20926_ (_12595_, _12390_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and _20927_ (_12596_, _12595_, _04856_);
  and _20928_ (_10374_, _12596_, _12594_);
  nor _20929_ (_12597_, _12431_, _05287_);
  or _20930_ (_12598_, _12395_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and _20931_ (_12599_, _12423_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and _20932_ (_12600_, _12599_, _12420_);
  and _20933_ (_12601_, _12407_, _12401_);
  and _20934_ (_12602_, _12601_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  nor _20935_ (_12603_, _12601_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  nor _20936_ (_12604_, _12603_, _12602_);
  or _20937_ (_12605_, _12604_, _12393_);
  or _20938_ (_12606_, _12605_, _12600_);
  nand _20939_ (_12607_, _12606_, _12598_);
  nor _20940_ (_12608_, _12607_, _12430_);
  or _20941_ (_12609_, _12608_, _12389_);
  or _20942_ (_12610_, _12609_, _12597_);
  or _20943_ (_12611_, _12390_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and _20944_ (_12612_, _12611_, _04856_);
  and _20945_ (_10416_, _12612_, _12610_);
  or _20946_ (_12613_, _12431_, _05718_);
  and _20947_ (_12614_, _12406_, _12401_);
  nor _20948_ (_12615_, _12614_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  nor _20949_ (_12616_, _12615_, _12601_);
  and _20950_ (_12617_, _12423_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and _20951_ (_12618_, _12617_, _12420_);
  or _20952_ (_12619_, _12618_, _12616_);
  and _20953_ (_12620_, _12619_, _12395_);
  and _20954_ (_12622_, _12393_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  or _20955_ (_12623_, _12622_, _12620_);
  or _20956_ (_12624_, _12623_, _12430_);
  and _20957_ (_12625_, _12624_, _12613_);
  or _20958_ (_12626_, _12625_, _12389_);
  not _20959_ (_12627_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  nand _20960_ (_12628_, _12389_, _12627_);
  and _20961_ (_12629_, _12628_, _04856_);
  and _20962_ (_10419_, _12629_, _12626_);
  or _20963_ (_12630_, _12395_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and _20964_ (_12631_, _12423_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and _20965_ (_12632_, _12631_, _12420_);
  not _20966_ (_12633_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  nand _20967_ (_12634_, _12405_, _12401_);
  and _20968_ (_12635_, _12634_, _12633_);
  nor _20969_ (_12636_, _12635_, _12614_);
  or _20970_ (_12637_, _12636_, _12393_);
  or _20971_ (_12638_, _12637_, _12632_);
  and _20972_ (_12639_, _12638_, _12630_);
  or _20973_ (_12640_, _12639_, _12430_);
  or _20974_ (_12641_, _12431_, _06410_);
  and _20975_ (_12642_, _12641_, _12640_);
  or _20976_ (_12643_, _12642_, _12389_);
  nand _20977_ (_12644_, _12389_, _12633_);
  and _20978_ (_12645_, _12644_, _04856_);
  and _20979_ (_10424_, _12645_, _12643_);
  and _20980_ (_12647_, _12404_, _12401_);
  or _20981_ (_12648_, _12647_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and _20982_ (_12649_, _12648_, _12634_);
  and _20983_ (_12650_, _12423_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and _20984_ (_12651_, _12650_, _12420_);
  or _20985_ (_12652_, _12651_, _12649_);
  and _20986_ (_12653_, _12652_, _12395_);
  and _20987_ (_12654_, _12393_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  or _20988_ (_12655_, _12654_, _12653_);
  or _20989_ (_12656_, _12655_, _12430_);
  nand _20990_ (_12657_, _12430_, _05669_);
  and _20991_ (_12658_, _12657_, _12656_);
  or _20992_ (_12659_, _12658_, _12389_);
  nand _20993_ (_12660_, _12389_, _08788_);
  and _20994_ (_12661_, _12660_, _04856_);
  and _20995_ (_10427_, _12661_, _12659_);
  and _20996_ (_12662_, _12423_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and _20997_ (_12663_, _12662_, _12420_);
  nand _20998_ (_12664_, _12403_, _12401_);
  and _20999_ (_12665_, _12664_, _08898_);
  nor _21000_ (_12666_, _12665_, _12647_);
  or _21001_ (_12667_, _12666_, _12393_);
  or _21002_ (_12668_, _12667_, _12663_);
  or _21003_ (_12669_, _12395_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  nand _21004_ (_12671_, _12669_, _12668_);
  nor _21005_ (_12672_, _12671_, _12430_);
  and _21006_ (_12674_, _12430_, _06705_);
  or _21007_ (_12675_, _12674_, _12389_);
  or _21008_ (_12676_, _12675_, _12672_);
  nand _21009_ (_12677_, _12389_, _08898_);
  and _21010_ (_12678_, _12677_, _04856_);
  and _21011_ (_10434_, _12678_, _12676_);
  and _21012_ (_12680_, _06721_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  or _21013_ (_12681_, _08197_, _06878_);
  and _21014_ (_12682_, _06594_, _05998_);
  or _21015_ (_12683_, _12682_, _06726_);
  and _21016_ (_12684_, _08198_, _05773_);
  or _21017_ (_12685_, _06625_, _12684_);
  or _21018_ (_12686_, _12685_, _12683_);
  or _21019_ (_12687_, _12686_, _12681_);
  or _21020_ (_12688_, _06865_, _06729_);
  and _21021_ (_12689_, _06624_, _06731_);
  and _21022_ (_12691_, _06745_, _06598_);
  or _21023_ (_12692_, _12691_, _12689_);
  or _21024_ (_12693_, _12692_, _12688_);
  and _21025_ (_12695_, _06857_, _06598_);
  or _21026_ (_12696_, _08193_, _12695_);
  and _21027_ (_12697_, _06598_, _06612_);
  or _21028_ (_12698_, _08246_, _06789_);
  or _21029_ (_12699_, _12698_, _12697_);
  or _21030_ (_12700_, _12699_, _12696_);
  and _21031_ (_12701_, _06857_, _06638_);
  or _21032_ (_12703_, _09075_, _06628_);
  or _21033_ (_12704_, _12703_, _12701_);
  or _21034_ (_12705_, _06835_, _06746_);
  or _21035_ (_12707_, _12705_, _12704_);
  or _21036_ (_12708_, _12707_, _12700_);
  or _21037_ (_12709_, _12708_, _12693_);
  or _21038_ (_12710_, _12709_, _12687_);
  and _21039_ (_12711_, _12710_, _06770_);
  or _21040_ (_10443_, _12711_, _12680_);
  and _21041_ (_12713_, _06125_, _05520_);
  and _21042_ (_12714_, _12713_, _12182_);
  not _21043_ (_12715_, _12714_);
  and _21044_ (_12716_, _12421_, _12221_);
  not _21045_ (_12717_, _12716_);
  and _21046_ (_12718_, _06494_, _06125_);
  and _21047_ (_12719_, _12718_, _12182_);
  nor _21048_ (_12720_, _12719_, _12717_);
  or _21049_ (_12721_, _12720_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  nand _21050_ (_12722_, _12720_, _08901_);
  and _21051_ (_12723_, _12722_, _12721_);
  and _21052_ (_12724_, _12723_, _12715_);
  and _21053_ (_12725_, _12714_, _06705_);
  or _21054_ (_12726_, _12725_, _12724_);
  and _21055_ (_10471_, _12726_, _04856_);
  or _21056_ (_12727_, _12720_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  not _21057_ (_12728_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  nand _21058_ (_12729_, _12720_, _12728_);
  and _21059_ (_12730_, _12729_, _12727_);
  or _21060_ (_12731_, _12730_, _12714_);
  nand _21061_ (_12732_, _12714_, _06032_);
  and _21062_ (_12733_, _12732_, _04856_);
  and _21063_ (_10473_, _12733_, _12731_);
  or _21064_ (_12734_, _12720_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  not _21065_ (_12735_, _12720_);
  or _21066_ (_12737_, _12735_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and _21067_ (_12738_, _12737_, _12734_);
  or _21068_ (_12739_, _12738_, _12714_);
  nand _21069_ (_12740_, _12714_, _06369_);
  and _21070_ (_12741_, _12740_, _04856_);
  and _21071_ (_10478_, _12741_, _12739_);
  and _21072_ (_12742_, _12735_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and _21073_ (_12743_, _12720_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or _21074_ (_12744_, _12743_, _12742_);
  and _21075_ (_12745_, _12744_, _12715_);
  and _21076_ (_12746_, _12714_, _06410_);
  or _21077_ (_12747_, _12746_, _12745_);
  and _21078_ (_10499_, _12747_, _04856_);
  nand _21079_ (_12748_, _12714_, _05287_);
  and _21080_ (_12749_, _12735_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and _21081_ (_12751_, _12720_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or _21082_ (_12752_, _12751_, _12749_);
  or _21083_ (_12753_, _12752_, _12714_);
  and _21084_ (_12754_, _12753_, _04856_);
  and _21085_ (_10507_, _12754_, _12748_);
  or _21086_ (_12755_, _12715_, _05718_);
  nor _21087_ (_12756_, _12720_, _12450_);
  and _21088_ (_12757_, _12720_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or _21089_ (_12758_, _12757_, _12756_);
  or _21090_ (_12759_, _12758_, _12714_);
  and _21091_ (_12760_, _12759_, _04856_);
  and _21092_ (_10514_, _12760_, _12755_);
  nor _21093_ (_12761_, _10231_, _10232_);
  and _21094_ (_12762_, _08067_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  and _21095_ (_12763_, _12762_, _10230_);
  or _21096_ (_12764_, _12763_, _12761_);
  and _21097_ (_12765_, _12764_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  and _21098_ (_12766_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], _09249_);
  nand _21099_ (_12767_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor _21100_ (_12768_, _12767_, _08087_);
  or _21101_ (_12769_, _12768_, _12766_);
  or _21102_ (_12770_, _12769_, _12765_);
  and _21103_ (_10531_, _12770_, _04856_);
  not _21104_ (_12771_, _12719_);
  or _21105_ (_12772_, _12771_, _06705_);
  and _21106_ (_12773_, _12717_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and _21107_ (_12774_, _12716_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or _21108_ (_12775_, _12774_, _12773_);
  or _21109_ (_12776_, _12775_, _12719_);
  and _21110_ (_12777_, _12776_, _12715_);
  and _21111_ (_12778_, _12777_, _12772_);
  and _21112_ (_12779_, _12714_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  or _21113_ (_12780_, _12779_, _12778_);
  and _21114_ (_10547_, _12780_, _04856_);
  nor _21115_ (_12781_, _12771_, _05287_);
  and _21116_ (_12782_, _12717_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and _21117_ (_12783_, _12716_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  nor _21118_ (_12784_, _12783_, _12782_);
  nor _21119_ (_12785_, _12784_, _12719_);
  or _21120_ (_12786_, _12785_, _12714_);
  or _21121_ (_12787_, _12786_, _12781_);
  or _21122_ (_12788_, _12715_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and _21123_ (_12789_, _12788_, _04856_);
  and _21124_ (_10549_, _12789_, _12787_);
  or _21125_ (_12790_, _12771_, _05718_);
  not _21126_ (_12791_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  nor _21127_ (_12792_, _12716_, _12791_);
  and _21128_ (_12793_, _12716_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or _21129_ (_12794_, _12793_, _12792_);
  or _21130_ (_12795_, _12794_, _12719_);
  and _21131_ (_12796_, _12795_, _12715_);
  and _21132_ (_12797_, _12796_, _12790_);
  and _21133_ (_12798_, _12714_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  or _21134_ (_12799_, _12798_, _12797_);
  and _21135_ (_10553_, _12799_, _04856_);
  or _21136_ (_12800_, _12771_, _06410_);
  and _21137_ (_12801_, _12717_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and _21138_ (_12802_, _12716_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or _21139_ (_12803_, _12802_, _12801_);
  or _21140_ (_12804_, _12803_, _12719_);
  and _21141_ (_12805_, _12804_, _12715_);
  and _21142_ (_12806_, _12805_, _12800_);
  and _21143_ (_12807_, _12714_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  or _21144_ (_12808_, _12807_, _12806_);
  and _21145_ (_10557_, _12808_, _04856_);
  nand _21146_ (_12809_, _12719_, _05669_);
  and _21147_ (_12810_, _12717_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and _21148_ (_12811_, _12716_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or _21149_ (_12812_, _12811_, _12810_);
  or _21150_ (_12813_, _12812_, _12719_);
  and _21151_ (_12814_, _12813_, _12715_);
  and _21152_ (_12815_, _12814_, _12809_);
  and _21153_ (_12816_, _12714_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  or _21154_ (_12817_, _12816_, _12815_);
  and _21155_ (_10566_, _12817_, _04856_);
  nor _21156_ (_12818_, _12761_, _09249_);
  or _21157_ (_12820_, _12818_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2]);
  or _21158_ (_12821_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _09249_);
  or _21159_ (_12822_, _12821_, _08087_);
  and _21160_ (_12823_, _12822_, _04856_);
  and _21161_ (_10761_, _12823_, _12820_);
  and _21162_ (_10850_, _05847_, _04856_);
  not _21163_ (_12824_, _05823_);
  and _21164_ (_12825_, _06612_, _12824_);
  nor _21165_ (_12826_, _12825_, _06610_);
  nand _21166_ (_12827_, _12826_, _12472_);
  nand _21167_ (_12828_, _12827_, _05959_);
  and _21168_ (_12829_, _05962_, _12532_);
  not _21169_ (_12830_, _12829_);
  and _21170_ (_12831_, _06822_, _05962_);
  and _21171_ (_12832_, _12831_, _05983_);
  nor _21172_ (_12833_, _12832_, _06847_);
  and _21173_ (_12834_, _12833_, _12830_);
  nand _21174_ (_12835_, _12834_, _12828_);
  or _21175_ (_12836_, _12835_, _07261_);
  and _21176_ (_12837_, _12834_, _12828_);
  nor _21177_ (_12838_, _05730_, _05177_);
  and _21178_ (_12839_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and _21179_ (_12840_, _05929_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and _21180_ (_12841_, _05742_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor _21181_ (_12842_, _12841_, _12840_);
  and _21182_ (_12843_, _05933_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and _21183_ (_12844_, _05935_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor _21184_ (_12845_, _12844_, _12843_);
  and _21185_ (_12846_, _12845_, _12842_);
  and _21186_ (_12847_, _05927_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and _21187_ (_12848_, _05758_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor _21188_ (_12849_, _12848_, _12847_);
  and _21189_ (_12850_, _12849_, _12846_);
  nor _21190_ (_12851_, _12850_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _21191_ (_12852_, _12851_, _12839_);
  nor _21192_ (_12853_, _12852_, _08257_);
  nor _21193_ (_12854_, _12853_, _12838_);
  or _21194_ (_12855_, _12854_, _12837_);
  and _21195_ (_12856_, _12855_, _12836_);
  or _21196_ (_12857_, _12856_, _05183_);
  nand _21197_ (_12858_, _12856_, _05183_);
  and _21198_ (_12859_, _12858_, _12857_);
  not _21199_ (_12860_, _07191_);
  and _21200_ (_12861_, _12837_, _12860_);
  nor _21201_ (_12862_, _05730_, _05060_);
  and _21202_ (_12863_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and _21203_ (_12864_, _05933_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and _21204_ (_12865_, _05758_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor _21205_ (_12866_, _12865_, _12864_);
  and _21206_ (_12867_, _05927_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and _21207_ (_12868_, _05935_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor _21208_ (_12869_, _12868_, _12867_);
  and _21209_ (_12870_, _05742_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  and _21210_ (_12871_, _05929_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nor _21211_ (_12872_, _12871_, _12870_);
  and _21212_ (_12873_, _12872_, _12869_);
  and _21213_ (_12874_, _12873_, _12866_);
  nor _21214_ (_12875_, _12874_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _21215_ (_12876_, _12875_, _12863_);
  nor _21216_ (_12877_, _12876_, _08257_);
  nor _21217_ (_12878_, _12877_, _12862_);
  not _21218_ (_12879_, _12878_);
  and _21219_ (_12880_, _12879_, _12835_);
  nor _21220_ (_12881_, _12880_, _12861_);
  not _21221_ (_12882_, _12881_);
  and _21222_ (_12883_, _12882_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  not _21223_ (_12884_, _12883_);
  not _21224_ (_12885_, _07142_);
  and _21225_ (_12886_, _12837_, _12885_);
  nor _21226_ (_12887_, _05730_, _05082_);
  and _21227_ (_12888_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and _21228_ (_12889_, _05929_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and _21229_ (_12890_, _05742_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor _21230_ (_12891_, _12890_, _12889_);
  and _21231_ (_12892_, _05933_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and _21232_ (_12893_, _05935_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor _21233_ (_12894_, _12893_, _12892_);
  and _21234_ (_12895_, _12894_, _12891_);
  and _21235_ (_12896_, _05927_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and _21236_ (_12897_, _05758_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor _21237_ (_12898_, _12897_, _12896_);
  and _21238_ (_12899_, _12898_, _12895_);
  nor _21239_ (_12900_, _12899_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _21240_ (_12901_, _12900_, _12888_);
  nor _21241_ (_12902_, _12901_, _08257_);
  nor _21242_ (_12903_, _12902_, _12887_);
  not _21243_ (_12904_, _12903_);
  and _21244_ (_12905_, _12904_, _12835_);
  nor _21245_ (_12906_, _12905_, _12886_);
  and _21246_ (_12907_, _12906_, _05087_);
  nor _21247_ (_12908_, _12906_, _05087_);
  or _21248_ (_12909_, _12835_, _07089_);
  nor _21249_ (_12910_, _05730_, _05154_);
  and _21250_ (_12911_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and _21251_ (_12912_, _05927_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and _21252_ (_12913_, _05742_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor _21253_ (_12914_, _12913_, _12912_);
  and _21254_ (_12915_, _05929_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and _21255_ (_12916_, _05758_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor _21256_ (_12917_, _12916_, _12915_);
  and _21257_ (_12918_, _05933_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and _21258_ (_12919_, _05935_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor _21259_ (_12920_, _12919_, _12918_);
  and _21260_ (_12921_, _12920_, _12917_);
  and _21261_ (_12922_, _12921_, _12914_);
  nor _21262_ (_12923_, _12922_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _21263_ (_12924_, _12923_, _12911_);
  nor _21264_ (_12925_, _12924_, _08257_);
  nor _21265_ (_12926_, _12925_, _12910_);
  or _21266_ (_12927_, _12926_, _12837_);
  and _21267_ (_12928_, _12927_, _12909_);
  or _21268_ (_12929_, _12928_, _05159_);
  not _21269_ (_12930_, _12929_);
  not _21270_ (_12931_, _07032_);
  or _21271_ (_12932_, _12835_, _12931_);
  nor _21272_ (_12933_, _05730_, _05135_);
  and _21273_ (_12934_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and _21274_ (_12935_, _05929_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and _21275_ (_12936_, _05742_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor _21276_ (_12937_, _12936_, _12935_);
  and _21277_ (_12938_, _05933_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and _21278_ (_12939_, _05935_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nor _21279_ (_12940_, _12939_, _12938_);
  and _21280_ (_12941_, _12940_, _12937_);
  and _21281_ (_12942_, _05927_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and _21282_ (_12943_, _05758_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor _21283_ (_12944_, _12943_, _12942_);
  and _21284_ (_12945_, _12944_, _12941_);
  nor _21285_ (_12946_, _12945_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _21286_ (_12947_, _12946_, _12934_);
  nor _21287_ (_12948_, _12947_, _08257_);
  nor _21288_ (_12949_, _12948_, _12933_);
  nand _21289_ (_12950_, _12949_, _12835_);
  and _21290_ (_12952_, _12950_, _12932_);
  nand _21291_ (_12953_, _12952_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  not _21292_ (_12954_, _06925_);
  and _21293_ (_12955_, _12837_, _12954_);
  nor _21294_ (_12956_, _05730_, _05106_);
  and _21295_ (_12957_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and _21296_ (_12958_, _05927_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and _21297_ (_12959_, _05742_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor _21298_ (_12960_, _12959_, _12958_);
  and _21299_ (_12961_, _05929_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and _21300_ (_12962_, _05758_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor _21301_ (_12963_, _12962_, _12961_);
  and _21302_ (_12964_, _05933_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and _21303_ (_12965_, _05935_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor _21304_ (_12966_, _12965_, _12964_);
  and _21305_ (_12967_, _12966_, _12963_);
  and _21306_ (_12968_, _12967_, _12960_);
  nor _21307_ (_12969_, _12968_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _21308_ (_12970_, _12969_, _12957_);
  nor _21309_ (_12971_, _12970_, _08257_);
  nor _21310_ (_12972_, _12971_, _12956_);
  not _21311_ (_12973_, _12972_);
  and _21312_ (_12974_, _12973_, _12835_);
  or _21313_ (_12975_, _12974_, _12955_);
  and _21314_ (_12976_, _12975_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  or _21315_ (_12977_, _12952_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and _21316_ (_12978_, _12977_, _12953_);
  and _21317_ (_12979_, _12978_, _12976_);
  not _21318_ (_12980_, _12979_);
  nand _21319_ (_12981_, _12980_, _12953_);
  nand _21320_ (_12982_, _12928_, _05159_);
  and _21321_ (_12983_, _12982_, _12929_);
  and _21322_ (_12984_, _12983_, _12981_);
  or _21323_ (_12985_, _12984_, _12930_);
  nor _21324_ (_12986_, _12985_, _12908_);
  nor _21325_ (_12987_, _12986_, _12907_);
  nor _21326_ (_12988_, _12882_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nor _21327_ (_12989_, _12988_, _12883_);
  nand _21328_ (_12990_, _12989_, _12987_);
  nand _21329_ (_12991_, _12990_, _12884_);
  and _21330_ (_12992_, _12991_, _12859_);
  not _21331_ (_12993_, _12992_);
  nand _21332_ (_12994_, _12993_, _12857_);
  not _21333_ (_12995_, _07294_);
  and _21334_ (_12996_, _12837_, _12995_);
  nor _21335_ (_12997_, _05730_, _05011_);
  and _21336_ (_12998_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and _21337_ (_12999_, _05929_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and _21338_ (_13000_, _05742_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor _21339_ (_13001_, _13000_, _12999_);
  and _21340_ (_13003_, _05933_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and _21341_ (_13004_, _05935_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor _21342_ (_13005_, _13004_, _13003_);
  and _21343_ (_13006_, _13005_, _13001_);
  and _21344_ (_13007_, _05927_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and _21345_ (_13008_, _05758_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor _21346_ (_13009_, _13008_, _13007_);
  and _21347_ (_13010_, _13009_, _13006_);
  nor _21348_ (_13011_, _13010_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _21349_ (_13012_, _13011_, _12998_);
  nor _21350_ (_13013_, _13012_, _08257_);
  nor _21351_ (_13014_, _13013_, _12997_);
  nor _21352_ (_13015_, _13014_, _12837_);
  nor _21353_ (_13016_, _13015_, _12996_);
  nor _21354_ (_13017_, _13016_, _05026_);
  and _21355_ (_13018_, _13016_, _05026_);
  nor _21356_ (_13019_, _13018_, _13017_);
  nand _21357_ (_13020_, _13019_, _12994_);
  or _21358_ (_13021_, _13019_, _12994_);
  and _21359_ (_13022_, _09088_, _05959_);
  nor _21360_ (_13023_, _13022_, _12534_);
  or _21361_ (_13024_, _13023_, _12835_);
  nor _21362_ (_13025_, _12521_, _08207_);
  and _21363_ (_13026_, _13025_, _12472_);
  and _21364_ (_13027_, _12527_, _12520_);
  and _21365_ (_13028_, _13027_, _13026_);
  nor _21366_ (_13029_, _13028_, _06647_);
  or _21367_ (_13030_, _13029_, _12832_);
  and _21368_ (_13031_, _13030_, _13024_);
  and _21369_ (_13032_, _13031_, _13021_);
  and _21370_ (_13033_, _13032_, _13020_);
  not _21371_ (_13034_, _06488_);
  nor _21372_ (_13035_, _13030_, _12835_);
  and _21373_ (_13036_, _13035_, _13023_);
  or _21374_ (_13037_, _13036_, _13022_);
  and _21375_ (_13038_, _13037_, _13034_);
  and _21376_ (_13039_, _05983_, _05962_);
  and _21377_ (_13040_, _13039_, _06822_);
  or _21378_ (_13041_, _13029_, _13040_);
  nor _21379_ (_13042_, _13041_, _13024_);
  and _21380_ (_13043_, _13042_, _12995_);
  and _21381_ (_13044_, _06847_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and _21382_ (_13045_, _13015_, _12534_);
  or _21383_ (_13046_, _13045_, _13044_);
  or _21384_ (_13047_, _13046_, _13043_);
  or _21385_ (_13048_, _13047_, _13038_);
  or _21386_ (_13049_, _13048_, _13033_);
  and _21387_ (_13050_, _13049_, _12547_);
  and _21388_ (_13051_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3], \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and _21389_ (_13052_, _13051_, _08368_);
  and _21390_ (_13053_, _13052_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and _21391_ (_13055_, _13053_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor _21392_ (_13056_, _13053_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or _21393_ (_13057_, _13056_, _13055_);
  nor _21394_ (_13058_, _13057_, _12547_);
  or _21395_ (_13059_, _13058_, _13050_);
  and _21396_ (_10866_, _13059_, _04856_);
  not _21397_ (_13060_, _07897_);
  and _21398_ (_13061_, _13037_, _13060_);
  nor _21399_ (_13062_, _12854_, _12830_);
  not _21400_ (_13063_, _07261_);
  and _21401_ (_13065_, _13042_, _13063_);
  and _21402_ (_13066_, _06847_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  or _21403_ (_13067_, _13066_, _13065_);
  or _21404_ (_13068_, _13067_, _13062_);
  or _21405_ (_13069_, _13068_, _13061_);
  and _21406_ (_13070_, _13041_, _13024_);
  nor _21407_ (_13071_, _12991_, _12859_);
  nor _21408_ (_13072_, _13071_, _12992_);
  and _21409_ (_13073_, _13072_, _13070_);
  or _21410_ (_13074_, _13073_, _13069_);
  and _21411_ (_13075_, _13074_, _12547_);
  nor _21412_ (_13076_, _13052_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  or _21413_ (_13077_, _13076_, _13053_);
  nor _21414_ (_13078_, _13077_, _12547_);
  or _21415_ (_13079_, _13078_, _13075_);
  and _21416_ (_10869_, _13079_, _04856_);
  nor _21417_ (_10883_, _13014_, rst);
  nor _21418_ (_13080_, _07774_, _06901_);
  and _21419_ (_13081_, _12829_, _12931_);
  or _21420_ (_13082_, _13081_, _13080_);
  and _21421_ (_13083_, _13042_, _05943_);
  and _21422_ (_13084_, _13036_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  or _21423_ (_13085_, _13084_, _13083_);
  or _21424_ (_13086_, _13085_, _13082_);
  not _21425_ (_13087_, _07380_);
  and _21426_ (_13088_, _12837_, _13087_);
  not _21427_ (_13089_, _08273_);
  and _21428_ (_13090_, _12835_, _13089_);
  nor _21429_ (_13091_, _13090_, _13088_);
  not _21430_ (_13092_, _13091_);
  nor _21431_ (_13093_, _13091_, _05327_);
  not _21432_ (_13094_, _13017_);
  and _21433_ (_13095_, _13091_, _05327_);
  nor _21434_ (_13096_, _13095_, _13094_);
  nor _21435_ (_13097_, _13096_, _13093_);
  nand _21436_ (_13098_, _12883_, _12859_);
  nand _21437_ (_13099_, _13098_, _12857_);
  nor _21438_ (_13100_, _13095_, _13093_);
  and _21439_ (_13101_, _13100_, _13019_);
  nand _21440_ (_13102_, _13101_, _13099_);
  and _21441_ (_13103_, _13102_, _13097_);
  and _21442_ (_13104_, _12989_, _12859_);
  and _21443_ (_13105_, _13101_, _13104_);
  nand _21444_ (_13106_, _13105_, _12987_);
  and _21445_ (_13107_, _13106_, _13103_);
  and _21446_ (_13108_, _13107_, _05111_);
  and _21447_ (_13109_, _13108_, _13092_);
  nor _21448_ (_13110_, _13107_, _05111_);
  and _21449_ (_13111_, _13110_, _13091_);
  nor _21450_ (_13112_, _13111_, _13109_);
  nand _21451_ (_13113_, _13112_, _05142_);
  or _21452_ (_13114_, _13112_, _05142_);
  and _21453_ (_13115_, _13114_, _13070_);
  and _21454_ (_13116_, _13115_, _13113_);
  or _21455_ (_13117_, _13116_, _13086_);
  nand _21456_ (_13118_, _13022_, _07743_);
  nand _21457_ (_13119_, _13118_, _12547_);
  or _21458_ (_13120_, _13119_, _13117_);
  and _21459_ (_13121_, _13055_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and _21460_ (_13122_, _13121_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor _21461_ (_13123_, _13122_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and _21462_ (_13124_, _13122_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  nor _21463_ (_13125_, _13124_, _13123_);
  or _21464_ (_13126_, _13125_, _12547_);
  and _21465_ (_13127_, _13126_, _04856_);
  and _21466_ (_10889_, _13127_, _13120_);
  and _21467_ (_13128_, _06688_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  and _21468_ (_13129_, _06370_, _05679_);
  or _21469_ (_13130_, _13129_, _13128_);
  and _21470_ (_10893_, _13130_, _04856_);
  and _21471_ (_13131_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and _21472_ (_13132_, _12165_, \oc8051_top_1.oc8051_rom1.data_o [24]);
  or _21473_ (_13133_, _13132_, _13131_);
  and _21474_ (_10902_, _13133_, _04856_);
  or _21475_ (_13134_, _08367_, \oc8051_top_1.oc8051_rom1.data_o [12]);
  nand _21476_ (_13135_, _08367_, _05861_);
  and _21477_ (_13136_, _13135_, _04856_);
  and _21478_ (_10908_, _13136_, _13134_);
  nor _21479_ (_13137_, _13121_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor _21480_ (_13138_, _13137_, _13122_);
  or _21481_ (_13139_, _13138_, _12547_);
  and _21482_ (_13140_, _13139_, _04856_);
  nor _21483_ (_13141_, _13107_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and _21484_ (_13142_, _13107_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor _21485_ (_13143_, _13142_, _13141_);
  nor _21486_ (_13144_, _13143_, _13092_);
  and _21487_ (_13145_, _13143_, _13092_);
  or _21488_ (_13146_, _13145_, _13144_);
  and _21489_ (_13147_, _13146_, _13031_);
  and _21490_ (_13148_, _13022_, _07676_);
  and _21491_ (_13149_, _13042_, _05895_);
  and _21492_ (_13150_, _12829_, _12954_);
  or _21493_ (_13151_, _13150_, _13149_);
  and _21494_ (_13152_, _13036_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  not _21495_ (_13153_, _07702_);
  and _21496_ (_13154_, _13153_, _06847_);
  or _21497_ (_13155_, _13154_, _13152_);
  or _21498_ (_13156_, _13155_, _13151_);
  nor _21499_ (_13157_, _13156_, _13148_);
  nand _21500_ (_13159_, _13157_, _12547_);
  or _21501_ (_13160_, _13159_, _13147_);
  and _21502_ (_10911_, _13160_, _13140_);
  and _21503_ (_13161_, _13020_, _13094_);
  nor _21504_ (_13162_, _13161_, _13100_);
  and _21505_ (_13163_, _13161_, _13100_);
  or _21506_ (_13164_, _13163_, _13162_);
  and _21507_ (_13166_, _13164_, _13031_);
  and _21508_ (_13167_, _13037_, _05641_);
  and _21509_ (_13169_, _12829_, _13089_);
  and _21510_ (_13170_, _13088_, _12534_);
  and _21511_ (_13171_, _06847_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  or _21512_ (_13172_, _13171_, _13170_);
  or _21513_ (_13173_, _13172_, _13169_);
  or _21514_ (_13174_, _13173_, _13167_);
  or _21515_ (_13175_, _13174_, _13166_);
  and _21516_ (_13176_, _13175_, _12547_);
  nor _21517_ (_13177_, _13055_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  or _21518_ (_13178_, _13177_, _13121_);
  nor _21519_ (_13179_, _13178_, _12547_);
  or _21520_ (_13180_, _13179_, _13176_);
  and _21521_ (_10919_, _13180_, _04856_);
  and _21522_ (_13181_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _04856_);
  and _21523_ (_13182_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _04856_);
  and _21524_ (_13183_, _13182_, _12206_);
  or _21525_ (_10992_, _13183_, _13181_);
  and _21526_ (_11042_, _05772_, _04856_);
  and _21527_ (_13184_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and _21528_ (_13185_, _12165_, \oc8051_top_1.oc8051_rom1.data_o [25]);
  or _21529_ (_13186_, _13185_, _13184_);
  and _21530_ (_11055_, _13186_, _04856_);
  and _21531_ (_13187_, _12371_, _05730_);
  nand _21532_ (_13189_, _13187_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor _21533_ (_13190_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , rst);
  or _21534_ (_13191_, _13187_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _21535_ (_13192_, _13191_, _13190_);
  and _21536_ (_11058_, _13192_, _13189_);
  or _21537_ (_13193_, _12375_, _12373_);
  and _21538_ (_13194_, _13193_, _12376_);
  or _21539_ (_13195_, _13194_, _08257_);
  or _21540_ (_13197_, _05730_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and _21541_ (_13198_, _13197_, _13190_);
  and _21542_ (_11089_, _13198_, _13195_);
  nor _21543_ (_11150_, _07089_, rst);
  nor _21544_ (_11174_, _07032_, rst);
  nand _21545_ (_13199_, _12171_, _06586_);
  or _21546_ (_13200_, _12171_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3]);
  and _21547_ (_13201_, _13200_, _04856_);
  and _21548_ (_11236_, _13201_, _13199_);
  nand _21549_ (_13202_, _12171_, _07702_);
  or _21550_ (_13204_, _12171_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  and _21551_ (_13206_, _13204_, _04856_);
  and _21552_ (_11247_, _13206_, _13202_);
  and _21553_ (_13207_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _04856_);
  and _21554_ (_13208_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _04856_);
  and _21555_ (_13209_, _13208_, _12206_);
  or _21556_ (_11312_, _13209_, _13207_);
  and _21557_ (_13210_, _12205_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  or _21558_ (_13211_, _13210_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  and _21559_ (_11327_, _13211_, _04856_);
  and _21560_ (_13212_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  and _21561_ (_13214_, _12165_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  or _21562_ (_13215_, _13214_, _13212_);
  and _21563_ (_11343_, _13215_, _04856_);
  or _21564_ (_13216_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  nand _21565_ (_13217_, _08367_, _05774_);
  and _21566_ (_13218_, _13217_, _04856_);
  and _21567_ (_11347_, _13218_, _13216_);
  and _21568_ (_13219_, _08277_, _05520_);
  nand _21569_ (_13220_, _13219_, _06088_);
  or _21570_ (_13221_, _13219_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and _21571_ (_13222_, _13221_, _06935_);
  and _21572_ (_13223_, _13222_, _13220_);
  or _21573_ (_13224_, _13223_, _06946_);
  and _21574_ (_11350_, _13224_, _04856_);
  or _21575_ (_13225_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  nand _21576_ (_13226_, _08367_, _05911_);
  and _21577_ (_13227_, _13226_, _04856_);
  and _21578_ (_11355_, _13227_, _13225_);
  or _21579_ (_13228_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  nand _21580_ (_13229_, _08367_, _05811_);
  and _21581_ (_13230_, _13229_, _04856_);
  and _21582_ (_11357_, _13230_, _13228_);
  or _21583_ (_13231_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  nand _21584_ (_13232_, _08367_, _05735_);
  and _21585_ (_13233_, _13232_, _04856_);
  and _21586_ (_11370_, _13233_, _13231_);
  and _21587_ (_13234_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  and _21588_ (_13235_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and _21589_ (_13236_, _13235_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor _21590_ (_13237_, _13235_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor _21591_ (_00001_, _13237_, _13236_);
  or _21592_ (_00002_, _00001_, _13234_);
  and _21593_ (_11406_, _00002_, _04856_);
  and _21594_ (_00003_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], _08359_);
  and _21595_ (_00004_, \oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or _21596_ (_00005_, _00004_, _00003_);
  and _21597_ (_11412_, _00005_, _04856_);
  nor _21598_ (_11426_, _12903_, rst);
  nor _21599_ (_11428_, _12972_, rst);
  and _21600_ (_00006_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6], \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  and _21601_ (_00007_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and _21602_ (_00008_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and _21603_ (_00009_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor _21604_ (_00010_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  nor _21605_ (_00011_, _00010_, _00008_);
  and _21606_ (_00012_, _00011_, _00009_);
  nor _21607_ (_00013_, _00012_, _00008_);
  not _21608_ (_00014_, _00013_);
  nor _21609_ (_00015_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor _21610_ (_00016_, _00015_, _00007_);
  and _21611_ (_00017_, _00016_, _00014_);
  nor _21612_ (_00018_, _00017_, _00007_);
  nor _21613_ (_00019_, _00018_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and _21614_ (_00020_, _00018_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor _21615_ (_00021_, _00020_, _00019_);
  not _21616_ (_00022_, _12361_);
  nor _21617_ (_00023_, _00011_, _00009_);
  nor _21618_ (_00024_, _00023_, _00012_);
  nand _21619_ (_00025_, _00024_, _00022_);
  nor _21620_ (_00026_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor _21621_ (_00027_, _00026_, _00009_);
  and _21622_ (_00028_, _00027_, _12371_);
  or _21623_ (_00029_, _00024_, _00022_);
  and _21624_ (_00030_, _00029_, _00025_);
  nand _21625_ (_00031_, _00030_, _00028_);
  nand _21626_ (_00032_, _00031_, _00025_);
  nor _21627_ (_00033_, _00016_, _00014_);
  nor _21628_ (_00034_, _00033_, _00017_);
  and _21629_ (_00035_, _00034_, _00032_);
  and _21630_ (_00036_, _00035_, _00021_);
  nor _21631_ (_00037_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3], \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or _21632_ (_00038_, _00037_, _13051_);
  nand _21633_ (_00039_, _00038_, _00019_);
  or _21634_ (_00040_, _00038_, _00019_);
  and _21635_ (_00042_, _00040_, _00039_);
  not _21636_ (_00043_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and _21637_ (_00044_, _00037_, _00043_);
  and _21638_ (_00045_, _00018_, _00044_);
  nand _21639_ (_00046_, _00018_, _00037_);
  and _21640_ (_00047_, _00046_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  or _21641_ (_00048_, _00047_, _00045_);
  and _21642_ (_00049_, _00048_, _00042_);
  and _21643_ (_00050_, _00049_, _00036_);
  not _21644_ (_00051_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor _21645_ (_00052_, _00045_, _00051_);
  and _21646_ (_00053_, _00045_, _00051_);
  or _21647_ (_00054_, _00053_, _00052_);
  and _21648_ (_00055_, _00054_, _00050_);
  nor _21649_ (_00056_, _00054_, _00050_);
  nor _21650_ (_00057_, _00056_, _00055_);
  or _21651_ (_00058_, _00057_, _06911_);
  not _21652_ (_00059_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _21653_ (_00060_, _06910_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and _21654_ (_00061_, _00060_, _00059_);
  and _21655_ (_00062_, _00061_, _00058_);
  or _21656_ (_00063_, _00062_, _00006_);
  and _21657_ (_11435_, _00063_, _04856_);
  and _21658_ (_00064_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor _21659_ (_00065_, _08367_, _05803_);
  or _21660_ (_00066_, _00065_, _00064_);
  and _21661_ (_11439_, _00066_, _04856_);
  and _21662_ (_00067_, _00042_, _00036_);
  or _21663_ (_00068_, _00048_, _00067_);
  nor _21664_ (_00069_, _00050_, _06911_);
  and _21665_ (_00070_, _00069_, _00068_);
  nor _21666_ (_00071_, _06910_, _05183_);
  or _21667_ (_00072_, _00071_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _21668_ (_00073_, _00072_, _00070_);
  or _21669_ (_00074_, _00059_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and _21670_ (_00075_, _00074_, _04856_);
  and _21671_ (_11443_, _00075_, _00073_);
  and _21672_ (_00076_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor _21673_ (_00077_, _08367_, _05754_);
  or _21674_ (_00078_, _00077_, _00076_);
  and _21675_ (_11451_, _00078_, _04856_);
  and _21676_ (_00079_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  nor _21677_ (_00080_, _08367_, _05850_);
  or _21678_ (_00081_, _00080_, _00079_);
  and _21679_ (_11464_, _00081_, _04856_);
  nor _21680_ (_00082_, _00042_, _00036_);
  nor _21681_ (_00083_, _00082_, _00067_);
  or _21682_ (_00084_, _00083_, _06911_);
  or _21683_ (_00085_, _06910_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _21684_ (_00086_, _00085_, _00059_);
  and _21685_ (_00087_, _00086_, _00084_);
  and _21686_ (_00088_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4], \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _21687_ (_00089_, _00088_, _00087_);
  and _21688_ (_11467_, _00089_, _04856_);
  and _21689_ (_00090_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  nor _21690_ (_00091_, _08367_, _05824_);
  or _21691_ (_00092_, _00091_, _00090_);
  and _21692_ (_11476_, _00092_, _04856_);
  and _21693_ (_00093_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3], \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  nor _21694_ (_00094_, _00035_, _00021_);
  nor _21695_ (_00095_, _00094_, _00036_);
  or _21696_ (_00096_, _00095_, _06911_);
  or _21697_ (_00097_, _06910_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and _21698_ (_00098_, _00097_, _00059_);
  and _21699_ (_00099_, _00098_, _00096_);
  or _21700_ (_00100_, _00099_, _00093_);
  and _21701_ (_11522_, _00100_, _04856_);
  and _21702_ (_00101_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  nor _21703_ (_00102_, _00034_, _00032_);
  nor _21704_ (_00103_, _00102_, _00035_);
  or _21705_ (_00104_, _00103_, _06911_);
  or _21706_ (_00105_, _06910_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and _21707_ (_00106_, _00105_, _00059_);
  and _21708_ (_00107_, _00106_, _00104_);
  or _21709_ (_00108_, _00107_, _00101_);
  and _21710_ (_11543_, _00108_, _04856_);
  or _21711_ (_00109_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  nand _21712_ (_00110_, _08367_, _05855_);
  and _21713_ (_00111_, _00110_, _04856_);
  and _21714_ (_11565_, _00111_, _00109_);
  and _21715_ (_00112_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], _08359_);
  and _21716_ (_00113_, \oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or _21717_ (_00114_, _00113_, _00112_);
  and _21718_ (_11579_, _00114_, _04856_);
  nor _21719_ (_11595_, _12878_, rst);
  and _21720_ (_00117_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  nor _21721_ (_00118_, _08367_, _05861_);
  or _21722_ (_00119_, _00118_, _00117_);
  and _21723_ (_11598_, _00119_, _04856_);
  and _21724_ (_00120_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  nor _21725_ (_00122_, _08367_, _05881_);
  or _21726_ (_00123_, _00122_, _00120_);
  and _21727_ (_11602_, _00123_, _04856_);
  and _21728_ (_00125_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13], \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  not _21729_ (_00127_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  not _21730_ (_00128_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  not _21731_ (_00129_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  not _21732_ (_00131_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor _21733_ (_00132_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8], \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  not _21734_ (_00134_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and _21735_ (_00135_, _00044_, _00051_);
  and _21736_ (_00136_, _00135_, _00134_);
  and _21737_ (_00138_, _00136_, _00132_);
  and _21738_ (_00139_, _00138_, _00131_);
  and _21739_ (_00141_, _00139_, _00018_);
  and _21740_ (_00142_, _00141_, _00129_);
  and _21741_ (_00143_, _00142_, _00128_);
  nor _21742_ (_00145_, _00143_, _00127_);
  and _21743_ (_00146_, _00143_, _00127_);
  nor _21744_ (_00147_, _00146_, _00145_);
  not _21745_ (_00148_, _00147_);
  nor _21746_ (_00149_, _00142_, _00128_);
  nor _21747_ (_00151_, _00149_, _00143_);
  not _21748_ (_00152_, _00151_);
  nor _21749_ (_00153_, _00141_, _00129_);
  nor _21750_ (_00154_, _00153_, _00142_);
  not _21751_ (_00155_, _00154_);
  and _21752_ (_00156_, _00138_, _00018_);
  nor _21753_ (_00158_, _00156_, _00131_);
  nor _21754_ (_00159_, _00158_, _00141_);
  not _21755_ (_00160_, _00159_);
  not _21756_ (_00161_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  not _21757_ (_00162_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and _21758_ (_00163_, _00136_, _00018_);
  and _21759_ (_00164_, _00163_, _00162_);
  nor _21760_ (_00166_, _00164_, _00161_);
  or _21761_ (_00167_, _00166_, _00156_);
  nor _21762_ (_00169_, _00163_, _00162_);
  nor _21763_ (_00171_, _00169_, _00164_);
  nor _21764_ (_00172_, _00053_, _00134_);
  nor _21765_ (_00173_, _00172_, _00163_);
  not _21766_ (_00174_, _00173_);
  and _21767_ (_00175_, _00174_, _00055_);
  not _21768_ (_00176_, _00175_);
  nor _21769_ (_00178_, _00176_, _00171_);
  and _21770_ (_00179_, _00178_, _00167_);
  and _21771_ (_00180_, _00179_, _00160_);
  and _21772_ (_00181_, _00180_, _00155_);
  and _21773_ (_00182_, _00181_, _00152_);
  and _21774_ (_00183_, _00182_, _00148_);
  nor _21775_ (_00184_, _00182_, _00148_);
  nor _21776_ (_00185_, _00184_, _00183_);
  or _21777_ (_00186_, _00185_, _06911_);
  or _21778_ (_00187_, _06910_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and _21779_ (_00188_, _00187_, _00059_);
  and _21780_ (_00189_, _00188_, _00186_);
  or _21781_ (_00190_, _00189_, _00125_);
  and _21782_ (_11605_, _00190_, _04856_);
  and _21783_ (_00191_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12], \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  nor _21784_ (_00192_, _00181_, _00152_);
  nor _21785_ (_00193_, _00192_, _00182_);
  or _21786_ (_00194_, _00193_, _06911_);
  or _21787_ (_00195_, _06910_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _21788_ (_00197_, _00195_, _00059_);
  and _21789_ (_00198_, _00197_, _00194_);
  or _21790_ (_00199_, _00198_, _00191_);
  and _21791_ (_11610_, _00199_, _04856_);
  nor _21792_ (_00200_, _00180_, _00155_);
  nor _21793_ (_00201_, _00200_, _00181_);
  or _21794_ (_00202_, _00201_, _06911_);
  or _21795_ (_00203_, _06910_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _21796_ (_00204_, _00203_, _00059_);
  and _21797_ (_00206_, _00204_, _00202_);
  and _21798_ (_00207_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11], \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _21799_ (_00208_, _00207_, _00206_);
  and _21800_ (_11616_, _00208_, _04856_);
  nor _21801_ (_00210_, _00179_, _00160_);
  nor _21802_ (_00211_, _00210_, _00180_);
  or _21803_ (_00212_, _00211_, _06911_);
  or _21804_ (_00213_, _06910_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and _21805_ (_00214_, _00213_, _00059_);
  and _21806_ (_00215_, _00214_, _00212_);
  and _21807_ (_00216_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10], \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _21808_ (_00217_, _00216_, _00215_);
  and _21809_ (_11618_, _00217_, _04856_);
  or _21810_ (_00218_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  nand _21811_ (_00219_, _08367_, _05808_);
  and _21812_ (_00220_, _00219_, _04856_);
  and _21813_ (_11620_, _00220_, _00218_);
  nor _21814_ (_00221_, _00178_, _00167_);
  nor _21815_ (_00222_, _00221_, _00179_);
  or _21816_ (_00223_, _00222_, _06911_);
  or _21817_ (_00224_, _06910_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and _21818_ (_00225_, _00224_, _00059_);
  and _21819_ (_00226_, _00225_, _00223_);
  and _21820_ (_00227_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  or _21821_ (_00228_, _00227_, _00226_);
  and _21822_ (_11624_, _00228_, _04856_);
  and _21823_ (_00229_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], _08359_);
  and _21824_ (_00230_, \oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or _21825_ (_00231_, _00230_, _00229_);
  and _21826_ (_11630_, _00231_, _04856_);
  nor _21827_ (_11638_, _12854_, rst);
  and _21828_ (_00232_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor _21829_ (_00233_, _08367_, _05884_);
  or _21830_ (_00234_, _00233_, _00232_);
  and _21831_ (_11641_, _00234_, _04856_);
  and _21832_ (_00235_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8], \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  and _21833_ (_00236_, _00176_, _00171_);
  nor _21834_ (_00237_, _00236_, _00178_);
  or _21835_ (_00238_, _00237_, _06911_);
  or _21836_ (_00239_, _06910_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and _21837_ (_00240_, _00239_, _00059_);
  and _21838_ (_00241_, _00240_, _00238_);
  or _21839_ (_00242_, _00241_, _00235_);
  and _21840_ (_11646_, _00242_, _04856_);
  and _21841_ (_00243_, \oc8051_top_1.oc8051_memory_interface1.cdata [5], _08359_);
  and _21842_ (_00244_, \oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or _21843_ (_00245_, _00244_, _00243_);
  and _21844_ (_11658_, _00245_, _04856_);
  not _21845_ (_00246_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  or _21846_ (_00247_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _00246_);
  or _21847_ (_00248_, _00247_, _08060_);
  nor _21848_ (_00249_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  and _21849_ (_00250_, _00249_, _00248_);
  or _21850_ (_00251_, _00250_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or _21851_ (_00252_, _00251_, _09259_);
  not _21852_ (_00253_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or _21853_ (_00254_, _04990_, _00253_);
  nand _21854_ (_00255_, _00254_, _09259_);
  or _21855_ (_00256_, _00255_, _07708_);
  and _21856_ (_00257_, _00256_, _00252_);
  or _21857_ (_00258_, _00257_, _09263_);
  nand _21858_ (_00259_, _09263_, _06369_);
  and _21859_ (_00260_, _00259_, _04856_);
  and _21860_ (_11698_, _00260_, _00258_);
  and _21861_ (_00261_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  nor _21862_ (_00262_, _08367_, _05749_);
  or _21863_ (_00263_, _00262_, _00261_);
  and _21864_ (_11704_, _00263_, _04856_);
  and _21865_ (_00264_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  nor _21866_ (_00265_, _08367_, _05805_);
  or _21867_ (_00266_, _00265_, _00264_);
  and _21868_ (_11710_, _00266_, _04856_);
  and _21869_ (_00267_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  nor _21870_ (_00268_, _08367_, _05782_);
  or _21871_ (_00269_, _00268_, _00267_);
  and _21872_ (_11715_, _00269_, _04856_);
  and _21873_ (_00270_, _08277_, _07855_);
  nand _21874_ (_00271_, _00270_, _06088_);
  or _21875_ (_00272_, _00270_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and _21876_ (_00273_, _00272_, _06935_);
  and _21877_ (_00274_, _00273_, _00271_);
  or _21878_ (_00275_, _00274_, _06937_);
  and _21879_ (_11718_, _00275_, _04856_);
  and _21880_ (_00276_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  nor _21881_ (_00277_, _08367_, _05909_);
  or _21882_ (_00278_, _00277_, _00276_);
  and _21883_ (_11720_, _00278_, _04856_);
  and _21884_ (_00279_, _06163_, _05510_);
  or _21885_ (_00280_, _00279_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and _21886_ (_00281_, _00280_, _04856_);
  nand _21887_ (_00282_, _00279_, _05287_);
  and _21888_ (_11723_, _00282_, _00281_);
  and _21889_ (_00283_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  and _21890_ (_00284_, _12165_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  or _21891_ (_00285_, _00284_, _00283_);
  and _21892_ (_11726_, _00285_, _04856_);
  or _21893_ (_00286_, _00279_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and _21894_ (_00287_, _00286_, _04856_);
  not _21895_ (_00288_, _00279_);
  or _21896_ (_00289_, _00288_, _05718_);
  and _21897_ (_11729_, _00289_, _00287_);
  and _21898_ (_00290_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  nor _21899_ (_00291_, _08367_, _05778_);
  or _21900_ (_00292_, _00291_, _00290_);
  and _21901_ (_11736_, _00292_, _04856_);
  and _21902_ (_00293_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor _21903_ (_00294_, _08367_, _05834_);
  or _21904_ (_00295_, _00294_, _00293_);
  and _21905_ (_11751_, _00295_, _04856_);
  nor _21906_ (_11754_, _07294_, rst);
  nor _21907_ (_11792_, _12926_, rst);
  nor _21908_ (_11801_, _12949_, rst);
  and _21909_ (_00296_, _06721_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  or _21910_ (_00297_, _06834_, _06733_);
  or _21911_ (_00298_, _12682_, _12695_);
  or _21912_ (_00299_, _00298_, _06866_);
  or _21913_ (_00300_, _00299_, _00297_);
  and _21914_ (_00301_, _06598_, _05950_);
  or _21915_ (_00302_, _09088_, _00301_);
  or _21916_ (_00303_, _00302_, _05988_);
  or _21917_ (_00304_, _06763_, _06799_);
  or _21918_ (_00305_, _00304_, _09097_);
  or _21919_ (_00306_, _00305_, _06756_);
  or _21920_ (_00308_, _06786_, _06760_);
  or _21921_ (_00309_, _00308_, _00306_);
  or _21922_ (_00310_, _00309_, _00303_);
  or _21923_ (_00311_, _09081_, _06740_);
  or _21924_ (_00312_, _00311_, _00310_);
  or _21925_ (_00313_, _00312_, _00300_);
  or _21926_ (_00314_, _05999_, _05962_);
  nor _21927_ (_00315_, rst, \oc8051_top_1.oc8051_sfr1.wait_data );
  and _21928_ (_00316_, _00315_, _00314_);
  and _21929_ (_00317_, _00316_, _00313_);
  or _21930_ (_11805_, _00317_, _00296_);
  or _21931_ (_00318_, _00279_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and _21932_ (_00319_, _00318_, _04856_);
  or _21933_ (_00320_, _00288_, _06410_);
  and _21934_ (_11825_, _00320_, _00319_);
  or _21935_ (_00321_, _00279_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  and _21936_ (_00322_, _00321_, _04856_);
  nand _21937_ (_00323_, _00279_, _05669_);
  and _21938_ (_11830_, _00323_, _00322_);
  and _21939_ (_00324_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], _08359_);
  and _21940_ (_00325_, \oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or _21941_ (_00326_, _00325_, _00324_);
  and _21942_ (_11848_, _00326_, _04856_);
  and _21943_ (_00327_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], _08359_);
  and _21944_ (_00328_, \oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or _21945_ (_00329_, _00328_, _00327_);
  and _21946_ (_11856_, _00329_, _04856_);
  and _21947_ (_00330_, _12429_, _05517_);
  and _21948_ (_00331_, _00330_, _05288_);
  and _21949_ (_00332_, _12718_, _05517_);
  and _21950_ (_00333_, _00332_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  not _21951_ (_00334_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _21952_ (_00335_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _00334_);
  and _21953_ (_00336_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _21954_ (_00337_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and _21955_ (_00338_, _00337_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _21956_ (_00339_, _00338_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and _21957_ (_00340_, _00339_, _00336_);
  and _21958_ (_00341_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and _21959_ (_00342_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  and _21960_ (_00343_, _00342_, _00341_);
  and _21961_ (_00344_, _00343_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  not _21962_ (_00345_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and _21963_ (_00346_, \oc8051_top_1.oc8051_sfr1.pres_ow , _00345_);
  not _21964_ (_00347_, t0_i);
  and _21965_ (_00348_, _00347_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and _21966_ (_00349_, _00348_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff );
  or _21967_ (_00350_, _00349_, _00346_);
  and _21968_ (_00351_, _00350_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and _21969_ (_00352_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and _21970_ (_00353_, _00352_, _00351_);
  and _21971_ (_00354_, _00353_, _00344_);
  and _21972_ (_00355_, _00354_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and _21973_ (_00356_, _00355_, _00340_);
  nor _21974_ (_00357_, _00356_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and _21975_ (_00358_, _00356_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nor _21976_ (_00359_, _00358_, _00357_);
  and _21977_ (_00360_, _00359_, _00335_);
  nor _21978_ (_00361_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _21979_ (_00362_, _00343_, _00351_);
  and _21980_ (_00363_, _00362_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and _21981_ (_00364_, _00363_, _00340_);
  nand _21982_ (_00365_, _00364_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or _21983_ (_00366_, _00364_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and _21984_ (_00367_, _00366_, _00365_);
  and _21985_ (_00368_, _00367_, _00361_);
  and _21986_ (_00369_, \oc8051_top_1.oc8051_sfr1.pres_ow , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and _21987_ (_00370_, _00369_, _00339_);
  and _21988_ (_00371_, _00370_, _00336_);
  and _21989_ (_00372_, _00371_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  nand _21990_ (_00373_, _00372_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or _21991_ (_00374_, _00372_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and _21992_ (_00375_, _00374_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _21993_ (_00376_, _00375_, _00373_);
  or _21994_ (_00377_, _00376_, _00368_);
  or _21995_ (_00378_, _00377_, _00360_);
  nor _21996_ (_00379_, _00332_, _00330_);
  and _21997_ (_00380_, _00379_, _00378_);
  or _21998_ (_00381_, _00380_, _00333_);
  or _21999_ (_00382_, _00381_, _00331_);
  and _22000_ (_11877_, _00382_, _04856_);
  and _22001_ (_00383_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], _08359_);
  and _22002_ (_00384_, \oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or _22003_ (_00385_, _00384_, _00383_);
  and _22004_ (_11883_, _00385_, _04856_);
  and _22005_ (_00386_, _00330_, _06410_);
  and _22006_ (_00387_, _00332_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _22007_ (_00388_, _00355_, _00339_);
  or _22008_ (_00389_, _00388_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _22009_ (_00390_, _00388_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  not _22010_ (_00391_, _00390_);
  and _22011_ (_00392_, _00391_, _00335_);
  and _22012_ (_00393_, _00392_, _00389_);
  and _22013_ (_00394_, _00339_, _00344_);
  and _22014_ (_00395_, _00394_, _00351_);
  nor _22015_ (_00396_, _00395_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _22016_ (_00397_, _00395_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nor _22017_ (_00398_, _00397_, _00396_);
  and _22018_ (_00399_, _00398_, _00361_);
  not _22019_ (_00400_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _22020_ (_00401_, _00370_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  nor _22021_ (_00402_, _00401_, _00400_);
  and _22022_ (_00403_, _00401_, _00400_);
  or _22023_ (_00404_, _00403_, _00402_);
  and _22024_ (_00405_, _00404_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  or _22025_ (_00406_, _00405_, _00399_);
  or _22026_ (_00407_, _00406_, _00393_);
  and _22027_ (_00408_, _00407_, _00379_);
  or _22028_ (_00409_, _00408_, _00387_);
  or _22029_ (_00410_, _00409_, _00386_);
  and _22030_ (_11888_, _00410_, _04856_);
  and _22031_ (_00411_, _00330_, _05718_);
  and _22032_ (_00412_, _00332_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _22033_ (_00413_, _07460_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  or _22034_ (_00414_, _00413_, _00335_);
  and _22035_ (_00415_, _00390_, _00334_);
  or _22036_ (_00416_, _00415_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nand _22037_ (_00417_, _00415_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _22038_ (_00418_, _00417_, _00416_);
  and _22039_ (_00419_, _00418_, _00414_);
  and _22040_ (_00420_, _00370_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or _22041_ (_00421_, _00420_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  not _22042_ (_00422_, _00371_);
  and _22043_ (_00423_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _22044_ (_00424_, _00423_, _00422_);
  and _22045_ (_00425_, _00424_, _00421_);
  nand _22046_ (_00426_, _00397_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  or _22047_ (_00427_, _00397_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _22048_ (_00428_, _00427_, _00426_);
  and _22049_ (_00429_, _00428_, _00361_);
  or _22050_ (_00430_, _00429_, _00425_);
  or _22051_ (_00431_, _00430_, _00419_);
  and _22052_ (_00432_, _00431_, _00379_);
  or _22053_ (_00433_, _00432_, _00412_);
  or _22054_ (_00434_, _00433_, _00411_);
  and _22055_ (_11891_, _00434_, _04856_);
  and _22056_ (_00435_, _00330_, _06705_);
  and _22057_ (_00436_, _00332_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _22058_ (_00437_, _00355_, _00338_);
  and _22059_ (_00438_, _00352_, _00344_);
  and _22060_ (_00439_, _00438_, _00351_);
  and _22061_ (_00440_, _00439_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and _22062_ (_00441_, _00440_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and _22063_ (_00442_, _00441_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  or _22064_ (_00443_, _00442_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nand _22065_ (_00444_, _00443_, _00335_);
  nor _22066_ (_00445_, _00444_, _00437_);
  and _22067_ (_00446_, _00363_, _00337_);
  or _22068_ (_00447_, _00446_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  not _22069_ (_00448_, _00361_);
  and _22070_ (_00449_, _00363_, _00338_);
  nor _22071_ (_00450_, _00449_, _00448_);
  and _22072_ (_00451_, _00450_, _00447_);
  and _22073_ (_00452_, _00369_, _00337_);
  and _22074_ (_00453_, _00452_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or _22075_ (_00454_, _00453_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nand _22076_ (_00455_, _00453_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _22077_ (_00456_, _00455_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _22078_ (_00457_, _00456_, _00454_);
  or _22079_ (_00458_, _00457_, _00451_);
  or _22080_ (_00459_, _00458_, _00445_);
  and _22081_ (_00460_, _00459_, _00379_);
  or _22082_ (_00461_, _00460_, _00436_);
  or _22083_ (_00462_, _00461_, _00435_);
  and _22084_ (_11897_, _00462_, _04856_);
  and _22085_ (_00463_, _00330_, _05670_);
  and _22086_ (_00464_, _00332_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and _22087_ (_00465_, _00437_, _00334_);
  or _22088_ (_00466_, _00465_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  not _22089_ (_00467_, _00388_);
  or _22090_ (_00468_, _00467_, _00413_);
  and _22091_ (_00469_, _00468_, _00414_);
  and _22092_ (_00470_, _00469_, _00466_);
  and _22093_ (_00471_, _00369_, _00338_);
  or _22094_ (_00472_, _00471_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  not _22095_ (_00473_, _00370_);
  and _22096_ (_00474_, _00423_, _00473_);
  and _22097_ (_00475_, _00474_, _00472_);
  not _22098_ (_00476_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  nor _22099_ (_00477_, _00449_, _00476_);
  and _22100_ (_00478_, _00449_, _00476_);
  or _22101_ (_00479_, _00478_, _00477_);
  and _22102_ (_00480_, _00479_, _00361_);
  or _22103_ (_00481_, _00480_, _00475_);
  or _22104_ (_00482_, _00481_, _00470_);
  and _22105_ (_00483_, _00482_, _00379_);
  or _22106_ (_00484_, _00483_, _00464_);
  or _22107_ (_00485_, _00484_, _00463_);
  and _22108_ (_11900_, _00485_, _04856_);
  not _22109_ (_00486_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  nor _22110_ (_00487_, _13234_, _00486_);
  nor _22111_ (_00488_, _00487_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and _22112_ (_00489_, _00487_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  or _22113_ (_00490_, _00489_, _00488_);
  nor _22114_ (_11904_, _00490_, rst);
  not _22115_ (_00491_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nand _22116_ (_00492_, _00355_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or _22117_ (_00493_, _00492_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  nand _22118_ (_00494_, _00493_, _00491_);
  not _22119_ (_00495_, _00442_);
  or _22120_ (_00496_, _00413_, _00495_);
  and _22121_ (_00497_, _00496_, _00414_);
  and _22122_ (_00499_, _00497_, _00494_);
  and _22123_ (_00500_, _00369_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or _22124_ (_00501_, _00500_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  not _22125_ (_00502_, _00452_);
  and _22126_ (_00503_, _00423_, _00502_);
  and _22127_ (_00504_, _00503_, _00501_);
  and _22128_ (_00505_, _00363_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or _22129_ (_00506_, _00505_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nor _22130_ (_00507_, _00446_, _00448_);
  and _22131_ (_00508_, _00507_, _00506_);
  or _22132_ (_00509_, _00508_, _00504_);
  or _22133_ (_00510_, _00509_, _00499_);
  and _22134_ (_00511_, _00510_, _00379_);
  and _22135_ (_00512_, _00332_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and _22136_ (_00513_, _00330_, _06033_);
  or _22137_ (_00514_, _00513_, _00512_);
  or _22138_ (_00515_, _00514_, _00511_);
  and _22139_ (_11907_, _00515_, _04856_);
  not _22140_ (_00516_, _00332_);
  or _22141_ (_00517_, _00516_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and _22142_ (_00518_, _00517_, _04856_);
  nand _22143_ (_00519_, _00330_, _06369_);
  and _22144_ (_00520_, _00440_, _00334_);
  or _22145_ (_00521_, _00520_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and _22146_ (_00522_, _00521_, _00493_);
  and _22147_ (_00523_, _00522_, _00414_);
  or _22148_ (_00524_, _00369_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand _22149_ (_00525_, _00524_, _00423_);
  nor _22150_ (_00526_, _00525_, _00500_);
  nor _22151_ (_00527_, _00363_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nor _22152_ (_00528_, _00527_, _00505_);
  and _22153_ (_00529_, _00528_, _00361_);
  or _22154_ (_00530_, _00529_, _00526_);
  or _22155_ (_00531_, _00530_, _00523_);
  or _22156_ (_00532_, _00531_, _00330_);
  and _22157_ (_00533_, _00532_, _00519_);
  or _22158_ (_00534_, _00533_, _00332_);
  and _22159_ (_11910_, _00534_, _00518_);
  and _22160_ (_00535_, _13234_, _00486_);
  nor _22161_ (_00536_, _00535_, _00487_);
  and _22162_ (_11914_, _00536_, _04856_);
  nand _22163_ (_00537_, _00279_, _06032_);
  or _22164_ (_00538_, _00279_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _22165_ (_00539_, _00538_, _04856_);
  and _22166_ (_11924_, _00539_, _00537_);
  or _22167_ (_00540_, _00288_, _06705_);
  or _22168_ (_00541_, _00279_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and _22169_ (_00542_, _00541_, _04856_);
  and _22170_ (_11927_, _00542_, _00540_);
  nor _22171_ (_00543_, _00279_, _07460_);
  and _22172_ (_00544_, _00279_, _06997_);
  or _22173_ (_00545_, _00544_, _00543_);
  and _22174_ (_11930_, _00545_, _04856_);
  and _22175_ (_00546_, _06721_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  and _22176_ (_00547_, _06612_, _05848_);
  or _22177_ (_00548_, _00547_, _09068_);
  or _22178_ (_00549_, _00548_, _09067_);
  or _22179_ (_00550_, _05999_, _05988_);
  or _22180_ (_00551_, _12689_, _06762_);
  or _22181_ (_00552_, _00551_, _00550_);
  or _22182_ (_00553_, _00552_, _06839_);
  or _22183_ (_00554_, _00553_, _00549_);
  not _22184_ (_00555_, _07509_);
  or _22185_ (_00556_, _08051_, _00555_);
  or _22186_ (_00557_, _12698_, _06760_);
  and _22187_ (_00558_, _06822_, _06598_);
  and _22188_ (_00559_, _06638_, _06635_);
  or _22189_ (_00560_, _00559_, _00558_);
  or _22190_ (_00561_, _00560_, _00557_);
  or _22191_ (_00562_, _00561_, _06727_);
  or _22192_ (_00563_, _00562_, _00556_);
  or _22193_ (_00564_, _00563_, _00554_);
  and _22194_ (_00565_, _00564_, _00316_);
  or _22195_ (_11945_, _00565_, _00546_);
  and _22196_ (_00566_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  nor _22197_ (_00567_, _08367_, _05904_);
  or _22198_ (_00568_, _00567_, _00566_);
  and _22199_ (_11979_, _00568_, _04856_);
  and _22200_ (_00569_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  and _22201_ (_00570_, _12165_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  or _22202_ (_00571_, _00570_, _00569_);
  and _22203_ (_11984_, _00571_, _04856_);
  or _22204_ (_00572_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  nand _22205_ (_00573_, _08367_, _05784_);
  and _22206_ (_00575_, _00573_, _04856_);
  and _22207_ (_11993_, _00575_, _00572_);
  or _22208_ (_00576_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  nand _22209_ (_00577_, _08367_, _05829_);
  and _22210_ (_00578_, _00577_, _04856_);
  and _22211_ (_11995_, _00578_, _00576_);
  and _22212_ (_00579_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  and _22213_ (_00580_, _12165_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  or _22214_ (_00581_, _00580_, _00579_);
  and _22215_ (_12001_, _00581_, _04856_);
  or _22216_ (_00582_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  nand _22217_ (_00583_, _08367_, _05875_);
  and _22218_ (_00584_, _00583_, _04856_);
  and _22219_ (_12006_, _00584_, _00582_);
  or _22220_ (_00585_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  nand _22221_ (_00586_, _08367_, _05826_);
  and _22222_ (_00587_, _00586_, _04856_);
  and _22223_ (_12011_, _00587_, _00585_);
  not _22224_ (_00588_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  not _22225_ (_00589_, t1_i);
  and _22226_ (_00590_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff , _00589_);
  nor _22227_ (_00591_, _00590_, _00588_);
  not _22228_ (_00592_, _00591_);
  not _22229_ (_00593_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and _22230_ (_00594_, _00593_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  nor _22231_ (_00595_, \oc8051_top_1.oc8051_sfr1.pres_ow , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  not _22232_ (_00596_, _00595_);
  and _22233_ (_00597_, _00596_, _00594_);
  and _22234_ (_00598_, _00597_, _00592_);
  and _22235_ (_00599_, _00598_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nor _22236_ (_00600_, _00599_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  and _22237_ (_00601_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  and _22238_ (_00602_, _00601_, _00598_);
  or _22239_ (_00603_, _00602_, _00600_);
  and _22240_ (_00604_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and _22241_ (_00605_, _12388_, _05517_);
  nor _22242_ (_00606_, _00605_, _00604_);
  nand _22243_ (_00607_, _00606_, _00603_);
  or _22244_ (_00608_, _00606_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  and _22245_ (_00609_, _00608_, _00607_);
  and _22246_ (_00610_, _12713_, _05517_);
  not _22247_ (_00611_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and _22248_ (_00612_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], _00611_);
  and _22249_ (_00613_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  and _22250_ (_00614_, _00613_, _00601_);
  and _22251_ (_00615_, _00614_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and _22252_ (_00616_, _00615_, _00598_);
  and _22253_ (_00617_, _00616_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and _22254_ (_00618_, _00617_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and _22255_ (_00619_, _00618_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and _22256_ (_00620_, _00619_, _00612_);
  nand _22257_ (_00621_, _00620_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nor _22258_ (_00622_, _00621_, _00605_);
  or _22259_ (_00623_, _00622_, _00610_);
  or _22260_ (_00624_, _00623_, _00609_);
  nand _22261_ (_00625_, _00610_, _06032_);
  and _22262_ (_00626_, _00625_, _04856_);
  and _22263_ (_12014_, _00626_, _00624_);
  and _22264_ (_00627_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and _22265_ (_00628_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and _22266_ (_00629_, _00628_, _00627_);
  and _22267_ (_00630_, _00629_, _00615_);
  nand _22268_ (_00631_, _00630_, _00612_);
  or _22269_ (_00632_, _00631_, _00605_);
  nand _22270_ (_00633_, _00632_, _00606_);
  and _22271_ (_00634_, _00633_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nor _22272_ (_00635_, _00598_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nor _22273_ (_00636_, _00635_, _00599_);
  and _22274_ (_00637_, _00636_, _00606_);
  or _22275_ (_00638_, _00637_, _00610_);
  or _22276_ (_00639_, _00638_, _00634_);
  nand _22277_ (_00640_, _00610_, _06369_);
  and _22278_ (_00641_, _00640_, _04856_);
  and _22279_ (_12017_, _00641_, _00639_);
  not _22280_ (_00642_, _00606_);
  and _22281_ (_00643_, _00642_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  and _22282_ (_00644_, _00620_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nor _22283_ (_00645_, _00602_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  and _22284_ (_00646_, _00602_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  or _22285_ (_00647_, _00646_, _00645_);
  nor _22286_ (_00648_, _00647_, _00604_);
  nor _22287_ (_00649_, _00648_, _00644_);
  nor _22288_ (_00650_, _00649_, _00605_);
  or _22289_ (_00651_, _00650_, _00610_);
  or _22290_ (_00652_, _00651_, _00643_);
  not _22291_ (_00653_, _00610_);
  or _22292_ (_00654_, _00653_, _06705_);
  and _22293_ (_00655_, _00654_, _04856_);
  and _22294_ (_12032_, _00655_, _00652_);
  or _22295_ (_00656_, _00653_, _06410_);
  and _22296_ (_00657_, _00642_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and _22297_ (_00658_, _00620_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and _22298_ (_00659_, _00613_, _00602_);
  or _22299_ (_00660_, _00659_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  nor _22300_ (_00661_, _00616_, _00604_);
  and _22301_ (_00662_, _00661_, _00660_);
  nor _22302_ (_00663_, _00662_, _00658_);
  nor _22303_ (_00664_, _00663_, _00605_);
  or _22304_ (_00665_, _00664_, _00657_);
  or _22305_ (_00666_, _00665_, _00610_);
  and _22306_ (_00667_, _00666_, _04856_);
  and _22307_ (_12035_, _00667_, _00656_);
  nor _22308_ (_00668_, _00646_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nor _22309_ (_00669_, _00668_, _00659_);
  and _22310_ (_00671_, _00669_, _00606_);
  nor _22311_ (_00672_, _00606_, _08808_);
  or _22312_ (_00673_, _00672_, _00671_);
  nand _22313_ (_00674_, _00620_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nor _22314_ (_00675_, _00674_, _00605_);
  or _22315_ (_00676_, _00675_, _00610_);
  or _22316_ (_00677_, _00676_, _00673_);
  nand _22317_ (_00678_, _00610_, _05669_);
  and _22318_ (_00679_, _00678_, _04856_);
  and _22319_ (_12038_, _00679_, _00677_);
  or _22320_ (_00680_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  nand _22321_ (_00681_, _08367_, _05745_);
  and _22322_ (_00682_, _00681_, _04856_);
  and _22323_ (_12040_, _00682_, _00680_);
  or _22324_ (_00683_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  nand _22325_ (_00684_, _08367_, _05879_);
  and _22326_ (_00685_, _00684_, _04856_);
  and _22327_ (_12042_, _00685_, _00683_);
  or _22328_ (_00686_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  nand _22329_ (_00687_, _08367_, _05852_);
  and _22330_ (_00688_, _00687_, _04856_);
  and _22331_ (_12049_, _00688_, _00686_);
  nand _22332_ (_00689_, _00610_, _05287_);
  not _22333_ (_00690_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and _22334_ (_00691_, _00690_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  nor _22335_ (_00692_, _00691_, _00612_);
  nor _22336_ (_00693_, _00605_, _00692_);
  not _22337_ (_00694_, _00693_);
  and _22338_ (_00695_, _00694_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nand _22339_ (_00696_, _00620_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nor _22340_ (_00697_, _00696_, _00605_);
  nor _22341_ (_00698_, _00617_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nor _22342_ (_00699_, _00698_, _00618_);
  and _22343_ (_00700_, _00699_, _00693_);
  or _22344_ (_00701_, _00700_, _00697_);
  or _22345_ (_00702_, _00701_, _00695_);
  or _22346_ (_00703_, _00702_, _00610_);
  and _22347_ (_00704_, _00703_, _04856_);
  and _22348_ (_12077_, _00704_, _00689_);
  or _22349_ (_00705_, _00653_, _05718_);
  not _22350_ (_00706_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  nor _22351_ (_00707_, _00693_, _00706_);
  and _22352_ (_00708_, _00620_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  not _22353_ (_00709_, _00692_);
  or _22354_ (_00710_, _00616_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  nand _22355_ (_00711_, _00710_, _00709_);
  nor _22356_ (_00712_, _00711_, _00617_);
  nor _22357_ (_00713_, _00712_, _00708_);
  nor _22358_ (_00714_, _00713_, _00605_);
  or _22359_ (_00715_, _00714_, _00707_);
  or _22360_ (_00716_, _00715_, _00610_);
  and _22361_ (_00717_, _00716_, _04856_);
  and _22362_ (_12082_, _00717_, _00705_);
  and _22363_ (_00718_, _12206_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  or _22364_ (_00719_, _00718_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and _22365_ (_12093_, _00719_, _04856_);
  nand _22366_ (_00720_, _00605_, _05287_);
  and _22367_ (_00721_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and _22368_ (_00722_, _00721_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and _22369_ (_00723_, _00615_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and _22370_ (_00724_, _00723_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and _22371_ (_00725_, _00724_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and _22372_ (_00726_, _00725_, _00598_);
  and _22373_ (_00727_, _00726_, _00722_);
  or _22374_ (_00728_, _00727_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nor _22375_ (_00729_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  not _22376_ (_00730_, _00729_);
  and _22377_ (_00731_, _00727_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nor _22378_ (_00732_, _00731_, _00730_);
  and _22379_ (_00733_, _00732_, _00728_);
  and _22380_ (_00734_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and _22381_ (_00735_, _00598_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and _22382_ (_00736_, _00630_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and _22383_ (_00737_, _00736_, _00735_);
  and _22384_ (_00738_, _00737_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and _22385_ (_00739_, _00738_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and _22386_ (_00740_, _00739_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and _22387_ (_00741_, _00740_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  or _22388_ (_00742_, _00740_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nand _22389_ (_00743_, _00742_, _00691_);
  nor _22390_ (_00744_, _00743_, _00741_);
  or _22391_ (_00745_, _00744_, _00734_);
  or _22392_ (_00746_, _00745_, _00733_);
  or _22393_ (_00747_, _00746_, _00605_);
  and _22394_ (_00748_, _00747_, _00720_);
  or _22395_ (_00749_, _00748_, _00610_);
  or _22396_ (_00750_, _00653_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and _22397_ (_00751_, _00750_, _04856_);
  and _22398_ (_12119_, _00751_, _00749_);
  nand _22399_ (_00752_, _00723_, _00598_);
  nor _22400_ (_00753_, _00752_, _00730_);
  and _22401_ (_00754_, _00691_, _00598_);
  and _22402_ (_00755_, _00754_, _00630_);
  or _22403_ (_00756_, _00755_, _00753_);
  and _22404_ (_00757_, _00756_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  or _22405_ (_00758_, _00757_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nor _22406_ (_00759_, _00726_, _00730_);
  or _22407_ (_00760_, _00759_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  or _22408_ (_00761_, _00737_, _00611_);
  nand _22409_ (_00762_, _00761_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  or _22410_ (_00763_, _00762_, _00760_);
  and _22411_ (_00764_, _00763_, _00758_);
  or _22412_ (_00765_, _00764_, _00605_);
  not _22413_ (_00766_, _00605_);
  or _22414_ (_00767_, _00766_, _06705_);
  and _22415_ (_00768_, _00767_, _00765_);
  or _22416_ (_00769_, _00768_, _00610_);
  or _22417_ (_00770_, _00653_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and _22418_ (_00771_, _00770_, _04856_);
  and _22419_ (_12128_, _00771_, _00769_);
  nand _22420_ (_00772_, _00605_, _05669_);
  or _22421_ (_00773_, _00737_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  not _22422_ (_00774_, _00691_);
  nor _22423_ (_00775_, _00738_, _00774_);
  and _22424_ (_00776_, _00775_, _00773_);
  and _22425_ (_00777_, _00726_, _00729_);
  or _22426_ (_00778_, _00777_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or _22427_ (_00779_, _00760_, _08812_);
  and _22428_ (_00780_, _00779_, _00778_);
  or _22429_ (_00781_, _00780_, _00776_);
  or _22430_ (_00782_, _00781_, _00605_);
  and _22431_ (_00783_, _00782_, _00772_);
  or _22432_ (_00784_, _00783_, _00610_);
  nand _22433_ (_00785_, _00610_, _08812_);
  and _22434_ (_00786_, _00785_, _04856_);
  and _22435_ (_12130_, _00786_, _00784_);
  or _22436_ (_00787_, _00766_, _06410_);
  or _22437_ (_00788_, _00738_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nor _22438_ (_00789_, _00739_, _00774_);
  and _22439_ (_00790_, _00789_, _00788_);
  and _22440_ (_00791_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and _22441_ (_00792_, _00726_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or _22442_ (_00793_, _00792_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and _22443_ (_00794_, _00792_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nor _22444_ (_00795_, _00794_, _00730_);
  and _22445_ (_00796_, _00795_, _00793_);
  or _22446_ (_00797_, _00796_, _00791_);
  or _22447_ (_00798_, _00797_, _00790_);
  or _22448_ (_00799_, _00798_, _00605_);
  and _22449_ (_00800_, _00799_, _00787_);
  or _22450_ (_00801_, _00800_, _00610_);
  or _22451_ (_00802_, _00653_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and _22452_ (_00803_, _00802_, _04856_);
  and _22453_ (_12135_, _00803_, _00801_);
  or _22454_ (_00804_, _00766_, _05718_);
  not _22455_ (_00805_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  nor _22456_ (_00806_, _00739_, _00611_);
  not _22457_ (_00807_, _00806_);
  nor _22458_ (_00808_, _00795_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and _22459_ (_00809_, _00808_, _00807_);
  and _22460_ (_00810_, _00809_, _00805_);
  nor _22461_ (_00811_, _00809_, _00805_);
  or _22462_ (_00812_, _00811_, _00810_);
  or _22463_ (_00813_, _00812_, _00605_);
  and _22464_ (_00814_, _00813_, _00804_);
  or _22465_ (_00815_, _00814_, _00610_);
  nand _22466_ (_00816_, _00610_, _00805_);
  and _22467_ (_00817_, _00816_, _04856_);
  and _22468_ (_12137_, _00817_, _00815_);
  or _22469_ (_00818_, _12818_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  or _22470_ (_00819_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _09249_);
  or _22471_ (_00820_, _00819_, _08087_);
  and _22472_ (_00821_, _00820_, _04856_);
  and _22473_ (_12141_, _00821_, _00818_);
  nor _22474_ (_00822_, _05669_, _06046_);
  and _22475_ (_00823_, _06046_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  or _22476_ (_00824_, _00823_, _05673_);
  or _22477_ (_00825_, _00824_, _00822_);
  or _22478_ (_00826_, _04861_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  and _22479_ (_00827_, _00826_, _04856_);
  and _22480_ (_12147_, _00827_, _00825_);
  nor _22481_ (_00828_, _00756_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nor _22482_ (_00829_, _00828_, _00757_);
  or _22483_ (_00830_, _00829_, _00605_);
  nand _22484_ (_00831_, _00605_, _06032_);
  and _22485_ (_00832_, _00831_, _00830_);
  or _22486_ (_00833_, _00832_, _00610_);
  not _22487_ (_00834_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nand _22488_ (_00835_, _00610_, _00834_);
  and _22489_ (_00836_, _00835_, _04856_);
  and _22490_ (_12151_, _00836_, _00833_);
  or _22491_ (_00837_, _06238_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  not _22492_ (_00838_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nand _22493_ (_00839_, _06238_, _00838_);
  and _22494_ (_00840_, _00839_, _04856_);
  and _22495_ (_12154_, _00840_, _00837_);
  nand _22496_ (_00841_, _00605_, _06369_);
  nand _22497_ (_00842_, _00629_, _00616_);
  and _22498_ (_00843_, _00842_, _00691_);
  or _22499_ (_00844_, _00619_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and _22500_ (_00845_, _00844_, _00843_);
  and _22501_ (_00846_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  or _22502_ (_00847_, _00616_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and _22503_ (_00848_, _00752_, _00729_);
  and _22504_ (_00849_, _00848_, _00847_);
  or _22505_ (_00850_, _00849_, _00846_);
  or _22506_ (_00851_, _00850_, _00845_);
  or _22507_ (_00852_, _00851_, _00605_);
  and _22508_ (_00853_, _00852_, _00841_);
  or _22509_ (_00854_, _00853_, _00610_);
  or _22510_ (_00855_, _00653_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and _22511_ (_00856_, _00855_, _04856_);
  and _22512_ (_12156_, _00856_, _00854_);
  and _22513_ (_00857_, _00330_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and _22514_ (_00858_, _00332_, _06997_);
  and _22515_ (_00859_, _00351_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  nor _22516_ (_00860_, _00351_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  nor _22517_ (_00861_, _00860_, _00859_);
  and _22518_ (_00862_, _00413_, _00441_);
  or _22519_ (_00863_, _00862_, _00861_);
  and _22520_ (_00864_, _00863_, _00379_);
  or _22521_ (_00866_, _00864_, _00858_);
  or _22522_ (_00867_, _00866_, _00857_);
  and _22523_ (_12163_, _00867_, _04856_);
  or _22524_ (_00868_, _00516_, _06705_);
  and _22525_ (_00869_, _00868_, _04856_);
  nor _22526_ (_00870_, _04984_, _04947_);
  and _22527_ (_00871_, _00870_, _04989_);
  and _22528_ (_00872_, _00871_, _05517_);
  and _22529_ (_00873_, _00872_, _05510_);
  and _22530_ (_00874_, _00341_, _00351_);
  nor _22531_ (_00875_, _00874_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  and _22532_ (_00876_, _00874_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  nor _22533_ (_00877_, _00876_, _00875_);
  and _22534_ (_00878_, _00413_, _00440_);
  and _22535_ (_00879_, _00878_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nor _22536_ (_00880_, _00879_, _00877_);
  nor _22537_ (_00881_, _00880_, _00873_);
  and _22538_ (_00882_, _00873_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  or _22539_ (_00883_, _00882_, _00881_);
  or _22540_ (_00884_, _00883_, _00332_);
  and _22541_ (_12169_, _00884_, _00869_);
  and _22542_ (_00885_, _00330_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  nor _22543_ (_00886_, _00876_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  nor _22544_ (_00887_, _00886_, _00362_);
  and _22545_ (_00888_, _00878_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  or _22546_ (_00889_, _00888_, _00887_);
  and _22547_ (_00890_, _00889_, _00379_);
  or _22548_ (_00891_, _00890_, _00885_);
  nor _22549_ (_00892_, _00516_, _05669_);
  or _22550_ (_00893_, _00892_, _00891_);
  and _22551_ (_12172_, _00893_, _04856_);
  and _22552_ (_00894_, _00330_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  nor _22553_ (_00895_, _00516_, _06032_);
  nor _22554_ (_00896_, _00859_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  nor _22555_ (_00897_, _00896_, _00874_);
  and _22556_ (_00898_, _00878_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  or _22557_ (_00899_, _00898_, _00897_);
  and _22558_ (_00900_, _00899_, _00379_);
  or _22559_ (_00901_, _00900_, _00895_);
  or _22560_ (_00902_, _00901_, _00894_);
  and _22561_ (_12173_, _00902_, _04856_);
  and _22562_ (_00903_, _00330_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and _22563_ (_00904_, _00363_, _00448_);
  and _22564_ (_00905_, _00904_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  nor _22565_ (_00906_, _00904_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  nor _22566_ (_00907_, _00906_, _00905_);
  and _22567_ (_00908_, _00878_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  or _22568_ (_00909_, _00908_, _00907_);
  and _22569_ (_00910_, _00909_, _00379_);
  or _22570_ (_00911_, _00910_, _00903_);
  and _22571_ (_00912_, _00332_, _05718_);
  or _22572_ (_00913_, _00912_, _00911_);
  and _22573_ (_12178_, _00913_, _04856_);
  and _22574_ (_00914_, _00330_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and _22575_ (_00915_, _00878_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nand _22576_ (_00916_, _00448_, _00439_);
  or _22577_ (_00917_, _00905_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and _22578_ (_00918_, _00917_, _00916_);
  or _22579_ (_00919_, _00918_, _00915_);
  and _22580_ (_00920_, _00919_, _00379_);
  or _22581_ (_00921_, _00920_, _00914_);
  nor _22582_ (_00922_, _00516_, _05287_);
  or _22583_ (_00923_, _00922_, _00921_);
  and _22584_ (_12181_, _00923_, _04856_);
  nor _22585_ (_00924_, _00362_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  nor _22586_ (_00925_, _00924_, _00363_);
  and _22587_ (_00926_, _00413_, _00355_);
  and _22588_ (_00927_, _00926_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nor _22589_ (_00928_, _00927_, _00925_);
  nor _22590_ (_00929_, _00928_, _00873_);
  and _22591_ (_00930_, _00873_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  or _22592_ (_00931_, _00930_, _00929_);
  and _22593_ (_00932_, _00931_, _00516_);
  and _22594_ (_00933_, _00332_, _06410_);
  or _22595_ (_00934_, _00933_, _00932_);
  and _22596_ (_12184_, _00934_, _04856_);
  and _22597_ (_12211_, _05963_, _04856_);
  or _22598_ (_00935_, _08367_, \oc8051_top_1.oc8051_rom1.data_o [11]);
  nand _22599_ (_00936_, _08367_, _05803_);
  and _22600_ (_00937_, _00936_, _04856_);
  and _22601_ (_12229_, _00937_, _00935_);
  or _22602_ (_00938_, _08367_, \oc8051_top_1.oc8051_rom1.data_o [4]);
  nand _22603_ (_00939_, _08367_, _05850_);
  and _22604_ (_00940_, _00939_, _04856_);
  and _22605_ (_12234_, _00940_, _00938_);
  and _22606_ (_00941_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and _22607_ (_00942_, _12165_, \oc8051_top_1.oc8051_rom1.data_o [23]);
  or _22608_ (_00943_, _00942_, _00941_);
  and _22609_ (_12239_, _00943_, _04856_);
  and _22610_ (_00944_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and _22611_ (_00945_, _12165_, \oc8051_top_1.oc8051_rom1.data_o [17]);
  or _22612_ (_00946_, _00945_, _00944_);
  and _22613_ (_12251_, _00946_, _04856_);
  nand _22614_ (_00947_, _12719_, _06369_);
  or _22615_ (_00948_, _12716_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  or _22616_ (_00949_, _12717_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and _22617_ (_00950_, _00949_, _00948_);
  or _22618_ (_00951_, _00950_, _12719_);
  and _22619_ (_00952_, _00951_, _00947_);
  or _22620_ (_00953_, _00952_, _12714_);
  or _22621_ (_00954_, _12715_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  and _22622_ (_00955_, _00954_, _04856_);
  and _22623_ (_12255_, _00955_, _00953_);
  and _22624_ (_00956_, _06238_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  not _22625_ (_00957_, _06238_);
  and _22626_ (_00958_, _00957_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  or _22627_ (_00959_, _00958_, _00956_);
  and _22628_ (_12267_, _00959_, _04856_);
  or _22629_ (_00960_, _06238_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nand _22630_ (_00961_, _06238_, _05295_);
  and _22631_ (_00962_, _00961_, _04856_);
  and _22632_ (_12274_, _00962_, _00960_);
  nand _22633_ (_00963_, _12171_, _06552_);
  or _22634_ (_00964_, _12171_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2]);
  and _22635_ (_00965_, _00964_, _04856_);
  and _22636_ (_12280_, _00965_, _00963_);
  nand _22637_ (_00966_, _12171_, _07774_);
  or _22638_ (_00967_, _12171_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1]);
  and _22639_ (_00968_, _00967_, _04856_);
  and _22640_ (_12300_, _00968_, _00966_);
  and _22641_ (_12303_, _07212_, _04856_);
  nor _22642_ (_12317_, _06925_, rst);
  not _22643_ (_00969_, _07815_);
  and _22644_ (_00970_, _13037_, _00969_);
  and _22645_ (_00971_, _12879_, _12829_);
  and _22646_ (_00972_, _06847_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and _22647_ (_00973_, _12861_, _12534_);
  or _22648_ (_00974_, _00973_, _00972_);
  or _22649_ (_00975_, _00974_, _00971_);
  or _22650_ (_00976_, _00975_, _00970_);
  or _22651_ (_00977_, _12989_, _12987_);
  and _22652_ (_00978_, _00977_, _12990_);
  and _22653_ (_00979_, _00978_, _13070_);
  or _22654_ (_00980_, _00979_, _00976_);
  and _22655_ (_00981_, _00980_, _12547_);
  nor _22656_ (_00982_, _08369_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or _22657_ (_00983_, _00982_, _13052_);
  nor _22658_ (_00984_, _00983_, _12547_);
  or _22659_ (_00985_, _00984_, _00981_);
  and _22660_ (_12338_, _00985_, _04856_);
  nand _22661_ (_00986_, _13108_, _05142_);
  or _22662_ (_00987_, _00986_, _13091_);
  nand _22663_ (_00988_, _13111_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and _22664_ (_00989_, _00988_, _00987_);
  nand _22665_ (_00990_, _00989_, _05157_);
  or _22666_ (_00991_, _00989_, _05157_);
  and _22667_ (_00992_, _00991_, _13031_);
  and _22668_ (_00993_, _00992_, _00990_);
  and _22669_ (_00994_, _13022_, _07598_);
  and _22670_ (_00995_, _13042_, _05919_);
  not _22671_ (_00996_, _07089_);
  and _22672_ (_00997_, _12829_, _00996_);
  or _22673_ (_00998_, _00997_, _00995_);
  and _22674_ (_00999_, _13036_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor _22675_ (_01000_, _06901_, _06552_);
  or _22676_ (_01001_, _01000_, _00999_);
  or _22677_ (_01002_, _01001_, _00998_);
  nor _22678_ (_01003_, _01002_, _00994_);
  nand _22679_ (_01004_, _01003_, _12547_);
  or _22680_ (_01005_, _01004_, _00993_);
  and _22681_ (_01006_, _13124_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor _22682_ (_01007_, _13124_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor _22683_ (_01008_, _01007_, _01006_);
  or _22684_ (_01009_, _01008_, _12547_);
  and _22685_ (_01010_, _01009_, _04856_);
  and _22686_ (_12343_, _01010_, _01005_);
  or _22687_ (_01011_, _12688_, _12683_);
  or _22688_ (_01012_, _05988_, _05949_);
  or _22689_ (_01013_, _06598_, _05965_);
  and _22690_ (_01014_, _01013_, _01012_);
  or _22691_ (_01015_, _01014_, _00548_);
  or _22692_ (_01016_, _01015_, _01011_);
  and _22693_ (_01017_, _06635_, _06730_);
  or _22694_ (_01018_, _08194_, _07508_);
  or _22695_ (_01019_, _01018_, _01017_);
  or _22696_ (_01021_, _06747_, _06724_);
  or _22697_ (_01022_, _01021_, _01019_);
  or _22698_ (_01024_, _01022_, _01016_);
  and _22699_ (_01025_, _01024_, _05730_);
  and _22700_ (_01026_, \oc8051_top_1.oc8051_decoder1.alu_op [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and _22701_ (_01027_, _06002_, _04859_);
  or _22702_ (_01028_, _01027_, _01026_);
  or _22703_ (_01029_, _01028_, _01025_);
  and _22704_ (_12372_, _01029_, _04856_);
  and _22705_ (_01030_, _05718_, _05675_);
  and _22706_ (_01032_, _06046_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  or _22707_ (_01033_, _01032_, _05673_);
  or _22708_ (_01034_, _01033_, _01030_);
  or _22709_ (_01035_, _04861_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  and _22710_ (_01036_, _01035_, _04856_);
  and _22711_ (_12445_, _01036_, _01034_);
  or _22712_ (_12482_, _07102_, rst);
  and _22713_ (_12485_, _07310_, _04856_);
  nor _22714_ (_12489_, _07274_, rst);
  and _22715_ (_12491_, _07223_, _04856_);
  nor _22716_ (_12493_, _07154_, rst);
  nand _22717_ (_12496_, _07067_, _04856_);
  nor _22718_ (_12621_, _07191_, rst);
  nor _22719_ (_12646_, _07142_, rst);
  and _22720_ (_01038_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _22721_ (_01039_, _00030_, _00028_);
  and _22722_ (_01041_, _01039_, _00031_);
  or _22723_ (_01042_, _01041_, _06911_);
  or _22724_ (_01043_, _06910_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and _22725_ (_01045_, _01043_, _00059_);
  and _22726_ (_01046_, _01045_, _01042_);
  or _22727_ (_01047_, _01046_, _01038_);
  and _22728_ (_12670_, _01047_, _04856_);
  not _22729_ (_01048_, _10587_);
  or _22730_ (_01049_, _01048_, _06410_);
  or _22731_ (_01050_, _10587_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  and _22732_ (_01052_, _01050_, _04856_);
  and _22733_ (_12673_, _01052_, _01049_);
  and _22734_ (_01053_, _12206_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  or _22735_ (_01054_, _01053_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and _22736_ (_12679_, _01054_, _04856_);
  nor _22737_ (_01055_, _05287_, _06046_);
  and _22738_ (_01056_, _06046_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  or _22739_ (_01057_, _01056_, _05673_);
  or _22740_ (_01058_, _01057_, _01055_);
  or _22741_ (_01059_, _04861_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  and _22742_ (_01060_, _01059_, _04856_);
  and _22743_ (_12690_, _01060_, _01058_);
  and _22744_ (_01061_, _12206_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  or _22745_ (_01062_, _01061_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  and _22746_ (_12694_, _01062_, _04856_);
  or _22747_ (_01063_, _00027_, _12371_);
  nor _22748_ (_01064_, _00028_, _06911_);
  and _22749_ (_01065_, _01064_, _01063_);
  nor _22750_ (_01067_, _06910_, _05109_);
  or _22751_ (_01068_, _01067_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _22752_ (_01069_, _01068_, _01065_);
  or _22753_ (_01070_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], _00059_);
  and _22754_ (_01071_, _01070_, _04856_);
  and _22755_ (_12702_, _01071_, _01069_);
  and _22756_ (_01072_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14], \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  not _22757_ (_01073_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor _22758_ (_01074_, _00146_, _01073_);
  and _22759_ (_01075_, _00146_, _01073_);
  or _22760_ (_01076_, _01075_, _01074_);
  nand _22761_ (_01077_, _01076_, _00183_);
  or _22762_ (_01078_, _01076_, _00183_);
  and _22763_ (_01079_, _01078_, _01077_);
  or _22764_ (_01080_, _01079_, _06911_);
  or _22765_ (_01081_, _06910_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and _22766_ (_01082_, _01081_, _00059_);
  and _22767_ (_01083_, _01082_, _01080_);
  or _22768_ (_01084_, _01083_, _01072_);
  and _22769_ (_12706_, _01084_, _04856_);
  and _22770_ (_01085_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7], \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  nor _22771_ (_01086_, _00174_, _00055_);
  nor _22772_ (_01087_, _01086_, _00175_);
  or _22773_ (_01088_, _01087_, _06911_);
  or _22774_ (_01089_, _06910_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and _22775_ (_01090_, _01089_, _00059_);
  and _22776_ (_01091_, _01090_, _01088_);
  or _22777_ (_01092_, _01091_, _01085_);
  and _22778_ (_12712_, _01092_, _04856_);
  nor _22779_ (_12736_, _07261_, rst);
  and _22780_ (_01093_, _12206_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  or _22781_ (_01094_, _01093_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and _22782_ (_12750_, _01094_, _04856_);
  and _22783_ (_12819_, _10047_, _06994_);
  nand _22784_ (_01095_, _07774_, _06498_);
  not _22785_ (_01096_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  nand _22786_ (_01097_, _06497_, _01096_);
  and _22787_ (_01098_, _01097_, _04856_);
  and _22788_ (_12951_, _01098_, _01095_);
  nor _22789_ (_01099_, _12257_, _08816_);
  or _22790_ (_01100_, _01099_, _07642_);
  and _22791_ (_01101_, _01100_, _09259_);
  and _22792_ (_01102_, _09259_, _04984_);
  nor _22793_ (_01103_, _01102_, _08816_);
  or _22794_ (_01104_, _01103_, _09263_);
  or _22795_ (_01105_, _01104_, _01101_);
  nand _22796_ (_01106_, _09263_, _05669_);
  and _22797_ (_01107_, _01106_, _04856_);
  and _22798_ (_13002_, _01107_, _01105_);
  nor _22799_ (_01108_, _07702_, _06497_);
  and _22800_ (_01109_, _06497_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  or _22801_ (_01111_, _01109_, _01108_);
  and _22802_ (_13064_, _01111_, _04856_);
  not _22803_ (_01113_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  nor _22804_ (_01114_, _08060_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and _22805_ (_01116_, _01114_, _01113_);
  nor _22806_ (_01117_, _01116_, _08922_);
  and _22807_ (_01118_, _01116_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  or _22808_ (_01119_, _01118_, _01117_);
  or _22809_ (_01120_, _01119_, _09259_);
  or _22810_ (_01121_, _06494_, _08922_);
  nand _22811_ (_01122_, _01121_, _09259_);
  or _22812_ (_01123_, _01122_, _07602_);
  and _22813_ (_01124_, _01123_, _01120_);
  or _22814_ (_01125_, _01124_, _09263_);
  or _22815_ (_01126_, _09264_, _06705_);
  and _22816_ (_01127_, _01126_, _04856_);
  and _22817_ (_13158_, _01127_, _01125_);
  nor _22818_ (_01128_, _01006_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and _22819_ (_01129_, _01006_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor _22820_ (_01130_, _01129_, _01128_);
  or _22821_ (_01131_, _01130_, _12547_);
  and _22822_ (_01132_, _01131_, _04856_);
  and _22823_ (_01133_, _13022_, _07640_);
  and _22824_ (_01134_, _12829_, _12885_);
  nor _22825_ (_01135_, _06901_, _06586_);
  or _22826_ (_01136_, _01135_, _01134_);
  and _22827_ (_01137_, \oc8051_top_1.oc8051_memory_interface1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and _22828_ (_01138_, _01137_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and _22829_ (_01139_, \oc8051_top_1.oc8051_memory_interface1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _22830_ (_01140_, _01139_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and _22831_ (_01141_, \oc8051_top_1.oc8051_memory_interface1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and _22832_ (_01142_, \oc8051_top_1.oc8051_memory_interface1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and _22833_ (_01143_, _01142_, _01141_);
  and _22834_ (_01144_, _01143_, _01140_);
  and _22835_ (_01145_, _01144_, _01138_);
  and _22836_ (_01146_, _01145_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor _22837_ (_01148_, _01145_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor _22838_ (_01149_, _01148_, _01146_);
  and _22839_ (_01150_, _01149_, _13042_);
  and _22840_ (_01151_, _13036_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  or _22841_ (_01152_, _01151_, _01150_);
  or _22842_ (_01153_, _01152_, _01136_);
  nor _22843_ (_01155_, _01153_, _01133_);
  nand _22844_ (_01156_, _01155_, _12547_);
  not _22845_ (_01157_, _01138_);
  nor _22846_ (_01159_, _01157_, _13107_);
  and _22847_ (_01160_, _01159_, _13091_);
  nor _22848_ (_01161_, _00986_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and _22849_ (_01162_, _01161_, _13092_);
  nor _22850_ (_01163_, _01162_, _01160_);
  nand _22851_ (_01165_, _01163_, _05089_);
  or _22852_ (_01166_, _01163_, _05089_);
  and _22853_ (_01167_, _01166_, _01165_);
  and _22854_ (_01168_, _01167_, _13070_);
  or _22855_ (_01169_, _01168_, _01156_);
  and _22856_ (_13165_, _01169_, _01132_);
  and _22857_ (_01170_, _09259_, _06091_);
  and _22858_ (_01171_, _01170_, _06144_);
  nor _22859_ (_01172_, _01170_, _00246_);
  or _22860_ (_01173_, _01172_, _09263_);
  or _22861_ (_01174_, _01173_, _01171_);
  or _22862_ (_01175_, _09264_, _05718_);
  and _22863_ (_01176_, _01175_, _04856_);
  and _22864_ (_13168_, _01176_, _01174_);
  nand _22865_ (_01177_, _01161_, _05089_);
  or _22866_ (_01178_, _01177_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor _22867_ (_01179_, _01178_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  or _22868_ (_01180_, _01179_, _13091_);
  and _22869_ (_01181_, _01159_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _22870_ (_01182_, _01181_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nand _22871_ (_01183_, _01182_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nand _22872_ (_01184_, _01183_, _13091_);
  and _22873_ (_01185_, _01184_, _01180_);
  nor _22874_ (_01186_, _01185_, _05022_);
  and _22875_ (_01187_, _01185_, _05022_);
  or _22876_ (_01188_, _01187_, _01186_);
  and _22877_ (_01189_, _01188_, _13031_);
  and _22878_ (_01190_, _13022_, _06452_);
  nor _22879_ (_01191_, _06901_, _06488_);
  and _22880_ (_01192_, _13036_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  and _22881_ (_01193_, _01146_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _22882_ (_01194_, _01193_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor _22883_ (_01195_, _01194_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and _22884_ (_01196_, _01194_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor _22885_ (_01197_, _01196_, _01195_);
  and _22886_ (_01198_, _01197_, _13042_);
  and _22887_ (_01199_, _12829_, _12995_);
  or _22888_ (_01200_, _01199_, _01198_);
  or _22889_ (_01201_, _01200_, _01192_);
  or _22890_ (_01202_, _01201_, _01191_);
  nor _22891_ (_01203_, _01202_, _01190_);
  nand _22892_ (_01204_, _01203_, _12547_);
  or _22893_ (_01205_, _01204_, _01189_);
  and _22894_ (_01206_, _01129_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and _22895_ (_01207_, _01206_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor _22896_ (_01208_, _01207_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  and _22897_ (_01209_, _01207_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor _22898_ (_01210_, _01209_, _01208_);
  or _22899_ (_01211_, _01210_, _12547_);
  and _22900_ (_01212_, _01211_, _04856_);
  and _22901_ (_13188_, _01212_, _01205_);
  and _22902_ (_01213_, _01178_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  or _22903_ (_01214_, _01213_, _01180_);
  or _22904_ (_01215_, _01182_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and _22905_ (_01216_, _01215_, _01183_);
  or _22906_ (_01217_, _01216_, _13092_);
  and _22907_ (_01218_, _01217_, _13031_);
  and _22908_ (_01219_, _01218_, _01214_);
  and _22909_ (_01220_, _13022_, _07924_);
  nor _22910_ (_01221_, _01193_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor _22911_ (_01222_, _01221_, _01194_);
  and _22912_ (_01223_, _01222_, _13042_);
  and _22913_ (_01224_, _13036_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or _22914_ (_01225_, _01224_, _01223_);
  and _22915_ (_01226_, _12829_, _13063_);
  nor _22916_ (_01227_, _07897_, _06901_);
  or _22917_ (_01228_, _01227_, _01226_);
  or _22918_ (_01229_, _01228_, _01225_);
  nor _22919_ (_01230_, _01229_, _01220_);
  nand _22920_ (_01231_, _01230_, _12547_);
  or _22921_ (_01232_, _01231_, _01219_);
  nor _22922_ (_01233_, _01206_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor _22923_ (_01234_, _01233_, _01207_);
  or _22924_ (_01235_, _01234_, _12547_);
  and _22925_ (_01236_, _01235_, _04856_);
  and _22926_ (_13196_, _01236_, _01232_);
  nand _22927_ (_01237_, _01177_, _13092_);
  or _22928_ (_01238_, _01181_, _13092_);
  nand _22929_ (_01239_, _01238_, _01237_);
  nand _22930_ (_01240_, _01239_, _05067_);
  or _22931_ (_01241_, _01239_, _05067_);
  and _22932_ (_01242_, _01241_, _13031_);
  and _22933_ (_01243_, _01242_, _01240_);
  and _22934_ (_01244_, _13022_, _07853_);
  nor _22935_ (_01245_, _07815_, _06901_);
  and _22936_ (_01246_, _12829_, _12860_);
  or _22937_ (_01247_, _01246_, _01245_);
  nor _22938_ (_01248_, _01146_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor _22939_ (_01249_, _01248_, _01193_);
  and _22940_ (_01250_, _01249_, _13042_);
  and _22941_ (_01251_, _13036_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  or _22942_ (_01252_, _01251_, _01250_);
  or _22943_ (_01253_, _01252_, _01247_);
  nor _22944_ (_01254_, _01253_, _01244_);
  nand _22945_ (_01255_, _01254_, _12547_);
  or _22946_ (_01256_, _01255_, _01243_);
  nor _22947_ (_01257_, _01129_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor _22948_ (_01258_, _01257_, _01206_);
  or _22949_ (_01259_, _01258_, _12547_);
  and _22950_ (_01260_, _01259_, _04856_);
  and _22951_ (_13203_, _01260_, _01256_);
  and _22952_ (_01261_, _09259_, _07857_);
  not _22953_ (_01262_, _09259_);
  or _22954_ (_01263_, _12246_, _01262_);
  or _22955_ (_01264_, _01263_, _01102_);
  and _22956_ (_01265_, _01264_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  or _22957_ (_01266_, _01265_, _09263_);
  or _22958_ (_01267_, _01266_, _01261_);
  or _22959_ (_01268_, _09264_, _06410_);
  and _22960_ (_01269_, _01268_, _04856_);
  and _22961_ (_13205_, _01269_, _01267_);
  and _22962_ (_01270_, _06370_, _05675_);
  nand _22963_ (_01271_, _05675_, _04861_);
  and _22964_ (_01272_, _01271_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  or _22965_ (_01273_, _01272_, _01270_);
  and _22966_ (_00041_, _01273_, _04856_);
  nand _22967_ (_01274_, _00332_, _06284_);
  nand _22968_ (_01275_, _00878_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or _22969_ (_01276_, _00916_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and _22970_ (_01277_, _01276_, _01275_);
  nor _22971_ (_01278_, _01277_, _00330_);
  or _22972_ (_01279_, _00916_, _00330_);
  and _22973_ (_01280_, _01279_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  or _22974_ (_01281_, _01280_, _01278_);
  or _22975_ (_01282_, _01281_, _00332_);
  and _22976_ (_01283_, _01282_, _04856_);
  and _22977_ (_00115_, _01283_, _01274_);
  nand _22978_ (_01284_, _00330_, _06284_);
  and _22979_ (_01285_, _00358_, _00334_);
  nand _22980_ (_01286_, _01285_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or _22981_ (_01287_, _01285_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and _22982_ (_01288_, _01287_, _01286_);
  and _22983_ (_01289_, _01288_, _00414_);
  and _22984_ (_01290_, _00369_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and _22985_ (_01291_, _01290_, _00340_);
  and _22986_ (_01292_, _01291_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or _22987_ (_01293_, _01291_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand _22988_ (_01294_, _01293_, _00423_);
  nor _22989_ (_01295_, _01294_, _01292_);
  and _22990_ (_01296_, _00344_, _00351_);
  and _22991_ (_01297_, _00340_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and _22992_ (_01298_, _01297_, _01296_);
  or _22993_ (_01299_, _01298_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and _22994_ (_01300_, _01297_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand _22995_ (_01301_, _01300_, _01296_);
  and _22996_ (_01302_, _01301_, _00361_);
  and _22997_ (_01303_, _01302_, _01299_);
  or _22998_ (_01304_, _01303_, _01295_);
  or _22999_ (_01305_, _01304_, _00330_);
  or _23000_ (_01306_, _01305_, _01289_);
  and _23001_ (_01307_, _01306_, _00516_);
  and _23002_ (_01308_, _01307_, _01284_);
  and _23003_ (_01309_, _00332_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or _23004_ (_01310_, _01309_, _01308_);
  and _23005_ (_00116_, _01310_, _04856_);
  and _23006_ (_01311_, _00610_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nand _23007_ (_01312_, _00605_, _06284_);
  or _23008_ (_01313_, _00741_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nand _23009_ (_01314_, _01313_, _00691_);
  and _23010_ (_01315_, _00741_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor _23011_ (_01316_, _01315_, _01314_);
  nand _23012_ (_01318_, _00690_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  or _23013_ (_01319_, _01318_, _00732_);
  and _23014_ (_01320_, _00731_, _00729_);
  or _23015_ (_01321_, _01320_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and _23016_ (_01322_, _01321_, _01319_);
  or _23017_ (_01323_, _01322_, _01316_);
  or _23018_ (_01324_, _01323_, _00605_);
  and _23019_ (_01325_, _01324_, _00653_);
  and _23020_ (_01326_, _01325_, _01312_);
  or _23021_ (_01327_, _01326_, _01311_);
  and _23022_ (_00121_, _01327_, _04856_);
  nor _23023_ (_01328_, _00351_, _06099_);
  or _23024_ (_01329_, _01300_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  or _23025_ (_01330_, _00361_, _00440_);
  nand _23026_ (_01331_, _01330_, _01329_);
  nor _23027_ (_01332_, _01331_, _01302_);
  or _23028_ (_01333_, _01332_, _01328_);
  and _23029_ (_01334_, _01333_, _04856_);
  and _23030_ (_00124_, _01334_, _00379_);
  not _23031_ (_01335_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  nor _23032_ (_01336_, _00598_, _01335_);
  or _23033_ (_01337_, _01336_, _01315_);
  and _23034_ (_01338_, _01337_, _00691_);
  and _23035_ (_01339_, _01320_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nand _23036_ (_01340_, _00598_, _00611_);
  nor _23037_ (_01341_, _00691_, _01335_);
  and _23038_ (_01342_, _01341_, _01340_);
  or _23039_ (_01343_, _01342_, _00620_);
  or _23040_ (_01344_, _01343_, _01339_);
  or _23041_ (_01345_, _01344_, _01338_);
  nor _23042_ (_01346_, _00605_, rst);
  and _23043_ (_01347_, _01346_, _00653_);
  and _23044_ (_00126_, _01347_, _01345_);
  or _23045_ (_01348_, _04989_, _06090_);
  not _23046_ (_01349_, _01348_);
  or _23047_ (_01350_, _01349_, _07855_);
  and _23048_ (_01351_, _06668_, _06930_);
  and _23049_ (_01352_, _01351_, _06670_);
  nand _23050_ (_01353_, _01352_, _01350_);
  and _23051_ (_01354_, _01353_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and _23052_ (_01355_, _01349_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  or _23053_ (_01356_, _01355_, _07857_);
  and _23054_ (_01357_, _01356_, _01352_);
  or _23055_ (_01358_, _01357_, _01354_);
  and _23056_ (_01359_, _01358_, _06093_);
  and _23057_ (_01360_, _08999_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and _23058_ (_01361_, _09122_, _06662_);
  nand _23059_ (_01362_, _01361_, _07815_);
  or _23060_ (_01363_, _01361_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and _23061_ (_01364_, _01363_, _05510_);
  and _23062_ (_01365_, _01364_, _01362_);
  or _23063_ (_01366_, _01365_, _01360_);
  or _23064_ (_01367_, _01366_, _01359_);
  and _23065_ (_00130_, _01367_, _04856_);
  nand _23066_ (_01368_, _00610_, _06284_);
  and _23067_ (_01369_, _00694_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and _23068_ (_01370_, _00620_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor _23069_ (_01371_, _00618_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  nor _23070_ (_01372_, _01371_, _00619_);
  and _23071_ (_01373_, _01372_, _00709_);
  nor _23072_ (_01374_, _01373_, _01370_);
  nor _23073_ (_01375_, _01374_, _00605_);
  or _23074_ (_01376_, _01375_, _01369_);
  or _23075_ (_01377_, _01376_, _00610_);
  and _23076_ (_01378_, _01377_, _04856_);
  and _23077_ (_00133_, _01378_, _01368_);
  not _23078_ (_01379_, _12547_);
  and _23079_ (_01380_, _13037_, _13153_);
  and _23080_ (_01381_, _06847_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and _23081_ (_01382_, _12973_, _12829_);
  and _23082_ (_01383_, _12955_, _12534_);
  or _23083_ (_01384_, _01383_, _01382_);
  or _23084_ (_01385_, _01384_, _01381_);
  or _23085_ (_01386_, _01385_, _01380_);
  nor _23086_ (_01387_, _12975_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor _23087_ (_01388_, _01387_, _12976_);
  and _23088_ (_01389_, _01388_, _13070_);
  or _23089_ (_01390_, _01389_, _01386_);
  or _23090_ (_01391_, _01390_, _01379_);
  or _23091_ (_01392_, _12547_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and _23092_ (_01393_, _01392_, _04856_);
  and _23093_ (_00137_, _01393_, _01391_);
  and _23094_ (_00140_, t1_i, _04856_);
  and _23095_ (_01394_, _01352_, _05520_);
  and _23096_ (_01395_, _01394_, _06088_);
  nor _23097_ (_01396_, _01394_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  or _23098_ (_01398_, _01396_, _06094_);
  nor _23099_ (_01399_, _01398_, _01395_);
  and _23100_ (_01400_, _08999_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  not _23101_ (_01401_, _01361_);
  and _23102_ (_01402_, _01401_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nor _23103_ (_01403_, _01401_, _06586_);
  or _23104_ (_01404_, _01403_, _01402_);
  and _23105_ (_01405_, _01404_, _05510_);
  or _23106_ (_01407_, _01405_, _01400_);
  or _23107_ (_01408_, _01407_, _01399_);
  and _23108_ (_00144_, _01408_, _04856_);
  and _23109_ (_00150_, t0_i, _04856_);
  not _23110_ (_01409_, _06586_);
  and _23111_ (_01410_, _13037_, _01409_);
  and _23112_ (_01411_, _12904_, _12829_);
  and _23113_ (_01413_, _12886_, _12534_);
  and _23114_ (_01414_, _06847_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  or _23115_ (_01416_, _01414_, _01413_);
  or _23116_ (_01417_, _01416_, _01411_);
  or _23117_ (_01418_, _01417_, _01410_);
  or _23118_ (_01419_, _12907_, _12908_);
  and _23119_ (_01420_, _01419_, _12985_);
  nor _23120_ (_01421_, _01419_, _12985_);
  or _23121_ (_01422_, _01421_, _01420_);
  and _23122_ (_01423_, _01422_, _13070_);
  or _23123_ (_01424_, _01423_, _01418_);
  or _23124_ (_01425_, _01424_, _01379_);
  or _23125_ (_01426_, _12547_, _08371_);
  and _23126_ (_01428_, _01426_, _04856_);
  and _23127_ (_00157_, _01428_, _01425_);
  or _23128_ (_01429_, _00279_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and _23129_ (_01430_, _01429_, _04856_);
  nand _23130_ (_01431_, _00279_, _06284_);
  and _23131_ (_00165_, _01431_, _01430_);
  and _23132_ (_01433_, _01352_, _06146_);
  nand _23133_ (_01434_, _01433_, _06088_);
  or _23134_ (_01435_, _01433_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and _23135_ (_01436_, _01435_, _06093_);
  and _23136_ (_01438_, _01436_, _01434_);
  and _23137_ (_01439_, _08999_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  nand _23138_ (_01440_, _01361_, _06488_);
  or _23139_ (_01441_, _01361_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and _23140_ (_01442_, _01441_, _05510_);
  and _23141_ (_01443_, _01442_, _01440_);
  or _23142_ (_01444_, _01443_, _01439_);
  or _23143_ (_01445_, _01444_, _01438_);
  and _23144_ (_00168_, _01445_, _04856_);
  not _23145_ (_01446_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 );
  nor _23146_ (_01447_, _00369_, _01446_);
  or _23147_ (_01448_, _01447_, _01292_);
  and _23148_ (_01449_, _00423_, _04856_);
  and _23149_ (_01450_, _01449_, _01448_);
  and _23150_ (_00170_, _01450_, _00379_);
  and _23151_ (_01451_, _06847_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  not _23152_ (_01452_, _06552_);
  and _23153_ (_01453_, _13037_, _01452_);
  nor _23154_ (_01454_, _12926_, _12830_);
  and _23155_ (_01455_, _13042_, _00996_);
  or _23156_ (_01456_, _01455_, _01454_);
  or _23157_ (_01457_, _01456_, _01453_);
  nor _23158_ (_01458_, _12983_, _12981_);
  nor _23159_ (_01459_, _01458_, _12984_);
  and _23160_ (_01460_, _01459_, _13070_);
  or _23161_ (_01461_, _01460_, _01457_);
  or _23162_ (_01462_, _01461_, _01451_);
  and _23163_ (_01463_, _01462_, _12547_);
  and _23164_ (_01464_, _01379_, _08387_);
  or _23165_ (_01465_, _01464_, _01463_);
  and _23166_ (_00177_, _01465_, _04856_);
  and _23167_ (_01466_, _12548_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  and _23168_ (_01467_, _12952_, _12534_);
  not _23169_ (_01468_, _07774_);
  and _23170_ (_01469_, _13037_, _01468_);
  or _23171_ (_01470_, _01469_, _01467_);
  nor _23172_ (_01471_, _12978_, _12976_);
  nor _23173_ (_01472_, _01471_, _12979_);
  and _23174_ (_01473_, _01472_, _13070_);
  or _23175_ (_01474_, _01473_, _01470_);
  and _23176_ (_01475_, _01474_, _12547_);
  or _23177_ (_01476_, _01475_, _01466_);
  and _23178_ (_00196_, _01476_, _04856_);
  and _23179_ (_01477_, _01352_, _04986_);
  nand _23180_ (_01478_, _01477_, _06088_);
  or _23181_ (_01479_, _01477_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and _23182_ (_01480_, _01479_, _06093_);
  and _23183_ (_01481_, _01480_, _01478_);
  and _23184_ (_01482_, _08999_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and _23185_ (_01483_, _01401_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  nor _23186_ (_01484_, _01401_, _07774_);
  or _23187_ (_01485_, _01484_, _01483_);
  and _23188_ (_01486_, _01485_, _05510_);
  or _23189_ (_01487_, _01486_, _01482_);
  or _23190_ (_01488_, _01487_, _01481_);
  and _23191_ (_00205_, _01488_, _04856_);
  or _23192_ (_01489_, _01401_, _06144_);
  or _23193_ (_01490_, _01361_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  and _23194_ (_01491_, _01490_, _06093_);
  and _23195_ (_01492_, _01491_, _01489_);
  and _23196_ (_01493_, _08999_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nand _23197_ (_01495_, _01361_, _07702_);
  and _23198_ (_01496_, _01495_, _05510_);
  and _23199_ (_01497_, _01496_, _01490_);
  or _23200_ (_01498_, _01497_, _01493_);
  or _23201_ (_01499_, _01498_, _01492_);
  and _23202_ (_00209_, _01499_, _04856_);
  nor _23203_ (_01500_, _06346_, rst);
  or _23204_ (_01501_, _06338_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  nand _23205_ (_01502_, _06338_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  and _23206_ (_01503_, _01502_, _01501_);
  and _23207_ (_00307_, _01503_, _01500_);
  and _23208_ (_01504_, _06721_, \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  or _23209_ (_01505_, _12825_, _06872_);
  or _23210_ (_01506_, _12697_, _08209_);
  or _23211_ (_01507_, _01506_, _01505_);
  or _23212_ (_01509_, _00298_, _06878_);
  or _23213_ (_01510_, _01509_, _01507_);
  or _23214_ (_01511_, _12693_, _08249_);
  or _23215_ (_01512_, _01511_, _01510_);
  and _23216_ (_01513_, _01512_, _06770_);
  or _23217_ (_00498_, _01513_, _01504_);
  and _23218_ (_01514_, _06410_, _05675_);
  and _23219_ (_01515_, _06046_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  or _23220_ (_01516_, _01515_, _05673_);
  or _23221_ (_01518_, _01516_, _01514_);
  or _23222_ (_01519_, _04861_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  and _23223_ (_01520_, _01519_, _04856_);
  and _23224_ (_00574_, _01520_, _01518_);
  and _23225_ (_01521_, _07176_, _07228_);
  and _23226_ (_01522_, _01521_, _07499_);
  and _23227_ (_01523_, _01522_, _06661_);
  nor _23228_ (_01524_, _01523_, _12477_);
  and _23229_ (_01525_, _07445_, _06410_);
  and _23230_ (_01526_, _07074_, _05288_);
  or _23231_ (_01527_, _01526_, _01525_);
  and _23232_ (_01528_, _01527_, _07406_);
  and _23233_ (_01529_, _07406_, _05718_);
  and _23234_ (_01530_, _07127_, _06033_);
  or _23235_ (_01531_, _01530_, _01529_);
  and _23236_ (_01532_, _01531_, _07461_);
  and _23237_ (_01533_, _07127_, _05670_);
  and _23238_ (_01534_, _07406_, _09282_);
  or _23239_ (_01535_, _01534_, _01533_);
  and _23240_ (_01536_, _01535_, _07452_);
  or _23241_ (_01537_, _01536_, _01532_);
  and _23242_ (_01538_, _07445_, _06997_);
  and _23243_ (_01539_, _07074_, _06705_);
  or _23244_ (_01540_, _01539_, _01538_);
  and _23245_ (_01541_, _01540_, _07127_);
  or _23246_ (_01542_, _01541_, _01537_);
  nor _23247_ (_01543_, _01542_, _01528_);
  nor _23248_ (_01544_, _01543_, _01524_);
  or _23249_ (_01545_, _07394_, _07228_);
  or _23250_ (_01546_, _01545_, _07402_);
  or _23251_ (_01548_, _07939_, _07406_);
  or _23252_ (_01549_, _07127_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and _23253_ (_01550_, _01549_, _07445_);
  and _23254_ (_01551_, _01550_, _01548_);
  and _23255_ (_01552_, _07127_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  and _23256_ (_01553_, _07406_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  or _23257_ (_01554_, _01553_, _01552_);
  and _23258_ (_01555_, _01554_, _07074_);
  or _23259_ (_01556_, _07127_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  or _23260_ (_01558_, _07406_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and _23261_ (_01560_, _01558_, _07461_);
  and _23262_ (_01561_, _01560_, _01556_);
  or _23263_ (_01562_, _07406_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  or _23264_ (_01564_, _07127_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  and _23265_ (_01565_, _01564_, _07452_);
  and _23266_ (_01566_, _01565_, _01562_);
  or _23267_ (_01567_, _01566_, _01561_);
  or _23268_ (_01568_, _01567_, _01555_);
  nor _23269_ (_01569_, _01568_, _01551_);
  nor _23270_ (_01571_, _01569_, _01546_);
  or _23271_ (_01572_, _07399_, _07398_);
  or _23272_ (_01573_, _07337_, _07176_);
  or _23273_ (_01574_, _01573_, _07400_);
  or _23274_ (_01575_, _01574_, _01572_);
  and _23275_ (_01576_, _07127_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and _23276_ (_01577_, _07406_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  or _23277_ (_01578_, _01577_, _01576_);
  and _23278_ (_01579_, _01578_, _07452_);
  or _23279_ (_01581_, _07127_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or _23280_ (_01582_, _07406_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and _23281_ (_01584_, _01582_, _07074_);
  and _23282_ (_01585_, _01584_, _01581_);
  and _23283_ (_01587_, _07406_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and _23284_ (_01588_, _07127_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  or _23285_ (_01589_, _01588_, _01587_);
  and _23286_ (_01590_, _01589_, _07445_);
  or _23287_ (_01591_, _07406_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or _23288_ (_01592_, _07127_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and _23289_ (_01594_, _01592_, _07461_);
  and _23290_ (_01595_, _01594_, _01591_);
  or _23291_ (_01596_, _01595_, _01590_);
  or _23292_ (_01598_, _01596_, _01585_);
  nor _23293_ (_01600_, _01598_, _01579_);
  nor _23294_ (_01601_, _01600_, _01575_);
  nand _23295_ (_01602_, _07482_, _07176_);
  and _23296_ (_01603_, _08841_, _07127_);
  or _23297_ (_01604_, _07531_, p1_in[7]);
  or _23298_ (_01605_, _07533_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and _23299_ (_01606_, _01605_, _01604_);
  and _23300_ (_01607_, _01606_, _07406_);
  or _23301_ (_01608_, _01607_, _01603_);
  and _23302_ (_01609_, _01608_, _07452_);
  or _23303_ (_01610_, _08940_, _07406_);
  or _23304_ (_01611_, _07531_, p1_in[6]);
  or _23305_ (_01612_, _07533_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and _23306_ (_01613_, _01612_, _01611_);
  or _23307_ (_01614_, _01613_, _07127_);
  and _23308_ (_01615_, _01614_, _07074_);
  and _23309_ (_01616_, _01615_, _01610_);
  or _23310_ (_01617_, _07531_, p1_in[4]);
  or _23311_ (_01618_, _07533_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and _23312_ (_01619_, _01618_, _01617_);
  and _23313_ (_01620_, _01619_, _07406_);
  and _23314_ (_01621_, _07555_, _07127_);
  or _23315_ (_01622_, _01621_, _01620_);
  and _23316_ (_01623_, _01622_, _07445_);
  nor _23317_ (_01624_, _07531_, p1_in[1]);
  not _23318_ (_01625_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and _23319_ (_01626_, _07531_, _01625_);
  nor _23320_ (_01627_, _01626_, _01624_);
  or _23321_ (_01628_, _01627_, _07406_);
  nor _23322_ (_01629_, _07531_, p1_in[5]);
  not _23323_ (_01630_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and _23324_ (_01631_, _07531_, _01630_);
  nor _23325_ (_01632_, _01631_, _01629_);
  or _23326_ (_01633_, _01632_, _07127_);
  and _23327_ (_01634_, _01633_, _07461_);
  and _23328_ (_01635_, _01634_, _01628_);
  or _23329_ (_01636_, _01635_, _01623_);
  or _23330_ (_01637_, _01636_, _01616_);
  nor _23331_ (_01638_, _01637_, _01609_);
  nor _23332_ (_01639_, _01638_, _01602_);
  and _23333_ (_01640_, _07394_, _07398_);
  and _23334_ (_01641_, _07127_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and _23335_ (_01642_, _07406_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  or _23336_ (_01643_, _01642_, _01641_);
  and _23337_ (_01645_, _01643_, _07461_);
  and _23338_ (_01646_, _07406_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and _23339_ (_01647_, _07127_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  or _23340_ (_01648_, _01647_, _01646_);
  and _23341_ (_01649_, _01648_, _07452_);
  or _23342_ (_01650_, _01649_, _01645_);
  and _23343_ (_01651_, _07406_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and _23344_ (_01652_, _07127_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  or _23345_ (_01653_, _01652_, _01651_);
  and _23346_ (_01654_, _01653_, _07445_);
  and _23347_ (_01655_, _07127_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and _23348_ (_01656_, _07406_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  or _23349_ (_01657_, _01656_, _01655_);
  and _23350_ (_01658_, _01657_, _07074_);
  or _23351_ (_01659_, _01658_, _01654_);
  or _23352_ (_01660_, _01659_, _01650_);
  and _23353_ (_01661_, _01660_, _07447_);
  and _23354_ (_01662_, _07127_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  and _23355_ (_01663_, _07406_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  or _23356_ (_01664_, _01663_, _01662_);
  and _23357_ (_01665_, _01664_, _07461_);
  and _23358_ (_01666_, _07406_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  and _23359_ (_01667_, _07127_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  or _23360_ (_01668_, _01667_, _01666_);
  and _23361_ (_01670_, _01668_, _07452_);
  or _23362_ (_01671_, _01670_, _01665_);
  and _23363_ (_01672_, _07406_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and _23364_ (_01673_, _07127_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or _23365_ (_01674_, _01673_, _01672_);
  and _23366_ (_01675_, _01674_, _07445_);
  and _23367_ (_01676_, _07127_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  and _23368_ (_01677_, _07406_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  or _23369_ (_01678_, _01677_, _01676_);
  and _23370_ (_01679_, _01678_, _07074_);
  or _23371_ (_01680_, _01679_, _01675_);
  or _23372_ (_01681_, _01680_, _01671_);
  and _23373_ (_01682_, _01681_, _07386_);
  or _23374_ (_01683_, _01682_, _01661_);
  and _23375_ (_01684_, _01683_, _01640_);
  or _23376_ (_01685_, _01684_, _01639_);
  or _23377_ (_01686_, _01685_, _01601_);
  or _23378_ (_01687_, _07401_, _07279_);
  or _23379_ (_01688_, _01545_, _01687_);
  and _23380_ (_01689_, _07127_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and _23381_ (_01690_, _07406_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  or _23382_ (_01691_, _01690_, _01689_);
  and _23383_ (_01692_, _01691_, _07452_);
  or _23384_ (_01693_, _07127_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  or _23385_ (_01694_, _07406_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and _23386_ (_01695_, _01694_, _07074_);
  and _23387_ (_01696_, _01695_, _01693_);
  and _23388_ (_01697_, _07406_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and _23389_ (_01698_, _07127_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  or _23390_ (_01699_, _01698_, _01697_);
  and _23391_ (_01700_, _01699_, _07445_);
  or _23392_ (_01701_, _07406_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  or _23393_ (_01702_, _07127_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and _23394_ (_01703_, _01702_, _07461_);
  and _23395_ (_01704_, _01703_, _01701_);
  or _23396_ (_01705_, _01704_, _01700_);
  or _23397_ (_01706_, _01705_, _01696_);
  nor _23398_ (_01707_, _01706_, _01692_);
  nor _23399_ (_01708_, _01707_, _01688_);
  or _23400_ (_01709_, _07991_, _04858_);
  and _23401_ (_01711_, _01688_, _01602_);
  nand _23402_ (_01712_, _07447_, _07176_);
  and _23403_ (_01713_, _01712_, _01575_);
  and _23404_ (_01714_, _01713_, _01711_);
  not _23405_ (_01715_, _01546_);
  nor _23406_ (_01716_, _01715_, _01522_);
  and _23407_ (_01717_, _01521_, _07386_);
  nand _23408_ (_01718_, _07385_, _07394_);
  nand _23409_ (_01719_, _01718_, \oc8051_top_1.oc8051_sfr1.bit_out );
  nor _23410_ (_01720_, _01719_, _01717_);
  and _23411_ (_01721_, _01720_, _01716_);
  nand _23412_ (_01722_, _01721_, _01714_);
  nand _23413_ (_01723_, _01722_, _01709_);
  or _23414_ (_01724_, _01723_, _01708_);
  and _23415_ (_01725_, _08836_, _07452_);
  nor _23416_ (_01726_, _07531_, p0_in[1]);
  not _23417_ (_01727_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and _23418_ (_01728_, _07531_, _01727_);
  nor _23419_ (_01729_, _01728_, _01726_);
  and _23420_ (_01730_, _01729_, _07461_);
  or _23421_ (_01731_, _01730_, _07406_);
  or _23422_ (_01732_, _01731_, _01725_);
  or _23423_ (_01733_, _07531_, p0_in[7]);
  or _23424_ (_01734_, _07533_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and _23425_ (_01735_, _01734_, _01733_);
  and _23426_ (_01736_, _01735_, _07452_);
  nor _23427_ (_01737_, _07531_, p0_in[5]);
  not _23428_ (_01738_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and _23429_ (_01739_, _07531_, _01738_);
  nor _23430_ (_01740_, _01739_, _01737_);
  and _23431_ (_01741_, _01740_, _07461_);
  or _23432_ (_01742_, _01741_, _07127_);
  or _23433_ (_01743_, _01742_, _01736_);
  and _23434_ (_01744_, _01743_, _01732_);
  or _23435_ (_01745_, _07531_, p0_in[6]);
  or _23436_ (_01746_, _07533_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and _23437_ (_01747_, _01746_, _01745_);
  and _23438_ (_01748_, _01747_, _07406_);
  and _23439_ (_01749_, _08944_, _07127_);
  or _23440_ (_01750_, _01749_, _01748_);
  and _23441_ (_01751_, _01750_, _07074_);
  or _23442_ (_01752_, _07531_, p0_in[4]);
  or _23443_ (_01753_, _07533_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and _23444_ (_01754_, _01753_, _01752_);
  and _23445_ (_01755_, _01754_, _07406_);
  and _23446_ (_01756_, _07550_, _07127_);
  or _23447_ (_01757_, _01756_, _01755_);
  and _23448_ (_01758_, _01757_, _07445_);
  or _23449_ (_01759_, _01758_, _01751_);
  or _23450_ (_01760_, _01759_, _01744_);
  and _23451_ (_01761_, _01760_, _01717_);
  and _23452_ (_01762_, _07127_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and _23453_ (_01763_, _07406_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or _23454_ (_01764_, _01763_, _01762_);
  and _23455_ (_01765_, _01764_, _07452_);
  or _23456_ (_01766_, _07127_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or _23457_ (_01767_, _07406_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and _23458_ (_01768_, _01767_, _07074_);
  and _23459_ (_01769_, _01768_, _01766_);
  and _23460_ (_01770_, _07406_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and _23461_ (_01771_, _07127_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or _23462_ (_01772_, _01771_, _01770_);
  and _23463_ (_01773_, _01772_, _07445_);
  or _23464_ (_01774_, _07406_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or _23465_ (_01775_, _07127_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and _23466_ (_01777_, _01775_, _07461_);
  and _23467_ (_01778_, _01777_, _01774_);
  or _23468_ (_01779_, _01778_, _01773_);
  or _23469_ (_01780_, _01779_, _01769_);
  or _23470_ (_01781_, _01780_, _01765_);
  and _23471_ (_01782_, _01781_, _01522_);
  or _23472_ (_01783_, _01782_, _01761_);
  or _23473_ (_01784_, _01783_, _01724_);
  or _23474_ (_01786_, _01784_, _01686_);
  and _23475_ (_01787_, _07406_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and _23476_ (_01788_, _07127_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  or _23477_ (_01789_, _01788_, _01787_);
  and _23478_ (_01790_, _01789_, _07445_);
  or _23479_ (_01792_, _07406_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or _23480_ (_01793_, _07127_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and _23481_ (_01795_, _01793_, _07461_);
  and _23482_ (_01797_, _01795_, _01792_);
  or _23483_ (_01798_, _01797_, _01790_);
  and _23484_ (_01800_, _07127_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and _23485_ (_01802_, _07406_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or _23486_ (_01804_, _01802_, _01800_);
  and _23487_ (_01806_, _01804_, _07074_);
  or _23488_ (_01807_, _07127_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or _23489_ (_01809_, _07406_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and _23490_ (_01810_, _01809_, _07452_);
  and _23491_ (_01811_, _01810_, _01807_);
  or _23492_ (_01813_, _01811_, _01806_);
  or _23493_ (_01814_, _01813_, _01798_);
  and _23494_ (_01815_, _01814_, _07387_);
  and _23495_ (_01816_, _07406_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  and _23496_ (_01818_, _07127_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  or _23497_ (_01819_, _01818_, _01816_);
  and _23498_ (_01820_, _01819_, _07445_);
  or _23499_ (_01821_, _07406_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  or _23500_ (_01822_, _07127_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and _23501_ (_01823_, _01822_, _07461_);
  and _23502_ (_01825_, _01823_, _01821_);
  or _23503_ (_01826_, _01825_, _01820_);
  and _23504_ (_01827_, _07127_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and _23505_ (_01828_, _07406_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  or _23506_ (_01830_, _01828_, _01827_);
  and _23507_ (_01831_, _01830_, _07074_);
  or _23508_ (_01832_, _07127_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  or _23509_ (_01833_, _07406_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and _23510_ (_01834_, _01833_, _07452_);
  and _23511_ (_01835_, _01834_, _01832_);
  or _23512_ (_01836_, _01835_, _01831_);
  or _23513_ (_01837_, _01836_, _01826_);
  and _23514_ (_01838_, _01837_, _07448_);
  or _23515_ (_01839_, _01838_, _01815_);
  and _23516_ (_01840_, _01839_, _07394_);
  and _23517_ (_01841_, _08953_, _07127_);
  or _23518_ (_01842_, _07531_, p2_in[6]);
  or _23519_ (_01843_, _07533_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and _23520_ (_01844_, _01843_, _01842_);
  and _23521_ (_01845_, _01844_, _07406_);
  or _23522_ (_01847_, _01845_, _01841_);
  and _23523_ (_01848_, _01847_, _07074_);
  nor _23524_ (_01850_, _07531_, p2_in[5]);
  not _23525_ (_01852_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and _23526_ (_01854_, _07531_, _01852_);
  nor _23527_ (_01855_, _01854_, _01850_);
  or _23528_ (_01857_, _01855_, _07127_);
  nor _23529_ (_01858_, _07531_, p2_in[1]);
  not _23530_ (_01860_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and _23531_ (_01861_, _07531_, _01860_);
  nor _23532_ (_01862_, _01861_, _01858_);
  or _23533_ (_01863_, _01862_, _07406_);
  and _23534_ (_01864_, _01863_, _07461_);
  and _23535_ (_01865_, _01864_, _01857_);
  or _23536_ (_01866_, _01865_, _01848_);
  or _23537_ (_01867_, _07531_, p2_in[4]);
  or _23538_ (_01868_, _07533_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and _23539_ (_01869_, _01868_, _01867_);
  and _23540_ (_01870_, _01869_, _07406_);
  and _23541_ (_01871_, _07536_, _07127_);
  or _23542_ (_01872_, _01871_, _01870_);
  and _23543_ (_01873_, _01872_, _07445_);
  or _23544_ (_01874_, _08847_, _07406_);
  or _23545_ (_01875_, _07531_, p2_in[7]);
  or _23546_ (_01876_, _07533_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and _23547_ (_01877_, _01876_, _01875_);
  or _23548_ (_01878_, _01877_, _07127_);
  and _23549_ (_01879_, _01878_, _07452_);
  and _23550_ (_01880_, _01879_, _01874_);
  or _23551_ (_01881_, _01880_, _01873_);
  or _23552_ (_01882_, _01881_, _01866_);
  and _23553_ (_01883_, _01882_, _07228_);
  nor _23554_ (_01885_, _07531_, p3_in[1]);
  not _23555_ (_01886_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and _23556_ (_01887_, _07531_, _01886_);
  nor _23557_ (_01888_, _01887_, _01885_);
  and _23558_ (_01889_, _01888_, _07127_);
  nor _23559_ (_01890_, _07531_, p3_in[5]);
  not _23560_ (_01891_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and _23561_ (_01892_, _07531_, _01891_);
  nor _23562_ (_01893_, _01892_, _01890_);
  and _23563_ (_01894_, _01893_, _07406_);
  or _23564_ (_01895_, _01894_, _01889_);
  and _23565_ (_01896_, _01895_, _07461_);
  or _23566_ (_01897_, _07531_, p3_in[4]);
  or _23567_ (_01898_, _07533_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and _23568_ (_01899_, _01898_, _01897_);
  or _23569_ (_01900_, _01899_, _07127_);
  or _23570_ (_01901_, _07544_, _07406_);
  and _23571_ (_01902_, _01901_, _07445_);
  and _23572_ (_01904_, _01902_, _01900_);
  or _23573_ (_01905_, _01904_, _01896_);
  or _23574_ (_01906_, _07531_, p3_in[6]);
  or _23575_ (_01907_, _07533_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and _23576_ (_01908_, _01907_, _01906_);
  and _23577_ (_01909_, _01908_, _07406_);
  and _23578_ (_01910_, _08949_, _07127_);
  or _23579_ (_01911_, _01910_, _01909_);
  and _23580_ (_01912_, _01911_, _07074_);
  or _23581_ (_01913_, _08852_, _07406_);
  or _23582_ (_01914_, _07531_, p3_in[7]);
  or _23583_ (_01915_, _07533_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and _23584_ (_01916_, _01915_, _01914_);
  or _23585_ (_01917_, _01916_, _07127_);
  and _23586_ (_01918_, _01917_, _07452_);
  and _23587_ (_01919_, _01918_, _01913_);
  or _23588_ (_01921_, _01919_, _01912_);
  or _23589_ (_01922_, _01921_, _01905_);
  and _23590_ (_01923_, _01922_, _07398_);
  nor _23591_ (_01925_, _01923_, _01883_);
  nor _23592_ (_01926_, _01925_, _01712_);
  or _23593_ (_01927_, _01926_, _01840_);
  or _23594_ (_01928_, _01927_, _01786_);
  or _23595_ (_01929_, _01928_, _01571_);
  or _23596_ (_01930_, _01709_, _06144_);
  and _23597_ (_01932_, _01930_, _01524_);
  and _23598_ (_01933_, _01932_, _01929_);
  or _23599_ (_01934_, _01933_, _01544_);
  and _23600_ (_00670_, _01934_, _04856_);
  and _23601_ (_01935_, _09254_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and _23602_ (_01936_, _01935_, _08063_);
  and _23603_ (_01937_, _09253_, _01936_);
  or _23604_ (_01938_, _01937_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0]);
  not _23605_ (_01939_, rxd_i);
  nand _23606_ (_01940_, _01937_, _01939_);
  and _23607_ (_01941_, _01940_, _04856_);
  and _23608_ (_00865_, _01941_, _01938_);
  or _23609_ (_01942_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  or _23610_ (_01944_, _01942_, _12219_);
  not _23611_ (_01945_, _06268_);
  nand _23612_ (_01946_, _01945_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  nand _23613_ (_01947_, _01946_, _12177_);
  or _23614_ (_01948_, _01947_, _06657_);
  and _23615_ (_01949_, _01948_, _01944_);
  or _23616_ (_01950_, _01949_, _12183_);
  nand _23617_ (_01951_, _12183_, _06284_);
  and _23618_ (_01952_, _01951_, _04856_);
  and _23619_ (_01020_, _01952_, _01950_);
  nor _23620_ (_01954_, _12453_, _12220_);
  not _23621_ (_01956_, _12391_);
  nor _23622_ (_01957_, _12393_, _01956_);
  and _23623_ (_01958_, _01957_, _12401_);
  and _23624_ (_01959_, _01958_, _12420_);
  and _23625_ (_01961_, _01959_, _12453_);
  or _23626_ (_01963_, _01961_, _01954_);
  and _23627_ (_01023_, _01963_, _04856_);
  and _23628_ (_01965_, _12401_, _01956_);
  and _23629_ (_01966_, _01965_, _12453_);
  not _23630_ (_01967_, _01966_);
  or _23631_ (_01968_, _01967_, _12420_);
  or _23632_ (_01969_, _01966_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  and _23633_ (_01970_, _01969_, _04856_);
  and _23634_ (_01031_, _01970_, _01968_);
  and _23635_ (_01971_, _05674_, _04861_);
  and _23636_ (_01972_, _01971_, _05718_);
  not _23637_ (_01973_, _01971_);
  and _23638_ (_01974_, _01973_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  or _23639_ (_01975_, _01974_, _01972_);
  and _23640_ (_01037_, _01975_, _04856_);
  nand _23641_ (_01976_, _12389_, _06284_);
  and _23642_ (_01977_, _12393_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  not _23643_ (_01978_, _01977_);
  and _23644_ (_01979_, _01978_, _12416_);
  nor _23645_ (_01980_, _01979_, _12430_);
  or _23646_ (_01981_, _01980_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  nand _23647_ (_01982_, _12422_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  and _23648_ (_01983_, _01982_, _12401_);
  nand _23649_ (_01984_, _01983_, _12420_);
  and _23650_ (_01985_, _01984_, _12395_);
  or _23651_ (_01986_, _01985_, _01977_);
  or _23652_ (_01987_, _01986_, _12430_);
  and _23653_ (_01988_, _01987_, _01981_);
  or _23654_ (_01989_, _01988_, _12389_);
  and _23655_ (_01990_, _01989_, _04856_);
  and _23656_ (_01040_, _01990_, _01976_);
  nand _23657_ (_01991_, _12430_, _06284_);
  and _23658_ (_01992_, _12393_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  nor _23659_ (_01993_, _12602_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  nor _23660_ (_01994_, _01993_, _12553_);
  and _23661_ (_01995_, _12423_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and _23662_ (_01996_, _01995_, _12420_);
  or _23663_ (_01997_, _01996_, _01994_);
  and _23664_ (_01998_, _01997_, _12395_);
  nor _23665_ (_01999_, _01998_, _01992_);
  nand _23666_ (_02000_, _01999_, _12431_);
  and _23667_ (_02001_, _02000_, _12390_);
  and _23668_ (_02002_, _02001_, _01991_);
  and _23669_ (_02003_, _12389_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or _23670_ (_02004_, _02003_, _02002_);
  and _23671_ (_01044_, _02004_, _04856_);
  or _23672_ (_02005_, _09251_, _08065_);
  or _23673_ (_02006_, _09253_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and _23674_ (_02007_, _02006_, _04856_);
  and _23675_ (_01051_, _02007_, _02005_);
  nand _23676_ (_02008_, _12714_, _06284_);
  and _23677_ (_02009_, _12735_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  and _23678_ (_02010_, _12720_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  or _23679_ (_02011_, _02010_, _02009_);
  or _23680_ (_02012_, _02011_, _12714_);
  and _23681_ (_02013_, _02012_, _04856_);
  and _23682_ (_01066_, _02013_, _02008_);
  nor _23683_ (_01110_, _07927_, rst);
  and _23684_ (_01112_, _07573_, _04856_);
  and _23685_ (_01115_, _07862_, _04856_);
  nor _23686_ (_01147_, _07712_, rst);
  and _23687_ (_02014_, _06238_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  not _23688_ (_02015_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nor _23689_ (_02017_, _06238_, _02015_);
  or _23690_ (_02018_, _02017_, _02014_);
  and _23691_ (_01154_, _02018_, _04856_);
  and _23692_ (_02019_, _06238_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  not _23693_ (_02020_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor _23694_ (_02021_, _06238_, _02020_);
  or _23695_ (_02023_, _02021_, _02019_);
  and _23696_ (_01158_, _02023_, _04856_);
  and _23697_ (_01317_, _07780_, _04856_);
  nand _23698_ (_02024_, _12719_, _06284_);
  and _23699_ (_02025_, _12717_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and _23700_ (_02026_, _12716_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or _23701_ (_02027_, _02026_, _02025_);
  or _23702_ (_02028_, _02027_, _12719_);
  and _23703_ (_02029_, _02028_, _12715_);
  and _23704_ (_02030_, _02029_, _02024_);
  and _23705_ (_02031_, _12714_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  or _23706_ (_02032_, _02031_, _02030_);
  and _23707_ (_01397_, _02032_, _04856_);
  and _23708_ (_01406_, t2ex_i, _04856_);
  nor _23709_ (_02033_, t2ex_i, rst);
  and _23710_ (_01412_, _02033_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r );
  nor _23711_ (_02034_, t2_i, rst);
  and _23712_ (_01415_, _02034_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r );
  or _23713_ (_02035_, _06238_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nand _23714_ (_02037_, _06238_, _05089_);
  and _23715_ (_02038_, _02037_, _04856_);
  and _23716_ (_01427_, _02038_, _02035_);
  and _23717_ (_02039_, _09282_, _05671_);
  and _23718_ (_02040_, _06696_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  or _23719_ (_02041_, _02040_, _02039_);
  and _23720_ (_01437_, _02041_, _04856_);
  and _23721_ (_01494_, t2_i, _04856_);
  and _23722_ (_02043_, _09251_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  not _23723_ (_02044_, _08062_);
  nor _23724_ (_02045_, _01935_, _02044_);
  or _23725_ (_02046_, _02045_, _02043_);
  and _23726_ (_02047_, _09254_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _23727_ (_02048_, _02047_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and _23728_ (_02050_, _02048_, _04856_);
  and _23729_ (_01508_, _02050_, _02046_);
  and _23730_ (_02051_, _08057_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  and _23731_ (_02052_, _08085_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  or _23732_ (_01557_, _02052_, _02051_);
  and _23733_ (_02053_, _06297_, _07855_);
  nand _23734_ (_02055_, _02053_, _06088_);
  or _23735_ (_02056_, _02053_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and _23736_ (_02057_, _02056_, _06305_);
  and _23737_ (_02058_, _02057_, _02055_);
  and _23738_ (_02059_, _06410_, _06304_);
  or _23739_ (_02060_, _02059_, _02058_);
  and _23740_ (_01559_, _02060_, _04856_);
  and _23741_ (_02061_, _06297_, _04986_);
  nand _23742_ (_02063_, _02061_, _06088_);
  or _23743_ (_02064_, _02061_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and _23744_ (_02065_, _02064_, _06305_);
  and _23745_ (_02066_, _02065_, _02063_);
  nor _23746_ (_02067_, _06305_, _06032_);
  or _23747_ (_02068_, _02067_, _02066_);
  and _23748_ (_01563_, _02068_, _04856_);
  and _23749_ (_02069_, _06270_, _07855_);
  or _23750_ (_02070_, _02069_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  and _23751_ (_02071_, _02070_, _06276_);
  nand _23752_ (_02073_, _02069_, _06088_);
  and _23753_ (_02074_, _02073_, _02071_);
  and _23754_ (_02075_, _06410_, _06275_);
  or _23755_ (_02076_, _02075_, _02074_);
  and _23756_ (_01570_, _02076_, _04856_);
  and _23757_ (_02077_, _06270_, _04986_);
  or _23758_ (_02078_, _02077_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and _23759_ (_02079_, _02078_, _06276_);
  nand _23760_ (_02080_, _02077_, _06088_);
  and _23761_ (_02081_, _02080_, _02079_);
  nor _23762_ (_02083_, _06276_, _06032_);
  or _23763_ (_02084_, _02083_, _02081_);
  and _23764_ (_01580_, _02084_, _04856_);
  and _23765_ (_02085_, _08085_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  or _23766_ (_01583_, _02085_, _08058_);
  or _23767_ (_02086_, _12716_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  not _23768_ (_02087_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  nand _23769_ (_02088_, _12716_, _02087_);
  and _23770_ (_02089_, _02088_, _02086_);
  or _23771_ (_02090_, _02089_, _12719_);
  nand _23772_ (_02092_, _12719_, _06032_);
  and _23773_ (_02093_, _02092_, _02090_);
  or _23774_ (_02094_, _02093_, _12714_);
  not _23775_ (_02095_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  nand _23776_ (_02096_, _12714_, _02095_);
  and _23777_ (_02097_, _02096_, _04856_);
  and _23778_ (_01586_, _02097_, _02094_);
  not _23779_ (_02098_, _06225_);
  nor _23780_ (_02099_, _02098_, _06202_);
  nand _23781_ (_02100_, _06249_, _02099_);
  and _23782_ (_02101_, _06249_, _06202_);
  or _23783_ (_02102_, _02101_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0]);
  and _23784_ (_02103_, _02102_, _04856_);
  and _23785_ (_01593_, _02103_, _02100_);
  nand _23786_ (_02104_, _06288_, _02099_);
  and _23787_ (_02105_, _06288_, _06202_);
  or _23788_ (_02106_, _02105_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0]);
  and _23789_ (_02107_, _02106_, _04856_);
  and _23790_ (_01597_, _02107_, _02104_);
  or _23791_ (_02108_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or _23792_ (_02109_, _02108_, _06206_);
  not _23793_ (_02110_, _06208_);
  or _23794_ (_02111_, _02110_, _06105_);
  not _23795_ (_02112_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  and _23796_ (_02113_, _06218_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or _23797_ (_02114_, _02113_, _02112_);
  and _23798_ (_02115_, _06216_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _23799_ (_02116_, _02115_, _06221_);
  nand _23800_ (_02117_, _02116_, _02114_);
  not _23801_ (_02118_, _06210_);
  or _23802_ (_02119_, _06222_, _06105_);
  and _23803_ (_02120_, _02119_, _02118_);
  and _23804_ (_02121_, _02120_, _02117_);
  and _23805_ (_02122_, _02108_, _06210_);
  or _23806_ (_02123_, _02122_, _06208_);
  or _23807_ (_02124_, _02123_, _02121_);
  and _23808_ (_02125_, _02124_, _02111_);
  or _23809_ (_02126_, _02125_, _06205_);
  nand _23810_ (_02127_, _02126_, _02109_);
  nand _23811_ (_02128_, _02127_, _02099_);
  and _23812_ (_02129_, _06194_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or _23813_ (_02130_, _02129_, _02112_);
  nor _23814_ (_02131_, _06190_, _06104_);
  nor _23815_ (_02132_, _02131_, _06198_);
  nand _23816_ (_02133_, _02132_, _02130_);
  or _23817_ (_02134_, _06199_, _06105_);
  and _23818_ (_02135_, _02134_, _02133_);
  or _23819_ (_02136_, _02135_, _06184_);
  not _23820_ (_02138_, _06182_);
  not _23821_ (_02139_, _06184_);
  or _23822_ (_02140_, _02108_, _02139_);
  and _23823_ (_02141_, _02140_, _02138_);
  and _23824_ (_02142_, _02141_, _02136_);
  and _23825_ (_02143_, _06182_, _06105_);
  or _23826_ (_02144_, _02143_, _06179_);
  or _23827_ (_02145_, _02144_, _02142_);
  or _23828_ (_02146_, _02108_, _06180_);
  and _23829_ (_02147_, _02146_, _02145_);
  or _23830_ (_02148_, _02147_, _06228_);
  and _23831_ (_02149_, _02148_, _02128_);
  or _23832_ (_02150_, _02149_, _06172_);
  nor _23833_ (_02151_, _06172_, _06226_);
  or _23834_ (_02152_, _02151_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  and _23835_ (_02153_, _02152_, _04856_);
  and _23836_ (_01599_, _02153_, _02150_);
  not _23837_ (_02154_, _05994_);
  and _23838_ (_02155_, _06859_, _02154_);
  or _23839_ (_02156_, _06872_, _06856_);
  or _23840_ (_02157_, _02156_, _06616_);
  or _23841_ (_02158_, _12685_, _06878_);
  or _23842_ (_02160_, _02158_, _12688_);
  or _23843_ (_02161_, _02160_, _02157_);
  and _23844_ (_02162_, _02161_, _05962_);
  or _23845_ (_02163_, _02162_, _02155_);
  and _23846_ (_01644_, _02163_, _04856_);
  and _23847_ (_02164_, _01973_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  and _23848_ (_02165_, _01971_, _06033_);
  or _23849_ (_02166_, _02165_, _02164_);
  and _23850_ (_01776_, _02166_, _04856_);
  and _23851_ (_02167_, _08057_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  and _23852_ (_02168_, _08085_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  or _23853_ (_01785_, _02168_, _02167_);
  and _23854_ (_02169_, _08057_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  and _23855_ (_02170_, _08085_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  or _23856_ (_01791_, _02170_, _02169_);
  and _23857_ (_02171_, _08085_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  and _23858_ (_02172_, _08057_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  or _23859_ (_01794_, _02172_, _02171_);
  nor _23860_ (_02173_, _06218_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nor _23861_ (_02174_, _02173_, _06216_);
  or _23862_ (_02175_, _02174_, _06221_);
  and _23863_ (_02176_, _02175_, _02118_);
  or _23864_ (_02177_, _02176_, _06208_);
  and _23865_ (_02178_, _02099_, _06206_);
  and _23866_ (_02179_, _02178_, _02177_);
  or _23867_ (_02180_, _06194_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and _23868_ (_02181_, _02180_, _06190_);
  or _23869_ (_02182_, _02181_, _06198_);
  and _23870_ (_02183_, _02182_, _02139_);
  or _23871_ (_02184_, _02183_, _06182_);
  and _23872_ (_02185_, _06202_, _06180_);
  and _23873_ (_02186_, _02185_, _02184_);
  or _23874_ (_02187_, _02186_, _06172_);
  or _23875_ (_02188_, _02187_, _02179_);
  nand _23876_ (_02189_, _06172_, _12199_);
  and _23877_ (_02190_, _02189_, _04856_);
  and _23878_ (_01796_, _02190_, _02188_);
  and _23879_ (_02191_, _06297_, _06091_);
  and _23880_ (_02192_, _02191_, _06088_);
  nor _23881_ (_02193_, _02191_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  or _23882_ (_02194_, _02193_, _02192_);
  nand _23883_ (_02195_, _02194_, _06305_);
  or _23884_ (_02196_, _06305_, _05718_);
  and _23885_ (_02197_, _02196_, _04856_);
  and _23886_ (_01799_, _02197_, _02195_);
  and _23887_ (_02199_, _06270_, _06091_);
  or _23888_ (_02200_, _02199_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and _23889_ (_02201_, _02200_, _06276_);
  nand _23890_ (_02202_, _02199_, _06088_);
  and _23891_ (_02203_, _02202_, _02201_);
  and _23892_ (_02204_, _06275_, _05718_);
  or _23893_ (_02205_, _02204_, _02203_);
  and _23894_ (_01801_, _02205_, _04856_);
  and _23895_ (_02206_, _06136_, _04990_);
  or _23896_ (_02207_, _02206_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and _23897_ (_02209_, _02207_, _06129_);
  nand _23898_ (_02210_, _02206_, _06088_);
  and _23899_ (_02211_, _02210_, _02209_);
  and _23900_ (_02212_, _06997_, _06127_);
  or _23901_ (_02213_, _02212_, _02211_);
  and _23902_ (_01803_, _02213_, _04856_);
  nand _23903_ (_02214_, _10587_, _05287_);
  or _23904_ (_02215_, _10587_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  and _23905_ (_02216_, _02215_, _04856_);
  and _23906_ (_01805_, _02216_, _02214_);
  or _23907_ (_02217_, _06235_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and _23908_ (_02218_, _02217_, _04856_);
  or _23909_ (_02219_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and _23910_ (_02220_, _02219_, _06180_);
  or _23911_ (_02221_, _02220_, _06186_);
  and _23912_ (_02222_, _06198_, _06110_);
  or _23913_ (_02223_, _02129_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  nand _23914_ (_02225_, _02223_, _02132_);
  nand _23915_ (_02226_, _02225_, _06185_);
  or _23916_ (_02227_, _02226_, _02222_);
  and _23917_ (_02228_, _02227_, _02221_);
  and _23918_ (_02229_, _06179_, _06110_);
  or _23919_ (_02230_, _02229_, _02228_);
  and _23920_ (_02231_, _02230_, _06202_);
  and _23921_ (_02232_, _02098_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and _23922_ (_02233_, _06205_, _06110_);
  and _23923_ (_02234_, _02219_, _06206_);
  or _23924_ (_02236_, _02234_, _06212_);
  or _23925_ (_02237_, _02113_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and _23926_ (_02238_, _02237_, _02116_);
  nand _23927_ (_02240_, _06221_, _06110_);
  nand _23928_ (_02241_, _02240_, _06211_);
  or _23929_ (_02242_, _02241_, _02238_);
  and _23930_ (_02243_, _02242_, _02236_);
  or _23931_ (_02244_, _02243_, _02233_);
  and _23932_ (_02245_, _02244_, _06225_);
  or _23933_ (_02246_, _02245_, _02232_);
  and _23934_ (_02247_, _02246_, _06228_);
  or _23935_ (_02248_, _02247_, _02231_);
  or _23936_ (_02249_, _02248_, _06172_);
  and _23937_ (_01808_, _02249_, _02218_);
  and _23938_ (_02250_, _06238_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  not _23939_ (_02251_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor _23940_ (_02252_, _06238_, _02251_);
  or _23941_ (_02253_, _02252_, _02250_);
  and _23942_ (_01812_, _02253_, _04856_);
  or _23943_ (_02254_, _06221_, _06210_);
  and _23944_ (_02255_, _06219_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or _23945_ (_02256_, _02255_, _02254_);
  and _23946_ (_02257_, _02256_, _02110_);
  and _23947_ (_02258_, _02257_, _02178_);
  or _23948_ (_02259_, _06198_, _06184_);
  and _23949_ (_02260_, _06196_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or _23950_ (_02261_, _02260_, _02259_);
  and _23951_ (_02262_, _02261_, _02138_);
  and _23952_ (_02263_, _02262_, _02185_);
  or _23953_ (_02264_, _02263_, _06172_);
  or _23954_ (_02265_, _02264_, _02258_);
  or _23955_ (_02266_, _06235_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and _23956_ (_02267_, _02266_, _04856_);
  and _23957_ (_01817_, _02267_, _02265_);
  and _23958_ (_02268_, _01973_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  and _23959_ (_02269_, _06370_, _05674_);
  or _23960_ (_02270_, _02269_, _02268_);
  and _23961_ (_01824_, _02270_, _04856_);
  and _23962_ (_02271_, _08057_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  and _23963_ (_02272_, _08085_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  or _23964_ (_01829_, _02272_, _02271_);
  and _23965_ (_02273_, _06172_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  or _23966_ (_02274_, _02273_, _02151_);
  and _23967_ (_01846_, _02274_, _04856_);
  and _23968_ (_01849_, _13181_, _06172_);
  and _23969_ (_02275_, _06172_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  or _23970_ (_02276_, _02275_, _02151_);
  and _23971_ (_01851_, _02276_, _04856_);
  and _23972_ (_01853_, _13207_, _06172_);
  and _23973_ (_02277_, _06222_, _06212_);
  nand _23974_ (_02278_, _02277_, _06203_);
  or _23975_ (_02279_, _02278_, _06219_);
  nor _23976_ (_02280_, _02279_, _06202_);
  and _23977_ (_02281_, _06172_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  or _23978_ (_02282_, _06172_, _06198_);
  nor _23979_ (_02283_, _02282_, _06177_);
  not _23980_ (_02284_, _06186_);
  nor _23981_ (_02285_, _06196_, _02284_);
  and _23982_ (_02286_, _02285_, _02283_);
  or _23983_ (_02287_, _02286_, _02281_);
  or _23984_ (_02288_, _02287_, _02280_);
  and _23985_ (_01856_, _02288_, _04856_);
  nand _23986_ (_02289_, _06288_, _06226_);
  nor _23987_ (_02290_, _06172_, _06202_);
  or _23988_ (_02291_, _02290_, _06104_);
  and _23989_ (_02292_, _02291_, _04856_);
  and _23990_ (_01859_, _02292_, _02289_);
  or _23991_ (_02293_, _12395_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and _23992_ (_02294_, _12423_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and _23993_ (_02295_, _02294_, _12420_);
  nand _23994_ (_02296_, _12412_, _12401_);
  and _23995_ (_02297_, _02296_, _08794_);
  nor _23996_ (_02298_, _02297_, _12440_);
  or _23997_ (_02299_, _02298_, _12393_);
  or _23998_ (_02300_, _02299_, _02295_);
  nand _23999_ (_02301_, _02300_, _02293_);
  nor _24000_ (_02302_, _02301_, _12430_);
  and _24001_ (_02303_, _12430_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or _24002_ (_02304_, _02303_, _12389_);
  or _24003_ (_02305_, _02304_, _02302_);
  nand _24004_ (_02306_, _12389_, _05669_);
  and _24005_ (_02307_, _02306_, _04856_);
  and _24006_ (_01884_, _02307_, _02305_);
  and _24007_ (_02308_, _09259_, _06268_);
  nand _24008_ (_02309_, _02308_, _06088_);
  or _24009_ (_02310_, _02308_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  and _24010_ (_02311_, _02310_, _09264_);
  and _24011_ (_02312_, _02311_, _02309_);
  nor _24012_ (_02313_, _09264_, _06284_);
  or _24013_ (_02314_, _02313_, _02312_);
  and _24014_ (_01903_, _02314_, _04856_);
  or _24015_ (_02315_, _09200_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  and _24016_ (_02316_, _02315_, _04856_);
  nand _24017_ (_02317_, _09200_, _06284_);
  and _24018_ (_01920_, _02317_, _02316_);
  and _24019_ (_02318_, _04856_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  and _24020_ (_02319_, _02318_, _09206_);
  and _24021_ (_02320_, _09217_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  nor _24022_ (_02321_, _09206_, rst);
  and _24023_ (_02322_, _02321_, _02320_);
  or _24024_ (_01924_, _02322_, _02319_);
  not _24025_ (_02323_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and _24026_ (_02324_, _02323_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _24027_ (_02325_, _02324_, _06179_);
  nor _24028_ (_02326_, _02325_, _06186_);
  nand _24029_ (_02327_, _06198_, _06109_);
  nor _24030_ (_02328_, _06190_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or _24031_ (_02329_, _02328_, _06198_);
  nand _24032_ (_02330_, _06194_, _06104_);
  and _24033_ (_02331_, _02330_, _02323_);
  or _24034_ (_02332_, _02331_, _02329_);
  and _24035_ (_02333_, _02332_, _06185_);
  and _24036_ (_02334_, _02333_, _02327_);
  or _24037_ (_02335_, _02334_, _02326_);
  nand _24038_ (_02336_, _06179_, _06109_);
  and _24039_ (_02337_, _02336_, _02335_);
  nand _24040_ (_02338_, _02337_, _06202_);
  nor _24041_ (_02339_, _02324_, _06205_);
  or _24042_ (_02341_, _02339_, _06212_);
  and _24043_ (_02342_, _06218_, _06104_);
  or _24044_ (_02343_, _02342_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and _24045_ (_02344_, _06216_, _06104_);
  nor _24046_ (_02345_, _02344_, _06221_);
  and _24047_ (_02346_, _02345_, _02343_);
  nand _24048_ (_02347_, _06221_, _06109_);
  nand _24049_ (_02348_, _02347_, _06211_);
  or _24050_ (_02349_, _02348_, _02346_);
  and _24051_ (_02350_, _02349_, _02341_);
  and _24052_ (_02351_, _06205_, _06109_);
  or _24053_ (_02352_, _02351_, _06202_);
  or _24054_ (_02353_, _02352_, _02098_);
  or _24055_ (_02354_, _02353_, _02350_);
  and _24056_ (_02355_, _02354_, _02338_);
  or _24057_ (_02356_, _02355_, _06172_);
  or _24058_ (_02357_, _02151_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and _24059_ (_02358_, _02357_, _04856_);
  and _24060_ (_01931_, _02358_, _02356_);
  not _24061_ (_02359_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  nor _24062_ (_02360_, _02151_, _02359_);
  or _24063_ (_02361_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _06104_);
  or _24064_ (_02362_, _02361_, _06180_);
  and _24065_ (_02363_, _02362_, _06202_);
  and _24066_ (_02364_, _02330_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  or _24067_ (_02365_, _02364_, _02329_);
  or _24068_ (_02366_, _06199_, _06103_);
  and _24069_ (_02367_, _02366_, _02365_);
  or _24070_ (_02368_, _02367_, _06184_);
  or _24071_ (_02369_, _02361_, _02139_);
  and _24072_ (_02370_, _02369_, _02138_);
  and _24073_ (_02371_, _02370_, _02368_);
  and _24074_ (_02372_, _06182_, _06103_);
  or _24075_ (_02373_, _02372_, _06179_);
  or _24076_ (_02374_, _02373_, _02371_);
  and _24077_ (_02375_, _02374_, _02363_);
  or _24078_ (_02376_, _02342_, _02359_);
  nand _24079_ (_02377_, _02376_, _02345_);
  or _24080_ (_02379_, _06222_, _06103_);
  and _24081_ (_02381_, _02379_, _02377_);
  or _24082_ (_02382_, _02381_, _06210_);
  or _24083_ (_02383_, _02361_, _02118_);
  and _24084_ (_02384_, _02383_, _02110_);
  and _24085_ (_02385_, _02384_, _02382_);
  and _24086_ (_02386_, _06208_, _06103_);
  or _24087_ (_02387_, _02386_, _06205_);
  or _24088_ (_02388_, _02387_, _02385_);
  or _24089_ (_02389_, _02361_, _06206_);
  and _24090_ (_02390_, _02389_, _02099_);
  and _24091_ (_02391_, _02390_, _02388_);
  or _24092_ (_02392_, _02391_, _02375_);
  and _24093_ (_02394_, _02392_, _06235_);
  or _24094_ (_02395_, _02394_, _02360_);
  and _24095_ (_01943_, _02395_, _04856_);
  and _24096_ (_01953_, _07173_, _04856_);
  and _24097_ (_01960_, _07124_, _04856_);
  and _24098_ (_01962_, _07053_, _04856_);
  and _24099_ (_01964_, _06991_, _04856_);
  and _24100_ (_02396_, _07855_, _06143_);
  or _24101_ (_02397_, _02396_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and _24102_ (_02398_, _02397_, _06129_);
  nand _24103_ (_02399_, _02396_, _06088_);
  and _24104_ (_02400_, _02399_, _02398_);
  and _24105_ (_02401_, _06410_, _06127_);
  or _24106_ (_02402_, _02401_, _02400_);
  and _24107_ (_02016_, _02402_, _04856_);
  and _24108_ (_02403_, _06494_, _06143_);
  or _24109_ (_02404_, _02403_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and _24110_ (_02405_, _02404_, _06129_);
  nand _24111_ (_02406_, _02403_, _06088_);
  and _24112_ (_02407_, _02406_, _02405_);
  and _24113_ (_02409_, _06705_, _06127_);
  or _24114_ (_02410_, _02409_, _02407_);
  and _24115_ (_02022_, _02410_, _04856_);
  and _24116_ (_02411_, _06270_, _04990_);
  or _24117_ (_02412_, _02411_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and _24118_ (_02413_, _02412_, _06276_);
  nand _24119_ (_02414_, _02411_, _06088_);
  and _24120_ (_02415_, _02414_, _02413_);
  and _24121_ (_02416_, _06997_, _06275_);
  or _24122_ (_02417_, _02416_, _02415_);
  and _24123_ (_02036_, _02417_, _04856_);
  and _24124_ (_02418_, _06269_, _06135_);
  and _24125_ (_02419_, _07642_, _02418_);
  nand _24126_ (_02420_, _02418_, _04984_);
  and _24127_ (_02421_, _02418_, _12258_);
  or _24128_ (_02422_, _02421_, _02420_);
  and _24129_ (_02423_, _02422_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  or _24130_ (_02425_, _02423_, _06275_);
  or _24131_ (_02426_, _02425_, _02419_);
  nand _24132_ (_02427_, _06275_, _05669_);
  and _24133_ (_02428_, _02427_, _04856_);
  and _24134_ (_02042_, _02428_, _02426_);
  not _24135_ (_02429_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  nor _24136_ (_02430_, _02421_, _02429_);
  or _24137_ (_02431_, _02430_, _06275_);
  and _24138_ (_02432_, _04985_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or _24139_ (_02433_, _02432_, _07602_);
  and _24140_ (_02434_, _02433_, _06270_);
  or _24141_ (_02435_, _02434_, _02431_);
  or _24142_ (_02436_, _06705_, _06276_);
  and _24143_ (_02437_, _02436_, _04856_);
  and _24144_ (_02049_, _02437_, _02435_);
  and _24145_ (_02439_, _06270_, _06146_);
  or _24146_ (_02440_, _02439_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and _24147_ (_02441_, _02440_, _06276_);
  nand _24148_ (_02442_, _02439_, _06088_);
  and _24149_ (_02443_, _02442_, _02441_);
  nor _24150_ (_02444_, _06276_, _05287_);
  or _24151_ (_02445_, _02444_, _02443_);
  and _24152_ (_02054_, _02445_, _04856_);
  and _24153_ (_02446_, _06297_, _04990_);
  and _24154_ (_02447_, _02446_, _06088_);
  nor _24155_ (_02448_, _02446_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  or _24156_ (_02449_, _02448_, _02447_);
  nand _24157_ (_02450_, _02449_, _06305_);
  nand _24158_ (_02451_, _06369_, _06304_);
  and _24159_ (_02453_, _02451_, _04856_);
  and _24160_ (_02062_, _02453_, _02450_);
  and _24161_ (_02455_, _06297_, _05520_);
  nand _24162_ (_02456_, _02455_, _06088_);
  or _24163_ (_02457_, _02455_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and _24164_ (_02458_, _02457_, _06305_);
  and _24165_ (_02459_, _02458_, _02456_);
  nor _24166_ (_02460_, _06305_, _05669_);
  or _24167_ (_02462_, _02460_, _02459_);
  and _24168_ (_02072_, _02462_, _04856_);
  and _24169_ (_02463_, _04985_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or _24170_ (_02464_, _02463_, _07602_);
  and _24171_ (_02465_, _02464_, _06297_);
  nand _24172_ (_02466_, _06297_, _12258_);
  and _24173_ (_02467_, _02466_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or _24174_ (_02468_, _02467_, _06304_);
  or _24175_ (_02469_, _02468_, _02465_);
  or _24176_ (_02470_, _06705_, _06305_);
  and _24177_ (_02471_, _02470_, _04856_);
  and _24178_ (_02082_, _02471_, _02469_);
  and _24179_ (_02472_, _06297_, _06146_);
  nand _24180_ (_02473_, _02472_, _06088_);
  or _24181_ (_02474_, _02472_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and _24182_ (_02475_, _02474_, _06305_);
  and _24183_ (_02476_, _02475_, _02473_);
  nor _24184_ (_02477_, _06305_, _05287_);
  or _24185_ (_02478_, _02477_, _02476_);
  and _24186_ (_02091_, _02478_, _04856_);
  and _24187_ (_02479_, _09212_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  and _24188_ (_02480_, _02479_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  and _24189_ (_02482_, _02480_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  or _24190_ (_02484_, _02482_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  nand _24191_ (_02485_, _02482_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  and _24192_ (_02487_, _02485_, _02484_);
  and _24193_ (_02137_, _02487_, _02321_);
  not _24194_ (_02488_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  and _24195_ (_02489_, _09215_, _02488_);
  and _24196_ (_02490_, _02489_, _09236_);
  nor _24197_ (_02491_, _09215_, _01113_);
  or _24198_ (_02492_, _02491_, _02490_);
  and _24199_ (_02493_, _02492_, _09212_);
  nand _24200_ (_02494_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  nor _24201_ (_02495_, _02494_, _09211_);
  nor _24202_ (_02496_, _02495_, _02493_);
  nor _24203_ (_02497_, _02496_, _09210_);
  or _24204_ (_02498_, _02497_, _09237_);
  and _24205_ (_02159_, _02498_, _02321_);
  nand _24206_ (_02499_, _02490_, _09211_);
  nand _24207_ (_02500_, _02499_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  nor _24208_ (_02501_, _02500_, _09237_);
  or _24209_ (_02502_, _02501_, _09206_);
  and _24210_ (_02198_, _02502_, _04856_);
  or _24211_ (_02504_, _12818_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1]);
  or _24212_ (_02505_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2], _09249_);
  or _24213_ (_02506_, _02505_, _08087_);
  and _24214_ (_02507_, _02506_, _04856_);
  and _24215_ (_02208_, _02507_, _02504_);
  nor _24216_ (_02508_, _02479_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  nor _24217_ (_02509_, _02508_, _02480_);
  and _24218_ (_02224_, _02509_, _02321_);
  or _24219_ (_02510_, _06238_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  nand _24220_ (_02511_, _06238_, _02015_);
  and _24221_ (_02513_, _02511_, _04856_);
  and _24222_ (_02235_, _02513_, _02510_);
  nor _24223_ (_02514_, _09212_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  nor _24224_ (_02515_, _02514_, _02479_);
  and _24225_ (_02239_, _02515_, _02321_);
  and _24226_ (_02340_, _06347_, _04856_);
  and _24227_ (_02516_, _06238_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  not _24228_ (_02517_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nor _24229_ (_02518_, _06238_, _02517_);
  or _24230_ (_02519_, _02518_, _02516_);
  and _24231_ (_02378_, _02519_, _04856_);
  and _24232_ (_02521_, _08037_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  and _24233_ (_02522_, _08790_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  and _24234_ (_02523_, _07411_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or _24235_ (_02524_, _02523_, _02522_);
  and _24236_ (_02525_, _07422_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and _24237_ (_02526_, _07429_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  or _24238_ (_02527_, _02526_, _02525_);
  or _24239_ (_02528_, _02527_, _02524_);
  and _24240_ (_02529_, _07437_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and _24241_ (_02530_, _07442_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  or _24242_ (_02531_, _02530_, _02529_);
  and _24243_ (_02532_, _07449_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and _24244_ (_02533_, _07455_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  or _24245_ (_02534_, _02533_, _02532_);
  or _24246_ (_02535_, _02534_, _02531_);
  or _24247_ (_02536_, _02535_, _02528_);
  and _24248_ (_02537_, _07466_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  nor _24249_ (_02538_, _07463_, _00593_);
  or _24250_ (_02539_, _02538_, _02537_);
  and _24251_ (_02540_, _07470_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and _24252_ (_02541_, _07473_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  or _24253_ (_02542_, _02541_, _02540_);
  or _24254_ (_02544_, _02542_, _02539_);
  not _24255_ (_02546_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  nor _24256_ (_02547_, _07486_, _02546_);
  and _24257_ (_02549_, _07484_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  or _24258_ (_02551_, _02549_, _02547_);
  and _24259_ (_02553_, _07477_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and _24260_ (_02554_, _07479_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or _24261_ (_02556_, _02554_, _02553_);
  or _24262_ (_02557_, _02556_, _02551_);
  or _24263_ (_02559_, _02557_, _02544_);
  or _24264_ (_02561_, _02559_, _02536_);
  and _24265_ (_02562_, _08028_, _07346_);
  and _24266_ (_02563_, _07500_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  or _24267_ (_02564_, _02563_, _02562_);
  and _24268_ (_02565_, _07389_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and _24269_ (_02566_, _07494_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or _24270_ (_02567_, _02566_, _02565_);
  or _24271_ (_02568_, _02567_, _02564_);
  and _24272_ (_02569_, _01877_, _07507_);
  and _24273_ (_02570_, _01916_, _07539_);
  or _24274_ (_02571_, _02570_, _02569_);
  and _24275_ (_02572_, _01735_, _07547_);
  and _24276_ (_02574_, _01606_, _07552_);
  or _24277_ (_02576_, _02574_, _02572_);
  or _24278_ (_02578_, _02576_, _02571_);
  or _24279_ (_02579_, _02578_, _02568_);
  and _24280_ (_02580_, _07943_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and _24281_ (_02581_, _07561_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or _24282_ (_02582_, _02581_, _02580_);
  or _24283_ (_02583_, _02582_, _02579_);
  or _24284_ (_02584_, _02583_, _02561_);
  and _24285_ (_02585_, _02584_, _08004_);
  or _24286_ (_02586_, _02585_, _07390_);
  or _24287_ (_02587_, _02586_, _02521_);
  or _24288_ (_02589_, _08786_, _05641_);
  and _24289_ (_02591_, _02589_, _04856_);
  and _24290_ (_02393_, _02591_, _02587_);
  nor _24291_ (_02593_, _02480_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  nor _24292_ (_02594_, _02593_, _02482_);
  and _24293_ (_02408_, _02594_, _02321_);
  nor _24294_ (_02595_, _07390_, rst);
  and _24295_ (_02424_, _02595_, _08787_);
  and _24296_ (_02596_, _09023_, _04987_);
  and _24297_ (_02597_, _02596_, _05510_);
  and _24298_ (_02598_, _02597_, _08070_);
  and _24299_ (_02599_, _02598_, _06705_);
  and _24300_ (_02600_, _09218_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  and _24301_ (_02601_, _09217_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  nor _24302_ (_02602_, _02601_, _02600_);
  nor _24303_ (_02603_, _02602_, _09206_);
  and _24304_ (_02604_, _02597_, _08060_);
  and _24305_ (_02605_, _02604_, _05670_);
  or _24306_ (_02606_, _02605_, _02603_);
  or _24307_ (_02607_, _02606_, _02599_);
  and _24308_ (_02438_, _02607_, _04856_);
  and _24309_ (_02608_, _08067_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  and _24310_ (_02609_, _02608_, _10230_);
  or _24311_ (_02610_, _02609_, _10232_);
  and _24312_ (_02611_, _08085_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  and _24313_ (_02612_, _02611_, _02610_);
  nand _24314_ (_02613_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9], _04856_);
  nor _24315_ (_02614_, _02613_, _12818_);
  or _24316_ (_02452_, _02614_, _02612_);
  and _24317_ (_02615_, _02604_, _06705_);
  and _24318_ (_02616_, _09218_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  and _24319_ (_02617_, _09217_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  nor _24320_ (_02618_, _02617_, _02616_);
  nor _24321_ (_02619_, _02618_, _09206_);
  and _24322_ (_02620_, _02598_, _06033_);
  or _24323_ (_02621_, _02620_, _02619_);
  or _24324_ (_02622_, _02621_, _02615_);
  and _24325_ (_02454_, _02622_, _04856_);
  and _24326_ (_02623_, _09218_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  and _24327_ (_02624_, _09217_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  nor _24328_ (_02626_, _02624_, _02623_);
  nor _24329_ (_02628_, _02626_, _09206_);
  and _24330_ (_02629_, _09223_, _05718_);
  or _24331_ (_02630_, _02629_, _02628_);
  and _24332_ (_02631_, _09207_, _05288_);
  or _24333_ (_02632_, _02631_, _02630_);
  and _24334_ (_02461_, _02632_, _04856_);
  not _24335_ (_02633_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  and _24336_ (_02634_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  not _24337_ (_02635_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and _24338_ (_02636_, _06316_, _02635_);
  nor _24339_ (_02638_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6], _02546_);
  or _24340_ (_02639_, _02638_, _02636_);
  nor _24341_ (_02640_, _02639_, _02634_);
  nand _24342_ (_02641_, _02640_, _02633_);
  nor _24343_ (_02642_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nor _24344_ (_02643_, _02642_, _02640_);
  nand _24345_ (_02644_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nand _24346_ (_02645_, _02644_, _02643_);
  and _24347_ (_02646_, _02645_, _04856_);
  and _24348_ (_02481_, _02646_, _02641_);
  and _24349_ (_02483_, _02643_, _04856_);
  not _24350_ (_02647_, _08082_);
  or _24351_ (_02648_, _08068_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  or _24352_ (_02649_, _02648_, _02044_);
  and _24353_ (_02650_, _02649_, _02647_);
  or _24354_ (_02651_, _02650_, rxd_i);
  and _24355_ (_02652_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1], rxd_i);
  nor _24356_ (_02653_, _02652_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0]);
  and _24357_ (_02654_, _02653_, _08067_);
  and _24358_ (_02656_, _02654_, _08062_);
  nor _24359_ (_02657_, _02656_, _10231_);
  and _24360_ (_02658_, _02657_, _02651_);
  or _24361_ (_02659_, _02658_, _09249_);
  not _24362_ (_02660_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  or _24363_ (_02661_, _08087_, _09249_);
  nand _24364_ (_02663_, _02661_, _02660_);
  and _24365_ (_02665_, _02663_, _04856_);
  and _24366_ (_02486_, _02665_, _02659_);
  and _24367_ (_02666_, _10232_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  and _24368_ (_02667_, _08077_, _08072_);
  or _24369_ (_02669_, _02667_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  or _24370_ (_02671_, _08077_, _08069_);
  and _24371_ (_02672_, _02671_, _02647_);
  and _24372_ (_02674_, _02672_, _02669_);
  or _24373_ (_02675_, _02674_, _02666_);
  and _24374_ (_02676_, _02675_, _08085_);
  or _24375_ (_02503_, _02676_, _02271_);
  not _24376_ (_02677_, _12761_);
  or _24377_ (_02678_, _02677_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  or _24378_ (_02679_, _08087_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  and _24379_ (_02680_, _02679_, _08085_);
  and _24380_ (_02681_, _02680_, _02678_);
  or _24381_ (_02520_, _02681_, _02167_);
  and _24382_ (_02682_, _09017_, _06146_);
  nand _24383_ (_02683_, _02682_, _06088_);
  or _24384_ (_02684_, _02682_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and _24385_ (_02685_, _02684_, _06093_);
  and _24386_ (_02686_, _02685_, _02683_);
  nand _24387_ (_02687_, _09024_, _05287_);
  or _24388_ (_02689_, _09024_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and _24389_ (_02690_, _02689_, _05510_);
  and _24390_ (_02692_, _02690_, _02687_);
  and _24391_ (_02694_, _08999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  or _24392_ (_02695_, _02694_, rst);
  or _24393_ (_02696_, _02695_, _02692_);
  or _24394_ (_02543_, _02696_, _02686_);
  and _24395_ (_02698_, _08988_, _07855_);
  nand _24396_ (_02699_, _02698_, _06088_);
  or _24397_ (_02700_, _02698_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and _24398_ (_02701_, _02700_, _06093_);
  and _24399_ (_02702_, _02701_, _02699_);
  not _24400_ (_02703_, _08994_);
  or _24401_ (_02704_, _02703_, _06410_);
  or _24402_ (_02705_, _08994_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and _24403_ (_02706_, _02705_, _05510_);
  and _24404_ (_02707_, _02706_, _02704_);
  and _24405_ (_02709_, _08999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or _24406_ (_02711_, _02709_, rst);
  or _24407_ (_02713_, _02711_, _02707_);
  or _24408_ (_02545_, _02713_, _02702_);
  not _24409_ (_02714_, _05631_);
  or _24410_ (_02715_, _06054_, _02714_);
  or _24411_ (_02716_, _05631_, _06053_);
  and _24412_ (_02717_, _02716_, _05583_);
  and _24413_ (_02718_, _02717_, _02715_);
  and _24414_ (_02719_, _05497_, ABINPUT001[0]);
  and _24415_ (_02721_, _05499_, ABINPUT000[0]);
  or _24416_ (_02722_, _02721_, _02719_);
  nand _24417_ (_02723_, _05431_, _05340_);
  and _24418_ (_02725_, _05433_, _05455_);
  and _24419_ (_02727_, _02725_, _02723_);
  or _24420_ (_02729_, _02727_, _02722_);
  or _24421_ (_02730_, _02729_, _02718_);
  and _24422_ (_02731_, _02730_, \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  not _24423_ (_02732_, \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  and _24424_ (_02733_, _02732_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or _24425_ (_02734_, _02733_, _08277_);
  or _24426_ (_02735_, _02734_, _02731_);
  not _24427_ (_02736_, _06494_);
  nand _24428_ (_02737_, _02736_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  nand _24429_ (_02738_, _02737_, _08277_);
  or _24430_ (_02739_, _02738_, _07602_);
  and _24431_ (_02741_, _02739_, _06935_);
  and _24432_ (_02742_, _02741_, _02735_);
  and _24433_ (_02743_, _06934_, _06705_);
  or _24434_ (_02744_, _02743_, _02742_);
  and _24435_ (_02548_, _02744_, _04856_);
  and _24436_ (_02745_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _24437_ (_02746_, _02745_, _12766_);
  and _24438_ (_02550_, _02746_, _04856_);
  and _24439_ (_02747_, _09132_, _07855_);
  nand _24440_ (_02748_, _02747_, _06088_);
  or _24441_ (_02750_, _02747_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and _24442_ (_02752_, _02750_, _06093_);
  and _24443_ (_02753_, _02752_, _02748_);
  and _24444_ (_02754_, _09138_, _06410_);
  and _24445_ (_02755_, _09139_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or _24446_ (_02757_, _02755_, _02754_);
  and _24447_ (_02758_, _02757_, _05510_);
  and _24448_ (_02759_, _08999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or _24449_ (_02760_, _02759_, rst);
  or _24450_ (_02761_, _02760_, _02758_);
  or _24451_ (_02552_, _02761_, _02753_);
  and _24452_ (_02762_, _09116_, _06494_);
  or _24453_ (_02764_, _02762_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and _24454_ (_02765_, _02764_, _06093_);
  nand _24455_ (_02766_, _02762_, _06088_);
  and _24456_ (_02767_, _02766_, _02765_);
  and _24457_ (_02769_, _09123_, _06705_);
  and _24458_ (_02770_, _09124_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or _24459_ (_02772_, _02770_, _02769_);
  and _24460_ (_02773_, _02772_, _05510_);
  and _24461_ (_02774_, _08999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or _24462_ (_02775_, _02774_, rst);
  or _24463_ (_02777_, _02775_, _02773_);
  or _24464_ (_02555_, _02777_, _02767_);
  and _24465_ (_02778_, _09116_, _06091_);
  or _24466_ (_02779_, _02778_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and _24467_ (_02780_, _02779_, _06093_);
  nand _24468_ (_02781_, _02778_, _06088_);
  and _24469_ (_02783_, _02781_, _02780_);
  and _24470_ (_02784_, _09123_, _05718_);
  nor _24471_ (_02785_, _09123_, _01891_);
  or _24472_ (_02786_, _02785_, _02784_);
  and _24473_ (_02788_, _02786_, _05510_);
  nor _24474_ (_02789_, _06092_, _01891_);
  or _24475_ (_02790_, _02789_, rst);
  or _24476_ (_02791_, _02790_, _02788_);
  or _24477_ (_02558_, _02791_, _02783_);
  or _24478_ (_02793_, _02045_, _09251_);
  and _24479_ (_02794_, _02793_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  or _24480_ (_02795_, _02794_, _01937_);
  and _24481_ (_02560_, _02795_, _04856_);
  and _24482_ (_02796_, _09017_, _05520_);
  nand _24483_ (_02797_, _02796_, _06088_);
  or _24484_ (_02799_, _02796_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and _24485_ (_02800_, _02799_, _06093_);
  and _24486_ (_02801_, _02800_, _02797_);
  nand _24487_ (_02802_, _09024_, _05669_);
  or _24488_ (_02803_, _09024_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and _24489_ (_02805_, _02803_, _05510_);
  and _24490_ (_02807_, _02805_, _02802_);
  nor _24491_ (_02808_, _06092_, _08839_);
  or _24492_ (_02810_, _02808_, rst);
  or _24493_ (_02811_, _02810_, _02807_);
  or _24494_ (_02573_, _02811_, _02801_);
  and _24495_ (_02812_, _08988_, _05520_);
  nand _24496_ (_02814_, _02812_, _06088_);
  or _24497_ (_02815_, _02812_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and _24498_ (_02817_, _02815_, _06093_);
  and _24499_ (_02818_, _02817_, _02814_);
  nand _24500_ (_02819_, _08994_, _05669_);
  or _24501_ (_02820_, _08994_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and _24502_ (_02821_, _02820_, _05510_);
  and _24503_ (_02822_, _02821_, _02819_);
  nor _24504_ (_02823_, _06092_, _08834_);
  or _24505_ (_02824_, _02823_, rst);
  or _24506_ (_02825_, _02824_, _02822_);
  or _24507_ (_02575_, _02825_, _02818_);
  and _24508_ (_02826_, _08988_, _06146_);
  nand _24509_ (_02827_, _02826_, _06088_);
  or _24510_ (_02828_, _02826_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and _24511_ (_02830_, _02828_, _06093_);
  and _24512_ (_02831_, _02830_, _02827_);
  nand _24513_ (_02832_, _08994_, _05287_);
  or _24514_ (_02834_, _08994_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and _24515_ (_02835_, _02834_, _05510_);
  and _24516_ (_02837_, _02835_, _02832_);
  and _24517_ (_02838_, _08999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  or _24518_ (_02840_, _02838_, rst);
  or _24519_ (_02841_, _02840_, _02837_);
  or _24520_ (_02577_, _02841_, _02831_);
  and _24521_ (_02842_, _09132_, _06146_);
  nand _24522_ (_02843_, _02842_, _06088_);
  or _24523_ (_02844_, _02842_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and _24524_ (_02845_, _02844_, _06093_);
  and _24525_ (_02846_, _02845_, _02843_);
  nor _24526_ (_02848_, _09139_, _05287_);
  and _24527_ (_02849_, _09139_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or _24528_ (_02850_, _02849_, _02848_);
  and _24529_ (_02851_, _02850_, _05510_);
  and _24530_ (_02852_, _08999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or _24531_ (_02853_, _02852_, rst);
  or _24532_ (_02854_, _02853_, _02851_);
  or _24533_ (_02588_, _02854_, _02846_);
  and _24534_ (_02855_, _09116_, _04990_);
  or _24535_ (_02856_, _02855_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and _24536_ (_02857_, _02856_, _06093_);
  nand _24537_ (_02858_, _02855_, _06088_);
  and _24538_ (_02859_, _02858_, _02857_);
  and _24539_ (_02861_, _09123_, _06997_);
  and _24540_ (_02862_, _09124_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  or _24541_ (_02863_, _02862_, _02861_);
  and _24542_ (_02865_, _02863_, _05510_);
  and _24543_ (_02866_, _08999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  or _24544_ (_02867_, _02866_, rst);
  or _24545_ (_02868_, _02867_, _02865_);
  or _24546_ (_02590_, _02868_, _02859_);
  and _24547_ (_02870_, _09116_, _07855_);
  or _24548_ (_02871_, _02870_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and _24549_ (_02872_, _02871_, _06093_);
  nand _24550_ (_02873_, _02870_, _06088_);
  and _24551_ (_02874_, _02873_, _02872_);
  and _24552_ (_02875_, _09123_, _06410_);
  and _24553_ (_02876_, _09124_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or _24554_ (_02878_, _02876_, _02875_);
  and _24555_ (_02879_, _02878_, _05510_);
  and _24556_ (_02880_, _08999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or _24557_ (_02881_, _02880_, rst);
  or _24558_ (_02882_, _02881_, _02879_);
  or _24559_ (_02592_, _02882_, _02874_);
  and _24560_ (_02884_, _09132_, _05520_);
  nand _24561_ (_02885_, _02884_, _06088_);
  or _24562_ (_02886_, _02884_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and _24563_ (_02888_, _02886_, _06093_);
  and _24564_ (_02889_, _02888_, _02885_);
  nor _24565_ (_02890_, _09139_, _05669_);
  nor _24566_ (_02891_, _09138_, _08845_);
  or _24567_ (_02892_, _02891_, _02890_);
  and _24568_ (_02893_, _02892_, _05510_);
  nor _24569_ (_02894_, _06092_, _08845_);
  or _24570_ (_02895_, _02894_, rst);
  or _24571_ (_02897_, _02895_, _02893_);
  or _24572_ (_02625_, _02897_, _02889_);
  and _24573_ (_02899_, _09132_, _06494_);
  nand _24574_ (_02900_, _02899_, _06088_);
  or _24575_ (_02901_, _02899_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and _24576_ (_02902_, _02901_, _06093_);
  and _24577_ (_02903_, _02902_, _02900_);
  and _24578_ (_02904_, _09138_, _06705_);
  and _24579_ (_02905_, _09139_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or _24580_ (_02907_, _02905_, _02904_);
  and _24581_ (_02908_, _02907_, _05510_);
  and _24582_ (_02909_, _08999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or _24583_ (_02910_, _02909_, rst);
  or _24584_ (_02912_, _02910_, _02908_);
  or _24585_ (_02627_, _02912_, _02903_);
  nand _24586_ (_02914_, _01352_, _12258_);
  and _24587_ (_02915_, _02914_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and _24588_ (_02916_, _04985_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or _24589_ (_02917_, _02916_, _07602_);
  and _24590_ (_02918_, _02917_, _01352_);
  or _24591_ (_02919_, _02918_, _02915_);
  and _24592_ (_02920_, _02919_, _06093_);
  and _24593_ (_02921_, _08999_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  nand _24594_ (_02922_, _01361_, _06552_);
  or _24595_ (_02924_, _01361_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and _24596_ (_02926_, _02924_, _05510_);
  and _24597_ (_02927_, _02926_, _02922_);
  or _24598_ (_02928_, _02927_, _02921_);
  or _24599_ (_02929_, _02928_, _02920_);
  and _24600_ (_02637_, _02929_, _04856_);
  and _24601_ (_02930_, _01352_, _06091_);
  nand _24602_ (_02931_, _02930_, _06088_);
  or _24603_ (_02932_, _02930_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and _24604_ (_02933_, _02932_, _06093_);
  and _24605_ (_02935_, _02933_, _02931_);
  and _24606_ (_02937_, _08999_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nand _24607_ (_02938_, _01361_, _07897_);
  or _24608_ (_02939_, _01361_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and _24609_ (_02940_, _02939_, _05510_);
  and _24610_ (_02942_, _02940_, _02938_);
  or _24611_ (_02943_, _02942_, _02937_);
  or _24612_ (_02944_, _02943_, _02935_);
  and _24613_ (_02655_, _02944_, _04856_);
  and _24614_ (_02945_, _09132_, _04986_);
  nand _24615_ (_02947_, _02945_, _06088_);
  or _24616_ (_02948_, _02945_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and _24617_ (_02949_, _02948_, _06093_);
  and _24618_ (_02951_, _02949_, _02947_);
  nor _24619_ (_02952_, _09139_, _06032_);
  nor _24620_ (_02953_, _09138_, _01860_);
  or _24621_ (_02955_, _02953_, _02952_);
  and _24622_ (_02956_, _02955_, _05510_);
  nor _24623_ (_02957_, _06092_, _01860_);
  or _24624_ (_02958_, _02957_, rst);
  or _24625_ (_02959_, _02958_, _02956_);
  or _24626_ (_02662_, _02959_, _02951_);
  and _24627_ (_02960_, _09132_, _04990_);
  nand _24628_ (_02961_, _02960_, _06088_);
  or _24629_ (_02963_, _02960_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and _24630_ (_02965_, _02963_, _06093_);
  and _24631_ (_02966_, _02965_, _02961_);
  and _24632_ (_02967_, _09138_, _06997_);
  and _24633_ (_02969_, _09139_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  or _24634_ (_02970_, _02969_, _02967_);
  and _24635_ (_02971_, _02970_, _05510_);
  and _24636_ (_02972_, _08999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  or _24637_ (_02973_, _02972_, rst);
  or _24638_ (_02974_, _02973_, _02971_);
  or _24639_ (_02664_, _02974_, _02966_);
  and _24640_ (_02975_, _09218_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  and _24641_ (_02976_, _09217_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  nor _24642_ (_02977_, _02976_, _02975_);
  nor _24643_ (_02978_, _02977_, _09206_);
  and _24644_ (_02979_, _09223_, _06410_);
  or _24645_ (_02980_, _02979_, _02978_);
  and _24646_ (_02981_, _09207_, _05718_);
  or _24647_ (_02982_, _02981_, _02980_);
  and _24648_ (_02668_, _02982_, _04856_);
  nand _24649_ (_02984_, _08988_, _12258_);
  and _24650_ (_02985_, _02984_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and _24651_ (_02986_, _04985_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or _24652_ (_02987_, _02986_, _07602_);
  and _24653_ (_02989_, _02987_, _08988_);
  or _24654_ (_02990_, _02989_, _02985_);
  and _24655_ (_02991_, _02990_, _06093_);
  or _24656_ (_02992_, _02703_, _06705_);
  or _24657_ (_02993_, _08994_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and _24658_ (_02994_, _02993_, _05510_);
  and _24659_ (_02995_, _02994_, _02992_);
  and _24660_ (_02996_, _08999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or _24661_ (_02997_, _02996_, rst);
  or _24662_ (_02998_, _02997_, _02995_);
  or _24663_ (_02670_, _02998_, _02991_);
  and _24664_ (_03000_, _05517_, _04999_);
  nand _24665_ (_03002_, _03000_, _06088_);
  or _24666_ (_03003_, _03000_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and _24667_ (_03004_, _03003_, _06093_);
  and _24668_ (_03005_, _03004_, _03002_);
  or _24669_ (_03006_, _08994_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  nand _24670_ (_03007_, _08994_, _06032_);
  and _24671_ (_03008_, _03007_, _05510_);
  and _24672_ (_03009_, _03008_, _03006_);
  nor _24673_ (_03010_, _06092_, _01727_);
  or _24674_ (_03011_, _03010_, rst);
  or _24675_ (_03012_, _03011_, _03009_);
  or _24676_ (_02673_, _03012_, _03005_);
  nand _24677_ (_03013_, _08988_, _04990_);
  or _24678_ (_03014_, _03013_, _06144_);
  or _24679_ (_03015_, _08994_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  and _24680_ (_03016_, _03015_, _06093_);
  and _24681_ (_03017_, _03016_, _03014_);
  nand _24682_ (_03018_, _08994_, _06369_);
  and _24683_ (_03019_, _03018_, _05510_);
  and _24684_ (_03020_, _03019_, _03015_);
  and _24685_ (_03021_, _08999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  or _24686_ (_03022_, _03021_, rst);
  or _24687_ (_03023_, _03022_, _03020_);
  or _24688_ (_02688_, _03023_, _03017_);
  and _24689_ (_03024_, _09017_, _04986_);
  nand _24690_ (_03025_, _03024_, _06088_);
  or _24691_ (_03026_, _03024_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and _24692_ (_03027_, _03026_, _06093_);
  and _24693_ (_03028_, _03027_, _03025_);
  or _24694_ (_03029_, _09024_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  nand _24695_ (_03030_, _09024_, _06032_);
  and _24696_ (_03031_, _03030_, _05510_);
  and _24697_ (_03032_, _03031_, _03029_);
  nor _24698_ (_03033_, _06092_, _01625_);
  or _24699_ (_03034_, _03033_, rst);
  or _24700_ (_03035_, _03034_, _03032_);
  or _24701_ (_02691_, _03035_, _03028_);
  nand _24702_ (_03037_, _09017_, _04990_);
  or _24703_ (_03038_, _03037_, _06144_);
  or _24704_ (_03039_, _09024_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and _24705_ (_03040_, _03039_, _06093_);
  and _24706_ (_03041_, _03040_, _03038_);
  nand _24707_ (_03042_, _09024_, _06369_);
  and _24708_ (_03043_, _03042_, _05510_);
  and _24709_ (_03044_, _03043_, _03039_);
  and _24710_ (_03045_, _08999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  or _24711_ (_03046_, _03045_, rst);
  or _24712_ (_03047_, _03046_, _03044_);
  or _24713_ (_02693_, _03047_, _03041_);
  and _24714_ (_03048_, _09017_, _06091_);
  nand _24715_ (_03049_, _03048_, _06088_);
  or _24716_ (_03050_, _03048_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and _24717_ (_03051_, _03050_, _06093_);
  and _24718_ (_03052_, _03051_, _03049_);
  not _24719_ (_03053_, _09024_);
  or _24720_ (_03054_, _03053_, _05718_);
  or _24721_ (_03055_, _09024_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and _24722_ (_03056_, _03055_, _05510_);
  and _24723_ (_03057_, _03056_, _03054_);
  nor _24724_ (_03058_, _06092_, _01630_);
  or _24725_ (_03059_, _03058_, rst);
  or _24726_ (_03060_, _03059_, _03057_);
  or _24727_ (_02697_, _03060_, _03052_);
  and _24728_ (_03061_, _09116_, _06146_);
  or _24729_ (_03063_, _03061_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and _24730_ (_03064_, _03063_, _06093_);
  nand _24731_ (_03065_, _03061_, _06088_);
  and _24732_ (_03066_, _03065_, _03064_);
  nor _24733_ (_03068_, _09124_, _05287_);
  and _24734_ (_03069_, _09124_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or _24735_ (_03070_, _03069_, _03068_);
  and _24736_ (_03071_, _03070_, _05510_);
  and _24737_ (_03072_, _08999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or _24738_ (_03073_, _03072_, rst);
  or _24739_ (_03075_, _03073_, _03071_);
  or _24740_ (_02708_, _03075_, _03066_);
  and _24741_ (_03076_, _09116_, _05520_);
  or _24742_ (_03077_, _03076_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and _24743_ (_03078_, _03077_, _06093_);
  nand _24744_ (_03079_, _03076_, _06088_);
  and _24745_ (_03080_, _03079_, _03078_);
  nor _24746_ (_03081_, _09124_, _05669_);
  nor _24747_ (_03082_, _09123_, _08850_);
  or _24748_ (_03083_, _03082_, _03081_);
  and _24749_ (_03084_, _03083_, _05510_);
  nor _24750_ (_03085_, _06092_, _08850_);
  or _24751_ (_03086_, _03085_, rst);
  or _24752_ (_03087_, _03086_, _03084_);
  or _24753_ (_02710_, _03087_, _03080_);
  nand _24754_ (_03088_, _09115_, _04933_);
  or _24755_ (_03089_, _03088_, _09132_);
  and _24756_ (_03090_, _03089_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  nor _24757_ (_03091_, _04986_, _01886_);
  or _24758_ (_03092_, _03091_, _07713_);
  and _24759_ (_03093_, _03092_, _09116_);
  or _24760_ (_03094_, _03093_, _03090_);
  and _24761_ (_03095_, _03094_, _06093_);
  nor _24762_ (_03096_, _09124_, _06032_);
  nor _24763_ (_03098_, _09123_, _01886_);
  or _24764_ (_03099_, _03098_, _03096_);
  and _24765_ (_03100_, _03099_, _05510_);
  nor _24766_ (_03101_, _06092_, _01886_);
  or _24767_ (_03103_, _03101_, rst);
  or _24768_ (_03104_, _03103_, _03100_);
  or _24769_ (_02712_, _03104_, _03095_);
  and _24770_ (_03105_, _08988_, _06091_);
  nand _24771_ (_03106_, _03105_, _06088_);
  or _24772_ (_03107_, _03105_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and _24773_ (_03108_, _03107_, _06093_);
  and _24774_ (_03109_, _03108_, _03106_);
  or _24775_ (_03110_, _02703_, _05718_);
  or _24776_ (_03111_, _08994_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and _24777_ (_03112_, _03111_, _05510_);
  and _24778_ (_03113_, _03112_, _03110_);
  nor _24779_ (_03114_, _06092_, _01738_);
  or _24780_ (_03115_, _03114_, rst);
  or _24781_ (_03116_, _03115_, _03113_);
  or _24782_ (_02720_, _03116_, _03109_);
  and _24783_ (_03117_, _09017_, _07855_);
  nand _24784_ (_03118_, _03117_, _06088_);
  or _24785_ (_03119_, _03117_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and _24786_ (_03120_, _03119_, _06093_);
  and _24787_ (_03121_, _03120_, _03118_);
  or _24788_ (_03122_, _03053_, _06410_);
  or _24789_ (_03123_, _09024_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and _24790_ (_03124_, _03123_, _05510_);
  and _24791_ (_03125_, _03124_, _03122_);
  and _24792_ (_03126_, _08999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  or _24793_ (_03127_, _03126_, rst);
  or _24794_ (_03128_, _03127_, _03125_);
  or _24795_ (_02724_, _03128_, _03121_);
  and _24796_ (_03129_, _09017_, _06494_);
  nand _24797_ (_03130_, _03129_, _06088_);
  or _24798_ (_03131_, _03129_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and _24799_ (_03132_, _03131_, _06093_);
  and _24800_ (_03133_, _03132_, _03130_);
  or _24801_ (_03134_, _03053_, _06705_);
  or _24802_ (_03135_, _09024_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and _24803_ (_03136_, _03135_, _05510_);
  and _24804_ (_03137_, _03136_, _03134_);
  and _24805_ (_03138_, _08999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  or _24806_ (_03139_, _03138_, rst);
  or _24807_ (_03140_, _03139_, _03137_);
  or _24808_ (_02726_, _03140_, _03133_);
  and _24809_ (_03141_, _09132_, _06091_);
  nand _24810_ (_03142_, _03141_, _06088_);
  or _24811_ (_03143_, _03141_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and _24812_ (_03144_, _03143_, _06093_);
  and _24813_ (_03145_, _03144_, _03142_);
  and _24814_ (_03146_, _09138_, _05718_);
  nor _24815_ (_03147_, _09138_, _01852_);
  or _24816_ (_03148_, _03147_, _03146_);
  and _24817_ (_03149_, _03148_, _05510_);
  nor _24818_ (_03150_, _06092_, _01852_);
  or _24819_ (_03151_, _03150_, rst);
  or _24820_ (_03152_, _03151_, _03149_);
  or _24821_ (_02728_, _03152_, _03145_);
  or _24822_ (_03154_, _08087_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  nand _24823_ (_03155_, _01114_, _08073_);
  or _24824_ (_03156_, _03155_, _08062_);
  nand _24825_ (_03157_, _03156_, _03154_);
  nand _24826_ (_02740_, _03157_, _08085_);
  and _24827_ (_03158_, _06238_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor _24828_ (_03159_, _06238_, _00838_);
  or _24829_ (_03160_, _03159_, _03158_);
  and _24830_ (_02749_, _03160_, _04856_);
  and _24831_ (_02751_, _07334_, _04856_);
  and _24832_ (_03161_, _09255_, _08064_);
  and _24833_ (_03162_, _09253_, _03161_);
  nand _24834_ (_03163_, _03162_, _01939_);
  or _24835_ (_03164_, _03162_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  and _24836_ (_03166_, _03164_, _04856_);
  and _24837_ (_02756_, _03166_, _03163_);
  and _24838_ (_02763_, _07346_, _04856_);
  and _24839_ (_03167_, _09218_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  and _24840_ (_03168_, _09217_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  or _24841_ (_03169_, _03168_, _03167_);
  and _24842_ (_03170_, _03169_, _02321_);
  or _24843_ (_03171_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3], _02546_);
  and _24844_ (_03172_, _03171_, _04856_);
  and _24845_ (_03173_, _03172_, _09223_);
  or _24846_ (_02768_, _03173_, _03170_);
  not _24847_ (_03174_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r );
  nor _24848_ (_03175_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , _08073_);
  not _24849_ (_03176_, _03175_);
  nor _24850_ (_03178_, _08060_, _09249_);
  and _24851_ (_03179_, _03178_, _03176_);
  and _24852_ (_03181_, _03179_, _02044_);
  nor _24853_ (_03183_, _03181_, _03174_);
  and _24854_ (_03184_, _03181_, rxd_i);
  or _24855_ (_03185_, _03184_, rst);
  or _24856_ (_02771_, _03185_, _03183_);
  and _24857_ (_02776_, _07246_, _04856_);
  or _24858_ (_03187_, _03174_, rxd_i);
  nand _24859_ (_03188_, _03187_, _08071_);
  or _24860_ (_03189_, _08072_, _08061_);
  and _24861_ (_03191_, _03189_, _03188_);
  or _24862_ (_03192_, _08081_, _08078_);
  or _24863_ (_03193_, _03192_, _03191_);
  and _24864_ (_02782_, _03193_, _08085_);
  not _24865_ (_03194_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  and _24866_ (_03196_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  not _24867_ (_03197_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and _24868_ (_03199_, _06316_, _03197_);
  or _24869_ (_03201_, _03199_, _02638_);
  nor _24870_ (_03203_, _03201_, _03196_);
  nand _24871_ (_03205_, _03203_, _03194_);
  nor _24872_ (_03206_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  nor _24873_ (_03207_, _03206_, _03203_);
  nand _24874_ (_03208_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  nand _24875_ (_03209_, _03208_, _03207_);
  and _24876_ (_03210_, _03209_, _04856_);
  and _24877_ (_02787_, _03210_, _03205_);
  and _24878_ (_03212_, _06041_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  and _24879_ (_03213_, _09282_, _06043_);
  or _24880_ (_03214_, _03213_, _03212_);
  and _24881_ (_02792_, _03214_, _04856_);
  nand _24882_ (_02798_, _07011_, _04856_);
  and _24883_ (_03215_, _09282_, _05719_);
  and _24884_ (_03216_, _05723_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  or _24885_ (_03217_, _03216_, _03215_);
  and _24886_ (_02804_, _03217_, _04856_);
  and _24887_ (_03218_, _06238_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and _24888_ (_03219_, _00957_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  or _24889_ (_03220_, _03219_, _03218_);
  and _24890_ (_02806_, _03220_, _04856_);
  or _24891_ (_03222_, _06238_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  not _24892_ (_03223_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  nand _24893_ (_03224_, _06238_, _03223_);
  and _24894_ (_03225_, _03224_, _04856_);
  and _24895_ (_02809_, _03225_, _03222_);
  or _24896_ (_03226_, _06238_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  not _24897_ (_03227_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  nand _24898_ (_03228_, _06238_, _03227_);
  and _24899_ (_03229_, _03228_, _04856_);
  and _24900_ (_02813_, _03229_, _03226_);
  and _24901_ (_03230_, _06238_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  not _24902_ (_03231_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _24903_ (_03232_, _06238_, _03231_);
  or _24904_ (_03233_, _03232_, _03230_);
  and _24905_ (_02816_, _03233_, _04856_);
  and _24906_ (_03234_, _06238_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor _24907_ (_03235_, _06238_, _06342_);
  or _24908_ (_03236_, _03235_, _03234_);
  and _24909_ (_02829_, _03236_, _04856_);
  and _24910_ (_03237_, _06238_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  not _24911_ (_03238_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  nor _24912_ (_03239_, _06238_, _03238_);
  or _24913_ (_03240_, _03239_, _03237_);
  and _24914_ (_02833_, _03240_, _04856_);
  and _24915_ (_03241_, _06238_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  not _24916_ (_03242_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor _24917_ (_03243_, _06238_, _03242_);
  or _24918_ (_03244_, _03243_, _03241_);
  and _24919_ (_02836_, _03244_, _04856_);
  nor _24920_ (_03245_, _06284_, _06046_);
  and _24921_ (_03246_, _06046_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  or _24922_ (_03247_, _03246_, _05673_);
  or _24923_ (_03248_, _03247_, _03245_);
  or _24924_ (_03250_, _04861_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  and _24925_ (_03251_, _03250_, _04856_);
  and _24926_ (_02839_, _03251_, _03248_);
  nand _24927_ (_03252_, _10587_, _06284_);
  or _24928_ (_03253_, _10587_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  and _24929_ (_03254_, _03253_, _04856_);
  and _24930_ (_02847_, _03254_, _03252_);
  nand _24931_ (_03255_, _09200_, _06032_);
  or _24932_ (_03256_, _09200_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  and _24933_ (_03257_, _03256_, _04856_);
  and _24934_ (_02860_, _03257_, _03255_);
  and _24935_ (_03258_, _01973_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  nor _24936_ (_03259_, _01973_, _06284_);
  or _24937_ (_03260_, _03259_, _03258_);
  and _24938_ (_02864_, _03260_, _04856_);
  nor _24939_ (_03261_, _01973_, _05287_);
  and _24940_ (_03262_, _01973_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  or _24941_ (_03263_, _03262_, _03261_);
  and _24942_ (_02869_, _03263_, _04856_);
  nor _24943_ (_03264_, _06688_, _06284_);
  and _24944_ (_03265_, _06688_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  or _24945_ (_03266_, _03265_, _03264_);
  and _24946_ (_02877_, _03266_, _04856_);
  nand _24947_ (_03267_, _09200_, _06369_);
  or _24948_ (_03268_, _09200_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  and _24949_ (_03269_, _03268_, _04856_);
  and _24950_ (_02883_, _03269_, _03267_);
  and _24951_ (_03270_, _09282_, _05009_);
  and _24952_ (_03271_, _05007_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  and _24953_ (_03272_, _04861_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  and _24954_ (_03273_, _03272_, _05005_);
  or _24955_ (_03274_, _03273_, _03271_);
  or _24956_ (_03275_, _03274_, _03270_);
  and _24957_ (_02887_, _03275_, _04856_);
  or _24958_ (_03276_, _06238_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  not _24959_ (_03277_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nand _24960_ (_03278_, _06238_, _03277_);
  and _24961_ (_03279_, _03278_, _04856_);
  and _24962_ (_02896_, _03279_, _03276_);
  and _24963_ (_03280_, _06238_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  not _24964_ (_03281_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nor _24965_ (_03282_, _06238_, _03281_);
  or _24966_ (_03283_, _03282_, _03280_);
  and _24967_ (_02898_, _03283_, _04856_);
  and _24968_ (_03284_, _06238_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor _24969_ (_03285_, _06238_, _03223_);
  or _24970_ (_03286_, _03285_, _03284_);
  and _24971_ (_02906_, _03286_, _04856_);
  or _24972_ (_03287_, _09200_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  and _24973_ (_03288_, _03287_, _04856_);
  or _24974_ (_03289_, _09203_, _05718_);
  and _24975_ (_02911_, _03289_, _03288_);
  and _24976_ (_03290_, _06238_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  not _24977_ (_03291_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _24978_ (_03292_, _06238_, _03291_);
  or _24979_ (_03293_, _03292_, _03290_);
  and _24980_ (_02913_, _03293_, _04856_);
  or _24981_ (_03294_, _09200_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  and _24982_ (_03295_, _03294_, _04856_);
  or _24983_ (_03296_, _09203_, _06410_);
  and _24984_ (_02923_, _03296_, _03295_);
  or _24985_ (_03297_, _02677_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  or _24986_ (_03298_, _08087_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  and _24987_ (_03299_, _03298_, _08085_);
  and _24988_ (_03300_, _03299_, _03297_);
  or _24989_ (_02925_, _03300_, _02169_);
  or _24990_ (_03301_, _09200_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  and _24991_ (_03302_, _03301_, _04856_);
  nand _24992_ (_03303_, _09200_, _05287_);
  and _24993_ (_02934_, _03303_, _03302_);
  or _24994_ (_03304_, _12818_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  or _24995_ (_03305_, _02661_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1]);
  and _24996_ (_03306_, _03305_, _04856_);
  and _24997_ (_02936_, _03306_, _03304_);
  nor _24998_ (_02941_, _06314_, rst);
  or _24999_ (_03307_, _06238_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  not _25000_ (_03308_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nand _25001_ (_03309_, _06238_, _03308_);
  and _25002_ (_03310_, _03309_, _04856_);
  and _25003_ (_02946_, _03310_, _03307_);
  and _25004_ (_03311_, _06238_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor _25005_ (_03312_, _06238_, _03277_);
  or _25006_ (_03313_, _03312_, _03311_);
  and _25007_ (_02950_, _03313_, _04856_);
  or _25008_ (_03314_, _06238_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  nand _25009_ (_03315_, _06238_, _02517_);
  and _25010_ (_03316_, _03315_, _04856_);
  and _25011_ (_02962_, _03316_, _03314_);
  and _25012_ (_03317_, _06238_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor _25013_ (_03318_, _06238_, _03308_);
  or _25014_ (_03319_, _03318_, _03317_);
  and _25015_ (_02964_, _03319_, _04856_);
  or _25016_ (_03320_, _05678_, _05673_);
  and _25017_ (_03321_, _03320_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  and _25018_ (_03322_, _04861_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  and _25019_ (_03323_, _03322_, _05677_);
  and _25020_ (_03324_, _01971_, _06705_);
  or _25021_ (_03325_, _03324_, _03323_);
  or _25022_ (_03326_, _03325_, _03321_);
  and _25023_ (_02968_, _03326_, _04856_);
  and _25024_ (_03327_, _03320_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  and _25025_ (_03328_, _04861_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  and _25026_ (_03329_, _03328_, _05677_);
  nor _25027_ (_03330_, _01973_, _05669_);
  or _25028_ (_03331_, _03330_, _03329_);
  or _25029_ (_03332_, _03331_, _03327_);
  and _25030_ (_02983_, _03332_, _04856_);
  and _25031_ (_02988_, _03207_, _04856_);
  and _25032_ (_03333_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _04856_);
  and _25033_ (_03334_, _03333_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nor _25034_ (_03335_, _01075_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and _25035_ (_03336_, _01075_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nor _25036_ (_03337_, _03336_, _03335_);
  and _25037_ (_03338_, _03337_, _01077_);
  nor _25038_ (_03339_, _03337_, _01077_);
  or _25039_ (_03340_, _03339_, _03338_);
  or _25040_ (_03341_, _03340_, _06911_);
  or _25041_ (_03342_, _06910_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and _25042_ (_03343_, _03342_, _13190_);
  and _25043_ (_03344_, _03343_, _03341_);
  or _25044_ (_03001_, _03344_, _03334_);
  or _25045_ (_03345_, _05919_, _06812_);
  or _25046_ (_03346_, _05729_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and _25047_ (_03347_, _03346_, _04856_);
  and _25048_ (_03062_, _03347_, _03345_);
  not _25049_ (_03348_, _00536_);
  and _25050_ (_03349_, _03348_, _00490_);
  or _25051_ (_03350_, _13236_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  and _25052_ (_03097_, _03350_, _04856_);
  and _25053_ (_03351_, _03097_, _00002_);
  and _25054_ (_03067_, _03351_, _03349_);
  and _25055_ (_03352_, _01973_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  and _25056_ (_03353_, _01971_, _06410_);
  or _25057_ (_03354_, _03353_, _03352_);
  and _25058_ (_03074_, _03354_, _04856_);
  or _25059_ (_03355_, _01048_, _05718_);
  or _25060_ (_03356_, _10587_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  and _25061_ (_03357_, _03356_, _04856_);
  and _25062_ (_03102_, _03357_, _03355_);
  and _25063_ (_03153_, _06816_, _04856_);
  and _25064_ (_03358_, _06705_, _05679_);
  and _25065_ (_03359_, _06688_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  or _25066_ (_03360_, _03359_, _03358_);
  or _25067_ (_03361_, _04861_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  and _25068_ (_03362_, _03361_, _04856_);
  and _25069_ (_03165_, _03362_, _03360_);
  and _25070_ (_03363_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and _25071_ (_03364_, _12165_, \oc8051_top_1.oc8051_rom1.data_o [30]);
  or _25072_ (_03365_, _03364_, _03363_);
  and _25073_ (_03177_, _03365_, _04856_);
  and _25074_ (_03366_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and _25075_ (_03367_, _12165_, \oc8051_top_1.oc8051_rom1.data_o [29]);
  or _25076_ (_03368_, _03367_, _03366_);
  and _25077_ (_03180_, _03368_, _04856_);
  and _25078_ (_03369_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and _25079_ (_03370_, _12165_, \oc8051_top_1.oc8051_rom1.data_o [28]);
  or _25080_ (_03371_, _03370_, _03369_);
  and _25081_ (_03182_, _03371_, _04856_);
  and _25082_ (_03372_, _06598_, _06001_);
  or _25083_ (_03373_, _03372_, _05956_);
  and _25084_ (_03374_, _03373_, _05962_);
  not _25085_ (_03375_, _12131_);
  and _25086_ (_03376_, _03375_, _05995_);
  or _25087_ (_03377_, _03376_, _05961_);
  or _25088_ (_03378_, _03377_, _03374_);
  or _25089_ (_03379_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2], _04859_);
  and _25090_ (_03380_, _03379_, _04856_);
  and _25091_ (_03186_, _03380_, _03378_);
  and _25092_ (_03381_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and _25093_ (_03382_, _12165_, \oc8051_top_1.oc8051_rom1.data_o [27]);
  or _25094_ (_03383_, _03382_, _03381_);
  and _25095_ (_03195_, _03383_, _04856_);
  not _25096_ (_03384_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nor _25097_ (_03385_, _01209_, _03384_);
  and _25098_ (_03386_, _01209_, _03384_);
  or _25099_ (_03388_, _03386_, _03385_);
  or _25100_ (_03389_, _03388_, _12547_);
  and _25101_ (_03390_, _03389_, _04856_);
  nor _25102_ (_03391_, _13091_, _05022_);
  and _25103_ (_03392_, _13091_, _05022_);
  nor _25104_ (_03393_, _03392_, _03391_);
  and _25105_ (_03394_, _03393_, _01185_);
  nand _25106_ (_03395_, _03394_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  or _25107_ (_03396_, _03394_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and _25108_ (_03397_, _03396_, _13031_);
  and _25109_ (_03398_, _03397_, _03395_);
  and _25110_ (_03399_, _13022_, _05507_);
  and _25111_ (_03400_, _06847_, _05641_);
  or _25112_ (_03401_, _01196_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nand _25113_ (_03402_, _01196_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and _25114_ (_03403_, _03402_, _03401_);
  and _25115_ (_03404_, _03403_, _13042_);
  and _25116_ (_03405_, _13036_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and _25117_ (_03406_, _12829_, _13087_);
  or _25118_ (_03407_, _03406_, _03405_);
  or _25119_ (_03408_, _03407_, _03404_);
  or _25120_ (_03409_, _03408_, _03400_);
  nor _25121_ (_03410_, _03409_, _03399_);
  nand _25122_ (_03411_, _03410_, _12547_);
  or _25123_ (_03412_, _03411_, _03398_);
  and _25124_ (_03198_, _03412_, _03390_);
  nor _25125_ (_03200_, _06938_, rst);
  and _25126_ (_03413_, \oc8051_top_1.oc8051_memory_interface1.cdata [7], _08359_);
  and _25127_ (_03414_, \oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or _25128_ (_03415_, _03414_, _03413_);
  and _25129_ (_03202_, _03415_, _04856_);
  nand _25130_ (_03416_, _05730_, _00059_);
  nand _25131_ (_03417_, _03416_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nand _25132_ (_03418_, _03417_, _12206_);
  and _25133_ (_03204_, _03418_, _04856_);
  and _25134_ (_03419_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and _25135_ (_03420_, _12165_, \oc8051_top_1.oc8051_rom1.data_o [26]);
  or _25136_ (_03421_, _03420_, _03419_);
  and _25137_ (_03211_, _03421_, _04856_);
  or _25138_ (_03422_, _06238_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nand _25139_ (_03423_, _06238_, _03238_);
  and _25140_ (_03424_, _03423_, _04856_);
  and _25141_ (_03249_, _03424_, _03422_);
  and _25142_ (_03425_, _06370_, _05000_);
  and _25143_ (_03426_, _05723_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  or _25144_ (_03427_, _03426_, _03425_);
  and _25145_ (_03387_, _03427_, _04856_);
  and _25146_ (_03428_, _01945_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or _25147_ (_03429_, _03428_, _06657_);
  and _25148_ (_03430_, _03429_, _08277_);
  or _25149_ (_03431_, _07949_, _06144_);
  nor _25150_ (_03432_, _07951_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor _25151_ (_03433_, _03432_, _08277_);
  and _25152_ (_03434_, _03433_, _03431_);
  or _25153_ (_03435_, _03434_, _06934_);
  or _25154_ (_03436_, _03435_, _03430_);
  nand _25155_ (_03437_, _06934_, _06284_);
  and _25156_ (_03438_, _03437_, _04856_);
  and _25157_ (_03471_, _03438_, _03436_);
  and _25158_ (_03439_, _06238_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and _25159_ (_03440_, _00957_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  or _25160_ (_03441_, _03440_, _03439_);
  and _25161_ (_03559_, _03441_, _04856_);
  or _25162_ (_03442_, _06757_, _06752_);
  or _25163_ (_03443_, _06787_, _06732_);
  or _25164_ (_03444_, _06777_, _06620_);
  and _25165_ (_03445_, _03444_, _06637_);
  or _25166_ (_03446_, _03445_, _03443_);
  or _25167_ (_03447_, _03446_, _03442_);
  and _25168_ (_03448_, _06777_, _05965_);
  or _25169_ (_03449_, _06835_, _03448_);
  or _25170_ (_03450_, _07508_, _06871_);
  or _25171_ (_03451_, _03450_, _03449_);
  and _25172_ (_03452_, _05998_, _05969_);
  or _25173_ (_03453_, _12689_, _08242_);
  or _25174_ (_03454_, _03453_, _03452_);
  or _25175_ (_03455_, _06786_, _06761_);
  or _25176_ (_03456_, _03455_, _03454_);
  or _25177_ (_03457_, _03456_, _03451_);
  or _25178_ (_03458_, _09071_, _08208_);
  or _25179_ (_03459_, _03458_, _09079_);
  or _25180_ (_03460_, _03459_, _09099_);
  or _25181_ (_03461_, _03460_, _03457_);
  or _25182_ (_03462_, _03461_, _03447_);
  and _25183_ (_03463_, _03462_, _05730_);
  and _25184_ (_03464_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _25185_ (_03465_, _03464_, _03376_);
  or _25186_ (_03466_, _03465_, _03463_);
  and _25187_ (_03577_, _03466_, _04856_);
  nor _25188_ (_03612_, _06947_, rst);
  or _25189_ (_03467_, _08367_, \oc8051_top_1.oc8051_rom1.data_o [13]);
  nand _25190_ (_03468_, _08367_, _05884_);
  and _25191_ (_03469_, _03468_, _04856_);
  and _25192_ (_03641_, _03469_, _03467_);
  and _25193_ (_03470_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and _25194_ (_03472_, _12165_, \oc8051_top_1.oc8051_rom1.data_o [16]);
  or _25195_ (_03473_, _03472_, _03470_);
  and _25196_ (_03643_, _03473_, _04856_);
  or _25197_ (_03474_, _08367_, \oc8051_top_1.oc8051_rom1.data_o [15]);
  nand _25198_ (_03475_, _08367_, _05904_);
  and _25199_ (_03476_, _03475_, _04856_);
  and _25200_ (_03647_, _03476_, _03474_);
  and _25201_ (_03477_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and _25202_ (_03478_, _12165_, \oc8051_top_1.oc8051_rom1.data_o [14]);
  or _25203_ (_03479_, _03478_, _03477_);
  and _25204_ (_03653_, _03479_, _04856_);
  and _25205_ (_03480_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and _25206_ (_03481_, _12165_, \oc8051_top_1.oc8051_rom1.data_o [18]);
  or _25207_ (_03482_, _03481_, _03480_);
  and _25208_ (_03677_, _03482_, _04856_);
  and _25209_ (_03483_, _06041_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  and _25210_ (_03484_, _06043_, _05718_);
  or _25211_ (_03485_, _03484_, _03483_);
  and _25212_ (_03698_, _03485_, _04856_);
  and _25213_ (_03486_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and _25214_ (_03487_, _12165_, \oc8051_top_1.oc8051_rom1.data_o [22]);
  or _25215_ (_03488_, _03487_, _03486_);
  and _25216_ (_03706_, _03488_, _04856_);
  and _25217_ (_03489_, _08037_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  nor _25218_ (_03490_, _07410_, _12633_);
  nor _25219_ (_03491_, _07404_, _02635_);
  or _25220_ (_03492_, _03491_, _03490_);
  and _25221_ (_03493_, _07429_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and _25222_ (_03494_, _07422_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  or _25223_ (_03495_, _03494_, _03493_);
  or _25224_ (_03496_, _03495_, _03492_);
  and _25225_ (_03497_, _07437_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and _25226_ (_03498_, _07442_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  or _25227_ (_03499_, _03498_, _03497_);
  and _25228_ (_03500_, _07449_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  and _25229_ (_03501_, _07455_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  or _25230_ (_03502_, _03501_, _03500_);
  or _25231_ (_03503_, _03502_, _03499_);
  or _25232_ (_03504_, _03503_, _03496_);
  and _25233_ (_03505_, _07466_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  nor _25234_ (_03506_, _07463_, _00611_);
  or _25235_ (_03507_, _03506_, _03505_);
  and _25236_ (_03508_, _07470_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and _25237_ (_03509_, _07473_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  or _25238_ (_03510_, _03509_, _03508_);
  or _25239_ (_03511_, _03510_, _03507_);
  nor _25240_ (_03512_, _07486_, _08073_);
  and _25241_ (_03513_, _07484_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  or _25242_ (_03514_, _03513_, _03512_);
  and _25243_ (_03515_, _07477_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _25244_ (_03516_, _07479_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  or _25245_ (_03517_, _03516_, _03515_);
  or _25246_ (_03518_, _03517_, _03514_);
  or _25247_ (_03519_, _03518_, _03511_);
  or _25248_ (_03520_, _03519_, _03504_);
  and _25249_ (_03521_, _07500_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and _25250_ (_03522_, _08028_, _07223_);
  or _25251_ (_03523_, _03522_, _03521_);
  and _25252_ (_03524_, _07494_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  and _25253_ (_03525_, _07389_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  or _25254_ (_03526_, _03525_, _03524_);
  or _25255_ (_03527_, _03526_, _03523_);
  and _25256_ (_03528_, _01899_, _07539_);
  and _25257_ (_03529_, _01869_, _07507_);
  or _25258_ (_03530_, _03529_, _03528_);
  and _25259_ (_03531_, _01754_, _07547_);
  and _25260_ (_03532_, _01619_, _07552_);
  or _25261_ (_03533_, _03532_, _03531_);
  or _25262_ (_03534_, _03533_, _03530_);
  or _25263_ (_03535_, _03534_, _03527_);
  and _25264_ (_03536_, _07943_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and _25265_ (_03537_, _07561_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  or _25266_ (_03538_, _03537_, _03536_);
  or _25267_ (_03539_, _03538_, _03535_);
  or _25268_ (_03540_, _03539_, _03520_);
  and _25269_ (_03541_, _03540_, _08004_);
  or _25270_ (_03542_, _03541_, _07390_);
  or _25271_ (_03543_, _03542_, _03489_);
  nand _25272_ (_03544_, _07390_, _07815_);
  and _25273_ (_03545_, _03544_, _04856_);
  and _25274_ (_03708_, _03545_, _03543_);
  and _25275_ (_03546_, _08037_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  nor _25276_ (_03547_, _07991_, _04904_);
  nand _25277_ (_03548_, _03547_, _04858_);
  nand _25278_ (_03549_, _07943_, _06661_);
  and _25279_ (_03550_, _07996_, _07997_);
  nand _25280_ (_03551_, _03550_, _06141_);
  and _25281_ (_03552_, _03551_, _03549_);
  and _25282_ (_03553_, _03552_, _03548_);
  nand _25283_ (_03554_, _03553_, _07958_);
  or _25284_ (_03555_, _07404_, _12397_);
  or _25285_ (_03556_, _07410_, _02087_);
  and _25286_ (_03557_, _03556_, _03555_);
  or _25287_ (_03558_, _07428_, _12728_);
  or _25288_ (_03560_, _07420_, _02095_);
  and _25289_ (_03561_, _03560_, _03558_);
  and _25290_ (_03562_, _03561_, _03557_);
  nand _25291_ (_03563_, _07437_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or _25292_ (_03564_, _07441_, _12549_);
  and _25293_ (_03565_, _03564_, _03563_);
  nand _25294_ (_03566_, _07449_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  nand _25295_ (_03567_, _07455_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and _25296_ (_03568_, _03567_, _03566_);
  and _25297_ (_03569_, _03568_, _03565_);
  and _25298_ (_03570_, _03569_, _03562_);
  or _25299_ (_03571_, _07463_, _00334_);
  nand _25300_ (_03572_, _07466_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  and _25301_ (_03573_, _03572_, _03571_);
  or _25302_ (_03574_, _07472_, _00834_);
  nand _25303_ (_03575_, _07470_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and _25304_ (_03576_, _03575_, _03574_);
  and _25305_ (_03578_, _03576_, _03573_);
  or _25306_ (_03579_, _07486_, _09271_);
  nand _25307_ (_03580_, _07484_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  and _25308_ (_03581_, _03580_, _03579_);
  nand _25309_ (_03582_, _07477_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nand _25310_ (_03583_, _07479_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  and _25311_ (_03584_, _03583_, _03582_);
  and _25312_ (_03585_, _03584_, _03581_);
  and _25313_ (_03586_, _03585_, _03578_);
  and _25314_ (_03587_, _03586_, _03570_);
  nand _25315_ (_03588_, _07500_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  or _25316_ (_03589_, _07503_, _07067_);
  and _25317_ (_03590_, _03589_, _03588_);
  or _25318_ (_03591_, _07953_, _08340_);
  or _25319_ (_03592_, _08025_, _01096_);
  and _25320_ (_03593_, _03592_, _03591_);
  and _25321_ (_03595_, _03593_, _03590_);
  nand _25322_ (_03596_, _01862_, _07507_);
  nand _25323_ (_03597_, _01888_, _07539_);
  and _25324_ (_03598_, _03597_, _03596_);
  nand _25325_ (_03599_, _01627_, _07552_);
  nand _25326_ (_03600_, _01729_, _07547_);
  and _25327_ (_03601_, _03600_, _03599_);
  and _25328_ (_03602_, _03601_, _03598_);
  and _25329_ (_03603_, _03602_, _03595_);
  nand _25330_ (_03604_, _07561_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  nand _25331_ (_03605_, _07943_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and _25332_ (_03606_, _03605_, _03604_);
  and _25333_ (_03607_, _03606_, _03603_);
  and _25334_ (_03608_, _03607_, _03587_);
  or _25335_ (_03609_, _03608_, _03554_);
  nand _25336_ (_03610_, _03609_, _08786_);
  or _25337_ (_03611_, _03610_, _03546_);
  nand _25338_ (_03613_, _07390_, _07774_);
  and _25339_ (_03614_, _03613_, _04856_);
  and _25340_ (_03712_, _03614_, _03611_);
  and _25341_ (_03615_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and _25342_ (_03616_, _12165_, \oc8051_top_1.oc8051_rom1.data_o [21]);
  or _25343_ (_03617_, _03616_, _03615_);
  and _25344_ (_03719_, _03617_, _04856_);
  and _25345_ (_03618_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and _25346_ (_03619_, _12165_, \oc8051_top_1.oc8051_rom1.data_o [20]);
  or _25347_ (_03620_, _03619_, _03618_);
  and _25348_ (_03721_, _03620_, _04856_);
  and _25349_ (_03621_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and _25350_ (_03622_, _12165_, \oc8051_top_1.oc8051_rom1.data_o [19]);
  or _25351_ (_03623_, _03622_, _03621_);
  and _25352_ (_03724_, _03623_, _04856_);
  or _25353_ (_03624_, _12720_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  nand _25354_ (_03625_, _12720_, _08794_);
  and _25355_ (_03626_, _03625_, _03624_);
  and _25356_ (_03627_, _03626_, _12715_);
  nor _25357_ (_03628_, _12715_, _05669_);
  or _25358_ (_03629_, _03628_, _03627_);
  and _25359_ (_03726_, _03629_, _04856_);
  or _25360_ (_03630_, _01048_, _06705_);
  or _25361_ (_03631_, _10587_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  and _25362_ (_03632_, _03631_, _04856_);
  and _25363_ (_03728_, _03632_, _03630_);
  and _25364_ (_03633_, _08037_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  or _25365_ (_03634_, _07404_, _03197_);
  or _25366_ (_03635_, _07410_, _12627_);
  and _25367_ (_03636_, _03635_, _03634_);
  or _25368_ (_03637_, _07420_, _12791_);
  or _25369_ (_03638_, _07428_, _12439_);
  and _25370_ (_03639_, _03638_, _03637_);
  and _25371_ (_03640_, _03639_, _03636_);
  nand _25372_ (_03642_, _07437_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or _25373_ (_03644_, _07441_, _12450_);
  and _25374_ (_03645_, _03644_, _03642_);
  nand _25375_ (_03646_, _07449_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  nand _25376_ (_03648_, _07455_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and _25377_ (_03649_, _03648_, _03646_);
  and _25378_ (_03650_, _03649_, _03645_);
  and _25379_ (_03651_, _03650_, _03640_);
  or _25380_ (_03652_, _07463_, _00690_);
  or _25381_ (_03654_, _07465_, _00706_);
  and _25382_ (_03655_, _03654_, _03652_);
  or _25383_ (_03656_, _07472_, _00805_);
  nand _25384_ (_03657_, _07470_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and _25385_ (_03658_, _03657_, _03656_);
  and _25386_ (_03659_, _03658_, _03655_);
  or _25387_ (_03660_, _07486_, _00246_);
  nand _25388_ (_03661_, _07484_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  and _25389_ (_03662_, _03661_, _03660_);
  nand _25390_ (_03663_, _07477_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nand _25391_ (_03664_, _07479_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  and _25392_ (_03665_, _03664_, _03663_);
  and _25393_ (_03666_, _03665_, _03662_);
  and _25394_ (_03667_, _03666_, _03659_);
  and _25395_ (_03668_, _03667_, _03651_);
  nand _25396_ (_03669_, _07500_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  or _25397_ (_03670_, _07503_, _07274_);
  and _25398_ (_03671_, _03670_, _03669_);
  or _25399_ (_03672_, _08025_, _08313_);
  or _25400_ (_03673_, _07953_, _08327_);
  and _25401_ (_03674_, _03673_, _03672_);
  and _25402_ (_03675_, _03674_, _03671_);
  nand _25403_ (_03676_, _01893_, _07539_);
  nand _25404_ (_03678_, _01855_, _07507_);
  and _25405_ (_03679_, _03678_, _03676_);
  nand _25406_ (_03680_, _01740_, _07547_);
  nand _25407_ (_03681_, _01632_, _07552_);
  and _25408_ (_03682_, _03681_, _03680_);
  and _25409_ (_03683_, _03682_, _03679_);
  and _25410_ (_03684_, _03683_, _03675_);
  nand _25411_ (_03685_, _07943_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nand _25412_ (_03686_, _07561_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and _25413_ (_03687_, _03686_, _03685_);
  and _25414_ (_03688_, _03687_, _03684_);
  and _25415_ (_03689_, _03688_, _03668_);
  or _25416_ (_03690_, _03689_, _03554_);
  nand _25417_ (_03691_, _03690_, _08786_);
  or _25418_ (_03692_, _03691_, _03633_);
  nand _25419_ (_03693_, _07390_, _07897_);
  and _25420_ (_03694_, _03693_, _04856_);
  and _25421_ (_03746_, _03694_, _03692_);
  nand _25422_ (_03695_, _10587_, _05669_);
  or _25423_ (_03696_, _10587_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  and _25424_ (_03697_, _03696_, _04856_);
  and _25425_ (_03751_, _03697_, _03695_);
  or _25426_ (_03699_, _08367_, \oc8051_top_1.oc8051_rom1.data_o [3]);
  nand _25427_ (_03700_, _08367_, _05805_);
  and _25428_ (_03701_, _03700_, _04856_);
  and _25429_ (_03754_, _03701_, _03699_);
  or _25430_ (_03702_, _08367_, \oc8051_top_1.oc8051_rom1.data_o [2]);
  nand _25431_ (_03703_, _08367_, _05782_);
  and _25432_ (_03704_, _03703_, _04856_);
  and _25433_ (_03756_, _03704_, _03702_);
  or _25434_ (_03705_, _08367_, \oc8051_top_1.oc8051_rom1.data_o [1]);
  nand _25435_ (_03707_, _08367_, _05824_);
  and _25436_ (_03709_, _03707_, _04856_);
  and _25437_ (_03760_, _03709_, _03705_);
  or _25438_ (_03710_, _08367_, \oc8051_top_1.oc8051_rom1.data_o [0]);
  nand _25439_ (_03711_, _08367_, _05749_);
  and _25440_ (_03713_, _03711_, _04856_);
  and _25441_ (_03763_, _03713_, _03710_);
  and _25442_ (_03714_, _08037_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  and _25443_ (_03715_, _07411_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  nor _25444_ (_03716_, _07404_, _12225_);
  or _25445_ (_03717_, _03716_, _03715_);
  and _25446_ (_03718_, _07422_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and _25447_ (_03720_, _07429_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or _25448_ (_03722_, _03720_, _03718_);
  or _25449_ (_03723_, _03722_, _03717_);
  and _25450_ (_03725_, _07437_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and _25451_ (_03727_, _07442_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  or _25452_ (_03729_, _03727_, _03725_);
  and _25453_ (_03730_, _07449_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and _25454_ (_03731_, _07455_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  or _25455_ (_03732_, _03731_, _03730_);
  or _25456_ (_03733_, _03732_, _03729_);
  or _25457_ (_03734_, _03733_, _03723_);
  nor _25458_ (_03735_, _07463_, _00588_);
  and _25459_ (_03736_, _07466_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  or _25460_ (_03737_, _03736_, _03735_);
  and _25461_ (_03738_, _07470_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and _25462_ (_03739_, _07473_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  or _25463_ (_03740_, _03739_, _03738_);
  or _25464_ (_03741_, _03740_, _03737_);
  and _25465_ (_03742_, _07487_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  and _25466_ (_03743_, _07484_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  or _25467_ (_03744_, _03743_, _03742_);
  and _25468_ (_03745_, _07477_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and _25469_ (_03747_, _07479_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  or _25470_ (_03748_, _03747_, _03745_);
  or _25471_ (_03749_, _03748_, _03744_);
  or _25472_ (_03750_, _03749_, _03741_);
  or _25473_ (_03752_, _03750_, _03734_);
  and _25474_ (_03753_, _08028_, _07310_);
  and _25475_ (_03755_, _07500_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  or _25476_ (_03757_, _03755_, _03753_);
  and _25477_ (_03758_, _07494_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  and _25478_ (_03759_, _07389_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  or _25479_ (_03761_, _03759_, _03758_);
  or _25480_ (_03762_, _03761_, _03757_);
  and _25481_ (_03764_, _01747_, _07547_);
  and _25482_ (_03766_, _01613_, _07552_);
  or _25483_ (_03767_, _03766_, _03764_);
  and _25484_ (_03768_, _01844_, _07507_);
  and _25485_ (_03769_, _01908_, _07539_);
  or _25486_ (_03770_, _03769_, _03768_);
  or _25487_ (_03771_, _03770_, _03767_);
  or _25488_ (_03772_, _03771_, _03762_);
  and _25489_ (_03773_, _07561_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and _25490_ (_03774_, _07943_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or _25491_ (_03775_, _03774_, _03773_);
  or _25492_ (_03776_, _03775_, _03772_);
  or _25493_ (_03777_, _03776_, _03752_);
  and _25494_ (_03778_, _03777_, _08004_);
  or _25495_ (_03780_, _03778_, _07390_);
  or _25496_ (_03781_, _03780_, _03714_);
  nand _25497_ (_03782_, _07390_, _06488_);
  and _25498_ (_03783_, _03782_, _04856_);
  and _25499_ (_03765_, _03783_, _03781_);
  nand _25500_ (_03784_, _12393_, _02095_);
  or _25501_ (_03785_, _12583_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and _25502_ (_03786_, _03785_, _12664_);
  or _25503_ (_03787_, _03786_, _12393_);
  and _25504_ (_03788_, _12423_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and _25505_ (_03790_, _03788_, _12420_);
  or _25506_ (_03792_, _03790_, _03787_);
  and _25507_ (_03793_, _03792_, _03784_);
  or _25508_ (_03794_, _03793_, _12430_);
  nand _25509_ (_03795_, _12430_, _06032_);
  and _25510_ (_03796_, _03795_, _03794_);
  or _25511_ (_03797_, _03796_, _12389_);
  nand _25512_ (_03799_, _12389_, _02087_);
  and _25513_ (_03800_, _03799_, _04856_);
  and _25514_ (_03779_, _03800_, _03797_);
  or _25515_ (_03802_, _08367_, \oc8051_top_1.oc8051_rom1.data_o [5]);
  nand _25516_ (_03804_, _08367_, _05881_);
  and _25517_ (_03806_, _03804_, _04856_);
  and _25518_ (_03789_, _03806_, _03802_);
  or _25519_ (_03807_, _08367_, \oc8051_top_1.oc8051_rom1.data_o [10]);
  nand _25520_ (_03808_, _08367_, _05778_);
  and _25521_ (_03809_, _03808_, _04856_);
  and _25522_ (_03791_, _03809_, _03807_);
  or _25523_ (_03810_, _08367_, \oc8051_top_1.oc8051_rom1.data_o [9]);
  nand _25524_ (_03811_, _08367_, _05834_);
  and _25525_ (_03812_, _03811_, _04856_);
  and _25526_ (_03798_, _03812_, _03810_);
  or _25527_ (_03813_, _08367_, \oc8051_top_1.oc8051_rom1.data_o [8]);
  nand _25528_ (_03814_, _08367_, _05754_);
  and _25529_ (_03815_, _03814_, _04856_);
  and _25530_ (_03801_, _03815_, _03813_);
  or _25531_ (_03816_, _08367_, \oc8051_top_1.oc8051_rom1.data_o [7]);
  nand _25532_ (_03817_, _08367_, _05909_);
  and _25533_ (_03818_, _03817_, _04856_);
  and _25534_ (_03803_, _03818_, _03816_);
  and _25535_ (_03819_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and _25536_ (_03820_, _12165_, \oc8051_top_1.oc8051_rom1.data_o [6]);
  or _25537_ (_03821_, _03820_, _03819_);
  and _25538_ (_03805_, _03821_, _04856_);
  and _25539_ (_03823_, _12423_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and _25540_ (_03824_, _03823_, _12420_);
  and _25541_ (_03825_, _12411_, _12401_);
  or _25542_ (_03826_, _03825_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and _25543_ (_03827_, _03826_, _02296_);
  or _25544_ (_03828_, _03827_, _12393_);
  or _25545_ (_03829_, _03828_, _03824_);
  or _25546_ (_03830_, _12395_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  nand _25547_ (_03831_, _03830_, _03829_);
  nor _25548_ (_03832_, _03831_, _12430_);
  and _25549_ (_03833_, _12430_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or _25550_ (_03834_, _03833_, _12389_);
  or _25551_ (_03835_, _03834_, _03832_);
  or _25552_ (_03836_, _12390_, _06705_);
  and _25553_ (_03837_, _03836_, _04856_);
  and _25554_ (_03822_, _03837_, _03835_);
  and _25555_ (_03838_, _06721_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  or _25556_ (_03839_, _08242_, _06736_);
  and _25557_ (_03840_, _06597_, _05848_);
  or _25558_ (_03841_, _07508_, _03840_);
  or _25559_ (_03842_, _03841_, _03839_);
  and _25560_ (_03843_, _03842_, _05773_);
  or _25561_ (_03844_, _12521_, _06763_);
  or _25562_ (_03845_, _03844_, _06750_);
  or _25563_ (_03846_, _03845_, _06889_);
  or _25564_ (_03847_, _03443_, _08212_);
  or _25565_ (_03848_, _03847_, _03846_);
  or _25566_ (_03849_, _06624_, _06612_);
  and _25567_ (_03850_, _03849_, _05998_);
  or _25568_ (_03851_, _08208_, _03850_);
  or _25569_ (_03852_, _03851_, _09083_);
  or _25570_ (_03853_, _03852_, _06758_);
  or _25571_ (_03854_, _03853_, _03848_);
  or _25572_ (_03855_, _03854_, _03843_);
  and _25573_ (_03856_, _03855_, _06770_);
  or _25574_ (_03857_, _03856_, _03838_);
  and _25575_ (_03858_, _12260_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or _25576_ (_03859_, _03858_, _12183_);
  and _25577_ (_03860_, _04985_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or _25578_ (_03862_, _03860_, _07602_);
  and _25579_ (_03863_, _03862_, _12177_);
  or _25580_ (_03864_, _03863_, _03859_);
  or _25581_ (_03866_, _12185_, _06705_);
  and _25582_ (_03867_, _03866_, _04856_);
  and _25583_ (_03861_, _03867_, _03864_);
  and _25584_ (_03868_, _06238_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nor _25585_ (_03869_, _06238_, _03227_);
  or _25586_ (_03870_, _03869_, _03868_);
  and _25587_ (_03865_, _03870_, _04856_);
  or _25588_ (_03871_, _01401_, _05641_);
  or _25589_ (_03872_, _01361_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and _25590_ (_03873_, _03872_, _05510_);
  and _25591_ (_03874_, _03873_, _03871_);
  and _25592_ (_03875_, _08999_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and _25593_ (_03876_, _01352_, _06268_);
  nand _25594_ (_03877_, _03876_, _06088_);
  or _25595_ (_03878_, _03876_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and _25596_ (_03879_, _03878_, _06093_);
  and _25597_ (_03880_, _03879_, _03877_);
  or _25598_ (_03881_, _03880_, _03875_);
  or _25599_ (_03882_, _03881_, _03874_);
  and _25600_ (_03916_, _03882_, _04856_);
  and _25601_ (_03883_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and _25602_ (_03884_, _03883_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  and _25603_ (_03885_, _03231_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and _25604_ (_03886_, _03885_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  nor _25605_ (_03887_, _03886_, _03884_);
  nor _25606_ (_03888_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and _25607_ (_03889_, _03888_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  and _25608_ (_03890_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _03281_);
  and _25609_ (_03891_, _03890_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  nor _25610_ (_03892_, _03891_, _03889_);
  and _25611_ (_03893_, _03892_, _03887_);
  and _25612_ (_03894_, _03893_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and _25613_ (_03895_, _03888_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  and _25614_ (_03896_, _03890_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  nor _25615_ (_03897_, _03896_, _03895_);
  and _25616_ (_03898_, _03883_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  and _25617_ (_03899_, _03885_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  nor _25618_ (_03900_, _03899_, _03898_);
  and _25619_ (_03901_, _03900_, _03897_);
  and _25620_ (_03902_, _03901_, _06261_);
  nor _25621_ (_03903_, _03902_, _03894_);
  nor _25622_ (_03904_, _03903_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  not _25623_ (_03905_, _03904_);
  and _25624_ (_03906_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _08439_);
  nor _25625_ (_03907_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [6]);
  nor _25626_ (_03908_, _03907_, _03906_);
  nor _25627_ (_03909_, _03908_, _06261_);
  nor _25628_ (_03910_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [2]);
  and _25629_ (_03911_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _09148_);
  nor _25630_ (_03912_, _03911_, _03910_);
  nor _25631_ (_03913_, _03912_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor _25632_ (_03914_, _03913_, _03909_);
  and _25633_ (_03915_, _03914_, _03885_);
  nor _25634_ (_03917_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [5]);
  and _25635_ (_03918_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _08363_);
  nor _25636_ (_03919_, _03918_, _03917_);
  nor _25637_ (_03920_, _03919_, _06261_);
  and _25638_ (_03921_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [9]);
  and _25639_ (_03922_, _06241_, \oc8051_symbolic_cxrom1.regvalid [1]);
  nor _25640_ (_03923_, _03922_, _03921_);
  and _25641_ (_03924_, _03923_, _06261_);
  nor _25642_ (_03925_, _03924_, _03920_);
  and _25643_ (_03926_, _03925_, _03890_);
  nor _25644_ (_03927_, _03926_, _03915_);
  nor _25645_ (_03928_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [7]);
  and _25646_ (_03929_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _08408_);
  nor _25647_ (_03930_, _03929_, _03928_);
  nor _25648_ (_03931_, _03930_, _06261_);
  nor _25649_ (_03932_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [3]);
  nor _25650_ (_03933_, _06241_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor _25651_ (_03934_, _03933_, _03932_);
  nor _25652_ (_03935_, _03934_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor _25653_ (_03936_, _03935_, _03931_);
  and _25654_ (_03937_, _03936_, _03883_);
  and _25655_ (_03938_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _09193_);
  nor _25656_ (_03939_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [4]);
  nor _25657_ (_03940_, _03939_, _03938_);
  nor _25658_ (_03941_, _03940_, _06261_);
  and _25659_ (_03942_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [8]);
  and _25660_ (_03943_, _06241_, \oc8051_symbolic_cxrom1.regvalid [0]);
  nor _25661_ (_03944_, _03943_, _03942_);
  and _25662_ (_03945_, _03944_, _06261_);
  nor _25663_ (_03946_, _03945_, _03941_);
  and _25664_ (_03947_, _03946_, _03888_);
  nor _25665_ (_03948_, _03947_, _03937_);
  and _25666_ (_03949_, _03948_, _03927_);
  and _25667_ (_03950_, _03885_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  and _25668_ (_03951_, _03883_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  nor _25669_ (_03952_, _03951_, _03950_);
  and _25670_ (_03953_, _03888_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  and _25671_ (_03954_, _03890_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  nor _25672_ (_03955_, _03954_, _03953_);
  and _25673_ (_03956_, _03955_, _03952_);
  and _25674_ (_03957_, _03956_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and _25675_ (_03958_, _03888_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  and _25676_ (_03959_, _03890_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  nor _25677_ (_03960_, _03959_, _03958_);
  and _25678_ (_03961_, _03883_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  and _25679_ (_03962_, _03885_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  nor _25680_ (_03963_, _03962_, _03961_);
  and _25681_ (_03964_, _03963_, _03960_);
  and _25682_ (_03965_, _03964_, _06261_);
  nor _25683_ (_03966_, _03965_, _03957_);
  nor _25684_ (_03967_, _03966_, _06241_);
  nor _25685_ (_03968_, _03967_, _03949_);
  and _25686_ (_03969_, _03968_, _03905_);
  nor _25687_ (_03970_, _03969_, _03308_);
  and _25688_ (_03971_, _03969_, _03308_);
  or _25689_ (_03972_, _03971_, _03970_);
  and _25690_ (_03973_, _03883_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  and _25691_ (_03974_, _03885_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  nor _25692_ (_03975_, _03974_, _03973_);
  and _25693_ (_03976_, _03888_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  and _25694_ (_03977_, _03890_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  nor _25695_ (_03978_, _03977_, _03976_);
  and _25696_ (_03979_, _03978_, _03975_);
  and _25697_ (_03980_, _03979_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and _25698_ (_03981_, _03888_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  and _25699_ (_03982_, _03890_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  nor _25700_ (_03983_, _03982_, _03981_);
  and _25701_ (_03984_, _03883_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  and _25702_ (_03985_, _03885_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  nor _25703_ (_03986_, _03985_, _03984_);
  and _25704_ (_03987_, _03986_, _03983_);
  and _25705_ (_03988_, _03987_, _06261_);
  nor _25706_ (_03989_, _03988_, _03980_);
  nor _25707_ (_03990_, _03989_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  not _25708_ (_03991_, _03990_);
  and _25709_ (_03992_, _03885_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  and _25710_ (_03993_, _03883_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  nor _25711_ (_03994_, _03993_, _03992_);
  and _25712_ (_03995_, _03888_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  and _25713_ (_03996_, _03890_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  nor _25714_ (_03997_, _03996_, _03995_);
  and _25715_ (_03998_, _03997_, _03994_);
  and _25716_ (_03999_, _03998_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and _25717_ (_04000_, _03888_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  and _25718_ (_04001_, _03890_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  nor _25719_ (_04002_, _04001_, _04000_);
  and _25720_ (_04003_, _03883_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  and _25721_ (_04004_, _03885_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  nor _25722_ (_04005_, _04004_, _04003_);
  and _25723_ (_04006_, _04005_, _04002_);
  and _25724_ (_04007_, _04006_, _06261_);
  nor _25725_ (_04008_, _04007_, _03999_);
  nor _25726_ (_04009_, _04008_, _06241_);
  nor _25727_ (_04010_, _04009_, _03949_);
  and _25728_ (_04011_, _04010_, _03991_);
  and _25729_ (_04012_, _04011_, _03277_);
  nor _25730_ (_04013_, _04011_, _03277_);
  or _25731_ (_04015_, _04013_, _04012_);
  or _25732_ (_04016_, _04015_, _03972_);
  and _25733_ (_04017_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  and _25734_ (_04018_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  and _25735_ (_04019_, _04018_, _04017_);
  and _25736_ (_04020_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  and _25737_ (_04021_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and _25738_ (_04022_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  and _25739_ (_04023_, _04022_, _04021_);
  and _25740_ (_04024_, _04023_, _04020_);
  and _25741_ (_04025_, _04024_, _04019_);
  and _25742_ (_04026_, _04025_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  nor _25743_ (_04027_, _04025_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  nor _25744_ (_04028_, _04027_, _04026_);
  nand _25745_ (_04029_, _04028_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  or _25746_ (_04030_, _04028_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and _25747_ (_04031_, _04030_, _04029_);
  and _25748_ (_04032_, _03890_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  nor _25749_ (_04033_, _04032_, _06261_);
  and _25750_ (_04034_, _03885_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  and _25751_ (_04035_, _03883_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  and _25752_ (_04036_, _03888_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  or _25753_ (_04037_, _04036_, _04035_);
  nor _25754_ (_04038_, _04037_, _04034_);
  and _25755_ (_04039_, _04038_, _04033_);
  and _25756_ (_04040_, _03883_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  and _25757_ (_04041_, _03885_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  nor _25758_ (_04042_, _04041_, _04040_);
  and _25759_ (_04043_, _03888_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  and _25760_ (_04044_, _03890_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  nor _25761_ (_04045_, _04044_, _04043_);
  and _25762_ (_04046_, _04045_, _04042_);
  and _25763_ (_04047_, _04046_, _06261_);
  nor _25764_ (_04048_, _04047_, _04039_);
  nor _25765_ (_04049_, _04048_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  not _25766_ (_04050_, _04049_);
  and _25767_ (_04051_, _03885_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  and _25768_ (_04052_, _03883_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  nor _25769_ (_04053_, _04052_, _04051_);
  and _25770_ (_04054_, _03888_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  and _25771_ (_04055_, _03890_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  nor _25772_ (_04056_, _04055_, _04054_);
  and _25773_ (_04057_, _04056_, _04053_);
  and _25774_ (_04058_, _04057_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and _25775_ (_04059_, _03888_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  and _25776_ (_04060_, _03890_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  nor _25777_ (_04061_, _04060_, _04059_);
  and _25778_ (_04062_, _03883_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  and _25779_ (_04063_, _03885_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  nor _25780_ (_04064_, _04063_, _04062_);
  and _25781_ (_04066_, _04064_, _04061_);
  and _25782_ (_04067_, _04066_, _06261_);
  nor _25783_ (_04068_, _04067_, _04058_);
  nor _25784_ (_04069_, _04068_, _06241_);
  nor _25785_ (_04070_, _04069_, _03949_);
  and _25786_ (_04071_, _04070_, _04050_);
  and _25787_ (_04072_, _04071_, _02517_);
  nor _25788_ (_04073_, _04071_, _02517_);
  or _25789_ (_04074_, _04073_, _04072_);
  or _25790_ (_04075_, _04074_, _04031_);
  or _25791_ (_04076_, _04075_, _04016_);
  and _25792_ (_04077_, _04026_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor _25793_ (_04078_, _04077_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  and _25794_ (_04079_, _04077_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  nor _25795_ (_04080_, _04079_, _04078_);
  nand _25796_ (_04081_, _04080_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  or _25797_ (_04082_, _04080_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and _25798_ (_04083_, _04082_, _04081_);
  nor _25799_ (_04084_, _04026_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor _25800_ (_04085_, _04084_, _04077_);
  and _25801_ (_04086_, _04085_, _06342_);
  nor _25802_ (_04087_, _04085_, _06342_);
  or _25803_ (_04088_, _04087_, _04086_);
  or _25804_ (_04089_, _04088_, _04083_);
  nor _25805_ (_04090_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  and _25806_ (_04091_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  nor _25807_ (_04092_, _04091_, _04090_);
  and _25808_ (_04093_, _04079_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  or _25809_ (_04094_, _04093_, _04092_);
  nand _25810_ (_04095_, _04093_, _04092_);
  and _25811_ (_04096_, _04095_, _04094_);
  nor _25812_ (_04097_, _04079_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor _25813_ (_04098_, _04097_, _04093_);
  and _25814_ (_04099_, _04098_, _00838_);
  nor _25815_ (_04100_, _04098_, _00838_);
  or _25816_ (_04101_, _04100_, _04099_);
  or _25817_ (_04102_, _04101_, _04096_);
  or _25818_ (_04103_, _04102_, _04089_);
  or _25819_ (_04104_, _04103_, _04076_);
  not _25820_ (_04105_, _03888_);
  and _25821_ (_04106_, _03883_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor _25822_ (_04107_, _04106_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and _25823_ (_04108_, _04106_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _25824_ (_04109_, _04108_, _04107_);
  and _25825_ (_04110_, _04109_, _08363_);
  not _25826_ (_04111_, _03917_);
  nor _25827_ (_04112_, _03883_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor _25828_ (_04113_, _04112_, _04106_);
  and _25829_ (_04114_, _04113_, _04111_);
  not _25830_ (_04115_, _04114_);
  nor _25831_ (_04116_, _04115_, _04110_);
  not _25832_ (_04117_, \oc8051_symbolic_cxrom1.regvalid [1]);
  nor _25833_ (_04118_, _04109_, _04117_);
  and _25834_ (_04119_, _04109_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor _25835_ (_04120_, _04119_, _04118_);
  nor _25836_ (_04121_, _04120_, _04113_);
  nor _25837_ (_04122_, _04121_, _04116_);
  nor _25838_ (_04123_, _04122_, _04105_);
  not _25839_ (_04124_, _04123_);
  not _25840_ (_04125_, _04113_);
  nor _25841_ (_04126_, _04109_, \oc8051_symbolic_cxrom1.regvalid [6]);
  not _25842_ (_04127_, _03890_);
  or _25843_ (_04128_, _03906_, _04127_);
  or _25844_ (_04129_, _04128_, _04126_);
  nor _25845_ (_04130_, _04109_, \oc8051_symbolic_cxrom1.regvalid [4]);
  not _25846_ (_04131_, _03883_);
  or _25847_ (_04132_, _03938_, _04131_);
  or _25848_ (_04133_, _04132_, _04130_);
  and _25849_ (_04134_, _04133_, _04129_);
  or _25850_ (_04135_, _04134_, _04125_);
  not _25851_ (_04136_, _04106_);
  not _25852_ (_04137_, \oc8051_symbolic_cxrom1.regvalid [0]);
  nor _25853_ (_04138_, _04109_, _04137_);
  and _25854_ (_04139_, _04109_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor _25855_ (_04140_, _04139_, _04138_);
  or _25856_ (_04141_, _04140_, _04136_);
  not _25857_ (_04142_, \oc8051_symbolic_cxrom1.regvalid [2]);
  nor _25858_ (_04143_, _04109_, _04142_);
  and _25859_ (_04144_, _04109_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor _25860_ (_04145_, _04144_, _04143_);
  nand _25861_ (_04146_, _04125_, _03890_);
  or _25862_ (_04147_, _04146_, _04145_);
  and _25863_ (_04148_, _04147_, _04141_);
  and _25864_ (_04149_, _04148_, _04135_);
  not _25865_ (_04150_, _03885_);
  and _25866_ (_04151_, _04109_, _08408_);
  not _25867_ (_04152_, _04151_);
  nor _25868_ (_04153_, _03928_, _04125_);
  and _25869_ (_04154_, _04153_, _04152_);
  nor _25870_ (_04155_, _04109_, _08399_);
  and _25871_ (_04156_, _04109_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor _25872_ (_04157_, _04156_, _04155_);
  nor _25873_ (_04158_, _04157_, _04113_);
  nor _25874_ (_04159_, _04158_, _04154_);
  nor _25875_ (_04160_, _04159_, _04150_);
  not _25876_ (_04161_, _04160_);
  and _25877_ (_04162_, _04161_, _04149_);
  and _25878_ (_04163_, _04162_, _04124_);
  and _25879_ (_04164_, _03890_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  and _25880_ (_04165_, _03883_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  nor _25881_ (_04166_, _04165_, _04164_);
  and _25882_ (_04167_, _03885_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  and _25883_ (_04168_, _03888_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  nor _25884_ (_04169_, _04168_, _04167_);
  and _25885_ (_04170_, _04169_, _04166_);
  and _25886_ (_04171_, _04170_, _04125_);
  not _25887_ (_04172_, _04109_);
  and _25888_ (_04173_, _03885_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  and _25889_ (_04174_, _03888_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  nor _25890_ (_04175_, _04174_, _04173_);
  and _25891_ (_04176_, _03890_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  and _25892_ (_04177_, _03883_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  nor _25893_ (_04178_, _04177_, _04176_);
  and _25894_ (_04179_, _04178_, _04175_);
  and _25895_ (_04180_, _04179_, _04113_);
  or _25896_ (_04181_, _04180_, _04172_);
  nor _25897_ (_04182_, _04181_, _04171_);
  and _25898_ (_04183_, _03885_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  and _25899_ (_04184_, _03890_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  nor _25900_ (_04185_, _04184_, _04183_);
  and _25901_ (_04186_, _03888_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  and _25902_ (_04187_, _03883_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  nor _25903_ (_04188_, _04187_, _04186_);
  and _25904_ (_04189_, _04188_, _04185_);
  nor _25905_ (_04190_, _04189_, _04113_);
  and _25906_ (_04191_, _03885_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  and _25907_ (_04192_, _03888_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  nor _25908_ (_04193_, _04192_, _04191_);
  and _25909_ (_04194_, _03890_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  and _25910_ (_04195_, _03883_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  nor _25911_ (_04196_, _04195_, _04194_);
  and _25912_ (_04197_, _04196_, _04193_);
  nor _25913_ (_04198_, _04197_, _04125_);
  or _25914_ (_04199_, _04198_, _04190_);
  and _25915_ (_04200_, _04199_, _04172_);
  nor _25916_ (_04201_, _04200_, _04182_);
  nor _25917_ (_04202_, _04201_, _04163_);
  nand _25918_ (_04203_, _04202_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  or _25919_ (_04204_, _04202_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and _25920_ (_04205_, _04204_, _04203_);
  and _25921_ (_04206_, _03890_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  and _25922_ (_04207_, _03883_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  nor _25923_ (_04208_, _04207_, _04206_);
  and _25924_ (_04209_, _03885_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  and _25925_ (_04210_, _03888_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  nor _25926_ (_04211_, _04210_, _04209_);
  and _25927_ (_04212_, _04211_, _04208_);
  and _25928_ (_04213_, _04212_, _04125_);
  and _25929_ (_04214_, _03890_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  and _25930_ (_04215_, _03883_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  nor _25931_ (_04216_, _04215_, _04214_);
  and _25932_ (_04217_, _03885_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  and _25933_ (_04218_, _03888_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  nor _25934_ (_04219_, _04218_, _04217_);
  and _25935_ (_04220_, _04219_, _04216_);
  and _25936_ (_04221_, _04220_, _04113_);
  or _25937_ (_04222_, _04221_, _04109_);
  nor _25938_ (_04223_, _04222_, _04213_);
  and _25939_ (_04224_, _03890_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and _25940_ (_04225_, _03883_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  nor _25941_ (_04226_, _04225_, _04224_);
  and _25942_ (_04227_, _03885_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and _25943_ (_04228_, _03888_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  nor _25944_ (_04229_, _04228_, _04227_);
  and _25945_ (_04230_, _04229_, _04226_);
  nor _25946_ (_04231_, _04230_, _04113_);
  and _25947_ (_04232_, _03890_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and _25948_ (_04233_, _03883_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  nor _25949_ (_04234_, _04233_, _04232_);
  and _25950_ (_04235_, _03885_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  and _25951_ (_04236_, _03888_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  nor _25952_ (_04237_, _04236_, _04235_);
  and _25953_ (_04238_, _04237_, _04234_);
  nor _25954_ (_04239_, _04238_, _04125_);
  or _25955_ (_04240_, _04239_, _04231_);
  and _25956_ (_04241_, _04240_, _04109_);
  nor _25957_ (_04242_, _04241_, _04223_);
  nor _25958_ (_04243_, _04242_, _04163_);
  and _25959_ (_04244_, _04243_, _03291_);
  nor _25960_ (_04245_, _04243_, _03291_);
  or _25961_ (_04246_, _04245_, _04244_);
  or _25962_ (_04247_, _04246_, _04205_);
  and _25963_ (_04248_, _03890_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  and _25964_ (_04249_, _03883_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  nor _25965_ (_04250_, _04249_, _04248_);
  and _25966_ (_04251_, _03885_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  and _25967_ (_04252_, _03888_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  nor _25968_ (_04253_, _04252_, _04251_);
  and _25969_ (_04254_, _04253_, _04250_);
  and _25970_ (_04255_, _04254_, _04125_);
  and _25971_ (_04256_, _03890_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  and _25972_ (_04257_, _03883_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  nor _25973_ (_04258_, _04257_, _04256_);
  and _25974_ (_04259_, _03885_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  and _25975_ (_04260_, _03888_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  nor _25976_ (_04261_, _04260_, _04259_);
  and _25977_ (_04262_, _04261_, _04258_);
  and _25978_ (_04263_, _04262_, _04113_);
  or _25979_ (_04264_, _04263_, _04109_);
  nor _25980_ (_04265_, _04264_, _04255_);
  and _25981_ (_04266_, _03890_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  and _25982_ (_04267_, _03885_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  nor _25983_ (_04268_, _04267_, _04266_);
  and _25984_ (_04269_, _03888_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  and _25985_ (_04270_, _03883_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  nor _25986_ (_04271_, _04270_, _04269_);
  and _25987_ (_04272_, _04271_, _04268_);
  and _25988_ (_04273_, _04272_, _04125_);
  and _25989_ (_04274_, _03885_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  and _25990_ (_04275_, _03883_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  nor _25991_ (_04276_, _04275_, _04274_);
  and _25992_ (_04277_, _03890_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  and _25993_ (_04278_, _03888_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  nor _25994_ (_04279_, _04278_, _04277_);
  and _25995_ (_04280_, _04279_, _04276_);
  and _25996_ (_04281_, _04280_, _04113_);
  or _25997_ (_04282_, _04281_, _04172_);
  nor _25998_ (_04283_, _04282_, _04273_);
  nor _25999_ (_04284_, _04283_, _04265_);
  nor _26000_ (_04285_, _04284_, _04163_);
  nand _26001_ (_04286_, _04285_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or _26002_ (_04287_, _04285_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _26003_ (_04288_, _04287_, _04286_);
  and _26004_ (_04289_, _03890_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  and _26005_ (_04290_, _03883_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  nor _26006_ (_04291_, _04290_, _04289_);
  and _26007_ (_04292_, _03885_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  and _26008_ (_04293_, _03888_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  nor _26009_ (_04294_, _04293_, _04292_);
  and _26010_ (_04295_, _04294_, _04291_);
  and _26011_ (_04296_, _04295_, _04125_);
  and _26012_ (_04297_, _03885_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  and _26013_ (_04298_, _03888_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  nor _26014_ (_04299_, _04298_, _04297_);
  and _26015_ (_04300_, _03890_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  and _26016_ (_04301_, _03883_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  nor _26017_ (_04302_, _04301_, _04300_);
  and _26018_ (_04303_, _04302_, _04299_);
  and _26019_ (_04304_, _04303_, _04113_);
  nor _26020_ (_04305_, _04304_, _04296_);
  nor _26021_ (_04306_, _04305_, _04172_);
  and _26022_ (_04307_, _03890_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  and _26023_ (_04308_, _03883_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  nor _26024_ (_04309_, _04308_, _04307_);
  and _26025_ (_04310_, _03885_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  and _26026_ (_04311_, _03888_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  nor _26027_ (_04312_, _04311_, _04310_);
  and _26028_ (_04313_, _04312_, _04309_);
  and _26029_ (_04314_, _04313_, _04125_);
  and _26030_ (_04315_, _03890_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  and _26031_ (_04316_, _03888_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  nor _26032_ (_04317_, _04316_, _04315_);
  and _26033_ (_04318_, _03885_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  and _26034_ (_04319_, _03883_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  nor _26035_ (_04320_, _04319_, _04318_);
  and _26036_ (_04321_, _04320_, _04317_);
  and _26037_ (_04322_, _04321_, _04113_);
  nor _26038_ (_04323_, _04322_, _04314_);
  nor _26039_ (_04324_, _04323_, _04109_);
  nor _26040_ (_04325_, _04324_, _04306_);
  not _26041_ (_04326_, _04325_);
  nor _26042_ (_04327_, _04326_, _04163_);
  nor _26043_ (_04328_, _04327_, _02251_);
  and _26044_ (_04329_, _04327_, _02251_);
  or _26045_ (_04330_, _04329_, _04328_);
  or _26046_ (_04331_, _04330_, _04288_);
  or _26047_ (_04332_, _04331_, _04247_);
  and _26048_ (_04333_, _03890_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  and _26049_ (_04334_, _03885_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  nor _26050_ (_04335_, _04334_, _04333_);
  and _26051_ (_04336_, _03888_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  and _26052_ (_04337_, _03883_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  nor _26053_ (_04338_, _04337_, _04336_);
  and _26054_ (_04339_, _04338_, _04335_);
  and _26055_ (_04340_, _04339_, _04125_);
  and _26056_ (_04341_, _03885_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  and _26057_ (_04342_, _03888_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  nor _26058_ (_04343_, _04342_, _04341_);
  and _26059_ (_04344_, _03890_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  and _26060_ (_04345_, _03883_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  nor _26061_ (_04346_, _04345_, _04344_);
  and _26062_ (_04347_, _04346_, _04343_);
  and _26063_ (_04348_, _04347_, _04113_);
  or _26064_ (_04349_, _04348_, _04109_);
  nor _26065_ (_04350_, _04349_, _04340_);
  and _26066_ (_04351_, _03890_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  and _26067_ (_04352_, _03885_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  nor _26068_ (_04353_, _04352_, _04351_);
  and _26069_ (_04354_, _03888_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  and _26070_ (_04355_, _03883_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  nor _26071_ (_04356_, _04355_, _04354_);
  and _26072_ (_04357_, _04356_, _04353_);
  and _26073_ (_04358_, _04357_, _04125_);
  and _26074_ (_04359_, _03890_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  and _26075_ (_04360_, _03883_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  nor _26076_ (_04361_, _04360_, _04359_);
  and _26077_ (_04362_, _03885_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  and _26078_ (_04363_, _03888_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  nor _26079_ (_04364_, _04363_, _04362_);
  and _26080_ (_04365_, _04364_, _04361_);
  and _26081_ (_04366_, _04365_, _04113_);
  or _26082_ (_04367_, _04366_, _04172_);
  nor _26083_ (_04368_, _04367_, _04358_);
  nor _26084_ (_04369_, _04368_, _04350_);
  nor _26085_ (_04370_, _04369_, _04163_);
  and _26086_ (_04371_, _04370_, _03227_);
  nor _26087_ (_04372_, _04370_, _03227_);
  or _26088_ (_04373_, _04372_, _04371_);
  and _26089_ (_04374_, _03890_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  and _26090_ (_04375_, _03883_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  nor _26091_ (_04376_, _04375_, _04374_);
  and _26092_ (_04377_, _03885_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  and _26093_ (_04378_, _03888_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  nor _26094_ (_04379_, _04378_, _04377_);
  and _26095_ (_04380_, _04379_, _04376_);
  and _26096_ (_04381_, _04380_, _04125_);
  and _26097_ (_04382_, _03885_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  and _26098_ (_04383_, _03888_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  nor _26099_ (_04384_, _04383_, _04382_);
  and _26100_ (_04385_, _03890_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  and _26101_ (_04386_, _03883_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  nor _26102_ (_04387_, _04386_, _04385_);
  and _26103_ (_04388_, _04387_, _04384_);
  and _26104_ (_04389_, _04388_, _04113_);
  or _26105_ (_04390_, _04389_, _04172_);
  nor _26106_ (_04391_, _04390_, _04381_);
  and _26107_ (_04392_, _03885_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  and _26108_ (_04393_, _03890_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  nor _26109_ (_04394_, _04393_, _04392_);
  and _26110_ (_04395_, _03888_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  and _26111_ (_04396_, _03883_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  nor _26112_ (_04397_, _04396_, _04395_);
  and _26113_ (_04398_, _04397_, _04394_);
  nor _26114_ (_04399_, _04398_, _04113_);
  and _26115_ (_04400_, _03890_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  and _26116_ (_04401_, _03883_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  nor _26117_ (_04402_, _04401_, _04400_);
  and _26118_ (_04403_, _03885_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  and _26119_ (_04404_, _03888_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  nor _26120_ (_04405_, _04404_, _04403_);
  and _26121_ (_04406_, _04405_, _04402_);
  nor _26122_ (_04407_, _04406_, _04125_);
  or _26123_ (_04408_, _04407_, _04399_);
  and _26124_ (_04409_, _04408_, _04172_);
  nor _26125_ (_04410_, _04409_, _04391_);
  nor _26126_ (_04411_, _04410_, _04163_);
  and _26127_ (_04412_, _04411_, _02015_);
  nor _26128_ (_04413_, _04411_, _02015_);
  or _26129_ (_04414_, _04413_, _04412_);
  or _26130_ (_04415_, _04414_, _04373_);
  and _26131_ (_04416_, _03890_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  and _26132_ (_04417_, _03883_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  nor _26133_ (_04418_, _04417_, _04416_);
  and _26134_ (_04419_, _03885_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  and _26135_ (_04420_, _03888_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  nor _26136_ (_04421_, _04420_, _04419_);
  and _26137_ (_04422_, _04421_, _04418_);
  and _26138_ (_04423_, _04422_, _04125_);
  and _26139_ (_04424_, _03885_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  and _26140_ (_04425_, _03888_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  nor _26141_ (_04426_, _04425_, _04424_);
  and _26142_ (_04427_, _03890_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  and _26143_ (_04428_, _03883_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  nor _26144_ (_04429_, _04428_, _04427_);
  and _26145_ (_04430_, _04429_, _04426_);
  and _26146_ (_04431_, _04430_, _04113_);
  or _26147_ (_04432_, _04431_, _04109_);
  nor _26148_ (_04433_, _04432_, _04423_);
  and _26149_ (_04434_, _03890_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  and _26150_ (_04435_, _03885_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  nor _26151_ (_04436_, _04435_, _04434_);
  and _26152_ (_04437_, _03888_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  and _26153_ (_04438_, _03883_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  nor _26154_ (_04439_, _04438_, _04437_);
  and _26155_ (_04440_, _04439_, _04436_);
  and _26156_ (_04441_, _04440_, _04125_);
  and _26157_ (_04442_, _03890_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  and _26158_ (_04443_, _03883_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  nor _26159_ (_04444_, _04443_, _04442_);
  and _26160_ (_04445_, _03885_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  and _26161_ (_04446_, _03888_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  nor _26162_ (_04447_, _04446_, _04445_);
  and _26163_ (_04448_, _04447_, _04444_);
  and _26164_ (_04449_, _04448_, _04113_);
  or _26165_ (_04450_, _04449_, _04172_);
  nor _26166_ (_04451_, _04450_, _04441_);
  nor _26167_ (_04452_, _04451_, _04433_);
  nor _26168_ (_04453_, _04452_, _04163_);
  and _26169_ (_04454_, _04453_, _03223_);
  nor _26170_ (_04455_, _04453_, _03223_);
  or _26171_ (_04456_, _04455_, _04454_);
  and _26172_ (_04457_, _03890_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  and _26173_ (_04458_, _03885_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  nor _26174_ (_04459_, _04458_, _04457_);
  and _26175_ (_04460_, _03888_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  and _26176_ (_04461_, _03883_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  nor _26177_ (_04462_, _04461_, _04460_);
  and _26178_ (_04463_, _04462_, _04459_);
  and _26179_ (_04464_, _04463_, _04125_);
  and _26180_ (_04465_, _03885_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  and _26181_ (_04466_, _03888_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  nor _26182_ (_04467_, _04466_, _04465_);
  and _26183_ (_04468_, _03890_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  and _26184_ (_04469_, _03883_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  nor _26185_ (_04470_, _04469_, _04468_);
  and _26186_ (_04471_, _04470_, _04467_);
  and _26187_ (_04472_, _04471_, _04113_);
  or _26188_ (_04473_, _04472_, _04109_);
  nor _26189_ (_04474_, _04473_, _04464_);
  and _26190_ (_04475_, _03890_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  and _26191_ (_04476_, _03885_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  nor _26192_ (_04477_, _04476_, _04475_);
  and _26193_ (_04478_, _03888_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  and _26194_ (_04479_, _03883_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  nor _26195_ (_04480_, _04479_, _04478_);
  and _26196_ (_04481_, _04480_, _04477_);
  and _26197_ (_04482_, _04481_, _04125_);
  and _26198_ (_04483_, _03885_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  and _26199_ (_04484_, _03883_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  nor _26200_ (_04485_, _04484_, _04483_);
  and _26201_ (_04486_, _03890_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  and _26202_ (_04487_, _03888_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  nor _26203_ (_04488_, _04487_, _04486_);
  and _26204_ (_04489_, _04488_, _04485_);
  and _26205_ (_04490_, _04489_, _04113_);
  or _26206_ (_04491_, _04490_, _04172_);
  nor _26207_ (_04492_, _04491_, _04482_);
  nor _26208_ (_04493_, _04492_, _04474_);
  nor _26209_ (_04494_, _04493_, _04163_);
  nor _26210_ (_04495_, _04494_, _03238_);
  and _26211_ (_04496_, _04494_, _03238_);
  or _26212_ (_04497_, _04496_, _04495_);
  or _26213_ (_04498_, _04497_, _04456_);
  or _26214_ (_04499_, _04498_, _04415_);
  or _26215_ (_04500_, _04499_, _04332_);
  or _26216_ (_04501_, _04500_, _04104_);
  nor _26217_ (_04502_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  or _26218_ (_04503_, _04502_, _02251_);
  not _26219_ (_04504_, _04503_);
  and _26220_ (_04505_, _04502_, _02251_);
  nor _26221_ (_04506_, _04505_, _04504_);
  nor _26222_ (_04507_, _04503_, _03242_);
  and _26223_ (_04508_, _04503_, _03242_);
  nor _26224_ (_04509_, _04508_, _04507_);
  and _26225_ (_04510_, _04509_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and _26226_ (_04511_, _03242_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or _26227_ (_04512_, _04511_, _04510_);
  and _26228_ (_04513_, _04512_, _04506_);
  not _26229_ (_04514_, _04506_);
  nor _26230_ (_04515_, _04509_, _04142_);
  and _26231_ (_04516_, _04509_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or _26232_ (_04517_, _04516_, _04515_);
  and _26233_ (_04518_, _04517_, _04514_);
  or _26234_ (_04519_, _04518_, _04513_);
  and _26235_ (_04520_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and _26236_ (_04521_, _04520_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  not _26237_ (_04522_, _04521_);
  and _26238_ (_04523_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  or _26239_ (_04524_, _04523_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and _26240_ (_04525_, _04524_, _04522_);
  not _26241_ (_04526_, _04525_);
  nor _26242_ (_04527_, _04521_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _26243_ (_04528_, _04521_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor _26244_ (_04529_, _04528_, _04527_);
  nor _26245_ (_04530_, _04529_, _04137_);
  and _26246_ (_04531_, _04529_, \oc8051_symbolic_cxrom1.regvalid [8]);
  or _26247_ (_04532_, _04531_, _04530_);
  and _26248_ (_04533_, _04532_, _04526_);
  or _26249_ (_04534_, _04529_, \oc8051_symbolic_cxrom1.regvalid [4]);
  or _26250_ (_04535_, _03242_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and _26251_ (_04536_, _04535_, _04525_);
  and _26252_ (_04537_, _04536_, _04534_);
  or _26253_ (_04538_, _04537_, _04533_);
  and _26254_ (_04539_, _04509_, \oc8051_symbolic_cxrom1.regvalid [13]);
  and _26255_ (_04540_, _03242_, \oc8051_symbolic_cxrom1.regvalid [5]);
  or _26256_ (_04541_, _04540_, _04514_);
  or _26257_ (_04542_, _04541_, _04539_);
  nand _26258_ (_04543_, _04509_, _08414_);
  or _26259_ (_04544_, _04509_, \oc8051_symbolic_cxrom1.regvalid [1]);
  and _26260_ (_04545_, _04544_, _04543_);
  or _26261_ (_04546_, _04545_, _04506_);
  and _26262_ (_04547_, _04546_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and _26263_ (_04548_, _04547_, _04542_);
  or _26264_ (_04549_, _03242_, \oc8051_symbolic_cxrom1.regvalid [15]);
  or _26265_ (_04550_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [7]);
  and _26266_ (_04551_, _04550_, _04549_);
  or _26267_ (_04552_, _04551_, _02251_);
  or _26268_ (_04553_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [3]);
  or _26269_ (_04554_, _03242_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and _26270_ (_04555_, _04554_, _04553_);
  or _26271_ (_04556_, _04555_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and _26272_ (_04557_, _04556_, _04552_);
  and _26273_ (_04558_, _04557_, _04548_);
  and _26274_ (_04559_, _04558_, _04538_);
  and _26275_ (_04560_, _04559_, _04519_);
  or _26276_ (_04561_, _04560_, _02020_);
  or _26277_ (_04562_, _04529_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or _26278_ (_04563_, _03242_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and _26279_ (_04564_, _04563_, _04525_);
  and _26280_ (_04565_, _04564_, _04562_);
  or _26281_ (_04566_, _04529_, \oc8051_symbolic_cxrom1.regvalid [2]);
  nand _26282_ (_04567_, _04529_, _09148_);
  and _26283_ (_04568_, _04567_, _04526_);
  and _26284_ (_04569_, _04568_, _04566_);
  or _26285_ (_04570_, _04569_, _04565_);
  or _26286_ (_04571_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [1]);
  or _26287_ (_04572_, _03242_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and _26288_ (_04573_, _04572_, _04571_);
  or _26289_ (_04574_, _04573_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and _26290_ (_04575_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [13]);
  or _26291_ (_04576_, _04575_, _04540_);
  or _26292_ (_04577_, _04576_, _02251_);
  and _26293_ (_04578_, _04577_, _04574_);
  and _26294_ (_04579_, _03242_, \oc8051_symbolic_cxrom1.regvalid [4]);
  and _26295_ (_04580_, _04509_, \oc8051_symbolic_cxrom1.regvalid [12]);
  or _26296_ (_04581_, _04580_, _04579_);
  and _26297_ (_04582_, _04581_, _04506_);
  nor _26298_ (_04583_, _04509_, _04137_);
  and _26299_ (_04584_, _04509_, \oc8051_symbolic_cxrom1.regvalid [8]);
  or _26300_ (_04585_, _04584_, _04583_);
  and _26301_ (_04586_, _04585_, _04514_);
  or _26302_ (_04587_, _04586_, _04582_);
  and _26303_ (_04588_, _04587_, _04578_);
  and _26304_ (_04589_, _04588_, _04570_);
  or _26305_ (_04590_, _04589_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  or _26306_ (_04591_, _04557_, _04548_);
  and _26307_ (_04592_, _04591_, _04590_);
  and _26308_ (_04593_, _04592_, _04561_);
  or _26309_ (_04594_, _04593_, _03291_);
  and _26310_ (_04595_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [14]);
  or _26311_ (_04596_, _04511_, _02251_);
  or _26312_ (_04597_, _04596_, _04595_);
  or _26313_ (_04598_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [2]);
  or _26314_ (_04599_, _03242_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and _26315_ (_04600_, _04599_, _04598_);
  or _26316_ (_04601_, _04600_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and _26317_ (_04602_, _04601_, _04597_);
  and _26318_ (_04603_, _04602_, _02020_);
  or _26319_ (_04604_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [8]);
  or _26320_ (_04605_, _03242_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and _26321_ (_04606_, _04605_, _04520_);
  and _26322_ (_04607_, _04606_, _04604_);
  and _26323_ (_04608_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], _02251_);
  and _26324_ (_04609_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [12]);
  or _26325_ (_04610_, _04609_, _04579_);
  and _26326_ (_04611_, _04610_, _04608_);
  or _26327_ (_04612_, _04611_, _04607_);
  or _26328_ (_04613_, _04612_, _04603_);
  or _26329_ (_04614_, _03242_, \oc8051_symbolic_cxrom1.regvalid [13]);
  or _26330_ (_04615_, _04529_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and _26331_ (_04616_, _04615_, _04614_);
  or _26332_ (_04617_, _04616_, _04526_);
  nand _26333_ (_04618_, _04529_, _08414_);
  or _26334_ (_04619_, _04529_, \oc8051_symbolic_cxrom1.regvalid [1]);
  and _26335_ (_04620_, _04619_, _04618_);
  or _26336_ (_04621_, _04620_, _04525_);
  and _26337_ (_04622_, _04621_, _04617_);
  nor _26338_ (_04623_, _04509_, _08399_);
  and _26339_ (_04624_, _04509_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or _26340_ (_04625_, _04624_, _04623_);
  or _26341_ (_04626_, _04625_, _04506_);
  and _26342_ (_04627_, _04509_, \oc8051_symbolic_cxrom1.regvalid [15]);
  nand _26343_ (_04628_, _03242_, \oc8051_symbolic_cxrom1.regvalid [7]);
  nand _26344_ (_04629_, _04628_, _04506_);
  or _26345_ (_04630_, _04629_, _04627_);
  or _26346_ (_04631_, _04610_, _02251_);
  or _26347_ (_04632_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [0]);
  or _26348_ (_04633_, _03242_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and _26349_ (_04634_, _04633_, _04632_);
  or _26350_ (_04635_, _04634_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and _26351_ (_04636_, _04635_, _02020_);
  and _26352_ (_04637_, _04636_, _04631_);
  and _26353_ (_04638_, _04637_, _04630_);
  and _26354_ (_04639_, _04638_, _04626_);
  and _26355_ (_04640_, _04639_, _04622_);
  nor _26356_ (_04641_, _04529_, _08399_);
  and _26357_ (_04642_, _04529_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or _26358_ (_04643_, _04642_, _04641_);
  or _26359_ (_04644_, _04643_, _04525_);
  or _26360_ (_04645_, _04529_, \oc8051_symbolic_cxrom1.regvalid [7]);
  and _26361_ (_04646_, _04645_, _04549_);
  or _26362_ (_04647_, _04646_, _04526_);
  and _26363_ (_04648_, _04647_, _04644_);
  and _26364_ (_04649_, _04602_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and _26365_ (_04650_, _04649_, _04542_);
  and _26366_ (_04651_, _04650_, _04546_);
  and _26367_ (_04652_, _04651_, _04648_);
  or _26368_ (_04653_, _04652_, _04640_);
  and _26369_ (_04654_, _04653_, _04613_);
  or _26370_ (_04655_, _04654_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _26371_ (_04656_, _03888_, _06261_);
  nor _26372_ (_04657_, _04656_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and _26373_ (_04658_, _04656_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _26374_ (_04659_, _04658_, _04657_);
  or _26375_ (_04660_, _04659_, \oc8051_symbolic_cxrom1.regvalid [7]);
  nand _26376_ (_04661_, _03888_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor _26377_ (_04662_, _04661_, _03929_);
  and _26378_ (_04663_, _04662_, _04660_);
  or _26379_ (_04664_, _04659_, \oc8051_symbolic_cxrom1.regvalid [3]);
  and _26380_ (_04665_, _03888_, _06261_);
  not _26381_ (_04666_, _04659_);
  or _26382_ (_04667_, _04666_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and _26383_ (_04668_, _04667_, _04665_);
  and _26384_ (_04669_, _04668_, _04664_);
  or _26385_ (_04670_, _04669_, _04663_);
  nand _26386_ (_04671_, _04659_, _08363_);
  nor _26387_ (_04672_, _04665_, _04656_);
  and _26388_ (_04673_, _04672_, _04111_);
  and _26389_ (_04674_, _04673_, _04671_);
  not _26390_ (_04675_, _04672_);
  nor _26391_ (_04676_, _04659_, _04117_);
  and _26392_ (_04677_, _04659_, \oc8051_symbolic_cxrom1.regvalid [9]);
  or _26393_ (_04678_, _04677_, _04676_);
  and _26394_ (_04679_, _04678_, _04675_);
  or _26395_ (_04680_, _04679_, _04674_);
  and _26396_ (_04681_, _04680_, _03885_);
  or _26397_ (_04682_, _04681_, _04670_);
  or _26398_ (_04683_, _04659_, \oc8051_symbolic_cxrom1.regvalid [6]);
  nor _26399_ (_04684_, _04675_, _03906_);
  and _26400_ (_04685_, _04684_, _04683_);
  and _26401_ (_04686_, _04659_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor _26402_ (_04687_, _04659_, _04142_);
  or _26403_ (_04688_, _04687_, _04686_);
  and _26404_ (_04689_, _04688_, _04675_);
  or _26405_ (_04690_, _04689_, _04685_);
  and _26406_ (_04691_, _04690_, _03883_);
  or _26407_ (_04692_, _04666_, \oc8051_symbolic_cxrom1.regvalid [8]);
  or _26408_ (_04693_, _04659_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and _26409_ (_04694_, _04693_, _04675_);
  and _26410_ (_04695_, _04694_, _04692_);
  or _26411_ (_04696_, _04659_, \oc8051_symbolic_cxrom1.regvalid [4]);
  nor _26412_ (_04697_, _04675_, _03938_);
  and _26413_ (_04698_, _04697_, _04696_);
  or _26414_ (_04699_, _04698_, _04695_);
  and _26415_ (_04700_, _04699_, _03890_);
  or _26416_ (_04701_, _04700_, _04691_);
  or _26417_ (_04702_, _04701_, _04682_);
  and _26418_ (_04703_, _03885_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  and _26419_ (_04704_, _03890_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  or _26420_ (_04705_, _04704_, _04703_);
  and _26421_ (_04706_, _03883_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  and _26422_ (_04707_, _03888_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  or _26423_ (_04708_, _04707_, _04706_);
  or _26424_ (_04709_, _04708_, _04705_);
  nand _26425_ (_04710_, _03888_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  or _26426_ (_04711_, \oc8051_symbolic_cxrom1.regarray[2] [3], \oc8051_symbolic_cxrom1.regarray[2] [2]);
  nand _26427_ (_04712_, _04711_, _03885_);
  and _26428_ (_04713_, _04712_, _04710_);
  nand _26429_ (_04714_, _03885_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  nand _26430_ (_04715_, _03890_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  and _26431_ (_04716_, _04715_, _04714_);
  and _26432_ (_04717_, _04716_, _04713_);
  nand _26433_ (_04718_, _03883_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  or _26434_ (_04719_, \oc8051_symbolic_cxrom1.regarray[0] [3], \oc8051_symbolic_cxrom1.regarray[0] [2]);
  nand _26435_ (_04720_, _04719_, _03888_);
  and _26436_ (_04721_, _04720_, _04718_);
  or _26437_ (_04722_, \oc8051_symbolic_cxrom1.regarray[3] [3], \oc8051_symbolic_cxrom1.regarray[3] [2]);
  nand _26438_ (_04723_, _04722_, _03883_);
  or _26439_ (_04724_, \oc8051_symbolic_cxrom1.regarray[1] [3], \oc8051_symbolic_cxrom1.regarray[1] [2]);
  nand _26440_ (_04725_, _04724_, _03890_);
  and _26441_ (_04726_, _04725_, _04723_);
  and _26442_ (_04727_, _04726_, _04721_);
  and _26443_ (_04728_, _04727_, _04717_);
  and _26444_ (_04729_, _04728_, _04709_);
  or _26445_ (_04730_, _04729_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and _26446_ (_04731_, _03883_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and _26447_ (_04732_, _03888_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  or _26448_ (_04733_, _04732_, _04731_);
  and _26449_ (_04734_, _03885_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and _26450_ (_04735_, _03890_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  or _26451_ (_04736_, _04735_, _04734_);
  or _26452_ (_04737_, _04736_, _04733_);
  nand _26453_ (_04738_, _03888_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  or _26454_ (_04739_, \oc8051_symbolic_cxrom1.regarray[10] [3], \oc8051_symbolic_cxrom1.regarray[10] [2]);
  nand _26455_ (_04740_, _04739_, _03885_);
  and _26456_ (_04741_, _04740_, _04738_);
  nand _26457_ (_04742_, _03885_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  nand _26458_ (_04743_, _03890_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  and _26459_ (_04744_, _04743_, _04742_);
  and _26460_ (_04745_, _04744_, _04741_);
  nand _26461_ (_04746_, _03883_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  or _26462_ (_04747_, \oc8051_symbolic_cxrom1.regarray[8] [3], \oc8051_symbolic_cxrom1.regarray[8] [2]);
  nand _26463_ (_04748_, _04747_, _03888_);
  and _26464_ (_04749_, _04748_, _04746_);
  or _26465_ (_04750_, \oc8051_symbolic_cxrom1.regarray[11] [3], \oc8051_symbolic_cxrom1.regarray[11] [2]);
  nand _26466_ (_04751_, _04750_, _03883_);
  or _26467_ (_04752_, \oc8051_symbolic_cxrom1.regarray[9] [3], \oc8051_symbolic_cxrom1.regarray[9] [2]);
  nand _26468_ (_04753_, _04752_, _03890_);
  and _26469_ (_04754_, _04753_, _04751_);
  and _26470_ (_04755_, _04754_, _04749_);
  and _26471_ (_04756_, _04755_, _04745_);
  and _26472_ (_04757_, _04756_, _04737_);
  or _26473_ (_04758_, _04757_, _06241_);
  and _26474_ (_04759_, _04758_, _06261_);
  and _26475_ (_04760_, _04759_, _04730_);
  and _26476_ (_04761_, _03885_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  and _26477_ (_04762_, _03890_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  or _26478_ (_04763_, _04762_, _04761_);
  and _26479_ (_04764_, _03883_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  and _26480_ (_04765_, _03888_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  or _26481_ (_04766_, _04765_, _04764_);
  or _26482_ (_04767_, _04766_, _04763_);
  nand _26483_ (_04768_, _03888_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  or _26484_ (_04769_, \oc8051_symbolic_cxrom1.regarray[6] [3], \oc8051_symbolic_cxrom1.regarray[6] [2]);
  nand _26485_ (_04770_, _04769_, _03885_);
  and _26486_ (_04771_, _04770_, _04768_);
  nand _26487_ (_04772_, _03885_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  nand _26488_ (_04773_, _03890_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  and _26489_ (_04774_, _04773_, _04772_);
  and _26490_ (_04775_, _04774_, _04771_);
  nand _26491_ (_04776_, _03883_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  or _26492_ (_04777_, \oc8051_symbolic_cxrom1.regarray[4] [3], \oc8051_symbolic_cxrom1.regarray[4] [2]);
  nand _26493_ (_04778_, _04777_, _03888_);
  and _26494_ (_04779_, _04778_, _04776_);
  or _26495_ (_04780_, \oc8051_symbolic_cxrom1.regarray[7] [3], \oc8051_symbolic_cxrom1.regarray[7] [2]);
  nand _26496_ (_04781_, _04780_, _03883_);
  or _26497_ (_04782_, \oc8051_symbolic_cxrom1.regarray[5] [3], \oc8051_symbolic_cxrom1.regarray[5] [2]);
  nand _26498_ (_04783_, _04782_, _03890_);
  and _26499_ (_04784_, _04783_, _04781_);
  and _26500_ (_04785_, _04784_, _04779_);
  and _26501_ (_04786_, _04785_, _04775_);
  and _26502_ (_04787_, _04786_, _04767_);
  or _26503_ (_04788_, _04787_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and _26504_ (_04789_, _03883_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  and _26505_ (_04790_, _03888_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  or _26506_ (_04791_, _04790_, _04789_);
  and _26507_ (_04792_, _03885_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and _26508_ (_04793_, _03890_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  or _26509_ (_04794_, _04793_, _04792_);
  or _26510_ (_04795_, _04794_, _04791_);
  nand _26511_ (_04796_, _03888_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  or _26512_ (_04797_, \oc8051_symbolic_cxrom1.regarray[14] [3], \oc8051_symbolic_cxrom1.regarray[14] [2]);
  nand _26513_ (_04798_, _04797_, _03885_);
  and _26514_ (_04799_, _04798_, _04796_);
  nand _26515_ (_04800_, _03885_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  nand _26516_ (_04801_, _03890_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  and _26517_ (_04802_, _04801_, _04800_);
  and _26518_ (_04803_, _04802_, _04799_);
  nand _26519_ (_04804_, _03883_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  or _26520_ (_04805_, \oc8051_symbolic_cxrom1.regarray[12] [3], \oc8051_symbolic_cxrom1.regarray[12] [2]);
  nand _26521_ (_04806_, _04805_, _03888_);
  and _26522_ (_04807_, _04806_, _04804_);
  or _26523_ (_04808_, \oc8051_symbolic_cxrom1.regarray[15] [3], \oc8051_symbolic_cxrom1.regarray[15] [2]);
  nand _26524_ (_04809_, _04808_, _03883_);
  or _26525_ (_04810_, \oc8051_symbolic_cxrom1.regarray[13] [3], \oc8051_symbolic_cxrom1.regarray[13] [2]);
  nand _26526_ (_04811_, _04810_, _03890_);
  and _26527_ (_04812_, _04811_, _04809_);
  and _26528_ (_04813_, _04812_, _04807_);
  and _26529_ (_04814_, _04813_, _04803_);
  and _26530_ (_04815_, _04814_, _04795_);
  or _26531_ (_04816_, _04815_, _06241_);
  and _26532_ (_04817_, _04816_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and _26533_ (_04818_, _04817_, _04788_);
  or _26534_ (_04819_, _04818_, _04760_);
  and _26535_ (_04820_, _03936_, _03890_);
  and _26536_ (_04821_, _03940_, _06261_);
  or _26537_ (_04822_, _06241_, \oc8051_symbolic_cxrom1.regvalid [0]);
  or _26538_ (_04823_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [8]);
  and _26539_ (_04824_, _04823_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and _26540_ (_04825_, _04824_, _04822_);
  or _26541_ (_04826_, _04825_, _04821_);
  and _26542_ (_04827_, _04826_, _03885_);
  or _26543_ (_04828_, _04827_, _04820_);
  and _26544_ (_04829_, _03914_, _03888_);
  and _26545_ (_04830_, _03919_, _06261_);
  or _26546_ (_04831_, _06241_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or _26547_ (_04832_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [9]);
  and _26548_ (_04833_, _04832_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and _26549_ (_04834_, _04833_, _04831_);
  or _26550_ (_04835_, _04834_, _04830_);
  and _26551_ (_04836_, _04835_, _03883_);
  or _26552_ (_04837_, _04836_, _04829_);
  or _26553_ (_04838_, _04837_, _04828_);
  nor _26554_ (_04839_, _00957_, first_instr);
  nand _26555_ (_04840_, _04839_, _04838_);
  nor _26556_ (_04841_, _04840_, _03949_);
  nand _26557_ (_04842_, _04841_, _04819_);
  nor _26558_ (_04843_, _04842_, _04163_);
  and _26559_ (_04844_, _04843_, _04702_);
  and _26560_ (_04845_, _04844_, _04655_);
  and _26561_ (_04846_, _04845_, _04594_);
  and _26562_ (property_invalid_ajmp, _04846_, _04501_);
  and _26563_ (_04847_, _00957_, first_instr);
  or _26564_ (_00000_, _04847_, rst);
  dff _26565_ (first_instr, _00000_, clk);
  dff _26566_ (\oc8051_symbolic_cxrom1.regarray[15] [0], _13248_, clk);
  dff _26567_ (\oc8051_symbolic_cxrom1.regarray[15] [1], _13249_, clk);
  dff _26568_ (\oc8051_symbolic_cxrom1.regarray[15] [2], _13250_, clk);
  dff _26569_ (\oc8051_symbolic_cxrom1.regarray[15] [3], _13251_, clk);
  dff _26570_ (\oc8051_symbolic_cxrom1.regarray[15] [4], _13252_, clk);
  dff _26571_ (\oc8051_symbolic_cxrom1.regarray[15] [5], _13253_, clk);
  dff _26572_ (\oc8051_symbolic_cxrom1.regarray[15] [6], _13254_, clk);
  dff _26573_ (\oc8051_symbolic_cxrom1.regarray[15] [7], _13255_, clk);
  dff _26574_ (\oc8051_symbolic_cxrom1.regarray[14] [0], _13246_, clk);
  dff _26575_ (\oc8051_symbolic_cxrom1.regarray[14] [1], _08691_, clk);
  dff _26576_ (\oc8051_symbolic_cxrom1.regarray[14] [2], _08694_, clk);
  dff _26577_ (\oc8051_symbolic_cxrom1.regarray[14] [3], _08697_, clk);
  dff _26578_ (\oc8051_symbolic_cxrom1.regarray[14] [4], _13247_, clk);
  dff _26579_ (\oc8051_symbolic_cxrom1.regarray[14] [5], _08702_, clk);
  dff _26580_ (\oc8051_symbolic_cxrom1.regarray[14] [6], _08705_, clk);
  dff _26581_ (\oc8051_symbolic_cxrom1.regarray[14] [7], _08709_, clk);
  dff _26582_ (\oc8051_symbolic_cxrom1.regarray[13] [0], _13238_, clk);
  dff _26583_ (\oc8051_symbolic_cxrom1.regarray[13] [1], _13239_, clk);
  dff _26584_ (\oc8051_symbolic_cxrom1.regarray[13] [2], _13240_, clk);
  dff _26585_ (\oc8051_symbolic_cxrom1.regarray[13] [3], _13241_, clk);
  dff _26586_ (\oc8051_symbolic_cxrom1.regarray[13] [4], _13242_, clk);
  dff _26587_ (\oc8051_symbolic_cxrom1.regarray[13] [5], _13243_, clk);
  dff _26588_ (\oc8051_symbolic_cxrom1.regarray[13] [6], _13244_, clk);
  dff _26589_ (\oc8051_symbolic_cxrom1.regarray[13] [7], _13245_, clk);
  dff _26590_ (\oc8051_symbolic_cxrom1.regarray[12] [0], _08492_, clk);
  dff _26591_ (\oc8051_symbolic_cxrom1.regarray[12] [1], _08497_, clk);
  dff _26592_ (\oc8051_symbolic_cxrom1.regarray[12] [2], _08499_, clk);
  dff _26593_ (\oc8051_symbolic_cxrom1.regarray[12] [3], _08501_, clk);
  dff _26594_ (\oc8051_symbolic_cxrom1.regarray[12] [4], _08504_, clk);
  dff _26595_ (\oc8051_symbolic_cxrom1.regarray[12] [5], _08508_, clk);
  dff _26596_ (\oc8051_symbolic_cxrom1.regarray[12] [6], _08510_, clk);
  dff _26597_ (\oc8051_symbolic_cxrom1.regarray[12] [7], _08513_, clk);
  dff _26598_ (\oc8051_symbolic_cxrom1.regarray[11] [0], _08374_, clk);
  dff _26599_ (\oc8051_symbolic_cxrom1.regarray[11] [1], _08379_, clk);
  dff _26600_ (\oc8051_symbolic_cxrom1.regarray[11] [2], _08384_, clk);
  dff _26601_ (\oc8051_symbolic_cxrom1.regarray[11] [3], _08388_, clk);
  dff _26602_ (\oc8051_symbolic_cxrom1.regarray[11] [4], _08391_, clk);
  dff _26603_ (\oc8051_symbolic_cxrom1.regarray[11] [5], _08395_, clk);
  dff _26604_ (\oc8051_symbolic_cxrom1.regarray[11] [6], _08400_, clk);
  dff _26605_ (\oc8051_symbolic_cxrom1.regarray[11] [7], _08402_, clk);
  dff _26606_ (\oc8051_symbolic_cxrom1.regarray[10] [0], _08293_, clk);
  dff _26607_ (\oc8051_symbolic_cxrom1.regarray[10] [1], _08297_, clk);
  dff _26608_ (\oc8051_symbolic_cxrom1.regarray[10] [2], _08299_, clk);
  dff _26609_ (\oc8051_symbolic_cxrom1.regarray[10] [3], _08300_, clk);
  dff _26610_ (\oc8051_symbolic_cxrom1.regarray[10] [4], _08301_, clk);
  dff _26611_ (\oc8051_symbolic_cxrom1.regarray[10] [5], _08302_, clk);
  dff _26612_ (\oc8051_symbolic_cxrom1.regarray[10] [6], _08303_, clk);
  dff _26613_ (\oc8051_symbolic_cxrom1.regarray[10] [7], _08307_, clk);
  dff _26614_ (\oc8051_symbolic_cxrom1.regarray[9] [0], _13261_, clk);
  dff _26615_ (\oc8051_symbolic_cxrom1.regarray[9] [1], _13262_, clk);
  dff _26616_ (\oc8051_symbolic_cxrom1.regarray[9] [2], _13263_, clk);
  dff _26617_ (\oc8051_symbolic_cxrom1.regarray[9] [3], _13264_, clk);
  dff _26618_ (\oc8051_symbolic_cxrom1.regarray[9] [4], _13265_, clk);
  dff _26619_ (\oc8051_symbolic_cxrom1.regarray[9] [5], _08227_, clk);
  dff _26620_ (\oc8051_symbolic_cxrom1.regarray[9] [6], _08230_, clk);
  dff _26621_ (\oc8051_symbolic_cxrom1.regarray[9] [7], _08234_, clk);
  dff _26622_ (\oc8051_symbolic_cxrom1.regarray[8] [0], _08129_, clk);
  dff _26623_ (\oc8051_symbolic_cxrom1.regarray[8] [1], _13256_, clk);
  dff _26624_ (\oc8051_symbolic_cxrom1.regarray[8] [2], _13257_, clk);
  dff _26625_ (\oc8051_symbolic_cxrom1.regarray[8] [3], _08141_, clk);
  dff _26626_ (\oc8051_symbolic_cxrom1.regarray[8] [4], _13258_, clk);
  dff _26627_ (\oc8051_symbolic_cxrom1.regarray[8] [5], _13259_, clk);
  dff _26628_ (\oc8051_symbolic_cxrom1.regarray[8] [6], _08148_, clk);
  dff _26629_ (\oc8051_symbolic_cxrom1.regarray[8] [7], _13260_, clk);
  dff _26630_ (\oc8051_symbolic_cxrom1.regarray[7] [0], _08020_, clk);
  dff _26631_ (\oc8051_symbolic_cxrom1.regarray[7] [1], _08023_, clk);
  dff _26632_ (\oc8051_symbolic_cxrom1.regarray[7] [2], _08026_, clk);
  dff _26633_ (\oc8051_symbolic_cxrom1.regarray[7] [3], _08030_, clk);
  dff _26634_ (\oc8051_symbolic_cxrom1.regarray[7] [4], _08035_, clk);
  dff _26635_ (\oc8051_symbolic_cxrom1.regarray[7] [5], _08039_, clk);
  dff _26636_ (\oc8051_symbolic_cxrom1.regarray[7] [6], _08042_, clk);
  dff _26637_ (\oc8051_symbolic_cxrom1.regarray[7] [7], _08045_, clk);
  dff _26638_ (\oc8051_symbolic_cxrom1.regarray[6] [0], _07923_, clk);
  dff _26639_ (\oc8051_symbolic_cxrom1.regarray[6] [1], _07926_, clk);
  dff _26640_ (\oc8051_symbolic_cxrom1.regarray[6] [2], _07930_, clk);
  dff _26641_ (\oc8051_symbolic_cxrom1.regarray[6] [3], _07934_, clk);
  dff _26642_ (\oc8051_symbolic_cxrom1.regarray[6] [4], _07938_, clk);
  dff _26643_ (\oc8051_symbolic_cxrom1.regarray[6] [5], _07941_, clk);
  dff _26644_ (\oc8051_symbolic_cxrom1.regarray[6] [6], _07946_, clk);
  dff _26645_ (\oc8051_symbolic_cxrom1.regarray[6] [7], _07950_, clk);
  dff _26646_ (\oc8051_symbolic_cxrom1.regarray[5] [0], _07827_, clk);
  dff _26647_ (\oc8051_symbolic_cxrom1.regarray[5] [1], _07830_, clk);
  dff _26648_ (\oc8051_symbolic_cxrom1.regarray[5] [2], _07834_, clk);
  dff _26649_ (\oc8051_symbolic_cxrom1.regarray[5] [3], _07839_, clk);
  dff _26650_ (\oc8051_symbolic_cxrom1.regarray[5] [4], _07844_, clk);
  dff _26651_ (\oc8051_symbolic_cxrom1.regarray[5] [5], _07849_, clk);
  dff _26652_ (\oc8051_symbolic_cxrom1.regarray[5] [6], _07852_, clk);
  dff _26653_ (\oc8051_symbolic_cxrom1.regarray[5] [7], _07856_, clk);
  dff _26654_ (\oc8051_symbolic_cxrom1.regarray[1] [0], _07413_, clk);
  dff _26655_ (\oc8051_symbolic_cxrom1.regarray[1] [1], _07416_, clk);
  dff _26656_ (\oc8051_symbolic_cxrom1.regarray[1] [2], _07419_, clk);
  dff _26657_ (\oc8051_symbolic_cxrom1.regarray[1] [3], _07421_, clk);
  dff _26658_ (\oc8051_symbolic_cxrom1.regarray[1] [4], _07423_, clk);
  dff _26659_ (\oc8051_symbolic_cxrom1.regarray[1] [5], _07427_, clk);
  dff _26660_ (\oc8051_symbolic_cxrom1.regarray[1] [6], _07431_, clk);
  dff _26661_ (\oc8051_symbolic_cxrom1.regarray[1] [7], _07434_, clk);
  dff _26662_ (\oc8051_symbolic_cxrom1.regarray[0] [0], _07298_, clk);
  dff _26663_ (\oc8051_symbolic_cxrom1.regarray[0] [1], _07302_, clk);
  dff _26664_ (\oc8051_symbolic_cxrom1.regarray[0] [2], _07307_, clk);
  dff _26665_ (\oc8051_symbolic_cxrom1.regarray[0] [3], _07313_, clk);
  dff _26666_ (\oc8051_symbolic_cxrom1.regarray[0] [4], _07318_, clk);
  dff _26667_ (\oc8051_symbolic_cxrom1.regarray[0] [5], _07324_, clk);
  dff _26668_ (\oc8051_symbolic_cxrom1.regarray[0] [6], _07329_, clk);
  dff _26669_ (\oc8051_symbolic_cxrom1.regarray[0] [7], _07332_, clk);
  dff _26670_ (\oc8051_symbolic_cxrom1.regarray[3] [0], _07608_, clk);
  dff _26671_ (\oc8051_symbolic_cxrom1.regarray[3] [1], _07611_, clk);
  dff _26672_ (\oc8051_symbolic_cxrom1.regarray[3] [2], _07615_, clk);
  dff _26673_ (\oc8051_symbolic_cxrom1.regarray[3] [3], _07618_, clk);
  dff _26674_ (\oc8051_symbolic_cxrom1.regarray[3] [4], _07623_, clk);
  dff _26675_ (\oc8051_symbolic_cxrom1.regarray[3] [5], _07627_, clk);
  dff _26676_ (\oc8051_symbolic_cxrom1.regarray[3] [6], _07630_, clk);
  dff _26677_ (\oc8051_symbolic_cxrom1.regarray[3] [7], _07635_, clk);
  dff _26678_ (\oc8051_symbolic_cxrom1.regarray[2] [0], _07517_, clk);
  dff _26679_ (\oc8051_symbolic_cxrom1.regarray[2] [1], _07520_, clk);
  dff _26680_ (\oc8051_symbolic_cxrom1.regarray[2] [2], _07524_, clk);
  dff _26681_ (\oc8051_symbolic_cxrom1.regarray[2] [3], _07529_, clk);
  dff _26682_ (\oc8051_symbolic_cxrom1.regarray[2] [4], _07534_, clk);
  dff _26683_ (\oc8051_symbolic_cxrom1.regarray[2] [5], _07537_, clk);
  dff _26684_ (\oc8051_symbolic_cxrom1.regarray[2] [6], _07540_, clk);
  dff _26685_ (\oc8051_symbolic_cxrom1.regarray[2] [7], _07543_, clk);
  dff _26686_ (\oc8051_symbolic_cxrom1.regarray[4] [0], _07728_, clk);
  dff _26687_ (\oc8051_symbolic_cxrom1.regarray[4] [1], _07731_, clk);
  dff _26688_ (\oc8051_symbolic_cxrom1.regarray[4] [2], _07734_, clk);
  dff _26689_ (\oc8051_symbolic_cxrom1.regarray[4] [3], _07738_, clk);
  dff _26690_ (\oc8051_symbolic_cxrom1.regarray[4] [4], _07742_, clk);
  dff _26691_ (\oc8051_symbolic_cxrom1.regarray[4] [5], _07745_, clk);
  dff _26692_ (\oc8051_symbolic_cxrom1.regarray[4] [6], _07747_, clk);
  dff _26693_ (\oc8051_symbolic_cxrom1.regarray[4] [7], _07750_, clk);
  dff _26694_ (\oc8051_symbolic_cxrom1.regvalid [0], _05859_, clk);
  dff _26695_ (\oc8051_symbolic_cxrom1.regvalid [1], _05887_, clk);
  dff _26696_ (\oc8051_symbolic_cxrom1.regvalid [2], _05931_, clk);
  dff _26697_ (\oc8051_symbolic_cxrom1.regvalid [3], _05981_, clk);
  dff _26698_ (\oc8051_symbolic_cxrom1.regvalid [4], _06031_, clk);
  dff _26699_ (\oc8051_symbolic_cxrom1.regvalid [5], _06085_, clk);
  dff _26700_ (\oc8051_symbolic_cxrom1.regvalid [6], _06158_, clk);
  dff _26701_ (\oc8051_symbolic_cxrom1.regvalid [7], _06239_, clk);
  dff _26702_ (\oc8051_symbolic_cxrom1.regvalid [8], _06315_, clk);
  dff _26703_ (\oc8051_symbolic_cxrom1.regvalid [9], _06394_, clk);
  dff _26704_ (\oc8051_symbolic_cxrom1.regvalid [10], _06484_, clk);
  dff _26705_ (\oc8051_symbolic_cxrom1.regvalid [11], _06577_, clk);
  dff _26706_ (\oc8051_symbolic_cxrom1.regvalid [12], _06683_, clk);
  dff _26707_ (\oc8051_symbolic_cxrom1.regvalid [13], _06785_, clk);
  dff _26708_ (\oc8051_symbolic_cxrom1.regvalid [14], _06896_, clk);
  dff _26709_ (\oc8051_symbolic_cxrom1.regvalid [15], _05809_, clk);
  dff _26710_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [0], _05508_, clk);
  dff _26711_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [1], _05511_, clk);
  dff _26712_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [2], _05514_, clk);
  dff _26713_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [3], _05516_, clk);
  dff _26714_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [4], _05518_, clk);
  dff _26715_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [5], _05521_, clk);
  dff _26716_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [6], _05523_, clk);
  dff _26717_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [7], _05358_, clk);
  dff _26718_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [0], _12317_, clk);
  dff _26719_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [1], _11174_, clk);
  dff _26720_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [2], _11150_, clk);
  dff _26721_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [4], _12621_, clk);
  dff _26722_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [5], _12736_, clk);
  dff _26723_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [6], _11754_, clk);
  dff _26724_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [7], _05361_, clk);
  dff _26725_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [0], _11428_, clk);
  dff _26726_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [3], _11426_, clk);
  dff _26727_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [4], _11595_, clk);
  dff _26728_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [5], _11638_, clk);
  dff _26729_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [6], _10883_, clk);
  dff _26730_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [7], _05364_, clk);
  dff _26731_ (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], _09788_, clk);
  dff _26732_ (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], _09822_, clk);
  dff _26733_ (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], _03153_, clk);
  dff _26734_ (\oc8051_top_1.oc8051_decoder1.mem_act [0], _09794_, clk);
  dff _26735_ (\oc8051_top_1.oc8051_decoder1.mem_act [1], _09820_, clk);
  dff _26736_ (\oc8051_top_1.oc8051_decoder1.mem_act [2], _05116_, clk);
  dff _26737_ (\oc8051_top_1.oc8051_decoder1.state [0], _09810_, clk);
  dff _26738_ (\oc8051_top_1.oc8051_decoder1.state [1], _05182_, clk);
  dff _26739_ (\oc8051_top_1.oc8051_decoder1.op [0], _09813_, clk);
  dff _26740_ (\oc8051_top_1.oc8051_decoder1.op [1], _09782_, clk);
  dff _26741_ (\oc8051_top_1.oc8051_decoder1.op [2], _09513_, clk);
  dff _26742_ (\oc8051_top_1.oc8051_decoder1.op [3], _09521_, clk);
  dff _26743_ (\oc8051_top_1.oc8051_decoder1.op [4], _09529_, clk);
  dff _26744_ (\oc8051_top_1.oc8051_decoder1.op [5], _09806_, clk);
  dff _26745_ (\oc8051_top_1.oc8051_decoder1.op [6], _09791_, clk);
  dff _26746_ (\oc8051_top_1.oc8051_decoder1.op [7], _03062_, clk);
  dff _26747_ (\oc8051_top_1.oc8051_decoder1.src_sel3 , _05222_, clk);
  dff _26748_ (\oc8051_top_1.oc8051_decoder1.wr_sfr [0], _03577_, clk);
  dff _26749_ (\oc8051_top_1.oc8051_decoder1.wr_sfr [1], _05127_, clk);
  dff _26750_ (\oc8051_top_1.oc8051_decoder1.src_sel2 [0], _03857_, clk);
  dff _26751_ (\oc8051_top_1.oc8051_decoder1.src_sel2 [1], _05136_, clk);
  dff _26752_ (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _03594_, clk);
  dff _26753_ (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _04891_, clk);
  dff _26754_ (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], _05200_, clk);
  dff _26755_ (\oc8051_top_1.oc8051_decoder1.src_sel1 [0], _06447_, clk);
  dff _26756_ (\oc8051_top_1.oc8051_decoder1.src_sel1 [1], _07107_, clk);
  dff _26757_ (\oc8051_top_1.oc8051_decoder1.src_sel1 [2], _03186_, clk);
  dff _26758_ (\oc8051_top_1.oc8051_decoder1.cy_sel [0], _10443_, clk);
  dff _26759_ (\oc8051_top_1.oc8051_decoder1.cy_sel [1], _05219_, clk);
  dff _26760_ (\oc8051_top_1.oc8051_decoder1.alu_op [0], _11805_, clk);
  dff _26761_ (\oc8051_top_1.oc8051_decoder1.alu_op [1], _11945_, clk);
  dff _26762_ (\oc8051_top_1.oc8051_decoder1.alu_op [2], _12372_, clk);
  dff _26763_ (\oc8051_top_1.oc8051_decoder1.alu_op [3], _05113_, clk);
  dff _26764_ (\oc8051_top_1.oc8051_decoder1.psw_set [0], _00498_, clk);
  dff _26765_ (\oc8051_top_1.oc8051_decoder1.psw_set [1], _05311_, clk);
  dff _26766_ (\oc8051_top_1.oc8051_decoder1.wr , _05302_, clk);
  dff _26767_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [0], _08362_, clk);
  dff _26768_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [1], _08582_, clk);
  dff _26769_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [2], _03728_, clk);
  dff _26770_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [3], _03751_, clk);
  dff _26771_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [4], _12673_, clk);
  dff _26772_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [5], _03102_, clk);
  dff _26773_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [6], _01805_, clk);
  dff _26774_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [7], _02847_, clk);
  dff _26775_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [0], _00041_, clk);
  dff _26776_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [1], _06640_, clk);
  dff _26777_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [2], _04854_, clk);
  dff _26778_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [3], _12147_, clk);
  dff _26779_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [4], _00574_, clk);
  dff _26780_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [5], _12445_, clk);
  dff _26781_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [6], _12690_, clk);
  dff _26782_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [7], _02839_, clk);
  dff _26783_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [0], _01824_, clk);
  dff _26784_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [1], _01776_, clk);
  dff _26785_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [2], _02968_, clk);
  dff _26786_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [3], _02983_, clk);
  dff _26787_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [4], _03074_, clk);
  dff _26788_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [5], _01037_, clk);
  dff _26789_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [6], _02869_, clk);
  dff _26790_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [7], _02864_, clk);
  dff _26791_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [0], _10893_, clk);
  dff _26792_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [1], _08283_, clk);
  dff _26793_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [2], _03165_, clk);
  dff _26794_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [3], _07837_, clk);
  dff _26795_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [4], _05251_, clk);
  dff _26796_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [5], _09073_, clk);
  dff _26797_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [6], _04065_, clk);
  dff _26798_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [7], _02877_, clk);
  dff _26799_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [0], _07842_, clk);
  dff _26800_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [1], _04849_, clk);
  dff _26801_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [2], _09492_, clk);
  dff _26802_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [3], _04850_, clk);
  dff _26803_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [4], _08879_, clk);
  dff _26804_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [5], _09831_, clk);
  dff _26805_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [6], _03190_, clk);
  dff _26806_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [7], _01437_, clk);
  dff _26807_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [0], _03387_, clk);
  dff _26808_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [1], _04970_, clk);
  dff _26809_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [2], _04855_, clk);
  dff _26810_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [3], _01669_, clk);
  dff _26811_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [4], _05203_, clk);
  dff _26812_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [5], _04852_, clk);
  dff _26813_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [6], _06909_, clk);
  dff _26814_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [7], _02804_, clk);
  dff _26815_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [0], _01432_, clk);
  dff _26816_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [1], _05235_, clk);
  dff _26817_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [2], _04853_, clk);
  dff _26818_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [3], _01710_, clk);
  dff _26819_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [4], _01517_, clk);
  dff _26820_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [5], _03698_, clk);
  dff _26821_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [6], _01955_, clk);
  dff _26822_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [7], _02792_, clk);
  dff _26823_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [0], _13213_, clk);
  dff _26824_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [1], _04983_, clk);
  dff _26825_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [2], _10214_, clk);
  dff _26826_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [3], _08279_, clk);
  dff _26827_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [4], _01547_, clk);
  dff _26828_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [5], _01164_, clk);
  dff _26829_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [6], _13054_, clk);
  dff _26830_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [7], _02887_, clk);
  dff _26831_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [0], _11042_, clk);
  dff _26832_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [1], _10850_, clk);
  dff _26833_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [2], _12211_, clk);
  dff _26834_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [3], _03612_, clk);
  dff _26835_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [4], _03200_, clk);
  dff _26836_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [0], _02913_, clk);
  dff _26837_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [1], _01158_, clk);
  dff _26838_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [2], _01812_, clk);
  dff _26839_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [3], _02836_, clk);
  dff _26840_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [4], _03865_, clk);
  dff _26841_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [5], _01154_, clk);
  dff _26842_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [6], _02833_, clk);
  dff _26843_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [7], _02906_, clk);
  dff _26844_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [8], _02950_, clk);
  dff _26845_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [9], _02964_, clk);
  dff _26846_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [10], _02378_, clk);
  dff _26847_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [11], _01427_, clk);
  dff _26848_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [12], _02829_, clk);
  dff _26849_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [13], _04851_, clk);
  dff _26850_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [14], _02749_, clk);
  dff _26851_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [15], _12274_, clk);
  dff _26852_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _02816_, clk);
  dff _26853_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _02898_, clk);
  dff _26854_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _09528_, clk);
  dff _26855_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _09192_, clk);
  dff _26856_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _02813_, clk);
  dff _26857_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _02235_, clk);
  dff _26858_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _03249_, clk);
  dff _26859_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _02809_, clk);
  dff _26860_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _02896_, clk);
  dff _26861_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _02946_, clk);
  dff _26862_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _02962_, clk);
  dff _26863_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _03559_, clk);
  dff _26864_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _12295_, clk);
  dff _26865_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _02806_, clk);
  dff _26866_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _12154_, clk);
  dff _26867_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _12267_, clk);
  dff _26868_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [0], _03763_, clk);
  dff _26869_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [1], _03760_, clk);
  dff _26870_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [2], _03756_, clk);
  dff _26871_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [3], _03754_, clk);
  dff _26872_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [4], _12234_, clk);
  dff _26873_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [5], _03789_, clk);
  dff _26874_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [6], _03805_, clk);
  dff _26875_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [7], _03803_, clk);
  dff _26876_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [8], _03801_, clk);
  dff _26877_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [9], _03798_, clk);
  dff _26878_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [10], _03791_, clk);
  dff _26879_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [11], _12229_, clk);
  dff _26880_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [12], _10908_, clk);
  dff _26881_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [13], _03641_, clk);
  dff _26882_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [14], _03653_, clk);
  dff _26883_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [15], _03647_, clk);
  dff _26884_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [16], _03643_, clk);
  dff _26885_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [17], _12251_, clk);
  dff _26886_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [18], _03677_, clk);
  dff _26887_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [19], _03724_, clk);
  dff _26888_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [20], _03721_, clk);
  dff _26889_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [21], _03719_, clk);
  dff _26890_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [22], _03706_, clk);
  dff _26891_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [23], _12239_, clk);
  dff _26892_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [24], _10902_, clk);
  dff _26893_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [25], _11055_, clk);
  dff _26894_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [26], _03211_, clk);
  dff _26895_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [27], _03195_, clk);
  dff _26896_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [28], _03182_, clk);
  dff _26897_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [29], _03180_, clk);
  dff _26898_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [30], _03177_, clk);
  dff _26899_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [31], _09996_, clk);
  dff _26900_ (\oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _10265_, clk);
  dff _26901_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [0], _01964_, clk);
  dff _26902_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [1], _01962_, clk);
  dff _26903_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [2], _01960_, clk);
  dff _26904_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [3], _01953_, clk);
  dff _26905_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [4], _12303_, clk);
  dff _26906_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [5], _02776_, clk);
  dff _26907_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [6], _02751_, clk);
  dff _26908_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [7], _10297_, clk);
  dff _26909_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [3], _12646_, clk);
  dff _26910_ (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _10310_, clk);
  dff _26911_ (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _10301_, clk);
  dff _26912_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [0], _00137_, clk);
  dff _26913_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [1], _00196_, clk);
  dff _26914_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _00177_, clk);
  dff _26915_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [3], _00157_, clk);
  dff _26916_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [4], _12338_, clk);
  dff _26917_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [5], _10869_, clk);
  dff _26918_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [6], _10866_, clk);
  dff _26919_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [7], _10919_, clk);
  dff _26920_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [8], _10911_, clk);
  dff _26921_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [9], _10889_, clk);
  dff _26922_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [10], _12343_, clk);
  dff _26923_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [11], _13165_, clk);
  dff _26924_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [12], _13203_, clk);
  dff _26925_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [13], _13196_, clk);
  dff _26926_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [14], _13188_, clk);
  dff _26927_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [15], _03198_, clk);
  dff _26928_ (\oc8051_top_1.oc8051_memory_interface1.pc [0], _12702_, clk);
  dff _26929_ (\oc8051_top_1.oc8051_memory_interface1.pc [1], _12670_, clk);
  dff _26930_ (\oc8051_top_1.oc8051_memory_interface1.pc [2], _11543_, clk);
  dff _26931_ (\oc8051_top_1.oc8051_memory_interface1.pc [3], _11522_, clk);
  dff _26932_ (\oc8051_top_1.oc8051_memory_interface1.pc [4], _11467_, clk);
  dff _26933_ (\oc8051_top_1.oc8051_memory_interface1.pc [5], _11443_, clk);
  dff _26934_ (\oc8051_top_1.oc8051_memory_interface1.pc [6], _11435_, clk);
  dff _26935_ (\oc8051_top_1.oc8051_memory_interface1.pc [7], _12712_, clk);
  dff _26936_ (\oc8051_top_1.oc8051_memory_interface1.pc [8], _11646_, clk);
  dff _26937_ (\oc8051_top_1.oc8051_memory_interface1.pc [9], _11624_, clk);
  dff _26938_ (\oc8051_top_1.oc8051_memory_interface1.pc [10], _11618_, clk);
  dff _26939_ (\oc8051_top_1.oc8051_memory_interface1.pc [11], _11616_, clk);
  dff _26940_ (\oc8051_top_1.oc8051_memory_interface1.pc [12], _11610_, clk);
  dff _26941_ (\oc8051_top_1.oc8051_memory_interface1.pc [13], _11605_, clk);
  dff _26942_ (\oc8051_top_1.oc8051_memory_interface1.pc [14], _12706_, clk);
  dff _26943_ (\oc8051_top_1.oc8051_memory_interface1.pc [15], _03001_, clk);
  dff _26944_ (\oc8051_top_1.oc8051_memory_interface1.int_ack , _10135_, clk);
  dff _26945_ (\oc8051_top_1.oc8051_memory_interface1.int_ack_t , _03204_, clk);
  dff _26946_ (\oc8051_top_1.oc8051_memory_interface1.int_ack_buff , _10114_, clk);
  dff _26947_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], _12694_, clk);
  dff _26948_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], _12679_, clk);
  dff _26949_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _10992_, clk);
  dff _26950_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], _12093_, clk);
  dff _26951_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _12750_, clk);
  dff _26952_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], _11327_, clk);
  dff _26953_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _11312_, clk);
  dff _26954_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _10174_, clk);
  dff _26955_ (\oc8051_top_1.oc8051_memory_interface1.op_pos [0], _11058_, clk);
  dff _26956_ (\oc8051_top_1.oc8051_memory_interface1.op_pos [1], _11089_, clk);
  dff _26957_ (\oc8051_top_1.oc8051_memory_interface1.op_pos [2], _10221_, clk);
  dff _26958_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [1], _11801_, clk);
  dff _26959_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [2], _11792_, clk);
  dff _26960_ (\oc8051_top_1.oc8051_memory_interface1.reti , _10190_, clk);
  dff _26961_ (\oc8051_top_1.oc8051_memory_interface1.cdata [0], _11856_, clk);
  dff _26962_ (\oc8051_top_1.oc8051_memory_interface1.cdata [1], _11848_, clk);
  dff _26963_ (\oc8051_top_1.oc8051_memory_interface1.cdata [2], _11412_, clk);
  dff _26964_ (\oc8051_top_1.oc8051_memory_interface1.cdata [3], _11579_, clk);
  dff _26965_ (\oc8051_top_1.oc8051_memory_interface1.cdata [4], _11630_, clk);
  dff _26966_ (\oc8051_top_1.oc8051_memory_interface1.cdata [5], _11658_, clk);
  dff _26967_ (\oc8051_top_1.oc8051_memory_interface1.cdata [6], _11883_, clk);
  dff _26968_ (\oc8051_top_1.oc8051_memory_interface1.cdata [7], _03202_, clk);
  dff _26969_ (\oc8051_top_1.oc8051_memory_interface1.cdone , _02999_, clk);
  dff _26970_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst , _03067_, clk);
  dff _26971_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], _11914_, clk);
  dff _26972_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], _11904_, clk);
  dff _26973_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], _11406_, clk);
  dff _26974_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], _03097_, clk);
  dff _26975_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [0], _11704_, clk);
  dff _26976_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [1], _11476_, clk);
  dff _26977_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [2], _11715_, clk);
  dff _26978_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [3], _11710_, clk);
  dff _26979_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [4], _11464_, clk);
  dff _26980_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [5], _11602_, clk);
  dff _26981_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [6], _11726_, clk);
  dff _26982_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [7], _11720_, clk);
  dff _26983_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [8], _11451_, clk);
  dff _26984_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [9], _11751_, clk);
  dff _26985_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [10], _11736_, clk);
  dff _26986_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [11], _11439_, clk);
  dff _26987_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [12], _11598_, clk);
  dff _26988_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [13], _11641_, clk);
  dff _26989_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [14], _11984_, clk);
  dff _26990_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [15], _11979_, clk);
  dff _26991_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [16], _11370_, clk);
  dff _26992_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [17], _11995_, clk);
  dff _26993_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [18], _11993_, clk);
  dff _26994_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [19], _11357_, clk);
  dff _26995_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [20], _11565_, clk);
  dff _26996_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [21], _12006_, clk);
  dff _26997_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [22], _12001_, clk);
  dff _26998_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [23], _11355_, clk);
  dff _26999_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [24], _12040_, clk);
  dff _27000_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [25], _12011_, clk);
  dff _27001_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [26], _11347_, clk);
  dff _27002_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [27], _11620_, clk);
  dff _27003_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [28], _12049_, clk);
  dff _27004_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [29], _12042_, clk);
  dff _27005_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [30], _11343_, clk);
  dff _27006_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [31], _09984_, clk);
  dff _27007_ (\oc8051_top_1.oc8051_memory_interface1.dmem_wait , _10072_, clk);
  dff _27008_ (\oc8051_top_1.oc8051_memory_interface1.istb_t , _10067_, clk);
  dff _27009_ (\oc8051_top_1.oc8051_memory_interface1.imem_wait , _10060_, clk);
  dff _27010_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _11247_, clk);
  dff _27011_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _12300_, clk);
  dff _27012_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _12280_, clk);
  dff _27013_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _11236_, clk);
  dff _27014_ (\oc8051_top_1.oc8051_memory_interface1.rd_ind , _10047_, clk);
  dff _27015_ (\oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0], clk);
  dff _27016_ (\oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1], clk);
  dff _27017_ (\oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2], clk);
  dff _27018_ (\oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3], clk);
  dff _27019_ (\oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4], clk);
  dff _27020_ (\oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5], clk);
  dff _27021_ (\oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6], clk);
  dff _27022_ (\oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7], clk);
  dff _27023_ (\oc8051_top_1.oc8051_rom1.data_o [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8], clk);
  dff _27024_ (\oc8051_top_1.oc8051_rom1.data_o [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9], clk);
  dff _27025_ (\oc8051_top_1.oc8051_rom1.data_o [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10], clk);
  dff _27026_ (\oc8051_top_1.oc8051_rom1.data_o [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11], clk);
  dff _27027_ (\oc8051_top_1.oc8051_rom1.data_o [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12], clk);
  dff _27028_ (\oc8051_top_1.oc8051_rom1.data_o [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13], clk);
  dff _27029_ (\oc8051_top_1.oc8051_rom1.data_o [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14], clk);
  dff _27030_ (\oc8051_top_1.oc8051_rom1.data_o [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15], clk);
  dff _27031_ (\oc8051_top_1.oc8051_rom1.data_o [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16], clk);
  dff _27032_ (\oc8051_top_1.oc8051_rom1.data_o [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17], clk);
  dff _27033_ (\oc8051_top_1.oc8051_rom1.data_o [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18], clk);
  dff _27034_ (\oc8051_top_1.oc8051_rom1.data_o [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19], clk);
  dff _27035_ (\oc8051_top_1.oc8051_rom1.data_o [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20], clk);
  dff _27036_ (\oc8051_top_1.oc8051_rom1.data_o [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21], clk);
  dff _27037_ (\oc8051_top_1.oc8051_rom1.data_o [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22], clk);
  dff _27038_ (\oc8051_top_1.oc8051_rom1.data_o [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23], clk);
  dff _27039_ (\oc8051_top_1.oc8051_rom1.data_o [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24], clk);
  dff _27040_ (\oc8051_top_1.oc8051_rom1.data_o [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25], clk);
  dff _27041_ (\oc8051_top_1.oc8051_rom1.data_o [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26], clk);
  dff _27042_ (\oc8051_top_1.oc8051_rom1.data_o [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27], clk);
  dff _27043_ (\oc8051_top_1.oc8051_rom1.data_o [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28], clk);
  dff _27044_ (\oc8051_top_1.oc8051_rom1.data_o [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29], clk);
  dff _27045_ (\oc8051_top_1.oc8051_rom1.data_o [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30], clk);
  dff _27046_ (\oc8051_top_1.oc8051_rom1.data_o [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31], clk);
  dff _27047_ (\oc8051_top_1.oc8051_sfr1.pres_ow , _02340_, clk);
  dff _27048_ (\oc8051_top_1.oc8051_sfr1.prescaler [0], _11844_, clk);
  dff _27049_ (\oc8051_top_1.oc8051_sfr1.prescaler [1], _11292_, clk);
  dff _27050_ (\oc8051_top_1.oc8051_sfr1.prescaler [2], _12580_, clk);
  dff _27051_ (\oc8051_top_1.oc8051_sfr1.prescaler [3], _00307_, clk);
  dff _27052_ (\oc8051_top_1.oc8051_sfr1.bit_out , _00670_, clk);
  dff _27053_ (\oc8051_top_1.oc8051_sfr1.wait_data , _02424_, clk);
  dff _27054_ (\oc8051_top_1.oc8051_sfr1.dat0 [0], _05133_, clk);
  dff _27055_ (\oc8051_top_1.oc8051_sfr1.dat0 [1], _03712_, clk);
  dff _27056_ (\oc8051_top_1.oc8051_sfr1.dat0 [2], _06111_, clk);
  dff _27057_ (\oc8051_top_1.oc8051_sfr1.dat0 [3], _05975_, clk);
  dff _27058_ (\oc8051_top_1.oc8051_sfr1.dat0 [4], _03708_, clk);
  dff _27059_ (\oc8051_top_1.oc8051_sfr1.dat0 [5], _03746_, clk);
  dff _27060_ (\oc8051_top_1.oc8051_sfr1.dat0 [6], _03765_, clk);
  dff _27061_ (\oc8051_top_1.oc8051_sfr1.dat0 [7], _02393_, clk);
  dff _27062_ (\oc8051_top_1.oc8051_sfr1.wr_bit_r , _01644_, clk);
  dff _27063_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], _01147_, clk);
  dff _27064_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], _01317_, clk);
  dff _27065_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], _06465_, clk);
  dff _27066_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3], _08881_, clk);
  dff _27067_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4], _01115_, clk);
  dff _27068_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], _01110_, clk);
  dff _27069_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], _01112_, clk);
  dff _27070_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], _04014_, clk);
  dff _27071_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0], _00209_, clk);
  dff _27072_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1], _00205_, clk);
  dff _27073_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2], _02637_, clk);
  dff _27074_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3], _00144_, clk);
  dff _27075_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4], _00130_, clk);
  dff _27076_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5], _02655_, clk);
  dff _27077_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6], _00168_, clk);
  dff _27078_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7], _03916_, clk);
  dff _27079_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], _05691_, clk);
  dff _27080_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], _05706_, clk);
  dff _27081_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], _05712_, clk);
  dff _27082_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], _05709_, clk);
  dff _27083_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], _05697_, clk);
  dff _27084_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], _05695_, clk);
  dff _27085_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], _02380_, clk);
  dff _27086_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7], _03221_, clk);
  dff _27087_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0], _13064_, clk);
  dff _27088_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1], _12951_, clk);
  dff _27089_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2], _02954_, clk);
  dff _27090_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3], _03036_, clk);
  dff _27091_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4], _05575_, clk);
  dff _27092_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5], _05566_, clk);
  dff _27093_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6], _02512_, clk);
  dff _27094_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7], _04848_, clk);
  dff _27095_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff , _10675_, clk);
  dff _27096_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], _01846_, clk);
  dff _27097_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], _01851_, clk);
  dff _27098_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _01849_, clk);
  dff _27099_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3], _01796_, clk);
  dff _27100_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4], _01817_, clk);
  dff _27101_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], _01856_, clk);
  dff _27102_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _01853_, clk);
  dff _27103_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _10459_, clk);
  dff _27104_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], _01859_, clk);
  dff _27105_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _09163_, clk);
  dff _27106_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc , _10162_, clk);
  dff _27107_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _01943_, clk);
  dff _27108_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _01931_, clk);
  dff _27109_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], _10318_, clk);
  dff _27110_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _01599_, clk);
  dff _27111_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _01808_, clk);
  dff _27112_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], _09318_, clk);
  dff _27113_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], _01597_, clk);
  dff _27114_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _01593_, clk);
  dff _27115_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , _10816_, clk);
  dff _27116_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , _08683_, clk);
  dff _27117_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , _08562_, clk);
  dff _27118_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , _10480_, clk);
  dff _27119_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0], _01803_, clk);
  dff _27120_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1], _02022_, clk);
  dff _27121_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2], _02016_, clk);
  dff _27122_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], _08584_, clk);
  dff _27123_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0], _02036_, clk);
  dff _27124_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], _01580_, clk);
  dff _27125_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], _02049_, clk);
  dff _27126_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3], _02042_, clk);
  dff _27127_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4], _01570_, clk);
  dff _27128_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5], _01801_, clk);
  dff _27129_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6], _02054_, clk);
  dff _27130_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _10217_, clk);
  dff _27131_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0], _02062_, clk);
  dff _27132_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1], _01563_, clk);
  dff _27133_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2], _02082_, clk);
  dff _27134_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3], _02072_, clk);
  dff _27135_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4], _01559_, clk);
  dff _27136_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5], _01799_, clk);
  dff _27137_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6], _02091_, clk);
  dff _27138_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7], _10339_, clk);
  dff _27139_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0], _02688_, clk);
  dff _27140_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1], _02673_, clk);
  dff _27141_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2], _02670_, clk);
  dff _27142_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3], _02575_, clk);
  dff _27143_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4], _02545_, clk);
  dff _27144_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5], _02720_, clk);
  dff _27145_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6], _02577_, clk);
  dff _27146_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7], _06167_, clk);
  dff _27147_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0], _02693_, clk);
  dff _27148_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1], _02691_, clk);
  dff _27149_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2], _02726_, clk);
  dff _27150_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3], _02573_, clk);
  dff _27151_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4], _02724_, clk);
  dff _27152_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5], _02697_, clk);
  dff _27153_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6], _02543_, clk);
  dff _27154_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7], _06247_, clk);
  dff _27155_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0], _02664_, clk);
  dff _27156_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1], _02662_, clk);
  dff _27157_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2], _02627_, clk);
  dff _27158_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3], _02625_, clk);
  dff _27159_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4], _02552_, clk);
  dff _27160_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5], _02728_, clk);
  dff _27161_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6], _02588_, clk);
  dff _27162_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7], _06472_, clk);
  dff _27163_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0], _02590_, clk);
  dff _27164_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1], _02712_, clk);
  dff _27165_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2], _02555_, clk);
  dff _27166_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3], _02710_, clk);
  dff _27167_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4], _02592_, clk);
  dff _27168_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5], _02558_, clk);
  dff _27169_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6], _02708_, clk);
  dff _27170_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7], _06467_, clk);
  dff _27171_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1], _09036_, clk);
  dff _27172_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], _02548_, clk);
  dff _27173_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3], _11350_, clk);
  dff _27174_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4], _11718_, clk);
  dff _27175_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5], _05539_, clk);
  dff _27176_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6], _05505_, clk);
  dff _27177_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], _03471_, clk);
  dff _27178_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], _02798_, clk);
  dff _27179_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], _12496_, clk);
  dff _27180_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2], _12482_, clk);
  dff _27181_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3], _12493_, clk);
  dff _27182_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4], _12491_, clk);
  dff _27183_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5], _12489_, clk);
  dff _27184_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6], _12485_, clk);
  dff _27185_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7], _02763_, clk);
  dff _27186_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop , _12819_, clk);
  dff _27187_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , _00150_, clk);
  dff _27188_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff , _00140_, clk);
  dff _27189_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0], _12017_, clk);
  dff _27190_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1], _12014_, clk);
  dff _27191_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2], _12032_, clk);
  dff _27192_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3], _12038_, clk);
  dff _27193_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4], _12035_, clk);
  dff _27194_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], _12082_, clk);
  dff _27195_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6], _12077_, clk);
  dff _27196_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7], _00133_, clk);
  dff _27197_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0], _12156_, clk);
  dff _27198_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1], _12151_, clk);
  dff _27199_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2], _12128_, clk);
  dff _27200_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3], _12130_, clk);
  dff _27201_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4], _12135_, clk);
  dff _27202_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5], _12137_, clk);
  dff _27203_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6], _12119_, clk);
  dff _27204_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7], _00121_, clk);
  dff _27205_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , _00126_, clk);
  dff _27206_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _00124_, clk);
  dff _27207_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0], _12163_, clk);
  dff _27208_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1], _12173_, clk);
  dff _27209_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2], _12169_, clk);
  dff _27210_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3], _12172_, clk);
  dff _27211_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4], _12184_, clk);
  dff _27212_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], _12178_, clk);
  dff _27213_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6], _12181_, clk);
  dff _27214_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7], _00115_, clk);
  dff _27215_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0], _11910_, clk);
  dff _27216_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1], _11907_, clk);
  dff _27217_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2], _11897_, clk);
  dff _27218_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3], _11900_, clk);
  dff _27219_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4], _11888_, clk);
  dff _27220_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5], _11891_, clk);
  dff _27221_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6], _11877_, clk);
  dff _27222_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7], _00116_, clk);
  dff _27223_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 , _00170_, clk);
  dff _27224_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _11930_, clk);
  dff _27225_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], _11924_, clk);
  dff _27226_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2], _11927_, clk);
  dff _27227_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3], _11830_, clk);
  dff _27228_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _11825_, clk);
  dff _27229_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], _11729_, clk);
  dff _27230_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6], _11723_, clk);
  dff _27231_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7], _00165_, clk);
  dff _27232_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r , _01494_, clk);
  dff _27233_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _01415_, clk);
  dff _27234_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , _01412_, clk);
  dff _27235_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r , _01406_, clk);
  dff _27236_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0], _12255_, clk);
  dff _27237_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1], _01586_, clk);
  dff _27238_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2], _10547_, clk);
  dff _27239_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3], _10566_, clk);
  dff _27240_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4], _10557_, clk);
  dff _27241_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5], _10553_, clk);
  dff _27242_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6], _10549_, clk);
  dff _27243_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7], _01397_, clk);
  dff _27244_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0], _10478_, clk);
  dff _27245_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1], _10473_, clk);
  dff _27246_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2], _10471_, clk);
  dff _27247_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3], _03726_, clk);
  dff _27248_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4], _10499_, clk);
  dff _27249_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5], _10514_, clk);
  dff _27250_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6], _10507_, clk);
  dff _27251_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7], _01066_, clk);
  dff _27252_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 , _01031_, clk);
  dff _27253_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0], _10374_, clk);
  dff _27254_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1], _03779_, clk);
  dff _27255_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2], _10434_, clk);
  dff _27256_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3], _10427_, clk);
  dff _27257_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4], _10424_, clk);
  dff _27258_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5], _10419_, clk);
  dff _27259_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6], _10416_, clk);
  dff _27260_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7], _01044_, clk);
  dff _27261_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0], _10344_, clk);
  dff _27262_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1], _10337_, clk);
  dff _27263_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2], _03822_, clk);
  dff _27264_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3], _01884_, clk);
  dff _27265_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4], _10257_, clk);
  dff _27266_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5], _10250_, clk);
  dff _27267_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6], _10247_, clk);
  dff _27268_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7], _01040_, clk);
  dff _27269_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set , _01023_, clk);
  dff _27270_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0], _10146_, clk);
  dff _27271_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1], _10143_, clk);
  dff _27272_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2], _03861_, clk);
  dff _27273_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3], _10208_, clk);
  dff _27274_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], _10202_, clk);
  dff _27275_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], _10199_, clk);
  dff _27276_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6], _10193_, clk);
  dff _27277_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], _01020_, clk);
  dff _27278_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0], _02936_, clk);
  dff _27279_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1], _02208_, clk);
  dff _27280_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2], _10761_, clk);
  dff _27281_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _08118_, clk);
  dff _27282_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _05143_, clk);
  dff _27283_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _12141_, clk);
  dff _27284_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _02925_, clk);
  dff _27285_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _02520_, clk);
  dff _27286_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8], _02503_, clk);
  dff _27287_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9], _02452_, clk);
  dff _27288_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], _10531_, clk);
  dff _27289_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _02486_, clk);
  dff _27290_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf , _02941_, clk);
  dff _27291_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , _02988_, clk);
  dff _27292_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , _02787_, clk);
  dff _27293_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive , _02782_, clk);
  dff _27294_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _02740_, clk);
  dff _27295_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r , _02771_, clk);
  dff _27296_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], _00865_, clk);
  dff _27297_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1], _02756_, clk);
  dff _27298_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], _01051_, clk);
  dff _27299_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], _06914_, clk);
  dff _27300_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _01508_, clk);
  dff _27301_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3], _02560_, clk);
  dff _27302_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0], _06954_, clk);
  dff _27303_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1], _01583_, clk);
  dff _27304_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2], _01557_, clk);
  dff _27305_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3], _01791_, clk);
  dff _27306_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4], _01785_, clk);
  dff _27307_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5], _01829_, clk);
  dff _27308_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6], _01794_, clk);
  dff _27309_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7], _02550_, clk);
  dff _27310_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr , _02483_, clk);
  dff _27311_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr , _02481_, clk);
  dff _27312_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans , _02198_, clk);
  dff _27313_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , _02159_, clk);
  dff _27314_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0], _02239_, clk);
  dff _27315_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1], _02224_, clk);
  dff _27316_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2], _02408_, clk);
  dff _27317_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3], _02137_, clk);
  dff _27318_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0], _06884_, clk);
  dff _27319_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1], _06945_, clk);
  dff _27320_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], _02454_, clk);
  dff _27321_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3], _02438_, clk);
  dff _27322_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4], _06881_, clk);
  dff _27323_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5], _02668_, clk);
  dff _27324_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6], _02461_, clk);
  dff _27325_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7], _06942_, clk);
  dff _27326_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8], _06975_, clk);
  dff _27327_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], _02768_, clk);
  dff _27328_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10], _01924_, clk);
  dff _27329_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0], _02883_, clk);
  dff _27330_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1], _02860_, clk);
  dff _27331_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2], _06874_, clk);
  dff _27332_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3], _06939_, clk);
  dff _27333_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4], _02923_, clk);
  dff _27334_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5], _02911_, clk);
  dff _27335_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6], _02934_, clk);
  dff _27336_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], _01920_, clk);
  dff _27337_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0], _11698_, clk);
  dff _27338_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], _06933_, clk);
  dff _27339_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2], _13158_, clk);
  dff _27340_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3], _13002_, clk);
  dff _27341_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], _13205_, clk);
  dff _27342_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5], _13168_, clk);
  dff _27343_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6], _06927_, clk);
  dff _27344_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], _01903_, clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_for_ajmp [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_out [0], \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_out [1], \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [0], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [3], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [4], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [5], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [6], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [7], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [0], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [1], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [2], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [3], \oc8051_top_1.oc8051_memory_interface1.imm_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [4], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [5], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [6], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [7], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [0], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [1], \oc8051_top_1.oc8051_memory_interface1.op3_buff [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [2], \oc8051_top_1.oc8051_memory_interface1.op3_buff [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [3], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [4], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [5], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [6], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [7], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [0], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [1], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [2], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [4], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [5], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [6], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [7], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [0], ABINPUT[1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [1], ABINPUT[2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [2], ABINPUT[3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [3], ABINPUT[4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [4], ABINPUT[5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [5], ABINPUT[6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [6], ABINPUT[7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [7], ABINPUT[8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.oc8051_memory_interface1.bit_in , ABINPUT[0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.rst , rst);
  buf(\oc8051_top_1.oc8051_memory_interface1.clk , clk);
  buf(\oc8051_top_1.oc8051_indi_addr1.wr_bit_r , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_indi_addr1.rst , rst);
  buf(\oc8051_top_1.oc8051_indi_addr1.clk , clk);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.oc8051_rom1.clk , clk);
  buf(\oc8051_top_1.oc8051_rom1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.oc8051_decoder1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.oc8051_sfr1.ip [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_decoder1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_sfr1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_decoder1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_alu_src_sel1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [3], \oc8051_top_1.oc8051_memory_interface1.imm_r [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3_r [1], \oc8051_top_1.oc8051_memory_interface1.op3_buff [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3_r [2], \oc8051_top_1.oc8051_memory_interface1.op3_buff [2]);
  buf(\oc8051_top_1.oc8051_sfr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.rst , rst);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_in , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_symbolic_cxrom1.clk , clk);
  buf(\oc8051_symbolic_cxrom1.rst , rst);
  buf(\oc8051_symbolic_cxrom1.word_in [0], word_in[0]);
  buf(\oc8051_symbolic_cxrom1.word_in [1], word_in[1]);
  buf(\oc8051_symbolic_cxrom1.word_in [2], word_in[2]);
  buf(\oc8051_symbolic_cxrom1.word_in [3], word_in[3]);
  buf(\oc8051_symbolic_cxrom1.word_in [4], word_in[4]);
  buf(\oc8051_symbolic_cxrom1.word_in [5], word_in[5]);
  buf(\oc8051_symbolic_cxrom1.word_in [6], word_in[6]);
  buf(\oc8051_symbolic_cxrom1.word_in [7], word_in[7]);
  buf(\oc8051_symbolic_cxrom1.word_in [8], word_in[8]);
  buf(\oc8051_symbolic_cxrom1.word_in [9], word_in[9]);
  buf(\oc8051_symbolic_cxrom1.word_in [10], word_in[10]);
  buf(\oc8051_symbolic_cxrom1.word_in [11], word_in[11]);
  buf(\oc8051_symbolic_cxrom1.word_in [12], word_in[12]);
  buf(\oc8051_symbolic_cxrom1.word_in [13], word_in[13]);
  buf(\oc8051_symbolic_cxrom1.word_in [14], word_in[14]);
  buf(\oc8051_symbolic_cxrom1.word_in [15], word_in[15]);
  buf(\oc8051_symbolic_cxrom1.word_in [16], word_in[16]);
  buf(\oc8051_symbolic_cxrom1.word_in [17], word_in[17]);
  buf(\oc8051_symbolic_cxrom1.word_in [18], word_in[18]);
  buf(\oc8051_symbolic_cxrom1.word_in [19], word_in[19]);
  buf(\oc8051_symbolic_cxrom1.word_in [20], word_in[20]);
  buf(\oc8051_symbolic_cxrom1.word_in [21], word_in[21]);
  buf(\oc8051_symbolic_cxrom1.word_in [22], word_in[22]);
  buf(\oc8051_symbolic_cxrom1.word_in [23], word_in[23]);
  buf(\oc8051_symbolic_cxrom1.word_in [24], word_in[24]);
  buf(\oc8051_symbolic_cxrom1.word_in [25], word_in[25]);
  buf(\oc8051_symbolic_cxrom1.word_in [26], word_in[26]);
  buf(\oc8051_symbolic_cxrom1.word_in [27], word_in[27]);
  buf(\oc8051_symbolic_cxrom1.word_in [28], word_in[28]);
  buf(\oc8051_symbolic_cxrom1.word_in [29], word_in[29]);
  buf(\oc8051_symbolic_cxrom1.word_in [30], word_in[30]);
  buf(\oc8051_symbolic_cxrom1.word_in [31], word_in[31]);
  buf(\oc8051_symbolic_cxrom1.pc1 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc1 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_symbolic_cxrom1.pc1 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_symbolic_cxrom1.pc1 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_symbolic_cxrom1.pc1 [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_symbolic_cxrom1.pc1 [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_symbolic_cxrom1.pc1 [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_symbolic_cxrom1.pc1 [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_symbolic_cxrom1.pc1 [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_symbolic_cxrom1.pc1 [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_symbolic_cxrom1.pc1 [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_symbolic_cxrom1.pc1 [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_symbolic_cxrom1.pc1 [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_symbolic_cxrom1.pc1 [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_symbolic_cxrom1.pc1 [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_symbolic_cxrom1.pc1 [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_symbolic_cxrom1.pc2 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_symbolic_cxrom1.pc2 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_symbolic_cxrom1.pc2 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_symbolic_cxrom1.pc2 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_symbolic_cxrom1.pc2 [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_symbolic_cxrom1.pc2 [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_symbolic_cxrom1.pc2 [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_symbolic_cxrom1.pc2 [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_symbolic_cxrom1.pc2 [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_symbolic_cxrom1.pc2 [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_symbolic_cxrom1.pc2 [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_symbolic_cxrom1.pc2 [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_symbolic_cxrom1.pc2 [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_symbolic_cxrom1.pc2 [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_symbolic_cxrom1.pc2 [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_symbolic_cxrom1.pc2 [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [0], word_in[0]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [1], word_in[1]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [2], word_in[2]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [3], word_in[3]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [4], word_in[4]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [5], word_in[5]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [6], word_in[6]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [7], word_in[7]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [0], word_in[8]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [1], word_in[9]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [2], word_in[10]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [3], word_in[11]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [4], word_in[12]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [5], word_in[13]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [6], word_in[14]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [7], word_in[15]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [0], word_in[16]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [1], word_in[17]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [2], word_in[18]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [3], word_in[19]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [4], word_in[20]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [5], word_in[21]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [6], word_in[22]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [7], word_in[23]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [0], word_in[24]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [1], word_in[25]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [2], word_in[26]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [3], word_in[27]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [4], word_in[28]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [5], word_in[29]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [6], word_in[30]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [7], word_in[31]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_symbolic_cxrom1.pc10 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc10 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_symbolic_cxrom1.pc10 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_symbolic_cxrom1.pc10 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_symbolic_cxrom1.pc12 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc12 [1], pc1_plus_2[1]);
  buf(\oc8051_symbolic_cxrom1.pc12 [2], pc1_plus_2[2]);
  buf(\oc8051_symbolic_cxrom1.pc12 [3], pc1_plus_2[3]);
  buf(\oc8051_symbolic_cxrom1.pc20 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_symbolic_cxrom1.pc20 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_symbolic_cxrom1.pc20 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_symbolic_cxrom1.pc20 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_symbolic_cxrom1.pc22 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.oc8051_comp1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_comp1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_comp1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_comp1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_comp1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_comp1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_comp1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_comp1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_comp1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [0], ABINPUT000[0]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [1], ABINPUT000[1]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [2], ABINPUT000[2]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [3], ABINPUT000[3]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [4], ABINPUT000[4]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [5], ABINPUT000[5]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [6], ABINPUT000[6]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [7], ABINPUT000[7]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [8], ABINPUT000[8]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [9], ABINPUT000[9]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [10], ABINPUT000[10]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [11], ABINPUT000[11]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [12], ABINPUT000[12]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [13], ABINPUT000[13]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [14], ABINPUT000[14]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [15], ABINPUT000[15]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [16], ABINPUT000[16]);
  buf(\oc8051_top_1.oc8051_alu1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_alu1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc1 [0], ABINPUT000[1]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc1 [1], ABINPUT000[2]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc1 [2], ABINPUT000[3]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc1 [3], ABINPUT000[4]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc1 [4], ABINPUT000[5]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc1 [5], ABINPUT000[6]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc1 [6], ABINPUT000[7]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc1 [7], ABINPUT000[8]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc2 [0], ABINPUT000[9]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc2 [1], ABINPUT000[10]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc2 [2], ABINPUT000[11]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc2 [3], ABINPUT000[12]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc2 [4], ABINPUT000[13]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc2 [5], ABINPUT000[14]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc2 [6], ABINPUT000[15]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc2 [7], ABINPUT000[16]);
  buf(\oc8051_top_1.oc8051_alu1.mulOv , ABINPUT000[0]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc1 [0], ABINPUT001[1]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc1 [1], ABINPUT001[2]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc1 [2], ABINPUT001[3]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc1 [3], ABINPUT001[4]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc1 [4], ABINPUT001[5]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc1 [5], ABINPUT001[6]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc1 [6], ABINPUT001[7]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc1 [7], ABINPUT001[8]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [0], ABINPUT001[9]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [1], ABINPUT001[10]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [2], ABINPUT001[11]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [3], ABINPUT001[12]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [4], ABINPUT001[13]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [5], ABINPUT001[14]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [6], ABINPUT001[15]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [7], ABINPUT001[16]);
  buf(\oc8051_top_1.oc8051_alu1.divOv , ABINPUT001[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [4], \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [5], \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.uart_int , \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.t2_int , \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [0], ABINPUT001[0]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [1], ABINPUT001[1]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [2], ABINPUT001[2]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [3], ABINPUT001[3]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [4], ABINPUT001[4]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [5], ABINPUT001[5]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [6], ABINPUT001[6]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [7], ABINPUT001[7]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [8], ABINPUT001[8]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [9], ABINPUT001[9]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [10], ABINPUT001[10]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [11], ABINPUT001[11]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [12], ABINPUT001[12]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [13], ABINPUT001[13]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [14], ABINPUT001[14]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [15], ABINPUT001[15]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [16], ABINPUT001[16]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [0], \oc8051_top_1.oc8051_sfr1.psw [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.p , \oc8051_top_1.oc8051_sfr1.psw [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk , clk);
  buf(\oc8051_top_1.ABINPUT000 [0], ABINPUT000[0]);
  buf(\oc8051_top_1.ABINPUT000 [1], ABINPUT000[1]);
  buf(\oc8051_top_1.ABINPUT000 [2], ABINPUT000[2]);
  buf(\oc8051_top_1.ABINPUT000 [3], ABINPUT000[3]);
  buf(\oc8051_top_1.ABINPUT000 [4], ABINPUT000[4]);
  buf(\oc8051_top_1.ABINPUT000 [5], ABINPUT000[5]);
  buf(\oc8051_top_1.ABINPUT000 [6], ABINPUT000[6]);
  buf(\oc8051_top_1.ABINPUT000 [7], ABINPUT000[7]);
  buf(\oc8051_top_1.ABINPUT000 [8], ABINPUT000[8]);
  buf(\oc8051_top_1.ABINPUT000 [9], ABINPUT000[9]);
  buf(\oc8051_top_1.ABINPUT000 [10], ABINPUT000[10]);
  buf(\oc8051_top_1.ABINPUT000 [11], ABINPUT000[11]);
  buf(\oc8051_top_1.ABINPUT000 [12], ABINPUT000[12]);
  buf(\oc8051_top_1.ABINPUT000 [13], ABINPUT000[13]);
  buf(\oc8051_top_1.ABINPUT000 [14], ABINPUT000[14]);
  buf(\oc8051_top_1.ABINPUT000 [15], ABINPUT000[15]);
  buf(\oc8051_top_1.ABINPUT000 [16], ABINPUT000[16]);
  buf(\oc8051_top_1.ABINPUT001 [0], ABINPUT001[0]);
  buf(\oc8051_top_1.ABINPUT001 [1], ABINPUT001[1]);
  buf(\oc8051_top_1.ABINPUT001 [2], ABINPUT001[2]);
  buf(\oc8051_top_1.ABINPUT001 [3], ABINPUT001[3]);
  buf(\oc8051_top_1.ABINPUT001 [4], ABINPUT001[4]);
  buf(\oc8051_top_1.ABINPUT001 [5], ABINPUT001[5]);
  buf(\oc8051_top_1.ABINPUT001 [6], ABINPUT001[6]);
  buf(\oc8051_top_1.ABINPUT001 [7], ABINPUT001[7]);
  buf(\oc8051_top_1.ABINPUT001 [8], ABINPUT001[8]);
  buf(\oc8051_top_1.ABINPUT001 [9], ABINPUT001[9]);
  buf(\oc8051_top_1.ABINPUT001 [10], ABINPUT001[10]);
  buf(\oc8051_top_1.ABINPUT001 [11], ABINPUT001[11]);
  buf(\oc8051_top_1.ABINPUT001 [12], ABINPUT001[12]);
  buf(\oc8051_top_1.ABINPUT001 [13], ABINPUT001[13]);
  buf(\oc8051_top_1.ABINPUT001 [14], ABINPUT001[14]);
  buf(\oc8051_top_1.ABINPUT001 [15], ABINPUT001[15]);
  buf(\oc8051_top_1.ABINPUT001 [16], ABINPUT001[16]);
  buf(\oc8051_top_1.ABINPUT [0], ABINPUT[0]);
  buf(\oc8051_top_1.ABINPUT [1], ABINPUT[1]);
  buf(\oc8051_top_1.ABINPUT [2], ABINPUT[2]);
  buf(\oc8051_top_1.ABINPUT [3], ABINPUT[3]);
  buf(\oc8051_top_1.ABINPUT [4], ABINPUT[4]);
  buf(\oc8051_top_1.ABINPUT [5], ABINPUT[5]);
  buf(\oc8051_top_1.ABINPUT [6], ABINPUT[6]);
  buf(\oc8051_top_1.ABINPUT [7], ABINPUT[7]);
  buf(\oc8051_top_1.ABINPUT [8], ABINPUT[8]);
  buf(\oc8051_top_1.wb_rst_i , rst);
  buf(\oc8051_top_1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.bit_data , ABINPUT[0]);
  buf(\oc8051_top_1.rd_ind , \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  buf(\oc8051_top_1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.wb_clk_i , clk);
  buf(\oc8051_top_1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.sfr_out [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.sfr_out [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.sfr_out [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.sfr_out [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.sfr_out [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.sfr_out [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.sfr_out [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.sfr_out [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.ram_data [0], ABINPUT[1]);
  buf(\oc8051_top_1.ram_data [1], ABINPUT[2]);
  buf(\oc8051_top_1.ram_data [2], ABINPUT[3]);
  buf(\oc8051_top_1.ram_data [3], ABINPUT[4]);
  buf(\oc8051_top_1.ram_data [4], ABINPUT[5]);
  buf(\oc8051_top_1.ram_data [5], ABINPUT[6]);
  buf(\oc8051_top_1.ram_data [6], ABINPUT[7]);
  buf(\oc8051_top_1.ram_data [7], ABINPUT[8]);
  buf(\oc8051_top_1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.src_sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.src_sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_top_1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_top_1.pc_log [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_top_1.pc_log [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_top_1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_top_1.pc_log [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_top_1.pc_log [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_top_1.pc_log [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_top_1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_top_1.pc_log [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_top_1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_top_1.pc_log [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_top_1.pc_log [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_top_1.pc_log [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_top_1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_top_1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.t2ex_i , t2ex_i);
  buf(\oc8051_top_1.t2_i , t2_i);
  buf(\oc8051_top_1.t1_i , t1_i);
  buf(\oc8051_top_1.t0_i , t0_i);
  buf(\oc8051_top_1.rxd_i , rxd_i);
  buf(\oc8051_top_1.p3_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.p3_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.p3_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.p3_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.p3_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.p3_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.p3_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.p3_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.p3_i [0], p3_in[0]);
  buf(\oc8051_top_1.p3_i [1], p3_in[1]);
  buf(\oc8051_top_1.p3_i [2], p3_in[2]);
  buf(\oc8051_top_1.p3_i [3], p3_in[3]);
  buf(\oc8051_top_1.p3_i [4], p3_in[4]);
  buf(\oc8051_top_1.p3_i [5], p3_in[5]);
  buf(\oc8051_top_1.p3_i [6], p3_in[6]);
  buf(\oc8051_top_1.p3_i [7], p3_in[7]);
  buf(\oc8051_top_1.p2_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.p2_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.p2_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.p2_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.p2_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.p2_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.p2_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.p2_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.p2_i [0], p2_in[0]);
  buf(\oc8051_top_1.p2_i [1], p2_in[1]);
  buf(\oc8051_top_1.p2_i [2], p2_in[2]);
  buf(\oc8051_top_1.p2_i [3], p2_in[3]);
  buf(\oc8051_top_1.p2_i [4], p2_in[4]);
  buf(\oc8051_top_1.p2_i [5], p2_in[5]);
  buf(\oc8051_top_1.p2_i [6], p2_in[6]);
  buf(\oc8051_top_1.p2_i [7], p2_in[7]);
  buf(\oc8051_top_1.p1_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.p1_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.p1_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.p1_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.p1_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.p1_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.p1_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.p1_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.p1_i [0], p1_in[0]);
  buf(\oc8051_top_1.p1_i [1], p1_in[1]);
  buf(\oc8051_top_1.p1_i [2], p1_in[2]);
  buf(\oc8051_top_1.p1_i [3], p1_in[3]);
  buf(\oc8051_top_1.p1_i [4], p1_in[4]);
  buf(\oc8051_top_1.p1_i [5], p1_in[5]);
  buf(\oc8051_top_1.p1_i [6], p1_in[6]);
  buf(\oc8051_top_1.p1_i [7], p1_in[7]);
  buf(\oc8051_top_1.p0_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.p0_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.p0_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.p0_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.p0_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.p0_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.p0_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.p0_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.p0_i [0], p0_in[0]);
  buf(\oc8051_top_1.p0_i [1], p0_in[1]);
  buf(\oc8051_top_1.p0_i [2], p0_in[2]);
  buf(\oc8051_top_1.p0_i [3], p0_in[3]);
  buf(\oc8051_top_1.p0_i [4], p0_in[4]);
  buf(\oc8051_top_1.p0_i [5], p0_in[5]);
  buf(\oc8051_top_1.p0_i [6], p0_in[6]);
  buf(\oc8051_top_1.p0_i [7], p0_in[7]);
  buf(\oc8051_top_1.cxrom_data_out [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.cxrom_data_out [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.cxrom_data_out [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.cxrom_data_out [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.cxrom_data_out [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.cxrom_data_out [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.cxrom_data_out [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.cxrom_data_out [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.cxrom_data_out [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.cxrom_data_out [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.cxrom_data_out [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.cxrom_data_out [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.cxrom_data_out [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.cxrom_data_out [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.cxrom_data_out [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.cxrom_data_out [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.cxrom_data_out [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.cxrom_data_out [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.cxrom_data_out [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.cxrom_data_out [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.cxrom_data_out [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.cxrom_data_out [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.cxrom_data_out [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.cxrom_data_out [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.cxrom_data_out [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.cxrom_data_out [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.cxrom_data_out [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.cxrom_data_out [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.cxrom_data_out [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.cxrom_data_out [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.cxrom_data_out [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.cxrom_data_out [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_top_1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_top_1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_top_1.pc_log_prev [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_top_1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_top_1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_top_1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_top_1.pc_log_prev [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_top_1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_top_1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_top_1.pc_log_prev [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_top_1.pc_log_prev [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_top_1.pc_log_prev [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_top_1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_top_1.pc_log_prev [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_top_1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(cy, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(pc1[0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(pc1[1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(pc1[2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(pc1[3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(pc1[4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(pc1[5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(pc1[6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(pc1[7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(pc1[8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(pc1[9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(pc1[10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(pc1[11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(pc1[12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(pc1[13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(pc1[14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(pc1[15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(pc2[0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(pc2[1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(pc2[2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(pc2[3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(pc2[4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(pc2[5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(pc2[6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(pc2[7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(pc2[8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(pc2[9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(pc2[10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(pc2[11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(pc2[12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(pc2[13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(pc2[14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(pc2[15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(cxrom_data_out[0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(cxrom_data_out[1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(cxrom_data_out[2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(cxrom_data_out[3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(cxrom_data_out[4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(cxrom_data_out[5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(cxrom_data_out[6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(cxrom_data_out[7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(cxrom_data_out[8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(cxrom_data_out[9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(cxrom_data_out[10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(cxrom_data_out[11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(cxrom_data_out[12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(cxrom_data_out[13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(cxrom_data_out[14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(cxrom_data_out[15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(cxrom_data_out[16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(cxrom_data_out[17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(cxrom_data_out[18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(cxrom_data_out[19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(cxrom_data_out[20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(cxrom_data_out[21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(cxrom_data_out[22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(cxrom_data_out[23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(cxrom_data_out[24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(cxrom_data_out[25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(cxrom_data_out[26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(cxrom_data_out[27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(cxrom_data_out[28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(cxrom_data_out[29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(cxrom_data_out[30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(cxrom_data_out[31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst , rst);
  buf(pc1_plus_2[0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk , clk);
  buf(p3_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(p3_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(p3_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(p3_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(p3_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(p3_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(p3_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(p3_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(p2_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(p2_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(p2_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(p2_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(p2_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(p2_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(p2_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(p2_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(p1_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(p1_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(p1_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(p1_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(p1_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(p1_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(p1_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(p1_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(p0_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(p0_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(p0_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(p0_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(p0_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(p0_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(p0_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(p0_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
endmodule
