
module oc8051_gm_top(clk, rst, word_in, p0_in, p1_in, p2_in, p3_in, property_invalid_rom_pc, ABINPUT);
  wire [7:0] _00000_;
  wire [7:0] _00001_;
  wire [7:0] _00002_;
  wire [7:0] _00003_;
  wire _00004_;
  wire _00005_;
  wire _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  wire _08001_;
  wire _08002_;
  wire _08003_;
  wire _08004_;
  wire _08005_;
  wire _08006_;
  wire _08007_;
  wire _08008_;
  wire _08009_;
  wire _08010_;
  wire _08011_;
  wire _08012_;
  wire _08013_;
  wire _08014_;
  wire _08015_;
  wire _08016_;
  wire _08017_;
  wire _08018_;
  wire _08019_;
  wire _08020_;
  wire _08021_;
  wire _08022_;
  wire _08023_;
  wire _08024_;
  wire _08025_;
  wire _08026_;
  wire _08027_;
  wire _08028_;
  wire _08029_;
  wire _08030_;
  wire _08031_;
  wire _08032_;
  wire _08033_;
  wire _08034_;
  wire _08035_;
  wire _08036_;
  wire _08037_;
  wire _08038_;
  wire _08039_;
  wire _08040_;
  wire _08041_;
  wire _08042_;
  wire _08043_;
  wire _08044_;
  wire _08045_;
  wire _08046_;
  wire _08047_;
  wire _08048_;
  wire _08049_;
  wire _08050_;
  wire _08051_;
  wire _08052_;
  wire _08053_;
  wire _08054_;
  wire _08055_;
  wire _08056_;
  wire _08057_;
  wire _08058_;
  wire _08059_;
  wire _08060_;
  wire _08061_;
  wire _08062_;
  wire _08063_;
  wire _08064_;
  wire _08065_;
  wire _08066_;
  wire _08067_;
  wire _08068_;
  wire _08069_;
  wire _08070_;
  wire _08071_;
  wire _08072_;
  wire _08073_;
  wire _08074_;
  wire _08075_;
  wire _08076_;
  wire _08077_;
  wire _08078_;
  wire _08079_;
  wire _08080_;
  wire _08081_;
  wire _08082_;
  wire _08083_;
  wire _08084_;
  wire _08085_;
  wire _08086_;
  wire _08087_;
  wire _08088_;
  wire _08089_;
  wire _08090_;
  wire _08091_;
  wire _08092_;
  wire _08093_;
  wire _08094_;
  wire _08095_;
  wire _08096_;
  wire _08097_;
  wire _08098_;
  wire _08099_;
  wire _08100_;
  wire _08101_;
  wire _08102_;
  wire _08103_;
  wire _08104_;
  wire _08105_;
  wire _08106_;
  wire _08107_;
  wire _08108_;
  wire _08109_;
  wire _08110_;
  wire _08111_;
  wire _08112_;
  wire _08113_;
  wire _08114_;
  wire _08115_;
  wire _08116_;
  wire _08117_;
  wire _08118_;
  wire _08119_;
  wire _08120_;
  wire _08121_;
  wire _08122_;
  wire _08123_;
  wire _08124_;
  wire _08125_;
  wire _08126_;
  wire _08127_;
  wire _08128_;
  wire _08129_;
  wire _08130_;
  wire _08131_;
  wire _08132_;
  wire _08133_;
  wire _08134_;
  wire _08135_;
  wire _08136_;
  wire _08137_;
  wire _08138_;
  wire _08139_;
  wire _08140_;
  wire _08141_;
  wire _08142_;
  wire _08143_;
  wire _08144_;
  wire _08145_;
  wire _08146_;
  wire _08147_;
  wire _08148_;
  wire _08149_;
  wire _08150_;
  wire _08151_;
  wire _08152_;
  wire _08153_;
  wire _08154_;
  wire _08155_;
  wire _08156_;
  wire _08157_;
  wire _08158_;
  wire _08159_;
  wire _08160_;
  wire _08161_;
  wire _08162_;
  wire _08163_;
  wire _08164_;
  wire _08165_;
  wire _08166_;
  wire _08167_;
  wire _08168_;
  wire _08169_;
  wire _08170_;
  wire _08171_;
  wire _08172_;
  wire _08173_;
  wire _08174_;
  wire _08175_;
  wire _08176_;
  wire _08177_;
  wire _08178_;
  wire _08179_;
  wire _08180_;
  wire _08181_;
  wire _08182_;
  wire _08183_;
  wire _08184_;
  wire _08185_;
  wire _08186_;
  wire _08187_;
  wire _08188_;
  wire _08189_;
  wire _08190_;
  wire _08191_;
  wire _08192_;
  wire _08193_;
  wire _08194_;
  wire _08195_;
  wire _08196_;
  wire _08197_;
  wire _08198_;
  wire _08199_;
  wire _08200_;
  wire _08201_;
  wire _08202_;
  wire _08203_;
  wire _08204_;
  wire _08205_;
  wire _08206_;
  wire _08207_;
  wire _08208_;
  wire _08209_;
  wire _08210_;
  wire _08211_;
  wire _08212_;
  wire _08213_;
  wire _08214_;
  wire _08215_;
  wire _08216_;
  wire _08217_;
  wire _08218_;
  wire _08219_;
  wire _08220_;
  wire _08221_;
  wire _08222_;
  wire _08223_;
  wire _08224_;
  wire _08225_;
  wire _08226_;
  wire _08227_;
  wire _08228_;
  wire _08229_;
  wire _08230_;
  wire _08231_;
  wire _08232_;
  wire _08233_;
  wire _08234_;
  wire _08235_;
  wire _08236_;
  wire _08237_;
  wire _08238_;
  wire _08239_;
  wire _08240_;
  wire _08241_;
  wire _08242_;
  wire _08243_;
  wire _08244_;
  wire _08245_;
  wire _08246_;
  wire _08247_;
  wire _08248_;
  wire _08249_;
  wire _08250_;
  wire _08251_;
  wire _08252_;
  wire _08253_;
  wire _08254_;
  wire _08255_;
  wire _08256_;
  wire _08257_;
  wire _08258_;
  wire _08259_;
  wire _08260_;
  wire _08261_;
  wire _08262_;
  wire _08263_;
  wire _08264_;
  wire _08265_;
  wire _08266_;
  wire _08267_;
  wire _08268_;
  wire _08269_;
  wire _08270_;
  wire _08271_;
  wire _08272_;
  wire _08273_;
  wire _08274_;
  wire _08275_;
  wire _08276_;
  wire _08277_;
  wire _08278_;
  wire _08279_;
  wire _08280_;
  wire _08281_;
  wire _08282_;
  wire _08283_;
  wire _08284_;
  wire _08285_;
  wire _08286_;
  wire _08287_;
  wire _08288_;
  wire _08289_;
  wire _08290_;
  wire _08291_;
  wire _08292_;
  wire _08293_;
  wire _08294_;
  wire _08295_;
  wire _08296_;
  wire _08297_;
  wire _08298_;
  wire _08299_;
  wire _08300_;
  wire _08301_;
  wire _08302_;
  wire _08303_;
  wire _08304_;
  wire _08305_;
  wire _08306_;
  wire _08307_;
  wire _08308_;
  wire _08309_;
  wire _08310_;
  wire _08311_;
  wire _08312_;
  wire _08313_;
  wire _08314_;
  wire _08315_;
  wire _08316_;
  wire _08317_;
  wire _08318_;
  wire _08319_;
  wire _08320_;
  wire _08321_;
  wire _08322_;
  wire _08323_;
  wire _08324_;
  wire _08325_;
  wire _08326_;
  wire _08327_;
  wire _08328_;
  wire _08329_;
  wire _08330_;
  wire _08331_;
  wire _08332_;
  wire _08333_;
  wire _08334_;
  wire _08335_;
  wire _08336_;
  wire _08337_;
  wire _08338_;
  wire _08339_;
  wire _08340_;
  wire _08341_;
  wire _08342_;
  wire _08343_;
  wire _08344_;
  wire _08345_;
  wire _08346_;
  wire _08347_;
  wire _08348_;
  wire _08349_;
  wire _08350_;
  wire _08351_;
  wire _08352_;
  wire _08353_;
  wire _08354_;
  wire _08355_;
  wire _08356_;
  wire _08357_;
  wire _08358_;
  wire _08359_;
  wire _08360_;
  wire _08361_;
  wire _08362_;
  wire _08363_;
  wire _08364_;
  wire _08365_;
  wire _08366_;
  wire _08367_;
  wire _08368_;
  wire _08369_;
  wire _08370_;
  wire _08371_;
  wire _08372_;
  wire _08373_;
  wire _08374_;
  wire _08375_;
  wire _08376_;
  wire _08377_;
  wire _08378_;
  wire _08379_;
  wire _08380_;
  wire _08381_;
  wire _08382_;
  wire _08383_;
  wire _08384_;
  wire _08385_;
  wire _08386_;
  wire _08387_;
  wire _08388_;
  wire _08389_;
  wire _08390_;
  wire _08391_;
  wire _08392_;
  wire _08393_;
  wire _08394_;
  wire _08395_;
  wire _08396_;
  wire _08397_;
  wire _08398_;
  wire _08399_;
  wire _08400_;
  wire _08401_;
  wire _08402_;
  wire _08403_;
  wire _08404_;
  wire _08405_;
  wire _08406_;
  wire _08407_;
  wire _08408_;
  wire _08409_;
  wire _08410_;
  wire _08411_;
  wire _08412_;
  wire _08413_;
  wire _08414_;
  wire _08415_;
  wire _08416_;
  wire _08417_;
  wire _08418_;
  wire _08419_;
  wire _08420_;
  wire _08421_;
  wire _08422_;
  wire _08423_;
  wire _08424_;
  wire _08425_;
  wire _08426_;
  wire _08427_;
  wire _08428_;
  wire _08429_;
  wire _08430_;
  wire _08431_;
  wire _08432_;
  wire _08433_;
  wire _08434_;
  wire _08435_;
  wire _08436_;
  wire _08437_;
  wire _08438_;
  wire _08439_;
  wire _08440_;
  wire _08441_;
  wire _08442_;
  wire _08443_;
  wire _08444_;
  wire _08445_;
  wire _08446_;
  wire _08447_;
  wire _08448_;
  wire _08449_;
  wire _08450_;
  wire _08451_;
  wire _08452_;
  wire _08453_;
  wire _08454_;
  wire _08455_;
  wire _08456_;
  wire _08457_;
  wire _08458_;
  wire _08459_;
  wire _08460_;
  wire _08461_;
  wire _08462_;
  wire _08463_;
  wire _08464_;
  wire _08465_;
  wire _08466_;
  wire _08467_;
  wire _08468_;
  wire _08469_;
  wire _08470_;
  wire _08471_;
  wire _08472_;
  wire _08473_;
  wire _08474_;
  wire _08475_;
  wire _08476_;
  wire _08477_;
  wire _08478_;
  wire _08479_;
  wire _08480_;
  wire _08481_;
  wire _08482_;
  wire _08483_;
  wire _08484_;
  wire _08485_;
  wire _08486_;
  wire _08487_;
  wire _08488_;
  wire _08489_;
  wire _08490_;
  wire _08491_;
  wire _08492_;
  wire _08493_;
  wire _08494_;
  wire _08495_;
  wire _08496_;
  wire _08497_;
  wire _08498_;
  wire _08499_;
  wire _08500_;
  wire _08501_;
  wire _08502_;
  wire _08503_;
  wire _08504_;
  wire _08505_;
  wire _08506_;
  wire _08507_;
  wire _08508_;
  wire _08509_;
  wire _08510_;
  wire _08511_;
  wire _08512_;
  wire _08513_;
  wire _08514_;
  wire _08515_;
  wire _08516_;
  wire _08517_;
  wire _08518_;
  wire _08519_;
  wire _08520_;
  wire _08521_;
  wire _08522_;
  wire _08523_;
  wire _08524_;
  wire _08525_;
  wire _08526_;
  wire _08527_;
  wire _08528_;
  wire _08529_;
  wire _08530_;
  wire _08531_;
  wire _08532_;
  wire _08533_;
  wire _08534_;
  wire _08535_;
  wire _08536_;
  wire _08537_;
  wire _08538_;
  wire _08539_;
  wire _08540_;
  wire _08541_;
  wire _08542_;
  wire _08543_;
  wire _08544_;
  wire _08545_;
  wire _08546_;
  wire _08547_;
  wire _08548_;
  wire _08549_;
  wire _08550_;
  wire _08551_;
  wire _08552_;
  wire _08553_;
  wire _08554_;
  wire _08555_;
  wire _08556_;
  wire _08557_;
  wire _08558_;
  wire _08559_;
  wire _08560_;
  wire _08561_;
  wire _08562_;
  wire _08563_;
  wire _08564_;
  wire _08565_;
  wire _08566_;
  wire _08567_;
  wire _08568_;
  wire _08569_;
  wire _08570_;
  wire _08571_;
  wire _08572_;
  wire _08573_;
  wire _08574_;
  wire _08575_;
  wire _08576_;
  wire _08577_;
  wire _08578_;
  wire _08579_;
  wire _08580_;
  wire _08581_;
  wire _08582_;
  wire _08583_;
  wire _08584_;
  wire _08585_;
  wire _08586_;
  wire _08587_;
  wire _08588_;
  wire _08589_;
  wire _08590_;
  wire _08591_;
  wire _08592_;
  wire _08593_;
  wire _08594_;
  wire _08595_;
  wire _08596_;
  wire _08597_;
  wire _08598_;
  wire _08599_;
  wire _08600_;
  wire _08601_;
  wire _08602_;
  wire _08603_;
  wire _08604_;
  wire _08605_;
  wire _08606_;
  wire _08607_;
  wire _08608_;
  wire _08609_;
  wire _08610_;
  wire _08611_;
  wire _08612_;
  wire _08613_;
  wire _08614_;
  wire _08615_;
  wire _08616_;
  wire _08617_;
  wire _08618_;
  wire _08619_;
  wire _08620_;
  wire _08621_;
  wire _08622_;
  wire _08623_;
  wire _08624_;
  wire _08625_;
  wire _08626_;
  wire _08627_;
  wire _08628_;
  wire _08629_;
  wire _08630_;
  wire _08631_;
  wire _08632_;
  wire _08633_;
  wire _08634_;
  wire _08635_;
  wire _08636_;
  wire _08637_;
  wire _08638_;
  wire _08639_;
  wire _08640_;
  wire _08641_;
  wire _08642_;
  wire _08643_;
  wire _08644_;
  wire _08645_;
  wire _08646_;
  wire _08647_;
  wire _08648_;
  wire _08649_;
  wire _08650_;
  wire _08651_;
  wire _08652_;
  wire _08653_;
  wire _08654_;
  wire _08655_;
  wire _08656_;
  wire _08657_;
  wire _08658_;
  wire _08659_;
  wire _08660_;
  wire _08661_;
  wire _08662_;
  wire _08663_;
  wire _08664_;
  wire _08665_;
  wire _08666_;
  wire _08667_;
  wire _08668_;
  wire _08669_;
  wire _08670_;
  wire _08671_;
  wire _08672_;
  wire _08673_;
  wire _08674_;
  wire _08675_;
  wire _08676_;
  wire _08677_;
  wire _08678_;
  wire _08679_;
  wire _08680_;
  wire _08681_;
  wire _08682_;
  wire _08683_;
  wire _08684_;
  wire _08685_;
  wire _08686_;
  wire _08687_;
  wire _08688_;
  wire _08689_;
  wire _08690_;
  wire _08691_;
  wire _08692_;
  wire _08693_;
  wire _08694_;
  wire _08695_;
  wire _08696_;
  wire _08697_;
  wire _08698_;
  wire _08699_;
  wire _08700_;
  wire _08701_;
  wire _08702_;
  wire _08703_;
  wire _08704_;
  wire _08705_;
  wire _08706_;
  wire _08707_;
  wire _08708_;
  wire _08709_;
  wire _08710_;
  wire _08711_;
  wire _08712_;
  wire _08713_;
  wire _08714_;
  wire _08715_;
  wire _08716_;
  wire _08717_;
  wire _08718_;
  wire _08719_;
  wire _08720_;
  wire _08721_;
  wire _08722_;
  wire _08723_;
  wire _08724_;
  wire _08725_;
  wire _08726_;
  wire _08727_;
  wire _08728_;
  wire _08729_;
  wire _08730_;
  wire _08731_;
  wire _08732_;
  wire _08733_;
  wire _08734_;
  wire _08735_;
  wire _08736_;
  wire _08737_;
  wire _08738_;
  wire _08739_;
  wire _08740_;
  wire _08741_;
  wire _08742_;
  wire _08743_;
  wire _08744_;
  wire _08745_;
  wire _08746_;
  wire _08747_;
  wire _08748_;
  wire _08749_;
  wire _08750_;
  wire _08751_;
  wire _08752_;
  wire _08753_;
  wire _08754_;
  wire _08755_;
  wire _08756_;
  wire _08757_;
  wire _08758_;
  wire _08759_;
  wire _08760_;
  wire _08761_;
  wire _08762_;
  wire _08763_;
  wire _08764_;
  wire _08765_;
  wire _08766_;
  wire _08767_;
  wire _08768_;
  wire _08769_;
  wire _08770_;
  wire _08771_;
  wire _08772_;
  wire _08773_;
  wire _08774_;
  wire _08775_;
  wire _08776_;
  wire _08777_;
  wire _08778_;
  wire _08779_;
  wire _08780_;
  wire _08781_;
  wire _08782_;
  wire _08783_;
  wire _08784_;
  wire _08785_;
  wire _08786_;
  wire _08787_;
  wire _08788_;
  wire _08789_;
  wire _08790_;
  wire _08791_;
  wire _08792_;
  wire _08793_;
  wire _08794_;
  wire _08795_;
  wire _08796_;
  wire _08797_;
  wire _08798_;
  wire _08799_;
  wire _08800_;
  wire _08801_;
  wire _08802_;
  wire _08803_;
  wire _08804_;
  wire _08805_;
  wire _08806_;
  wire _08807_;
  wire _08808_;
  wire _08809_;
  wire _08810_;
  wire _08811_;
  wire _08812_;
  wire _08813_;
  wire _08814_;
  wire _08815_;
  wire _08816_;
  wire _08817_;
  wire _08818_;
  wire _08819_;
  wire _08820_;
  wire _08821_;
  wire _08822_;
  wire _08823_;
  wire _08824_;
  wire _08825_;
  wire _08826_;
  wire _08827_;
  wire _08828_;
  wire _08829_;
  wire _08830_;
  wire _08831_;
  wire _08832_;
  wire _08833_;
  wire _08834_;
  wire _08835_;
  wire _08836_;
  wire _08837_;
  wire _08838_;
  wire _08839_;
  wire _08840_;
  wire _08841_;
  wire _08842_;
  wire _08843_;
  wire _08844_;
  wire _08845_;
  wire _08846_;
  wire _08847_;
  wire _08848_;
  wire _08849_;
  wire _08850_;
  wire _08851_;
  wire _08852_;
  wire _08853_;
  wire _08854_;
  wire _08855_;
  wire _08856_;
  wire _08857_;
  wire _08858_;
  wire _08859_;
  wire _08860_;
  wire _08861_;
  wire _08862_;
  wire _08863_;
  wire _08864_;
  wire _08865_;
  wire _08866_;
  wire _08867_;
  wire _08868_;
  wire _08869_;
  wire _08870_;
  wire _08871_;
  wire _08872_;
  wire _08873_;
  wire _08874_;
  wire _08875_;
  wire _08876_;
  wire _08877_;
  wire _08878_;
  wire _08879_;
  wire _08880_;
  wire _08881_;
  wire _08882_;
  wire _08883_;
  wire _08884_;
  wire _08885_;
  wire _08886_;
  wire _08887_;
  wire _08888_;
  wire _08889_;
  wire _08890_;
  wire _08891_;
  wire _08892_;
  wire _08893_;
  wire _08894_;
  wire _08895_;
  wire _08896_;
  wire _08897_;
  wire _08898_;
  wire _08899_;
  wire _08900_;
  wire _08901_;
  wire _08902_;
  wire _08903_;
  wire _08904_;
  wire _08905_;
  wire _08906_;
  wire _08907_;
  wire _08908_;
  wire _08909_;
  wire _08910_;
  wire _08911_;
  wire _08912_;
  wire _08913_;
  wire _08914_;
  wire _08915_;
  wire _08916_;
  wire _08917_;
  wire _08918_;
  wire _08919_;
  wire _08920_;
  wire _08921_;
  wire _08922_;
  wire _08923_;
  wire _08924_;
  wire _08925_;
  wire _08926_;
  wire _08927_;
  wire _08928_;
  wire _08929_;
  wire _08930_;
  wire _08931_;
  wire _08932_;
  wire _08933_;
  wire _08934_;
  wire _08935_;
  wire _08936_;
  wire _08937_;
  wire _08938_;
  wire _08939_;
  wire _08940_;
  wire _08941_;
  wire _08942_;
  wire _08943_;
  wire _08944_;
  wire _08945_;
  wire _08946_;
  wire _08947_;
  wire _08948_;
  wire _08949_;
  wire _08950_;
  wire _08951_;
  wire _08952_;
  wire _08953_;
  wire _08954_;
  wire _08955_;
  wire _08956_;
  wire _08957_;
  wire _08958_;
  wire _08959_;
  wire _08960_;
  wire _08961_;
  wire _08962_;
  wire _08963_;
  wire _08964_;
  wire _08965_;
  wire _08966_;
  wire _08967_;
  wire _08968_;
  wire _08969_;
  wire _08970_;
  wire _08971_;
  wire _08972_;
  wire _08973_;
  wire _08974_;
  wire _08975_;
  wire _08976_;
  wire _08977_;
  wire _08978_;
  wire _08979_;
  wire _08980_;
  wire _08981_;
  wire _08982_;
  wire _08983_;
  wire _08984_;
  wire _08985_;
  wire _08986_;
  wire _08987_;
  wire _08988_;
  wire _08989_;
  wire _08990_;
  wire _08991_;
  wire _08992_;
  wire _08993_;
  wire _08994_;
  wire _08995_;
  wire _08996_;
  wire _08997_;
  wire _08998_;
  wire _08999_;
  wire _09000_;
  wire _09001_;
  wire _09002_;
  wire _09003_;
  wire _09004_;
  wire _09005_;
  wire _09006_;
  wire _09007_;
  wire _09008_;
  wire _09009_;
  wire _09010_;
  wire _09011_;
  wire _09012_;
  wire _09013_;
  wire _09014_;
  wire _09015_;
  wire _09016_;
  wire _09017_;
  wire _09018_;
  wire _09019_;
  wire _09020_;
  wire _09021_;
  wire _09022_;
  wire _09023_;
  wire _09024_;
  wire _09025_;
  wire _09026_;
  wire _09027_;
  wire _09028_;
  wire _09029_;
  wire _09030_;
  wire _09031_;
  wire _09032_;
  wire _09033_;
  wire _09034_;
  wire _09035_;
  wire _09036_;
  wire _09037_;
  wire _09038_;
  wire _09039_;
  wire _09040_;
  wire _09041_;
  wire _09042_;
  wire _09043_;
  wire _09044_;
  wire _09045_;
  wire _09046_;
  wire _09047_;
  wire _09048_;
  wire _09049_;
  wire _09050_;
  wire _09051_;
  wire _09052_;
  wire _09053_;
  wire _09054_;
  wire _09055_;
  wire _09056_;
  wire _09057_;
  wire _09058_;
  wire _09059_;
  wire _09060_;
  wire _09061_;
  wire _09062_;
  wire _09063_;
  wire _09064_;
  wire _09065_;
  wire _09066_;
  wire _09067_;
  wire _09068_;
  wire _09069_;
  wire _09070_;
  wire _09071_;
  wire _09072_;
  wire _09073_;
  wire _09074_;
  wire _09075_;
  wire _09076_;
  wire _09077_;
  wire _09078_;
  wire _09079_;
  wire _09080_;
  wire _09081_;
  wire _09082_;
  wire _09083_;
  wire _09084_;
  wire _09085_;
  wire _09086_;
  wire _09087_;
  wire _09088_;
  wire _09089_;
  wire _09090_;
  wire _09091_;
  wire _09092_;
  wire _09093_;
  wire _09094_;
  wire _09095_;
  wire _09096_;
  wire _09097_;
  wire _09098_;
  wire _09099_;
  wire _09100_;
  wire _09101_;
  wire _09102_;
  wire _09103_;
  wire _09104_;
  wire _09105_;
  wire _09106_;
  wire _09107_;
  wire _09108_;
  wire _09109_;
  wire _09110_;
  wire _09111_;
  wire _09112_;
  wire _09113_;
  wire _09114_;
  wire _09115_;
  wire _09116_;
  wire _09117_;
  wire _09118_;
  wire _09119_;
  wire _09120_;
  wire _09121_;
  wire _09122_;
  wire _09123_;
  wire _09124_;
  wire _09125_;
  wire _09126_;
  wire _09127_;
  wire _09128_;
  wire _09129_;
  wire _09130_;
  wire _09131_;
  wire _09132_;
  wire _09133_;
  wire _09134_;
  wire _09135_;
  wire _09136_;
  wire _09137_;
  wire _09138_;
  wire _09139_;
  wire _09140_;
  wire _09141_;
  wire _09142_;
  wire _09143_;
  wire _09144_;
  wire _09145_;
  wire _09146_;
  wire _09147_;
  wire _09148_;
  wire _09149_;
  wire _09150_;
  wire _09151_;
  wire _09152_;
  wire _09153_;
  wire _09154_;
  wire _09155_;
  wire _09156_;
  wire _09157_;
  wire _09158_;
  wire _09159_;
  wire _09160_;
  wire _09161_;
  wire _09162_;
  wire _09163_;
  wire _09164_;
  wire _09165_;
  wire _09166_;
  wire _09167_;
  wire _09168_;
  wire _09169_;
  wire _09170_;
  wire _09171_;
  wire _09172_;
  wire _09173_;
  wire _09174_;
  wire _09175_;
  wire _09176_;
  wire _09177_;
  wire _09178_;
  wire _09179_;
  wire _09180_;
  wire _09181_;
  wire _09182_;
  wire _09183_;
  wire _09184_;
  wire _09185_;
  wire _09186_;
  wire _09187_;
  wire _09188_;
  wire _09189_;
  wire _09190_;
  wire _09191_;
  wire _09192_;
  wire _09193_;
  wire _09194_;
  wire _09195_;
  wire _09196_;
  wire _09197_;
  wire _09198_;
  wire _09199_;
  wire _09200_;
  wire _09201_;
  wire _09202_;
  wire _09203_;
  wire _09204_;
  wire _09205_;
  wire _09206_;
  wire _09207_;
  wire _09208_;
  wire _09209_;
  wire _09210_;
  wire _09211_;
  wire _09212_;
  wire _09213_;
  wire _09214_;
  wire _09215_;
  wire _09216_;
  wire _09217_;
  wire _09218_;
  wire _09219_;
  wire _09220_;
  wire _09221_;
  wire _09222_;
  wire _09223_;
  wire _09224_;
  wire _09225_;
  wire _09226_;
  wire _09227_;
  wire _09228_;
  wire _09229_;
  wire _09230_;
  wire _09231_;
  wire _09232_;
  wire _09233_;
  wire _09234_;
  wire _09235_;
  wire _09236_;
  wire _09237_;
  wire _09238_;
  wire _09239_;
  wire _09240_;
  wire _09241_;
  wire _09242_;
  wire _09243_;
  wire _09244_;
  wire _09245_;
  wire _09246_;
  wire _09247_;
  wire _09248_;
  wire _09249_;
  wire _09250_;
  wire _09251_;
  wire _09252_;
  wire _09253_;
  wire _09254_;
  wire _09255_;
  wire _09256_;
  wire _09257_;
  wire _09258_;
  wire _09259_;
  wire _09260_;
  wire _09261_;
  wire _09262_;
  wire _09263_;
  wire _09264_;
  wire _09265_;
  wire _09266_;
  wire _09267_;
  wire _09268_;
  wire _09269_;
  wire _09270_;
  wire _09271_;
  wire _09272_;
  wire _09273_;
  wire _09274_;
  wire _09275_;
  wire _09276_;
  wire _09277_;
  wire _09278_;
  wire _09279_;
  wire _09280_;
  wire _09281_;
  wire _09282_;
  wire _09283_;
  wire _09284_;
  wire _09285_;
  wire _09286_;
  wire _09287_;
  wire _09288_;
  wire _09289_;
  wire _09290_;
  wire _09291_;
  wire _09292_;
  wire _09293_;
  wire _09294_;
  wire _09295_;
  wire _09296_;
  wire _09297_;
  wire _09298_;
  wire _09299_;
  wire _09300_;
  wire _09301_;
  wire _09302_;
  wire _09303_;
  wire _09304_;
  wire _09305_;
  wire _09306_;
  wire _09307_;
  wire _09308_;
  wire _09309_;
  wire _09310_;
  wire _09311_;
  wire _09312_;
  wire _09313_;
  wire _09314_;
  wire _09315_;
  wire _09316_;
  wire _09317_;
  wire _09318_;
  wire _09319_;
  wire _09320_;
  wire _09321_;
  wire _09322_;
  wire _09323_;
  wire _09324_;
  wire _09325_;
  wire _09326_;
  wire _09327_;
  wire _09328_;
  wire _09329_;
  wire _09330_;
  wire _09331_;
  wire _09332_;
  wire _09333_;
  wire _09334_;
  wire _09335_;
  wire _09336_;
  wire _09337_;
  wire _09338_;
  wire _09339_;
  wire _09340_;
  wire _09341_;
  wire _09342_;
  wire _09343_;
  wire _09344_;
  wire _09345_;
  wire _09346_;
  wire _09347_;
  wire _09348_;
  wire _09349_;
  wire _09350_;
  wire _09351_;
  wire _09352_;
  wire _09353_;
  wire _09354_;
  wire _09355_;
  wire _09356_;
  wire _09357_;
  wire _09358_;
  wire _09359_;
  wire _09360_;
  wire _09361_;
  wire _09362_;
  wire _09363_;
  wire _09364_;
  wire _09365_;
  wire _09366_;
  wire _09367_;
  wire _09368_;
  wire _09369_;
  wire _09370_;
  wire _09371_;
  wire _09372_;
  wire _09373_;
  wire _09374_;
  wire _09375_;
  wire _09376_;
  wire _09377_;
  wire _09378_;
  wire _09379_;
  wire _09380_;
  wire _09381_;
  wire _09382_;
  wire _09383_;
  wire _09384_;
  wire _09385_;
  wire _09386_;
  wire _09387_;
  wire _09388_;
  wire _09389_;
  wire _09390_;
  wire _09391_;
  wire _09392_;
  wire _09393_;
  wire _09394_;
  wire _09395_;
  wire _09396_;
  wire _09397_;
  wire _09398_;
  wire _09399_;
  wire _09400_;
  wire _09401_;
  wire _09402_;
  wire _09403_;
  wire _09404_;
  wire _09405_;
  wire _09406_;
  wire _09407_;
  wire _09408_;
  wire _09409_;
  wire _09410_;
  wire _09411_;
  wire _09412_;
  wire _09413_;
  wire _09414_;
  wire _09415_;
  wire _09416_;
  wire _09417_;
  wire _09418_;
  wire _09419_;
  wire _09420_;
  wire _09421_;
  wire _09422_;
  wire _09423_;
  wire _09424_;
  wire _09425_;
  wire _09426_;
  wire _09427_;
  wire _09428_;
  wire _09429_;
  wire _09430_;
  wire _09431_;
  wire _09432_;
  wire _09433_;
  wire _09434_;
  wire _09435_;
  wire _09436_;
  wire _09437_;
  wire _09438_;
  wire _09439_;
  wire _09440_;
  wire _09441_;
  wire _09442_;
  wire _09443_;
  wire _09444_;
  wire _09445_;
  wire _09446_;
  wire _09447_;
  wire _09448_;
  wire _09449_;
  wire _09450_;
  wire _09451_;
  wire _09452_;
  wire _09453_;
  wire _09454_;
  wire _09455_;
  wire _09456_;
  wire _09457_;
  wire _09458_;
  wire _09459_;
  wire _09460_;
  wire _09461_;
  wire _09462_;
  wire _09463_;
  wire _09464_;
  wire _09465_;
  wire _09466_;
  wire _09467_;
  wire _09468_;
  wire _09469_;
  wire _09470_;
  wire _09471_;
  wire _09472_;
  wire _09473_;
  wire _09474_;
  wire _09475_;
  wire _09476_;
  wire _09477_;
  wire _09478_;
  wire _09479_;
  wire _09480_;
  wire _09481_;
  wire _09482_;
  wire _09483_;
  wire _09484_;
  wire _09485_;
  wire _09486_;
  wire _09487_;
  wire _09488_;
  wire _09489_;
  wire _09490_;
  wire _09491_;
  wire _09492_;
  wire _09493_;
  wire _09494_;
  wire _09495_;
  wire _09496_;
  wire _09497_;
  wire _09498_;
  wire _09499_;
  wire _09500_;
  wire _09501_;
  wire _09502_;
  wire _09503_;
  wire _09504_;
  wire _09505_;
  wire _09506_;
  wire _09507_;
  wire _09508_;
  wire _09509_;
  wire _09510_;
  wire _09511_;
  wire _09512_;
  wire _09513_;
  wire _09514_;
  wire _09515_;
  wire _09516_;
  wire _09517_;
  wire _09518_;
  wire _09519_;
  wire _09520_;
  wire _09521_;
  wire _09522_;
  wire _09523_;
  wire _09524_;
  wire _09525_;
  wire _09526_;
  wire _09527_;
  wire _09528_;
  wire _09529_;
  wire _09530_;
  wire _09531_;
  wire _09532_;
  wire _09533_;
  wire _09534_;
  wire _09535_;
  wire _09536_;
  wire _09537_;
  wire _09538_;
  wire _09539_;
  wire _09540_;
  wire _09541_;
  wire _09542_;
  wire _09543_;
  wire _09544_;
  wire _09545_;
  wire _09546_;
  wire _09547_;
  wire _09548_;
  wire _09549_;
  wire _09550_;
  wire _09551_;
  wire _09552_;
  wire _09553_;
  wire _09554_;
  wire _09555_;
  wire _09556_;
  wire _09557_;
  wire _09558_;
  wire _09559_;
  wire _09560_;
  wire _09561_;
  wire _09562_;
  wire _09563_;
  wire _09564_;
  wire _09565_;
  wire _09566_;
  wire _09567_;
  wire _09568_;
  wire _09569_;
  wire _09570_;
  wire _09571_;
  wire _09572_;
  wire _09573_;
  wire _09574_;
  wire _09575_;
  wire _09576_;
  wire _09577_;
  wire _09578_;
  wire _09579_;
  wire _09580_;
  wire _09581_;
  wire _09582_;
  wire _09583_;
  wire _09584_;
  wire _09585_;
  wire _09586_;
  wire _09587_;
  wire _09588_;
  wire _09589_;
  wire _09590_;
  wire _09591_;
  wire _09592_;
  wire _09593_;
  wire _09594_;
  wire _09595_;
  wire _09596_;
  wire _09597_;
  wire _09598_;
  wire _09599_;
  wire _09600_;
  wire _09601_;
  wire _09602_;
  wire _09603_;
  wire _09604_;
  wire _09605_;
  wire _09606_;
  wire _09607_;
  wire _09608_;
  wire _09609_;
  wire _09610_;
  wire _09611_;
  wire _09612_;
  wire _09613_;
  wire _09614_;
  wire _09615_;
  wire _09616_;
  wire _09617_;
  wire _09618_;
  wire _09619_;
  wire _09620_;
  wire _09621_;
  wire _09622_;
  wire _09623_;
  wire _09624_;
  wire _09625_;
  wire _09626_;
  wire _09627_;
  wire _09628_;
  wire _09629_;
  wire _09630_;
  wire _09631_;
  wire _09632_;
  wire _09633_;
  wire _09634_;
  wire _09635_;
  wire _09636_;
  wire _09637_;
  wire _09638_;
  wire _09639_;
  wire _09640_;
  wire _09641_;
  wire _09642_;
  wire _09643_;
  wire _09644_;
  wire _09645_;
  wire _09646_;
  wire _09647_;
  wire _09648_;
  wire _09649_;
  wire _09650_;
  wire _09651_;
  wire _09652_;
  wire _09653_;
  wire _09654_;
  wire _09655_;
  wire _09656_;
  wire _09657_;
  wire _09658_;
  wire _09659_;
  wire _09660_;
  wire _09661_;
  wire _09662_;
  wire _09663_;
  wire _09664_;
  wire _09665_;
  wire _09666_;
  wire _09667_;
  wire _09668_;
  wire _09669_;
  wire _09670_;
  wire _09671_;
  wire _09672_;
  wire _09673_;
  wire _09674_;
  wire _09675_;
  wire _09676_;
  wire _09677_;
  wire _09678_;
  wire _09679_;
  wire _09680_;
  wire _09681_;
  wire _09682_;
  wire _09683_;
  wire _09684_;
  wire _09685_;
  wire _09686_;
  wire _09687_;
  wire _09688_;
  wire _09689_;
  wire _09690_;
  wire _09691_;
  wire _09692_;
  wire _09693_;
  wire _09694_;
  wire _09695_;
  wire _09696_;
  wire _09697_;
  wire _09698_;
  wire _09699_;
  wire _09700_;
  wire _09701_;
  wire _09702_;
  wire _09703_;
  wire _09704_;
  wire _09705_;
  wire _09706_;
  wire _09707_;
  wire _09708_;
  wire _09709_;
  wire _09710_;
  wire _09711_;
  wire _09712_;
  wire _09713_;
  wire _09714_;
  wire _09715_;
  wire _09716_;
  wire _09717_;
  wire _09718_;
  wire _09719_;
  wire _09720_;
  wire _09721_;
  wire _09722_;
  wire _09723_;
  wire _09724_;
  wire _09725_;
  wire _09726_;
  wire _09727_;
  wire _09728_;
  wire _09729_;
  wire _09730_;
  wire _09731_;
  wire _09732_;
  wire _09733_;
  wire _09734_;
  wire _09735_;
  wire _09736_;
  wire _09737_;
  wire _09738_;
  wire _09739_;
  wire _09740_;
  wire _09741_;
  wire _09742_;
  wire _09743_;
  wire _09744_;
  wire _09745_;
  wire _09746_;
  wire _09747_;
  wire _09748_;
  wire _09749_;
  wire _09750_;
  wire _09751_;
  wire _09752_;
  wire _09753_;
  wire _09754_;
  wire _09755_;
  wire _09756_;
  wire _09757_;
  wire _09758_;
  wire _09759_;
  wire _09760_;
  wire _09761_;
  wire _09762_;
  wire _09763_;
  wire _09764_;
  wire _09765_;
  wire _09766_;
  wire _09767_;
  wire _09768_;
  wire _09769_;
  wire _09770_;
  wire _09771_;
  wire _09772_;
  wire _09773_;
  wire _09774_;
  wire _09775_;
  wire _09776_;
  wire _09777_;
  wire _09778_;
  wire _09779_;
  wire _09780_;
  wire _09781_;
  wire _09782_;
  wire _09783_;
  wire _09784_;
  wire _09785_;
  wire _09786_;
  wire _09787_;
  wire _09788_;
  wire _09789_;
  wire _09790_;
  wire _09791_;
  wire _09792_;
  wire _09793_;
  wire _09794_;
  wire _09795_;
  wire _09796_;
  wire _09797_;
  wire _09798_;
  wire _09799_;
  wire _09800_;
  wire _09801_;
  wire _09802_;
  wire _09803_;
  wire _09804_;
  wire _09805_;
  wire _09806_;
  wire _09807_;
  wire _09808_;
  wire _09809_;
  wire _09810_;
  wire _09811_;
  wire _09812_;
  wire _09813_;
  wire _09814_;
  wire _09815_;
  wire _09816_;
  wire _09817_;
  wire _09818_;
  wire _09819_;
  wire _09820_;
  wire _09821_;
  wire _09822_;
  wire _09823_;
  wire _09824_;
  wire _09825_;
  wire _09826_;
  wire _09827_;
  wire _09828_;
  wire _09829_;
  wire _09830_;
  wire _09831_;
  wire _09832_;
  wire _09833_;
  wire _09834_;
  wire _09835_;
  wire _09836_;
  wire _09837_;
  wire _09838_;
  wire _09839_;
  wire _09840_;
  wire _09841_;
  wire _09842_;
  wire _09843_;
  wire _09844_;
  wire _09845_;
  wire _09846_;
  wire _09847_;
  wire _09848_;
  wire _09849_;
  wire _09850_;
  wire _09851_;
  wire _09852_;
  wire _09853_;
  wire _09854_;
  wire _09855_;
  wire _09856_;
  wire _09857_;
  wire _09858_;
  wire _09859_;
  wire _09860_;
  wire _09861_;
  wire _09862_;
  wire _09863_;
  wire _09864_;
  wire _09865_;
  wire _09866_;
  wire _09867_;
  wire _09868_;
  wire _09869_;
  wire _09870_;
  wire _09871_;
  wire _09872_;
  wire _09873_;
  wire _09874_;
  wire _09875_;
  wire _09876_;
  wire _09877_;
  wire _09878_;
  wire _09879_;
  wire _09880_;
  wire _09881_;
  wire _09882_;
  wire _09883_;
  wire _09884_;
  wire _09885_;
  wire _09886_;
  wire _09887_;
  wire _09888_;
  wire _09889_;
  wire _09890_;
  wire _09891_;
  wire _09892_;
  wire _09893_;
  wire _09894_;
  wire _09895_;
  wire _09896_;
  wire _09897_;
  wire _09898_;
  wire _09899_;
  wire _09900_;
  wire _09901_;
  wire _09902_;
  wire _09903_;
  wire _09904_;
  wire _09905_;
  wire _09906_;
  wire _09907_;
  wire _09908_;
  wire _09909_;
  wire _09910_;
  wire _09911_;
  wire _09912_;
  wire _09913_;
  wire _09914_;
  wire _09915_;
  wire _09916_;
  wire _09917_;
  wire _09918_;
  wire _09919_;
  wire _09920_;
  wire _09921_;
  wire _09922_;
  wire _09923_;
  wire _09924_;
  wire _09925_;
  wire _09926_;
  wire _09927_;
  wire _09928_;
  wire _09929_;
  wire _09930_;
  wire _09931_;
  wire _09932_;
  wire _09933_;
  wire _09934_;
  wire _09935_;
  wire _09936_;
  wire _09937_;
  wire _09938_;
  wire _09939_;
  wire _09940_;
  wire _09941_;
  wire _09942_;
  wire _09943_;
  wire _09944_;
  wire _09945_;
  wire _09946_;
  wire _09947_;
  wire _09948_;
  wire _09949_;
  wire _09950_;
  wire _09951_;
  wire _09952_;
  wire _09953_;
  wire _09954_;
  wire _09955_;
  wire _09956_;
  wire _09957_;
  wire _09958_;
  wire _09959_;
  wire _09960_;
  wire _09961_;
  wire _09962_;
  wire _09963_;
  wire _09964_;
  wire _09965_;
  wire _09966_;
  wire _09967_;
  wire _09968_;
  wire _09969_;
  wire _09970_;
  wire _09971_;
  wire _09972_;
  wire _09973_;
  wire _09974_;
  wire _09975_;
  wire _09976_;
  wire _09977_;
  wire _09978_;
  wire _09979_;
  wire _09980_;
  wire _09981_;
  wire _09982_;
  wire _09983_;
  wire _09984_;
  wire _09985_;
  wire _09986_;
  wire _09987_;
  wire _09988_;
  wire _09989_;
  wire _09990_;
  wire _09991_;
  wire _09992_;
  wire _09993_;
  wire _09994_;
  wire _09995_;
  wire _09996_;
  wire _09997_;
  wire _09998_;
  wire _09999_;
  wire _10000_;
  wire _10001_;
  wire _10002_;
  wire _10003_;
  wire _10004_;
  wire _10005_;
  wire _10006_;
  wire _10007_;
  wire _10008_;
  wire _10009_;
  wire _10010_;
  wire _10011_;
  wire _10012_;
  wire _10013_;
  wire _10014_;
  wire _10015_;
  wire _10016_;
  wire _10017_;
  wire _10018_;
  wire _10019_;
  wire _10020_;
  wire _10021_;
  wire _10022_;
  wire _10023_;
  wire _10024_;
  wire _10025_;
  wire _10026_;
  wire _10027_;
  wire _10028_;
  wire _10029_;
  wire _10030_;
  wire _10031_;
  wire _10032_;
  wire _10033_;
  wire _10034_;
  wire _10035_;
  wire _10036_;
  wire _10037_;
  wire _10038_;
  wire _10039_;
  wire _10040_;
  wire _10041_;
  wire _10042_;
  wire _10043_;
  wire _10044_;
  wire _10045_;
  wire _10046_;
  wire _10047_;
  wire _10048_;
  wire _10049_;
  wire _10050_;
  wire _10051_;
  wire _10052_;
  wire _10053_;
  wire _10054_;
  wire _10055_;
  wire _10056_;
  wire _10057_;
  wire _10058_;
  wire _10059_;
  wire _10060_;
  wire _10061_;
  wire _10062_;
  wire _10063_;
  wire _10064_;
  wire _10065_;
  wire _10066_;
  wire _10067_;
  wire _10068_;
  wire _10069_;
  wire _10070_;
  wire _10071_;
  wire _10072_;
  wire _10073_;
  wire _10074_;
  wire _10075_;
  wire _10076_;
  wire _10077_;
  wire _10078_;
  wire _10079_;
  wire _10080_;
  wire _10081_;
  wire _10082_;
  wire _10083_;
  wire _10084_;
  wire _10085_;
  wire _10086_;
  wire _10087_;
  wire _10088_;
  wire _10089_;
  wire _10090_;
  wire _10091_;
  wire _10092_;
  wire _10093_;
  wire _10094_;
  wire _10095_;
  wire _10096_;
  wire _10097_;
  wire _10098_;
  wire _10099_;
  wire _10100_;
  wire _10101_;
  wire _10102_;
  wire _10103_;
  wire _10104_;
  wire _10105_;
  wire _10106_;
  wire _10107_;
  wire _10108_;
  wire _10109_;
  wire _10110_;
  wire _10111_;
  wire _10112_;
  wire _10113_;
  wire _10114_;
  wire _10115_;
  wire _10116_;
  wire _10117_;
  wire _10118_;
  wire _10119_;
  wire _10120_;
  wire _10121_;
  wire _10122_;
  wire _10123_;
  wire _10124_;
  wire _10125_;
  wire _10126_;
  wire _10127_;
  wire _10128_;
  wire _10129_;
  wire _10130_;
  wire _10131_;
  wire _10132_;
  wire _10133_;
  wire _10134_;
  wire _10135_;
  wire _10136_;
  wire _10137_;
  wire _10138_;
  wire _10139_;
  wire _10140_;
  wire _10141_;
  wire _10142_;
  wire _10143_;
  wire _10144_;
  wire _10145_;
  wire _10146_;
  wire _10147_;
  wire _10148_;
  wire _10149_;
  wire _10150_;
  wire _10151_;
  wire _10152_;
  wire _10153_;
  wire _10154_;
  wire _10155_;
  wire _10156_;
  wire _10157_;
  wire _10158_;
  wire _10159_;
  wire _10160_;
  wire _10161_;
  wire _10162_;
  wire _10163_;
  wire _10164_;
  wire _10165_;
  wire _10166_;
  wire _10167_;
  wire _10168_;
  wire _10169_;
  wire _10170_;
  wire _10171_;
  wire _10172_;
  wire _10173_;
  wire _10174_;
  wire _10175_;
  wire _10176_;
  wire _10177_;
  wire _10178_;
  wire _10179_;
  wire _10180_;
  wire _10181_;
  wire _10182_;
  wire _10183_;
  wire _10184_;
  wire _10185_;
  wire _10186_;
  wire _10187_;
  wire _10188_;
  wire _10189_;
  wire _10190_;
  wire _10191_;
  wire _10192_;
  wire _10193_;
  wire _10194_;
  wire _10195_;
  wire _10196_;
  wire _10197_;
  wire _10198_;
  wire _10199_;
  wire _10200_;
  wire _10201_;
  wire _10202_;
  wire _10203_;
  wire _10204_;
  wire _10205_;
  wire _10206_;
  wire _10207_;
  wire _10208_;
  wire _10209_;
  wire _10210_;
  wire _10211_;
  wire _10212_;
  wire _10213_;
  wire _10214_;
  wire _10215_;
  wire _10216_;
  wire _10217_;
  wire _10218_;
  wire _10219_;
  wire _10220_;
  wire _10221_;
  wire _10222_;
  wire _10223_;
  wire _10224_;
  wire _10225_;
  wire _10226_;
  wire _10227_;
  wire _10228_;
  wire _10229_;
  wire _10230_;
  wire _10231_;
  wire _10232_;
  wire _10233_;
  wire _10234_;
  wire _10235_;
  wire _10236_;
  wire _10237_;
  wire _10238_;
  wire _10239_;
  wire _10240_;
  wire _10241_;
  wire _10242_;
  wire _10243_;
  wire _10244_;
  wire _10245_;
  wire _10246_;
  wire _10247_;
  wire _10248_;
  wire _10249_;
  wire _10250_;
  wire _10251_;
  wire _10252_;
  wire _10253_;
  wire _10254_;
  wire _10255_;
  wire _10256_;
  wire _10257_;
  wire _10258_;
  wire _10259_;
  wire _10260_;
  wire _10261_;
  wire _10262_;
  wire _10263_;
  wire _10264_;
  wire _10265_;
  wire _10266_;
  wire _10267_;
  wire _10268_;
  wire _10269_;
  wire _10270_;
  wire _10271_;
  wire _10272_;
  wire _10273_;
  wire _10274_;
  wire _10275_;
  wire _10276_;
  wire _10277_;
  wire _10278_;
  wire _10279_;
  wire _10280_;
  wire _10281_;
  wire _10282_;
  wire _10283_;
  wire _10284_;
  wire _10285_;
  wire _10286_;
  wire _10287_;
  wire _10288_;
  wire _10289_;
  wire _10290_;
  wire _10291_;
  wire _10292_;
  wire _10293_;
  wire _10294_;
  wire _10295_;
  wire _10296_;
  wire _10297_;
  wire _10298_;
  wire _10299_;
  wire _10300_;
  wire _10301_;
  wire _10302_;
  wire _10303_;
  wire _10304_;
  wire _10305_;
  wire _10306_;
  wire _10307_;
  wire _10308_;
  wire _10309_;
  wire _10310_;
  wire _10311_;
  wire _10312_;
  wire _10313_;
  wire _10314_;
  wire _10315_;
  wire _10316_;
  wire _10317_;
  wire _10318_;
  wire _10319_;
  wire _10320_;
  wire _10321_;
  wire _10322_;
  wire _10323_;
  wire _10324_;
  wire _10325_;
  wire _10326_;
  wire _10327_;
  wire _10328_;
  wire _10329_;
  wire _10330_;
  wire _10331_;
  wire _10332_;
  wire _10333_;
  wire _10334_;
  wire _10335_;
  wire _10336_;
  wire _10337_;
  wire _10338_;
  wire _10339_;
  wire _10340_;
  wire _10341_;
  wire _10342_;
  wire _10343_;
  wire _10344_;
  wire _10345_;
  wire _10346_;
  wire _10347_;
  wire _10348_;
  wire _10349_;
  wire _10350_;
  wire _10351_;
  wire _10352_;
  wire _10353_;
  wire _10354_;
  wire _10355_;
  wire _10356_;
  wire _10357_;
  wire _10358_;
  wire _10359_;
  wire _10360_;
  wire _10361_;
  wire _10362_;
  wire _10363_;
  wire _10364_;
  wire _10365_;
  wire _10366_;
  wire _10367_;
  wire _10368_;
  wire _10369_;
  wire _10370_;
  wire _10371_;
  wire _10372_;
  wire _10373_;
  wire _10374_;
  wire _10375_;
  wire _10376_;
  wire _10377_;
  wire _10378_;
  wire _10379_;
  wire _10380_;
  wire _10381_;
  wire _10382_;
  wire _10383_;
  wire _10384_;
  wire _10385_;
  wire _10386_;
  wire _10387_;
  wire _10388_;
  wire _10389_;
  wire _10390_;
  wire _10391_;
  wire _10392_;
  wire _10393_;
  wire _10394_;
  wire _10395_;
  wire _10396_;
  wire _10397_;
  wire _10398_;
  wire _10399_;
  wire _10400_;
  wire _10401_;
  wire _10402_;
  wire _10403_;
  wire _10404_;
  wire _10405_;
  wire _10406_;
  wire _10407_;
  wire _10408_;
  wire _10409_;
  wire _10410_;
  wire _10411_;
  wire _10412_;
  wire _10413_;
  wire _10414_;
  wire _10415_;
  wire _10416_;
  wire _10417_;
  wire _10418_;
  wire _10419_;
  wire _10420_;
  wire _10421_;
  wire _10422_;
  wire _10423_;
  wire _10424_;
  wire _10425_;
  wire _10426_;
  wire _10427_;
  wire _10428_;
  wire _10429_;
  wire _10430_;
  wire _10431_;
  wire _10432_;
  wire _10433_;
  wire _10434_;
  wire _10435_;
  wire _10436_;
  wire _10437_;
  wire _10438_;
  wire _10439_;
  wire _10440_;
  wire _10441_;
  wire _10442_;
  wire _10443_;
  wire _10444_;
  wire _10445_;
  wire _10446_;
  wire _10447_;
  wire _10448_;
  wire _10449_;
  wire _10450_;
  wire _10451_;
  wire _10452_;
  wire _10453_;
  wire _10454_;
  wire _10455_;
  wire _10456_;
  wire _10457_;
  wire _10458_;
  wire _10459_;
  wire _10460_;
  wire _10461_;
  wire _10462_;
  wire _10463_;
  wire _10464_;
  wire _10465_;
  wire _10466_;
  wire _10467_;
  wire _10468_;
  wire _10469_;
  wire _10470_;
  wire _10471_;
  wire _10472_;
  wire _10473_;
  wire _10474_;
  wire _10475_;
  wire _10476_;
  wire _10477_;
  wire _10478_;
  wire _10479_;
  wire _10480_;
  wire _10481_;
  wire _10482_;
  wire _10483_;
  wire _10484_;
  wire _10485_;
  wire _10486_;
  wire _10487_;
  wire _10488_;
  wire _10489_;
  wire _10490_;
  wire _10491_;
  wire _10492_;
  wire _10493_;
  wire _10494_;
  wire _10495_;
  wire _10496_;
  wire _10497_;
  wire _10498_;
  wire _10499_;
  wire _10500_;
  wire _10501_;
  wire _10502_;
  wire _10503_;
  wire _10504_;
  wire _10505_;
  wire _10506_;
  wire _10507_;
  wire _10508_;
  wire _10509_;
  wire _10510_;
  wire _10511_;
  wire _10512_;
  wire _10513_;
  wire _10514_;
  wire _10515_;
  wire _10516_;
  wire _10517_;
  wire _10518_;
  wire _10519_;
  wire _10520_;
  wire _10521_;
  wire _10522_;
  wire _10523_;
  wire _10524_;
  wire _10525_;
  wire _10526_;
  wire _10527_;
  wire _10528_;
  wire _10529_;
  wire _10530_;
  wire _10531_;
  wire _10532_;
  wire _10533_;
  wire _10534_;
  wire _10535_;
  wire _10536_;
  wire _10537_;
  wire _10538_;
  wire _10539_;
  wire _10540_;
  wire _10541_;
  wire _10542_;
  wire _10543_;
  wire _10544_;
  wire _10545_;
  wire _10546_;
  wire _10547_;
  wire _10548_;
  wire _10549_;
  wire _10550_;
  wire _10551_;
  wire _10552_;
  wire _10553_;
  wire _10554_;
  wire _10555_;
  wire _10556_;
  wire _10557_;
  wire _10558_;
  wire _10559_;
  wire _10560_;
  wire _10561_;
  wire _10562_;
  wire _10563_;
  wire _10564_;
  wire _10565_;
  wire _10566_;
  wire _10567_;
  wire _10568_;
  wire _10569_;
  wire _10570_;
  wire _10571_;
  wire _10572_;
  wire _10573_;
  wire _10574_;
  wire _10575_;
  wire _10576_;
  wire _10577_;
  wire _10578_;
  wire _10579_;
  wire _10580_;
  wire _10581_;
  wire _10582_;
  wire _10583_;
  wire _10584_;
  wire _10585_;
  wire _10586_;
  wire _10587_;
  wire _10588_;
  wire _10589_;
  wire _10590_;
  wire _10591_;
  wire _10592_;
  wire _10593_;
  wire _10594_;
  wire _10595_;
  wire _10596_;
  wire _10597_;
  wire _10598_;
  wire _10599_;
  wire _10600_;
  wire _10601_;
  wire _10602_;
  wire _10603_;
  wire _10604_;
  wire _10605_;
  wire _10606_;
  wire _10607_;
  wire _10608_;
  wire _10609_;
  wire _10610_;
  wire _10611_;
  wire _10612_;
  wire _10613_;
  wire _10614_;
  wire _10615_;
  wire _10616_;
  wire _10617_;
  wire _10618_;
  wire _10619_;
  wire _10620_;
  wire _10621_;
  wire _10622_;
  wire _10623_;
  wire _10624_;
  wire _10625_;
  wire _10626_;
  wire _10627_;
  wire _10628_;
  wire _10629_;
  wire _10630_;
  wire _10631_;
  wire _10632_;
  wire _10633_;
  wire _10634_;
  wire _10635_;
  wire _10636_;
  wire _10637_;
  wire _10638_;
  wire _10639_;
  wire _10640_;
  wire _10641_;
  wire _10642_;
  wire _10643_;
  wire _10644_;
  wire _10645_;
  wire _10646_;
  wire _10647_;
  wire _10648_;
  wire _10649_;
  wire _10650_;
  wire _10651_;
  wire _10652_;
  wire _10653_;
  wire _10654_;
  wire _10655_;
  wire _10656_;
  wire _10657_;
  wire _10658_;
  wire _10659_;
  wire _10660_;
  wire _10661_;
  wire _10662_;
  wire _10663_;
  wire _10664_;
  wire _10665_;
  wire _10666_;
  wire _10667_;
  wire _10668_;
  wire _10669_;
  wire _10670_;
  wire _10671_;
  wire _10672_;
  wire _10673_;
  wire _10674_;
  wire _10675_;
  wire _10676_;
  wire _10677_;
  wire _10678_;
  wire _10679_;
  wire _10680_;
  wire _10681_;
  wire _10682_;
  wire _10683_;
  wire _10684_;
  wire _10685_;
  wire _10686_;
  wire _10687_;
  wire _10688_;
  wire _10689_;
  wire _10690_;
  wire _10691_;
  wire _10692_;
  wire _10693_;
  wire _10694_;
  wire _10695_;
  wire _10696_;
  wire _10697_;
  wire _10698_;
  wire _10699_;
  wire _10700_;
  wire _10701_;
  wire _10702_;
  wire _10703_;
  wire _10704_;
  wire _10705_;
  wire _10706_;
  wire _10707_;
  wire _10708_;
  wire _10709_;
  wire _10710_;
  wire _10711_;
  wire _10712_;
  wire _10713_;
  wire _10714_;
  wire _10715_;
  wire _10716_;
  wire _10717_;
  wire _10718_;
  wire _10719_;
  wire _10720_;
  wire _10721_;
  wire _10722_;
  wire _10723_;
  wire _10724_;
  wire _10725_;
  wire _10726_;
  wire _10727_;
  wire _10728_;
  wire _10729_;
  wire _10730_;
  wire _10731_;
  wire _10732_;
  wire _10733_;
  wire _10734_;
  wire _10735_;
  wire _10736_;
  wire _10737_;
  wire _10738_;
  wire _10739_;
  wire _10740_;
  wire _10741_;
  wire _10742_;
  wire _10743_;
  wire _10744_;
  wire _10745_;
  wire _10746_;
  wire _10747_;
  wire _10748_;
  wire _10749_;
  wire _10750_;
  wire _10751_;
  wire _10752_;
  wire _10753_;
  wire _10754_;
  wire _10755_;
  wire _10756_;
  wire _10757_;
  wire _10758_;
  wire _10759_;
  wire _10760_;
  wire _10761_;
  wire _10762_;
  wire _10763_;
  wire _10764_;
  wire _10765_;
  wire _10766_;
  wire _10767_;
  wire _10768_;
  wire _10769_;
  wire _10770_;
  wire _10771_;
  wire _10772_;
  wire _10773_;
  wire _10774_;
  wire _10775_;
  wire _10776_;
  wire _10777_;
  wire _10778_;
  wire _10779_;
  wire _10780_;
  wire _10781_;
  wire _10782_;
  wire _10783_;
  wire _10784_;
  wire _10785_;
  wire _10786_;
  wire _10787_;
  wire _10788_;
  wire _10789_;
  wire _10790_;
  wire _10791_;
  wire _10792_;
  wire _10793_;
  wire _10794_;
  wire _10795_;
  wire _10796_;
  wire _10797_;
  wire _10798_;
  wire _10799_;
  wire _10800_;
  wire _10801_;
  wire _10802_;
  wire _10803_;
  wire _10804_;
  wire _10805_;
  wire _10806_;
  wire _10807_;
  wire _10808_;
  wire _10809_;
  wire _10810_;
  wire _10811_;
  wire _10812_;
  wire _10813_;
  wire _10814_;
  wire _10815_;
  wire _10816_;
  wire _10817_;
  wire _10818_;
  wire _10819_;
  wire _10820_;
  wire _10821_;
  wire _10822_;
  wire _10823_;
  wire _10824_;
  wire _10825_;
  wire _10826_;
  wire _10827_;
  wire _10828_;
  wire _10829_;
  wire _10830_;
  wire _10831_;
  wire _10832_;
  wire _10833_;
  wire _10834_;
  wire _10835_;
  wire _10836_;
  wire _10837_;
  wire _10838_;
  wire _10839_;
  wire _10840_;
  wire _10841_;
  wire _10842_;
  wire _10843_;
  wire _10844_;
  wire _10845_;
  wire _10846_;
  wire _10847_;
  wire _10848_;
  wire _10849_;
  wire _10850_;
  wire _10851_;
  wire _10852_;
  wire _10853_;
  wire _10854_;
  wire _10855_;
  wire _10856_;
  wire _10857_;
  wire _10858_;
  wire _10859_;
  wire _10860_;
  wire _10861_;
  wire _10862_;
  wire _10863_;
  wire _10864_;
  wire _10865_;
  wire _10866_;
  wire _10867_;
  wire _10868_;
  wire _10869_;
  wire _10870_;
  wire _10871_;
  wire _10872_;
  wire _10873_;
  wire _10874_;
  wire _10875_;
  wire _10876_;
  wire _10877_;
  wire _10878_;
  wire _10879_;
  wire _10880_;
  wire _10881_;
  wire _10882_;
  wire _10883_;
  wire _10884_;
  wire _10885_;
  wire _10886_;
  wire _10887_;
  wire _10888_;
  wire _10889_;
  wire _10890_;
  wire _10891_;
  wire _10892_;
  wire _10893_;
  wire _10894_;
  wire _10895_;
  wire _10896_;
  wire _10897_;
  wire _10898_;
  wire _10899_;
  wire _10900_;
  wire _10901_;
  wire _10902_;
  wire _10903_;
  wire _10904_;
  wire _10905_;
  wire _10906_;
  wire _10907_;
  wire _10908_;
  wire _10909_;
  wire _10910_;
  wire _10911_;
  wire _10912_;
  wire _10913_;
  wire _10914_;
  wire _10915_;
  wire _10916_;
  wire _10917_;
  wire _10918_;
  wire _10919_;
  wire _10920_;
  wire _10921_;
  wire _10922_;
  wire _10923_;
  wire _10924_;
  wire _10925_;
  wire _10926_;
  wire _10927_;
  wire _10928_;
  wire _10929_;
  wire _10930_;
  wire _10931_;
  wire _10932_;
  wire _10933_;
  wire _10934_;
  wire _10935_;
  wire _10936_;
  wire _10937_;
  wire _10938_;
  wire _10939_;
  wire _10940_;
  wire _10941_;
  wire _10942_;
  wire _10943_;
  wire _10944_;
  wire _10945_;
  wire _10946_;
  wire _10947_;
  wire _10948_;
  wire _10949_;
  wire _10950_;
  wire _10951_;
  wire _10952_;
  wire _10953_;
  wire _10954_;
  wire _10955_;
  wire _10956_;
  wire _10957_;
  wire _10958_;
  wire _10959_;
  wire _10960_;
  wire _10961_;
  wire _10962_;
  wire _10963_;
  wire _10964_;
  wire _10965_;
  wire _10966_;
  wire _10967_;
  wire _10968_;
  wire _10969_;
  wire _10970_;
  wire _10971_;
  wire _10972_;
  wire _10973_;
  wire _10974_;
  wire _10975_;
  wire _10976_;
  wire _10977_;
  wire _10978_;
  wire _10979_;
  wire _10980_;
  wire _10981_;
  wire _10982_;
  wire _10983_;
  wire _10984_;
  wire _10985_;
  wire _10986_;
  wire _10987_;
  wire _10988_;
  wire _10989_;
  wire _10990_;
  wire _10991_;
  wire _10992_;
  wire _10993_;
  wire _10994_;
  wire _10995_;
  wire _10996_;
  wire _10997_;
  wire _10998_;
  wire _10999_;
  wire _11000_;
  wire _11001_;
  wire _11002_;
  wire _11003_;
  wire _11004_;
  wire _11005_;
  wire _11006_;
  wire _11007_;
  wire _11008_;
  wire _11009_;
  wire _11010_;
  wire _11011_;
  wire _11012_;
  wire _11013_;
  wire _11014_;
  wire _11015_;
  wire _11016_;
  wire _11017_;
  wire _11018_;
  wire _11019_;
  wire _11020_;
  wire _11021_;
  wire _11022_;
  wire _11023_;
  wire _11024_;
  wire _11025_;
  wire _11026_;
  wire _11027_;
  wire _11028_;
  wire _11029_;
  wire _11030_;
  wire _11031_;
  wire _11032_;
  wire _11033_;
  wire _11034_;
  wire _11035_;
  wire _11036_;
  wire _11037_;
  wire _11038_;
  wire _11039_;
  wire _11040_;
  wire _11041_;
  wire _11042_;
  wire _11043_;
  wire _11044_;
  wire _11045_;
  wire _11046_;
  wire _11047_;
  wire _11048_;
  wire _11049_;
  wire _11050_;
  wire _11051_;
  wire _11052_;
  wire _11053_;
  wire _11054_;
  wire _11055_;
  wire _11056_;
  wire _11057_;
  wire _11058_;
  wire _11059_;
  wire _11060_;
  wire _11061_;
  wire _11062_;
  wire _11063_;
  wire _11064_;
  wire _11065_;
  wire _11066_;
  wire _11067_;
  wire _11068_;
  wire _11069_;
  wire _11070_;
  wire _11071_;
  wire _11072_;
  wire _11073_;
  wire _11074_;
  wire _11075_;
  wire _11076_;
  wire _11077_;
  wire _11078_;
  wire _11079_;
  wire _11080_;
  wire _11081_;
  wire _11082_;
  wire _11083_;
  wire _11084_;
  wire _11085_;
  wire _11086_;
  wire _11087_;
  wire _11088_;
  wire _11089_;
  wire _11090_;
  wire _11091_;
  wire _11092_;
  wire _11093_;
  wire _11094_;
  wire _11095_;
  wire _11096_;
  wire _11097_;
  wire _11098_;
  wire _11099_;
  wire _11100_;
  wire _11101_;
  wire _11102_;
  wire _11103_;
  wire _11104_;
  wire _11105_;
  wire _11106_;
  wire _11107_;
  wire _11108_;
  wire _11109_;
  wire _11110_;
  wire _11111_;
  wire _11112_;
  wire _11113_;
  wire _11114_;
  wire _11115_;
  wire _11116_;
  wire _11117_;
  wire _11118_;
  wire _11119_;
  wire _11120_;
  wire _11121_;
  wire _11122_;
  wire _11123_;
  wire _11124_;
  wire _11125_;
  wire _11126_;
  wire _11127_;
  wire _11128_;
  wire _11129_;
  wire _11130_;
  wire _11131_;
  wire _11132_;
  wire _11133_;
  wire _11134_;
  wire _11135_;
  wire _11136_;
  wire _11137_;
  wire _11138_;
  wire _11139_;
  wire _11140_;
  wire _11141_;
  wire _11142_;
  wire _11143_;
  wire _11144_;
  wire _11145_;
  wire _11146_;
  wire _11147_;
  wire _11148_;
  wire _11149_;
  wire _11150_;
  wire _11151_;
  wire _11152_;
  wire _11153_;
  wire _11154_;
  wire _11155_;
  wire _11156_;
  wire _11157_;
  wire _11158_;
  wire _11159_;
  wire _11160_;
  wire _11161_;
  wire _11162_;
  wire _11163_;
  wire _11164_;
  wire _11165_;
  wire _11166_;
  wire _11167_;
  wire _11168_;
  wire _11169_;
  wire _11170_;
  wire _11171_;
  wire _11172_;
  wire _11173_;
  wire _11174_;
  wire _11175_;
  wire _11176_;
  wire _11177_;
  wire _11178_;
  wire _11179_;
  wire _11180_;
  wire _11181_;
  wire _11182_;
  wire _11183_;
  wire _11184_;
  wire _11185_;
  wire _11186_;
  wire _11187_;
  wire _11188_;
  wire _11189_;
  wire _11190_;
  wire _11191_;
  wire _11192_;
  wire _11193_;
  wire _11194_;
  wire _11195_;
  wire _11196_;
  wire _11197_;
  wire _11198_;
  wire _11199_;
  wire _11200_;
  wire _11201_;
  wire _11202_;
  wire _11203_;
  wire _11204_;
  wire _11205_;
  wire _11206_;
  wire _11207_;
  wire _11208_;
  wire _11209_;
  wire _11210_;
  wire _11211_;
  wire _11212_;
  wire _11213_;
  wire _11214_;
  wire _11215_;
  wire _11216_;
  wire _11217_;
  wire _11218_;
  wire _11219_;
  wire _11220_;
  wire _11221_;
  wire _11222_;
  wire _11223_;
  wire _11224_;
  wire _11225_;
  wire _11226_;
  wire _11227_;
  wire _11228_;
  wire _11229_;
  wire _11230_;
  wire _11231_;
  wire _11232_;
  wire _11233_;
  wire _11234_;
  wire _11235_;
  wire _11236_;
  wire _11237_;
  wire _11238_;
  wire _11239_;
  wire _11240_;
  wire _11241_;
  wire _11242_;
  wire _11243_;
  wire _11244_;
  wire _11245_;
  wire _11246_;
  wire _11247_;
  wire _11248_;
  wire _11249_;
  wire _11250_;
  wire _11251_;
  wire _11252_;
  wire _11253_;
  wire _11254_;
  wire _11255_;
  wire _11256_;
  wire _11257_;
  wire _11258_;
  wire _11259_;
  wire _11260_;
  wire _11261_;
  wire _11262_;
  wire _11263_;
  wire _11264_;
  wire _11265_;
  wire _11266_;
  wire _11267_;
  wire _11268_;
  wire _11269_;
  wire _11270_;
  wire _11271_;
  wire _11272_;
  wire _11273_;
  wire _11274_;
  wire _11275_;
  wire _11276_;
  wire _11277_;
  wire _11278_;
  wire _11279_;
  wire _11280_;
  wire _11281_;
  wire _11282_;
  wire _11283_;
  wire _11284_;
  wire _11285_;
  wire _11286_;
  wire _11287_;
  wire _11288_;
  wire _11289_;
  wire _11290_;
  wire _11291_;
  wire _11292_;
  wire _11293_;
  wire _11294_;
  wire _11295_;
  wire _11296_;
  wire _11297_;
  wire _11298_;
  wire _11299_;
  wire _11300_;
  wire _11301_;
  wire _11302_;
  wire _11303_;
  wire _11304_;
  wire _11305_;
  wire _11306_;
  wire _11307_;
  wire _11308_;
  wire _11309_;
  wire _11310_;
  wire _11311_;
  wire _11312_;
  wire _11313_;
  wire _11314_;
  wire _11315_;
  wire _11316_;
  wire _11317_;
  wire _11318_;
  wire _11319_;
  wire _11320_;
  wire _11321_;
  wire _11322_;
  wire _11323_;
  wire _11324_;
  wire _11325_;
  wire _11326_;
  wire _11327_;
  wire _11328_;
  wire _11329_;
  wire _11330_;
  wire _11331_;
  wire _11332_;
  wire _11333_;
  wire _11334_;
  wire _11335_;
  wire _11336_;
  wire _11337_;
  wire _11338_;
  wire _11339_;
  wire _11340_;
  wire _11341_;
  wire _11342_;
  wire _11343_;
  wire _11344_;
  wire _11345_;
  wire _11346_;
  wire _11347_;
  wire _11348_;
  wire _11349_;
  wire _11350_;
  wire _11351_;
  wire _11352_;
  wire _11353_;
  wire _11354_;
  wire _11355_;
  wire _11356_;
  wire _11357_;
  wire _11358_;
  wire _11359_;
  wire _11360_;
  wire _11361_;
  wire _11362_;
  wire _11363_;
  wire _11364_;
  wire _11365_;
  wire _11366_;
  wire _11367_;
  wire _11368_;
  wire _11369_;
  wire _11370_;
  wire _11371_;
  wire _11372_;
  wire _11373_;
  wire _11374_;
  wire _11375_;
  wire _11376_;
  wire _11377_;
  wire _11378_;
  wire _11379_;
  wire _11380_;
  wire _11381_;
  wire _11382_;
  wire _11383_;
  wire _11384_;
  wire _11385_;
  wire _11386_;
  wire _11387_;
  wire _11388_;
  wire _11389_;
  wire _11390_;
  wire _11391_;
  wire _11392_;
  wire _11393_;
  wire _11394_;
  wire _11395_;
  wire _11396_;
  wire _11397_;
  wire _11398_;
  wire _11399_;
  wire _11400_;
  wire _11401_;
  wire _11402_;
  wire _11403_;
  wire _11404_;
  wire _11405_;
  wire _11406_;
  wire _11407_;
  wire _11408_;
  wire _11409_;
  wire _11410_;
  wire _11411_;
  wire _11412_;
  wire _11413_;
  wire _11414_;
  wire _11415_;
  wire _11416_;
  wire _11417_;
  wire _11418_;
  wire _11419_;
  wire _11420_;
  wire _11421_;
  wire _11422_;
  wire _11423_;
  wire _11424_;
  wire _11425_;
  wire _11426_;
  wire _11427_;
  wire _11428_;
  wire _11429_;
  wire _11430_;
  wire _11431_;
  wire _11432_;
  wire _11433_;
  wire _11434_;
  wire _11435_;
  wire _11436_;
  wire _11437_;
  wire _11438_;
  wire _11439_;
  wire _11440_;
  wire _11441_;
  wire _11442_;
  wire _11443_;
  wire _11444_;
  wire _11445_;
  wire _11446_;
  wire _11447_;
  wire _11448_;
  wire _11449_;
  wire _11450_;
  wire _11451_;
  wire _11452_;
  wire _11453_;
  wire _11454_;
  wire _11455_;
  wire _11456_;
  wire _11457_;
  wire _11458_;
  wire _11459_;
  wire _11460_;
  wire _11461_;
  wire _11462_;
  wire _11463_;
  wire _11464_;
  wire _11465_;
  wire _11466_;
  wire _11467_;
  wire _11468_;
  wire _11469_;
  wire _11470_;
  wire _11471_;
  wire _11472_;
  wire _11473_;
  wire _11474_;
  wire _11475_;
  wire _11476_;
  wire _11477_;
  wire _11478_;
  wire _11479_;
  wire _11480_;
  wire _11481_;
  wire _11482_;
  wire _11483_;
  wire _11484_;
  wire _11485_;
  wire _11486_;
  wire _11487_;
  wire _11488_;
  wire _11489_;
  wire _11490_;
  wire _11491_;
  wire _11492_;
  wire _11493_;
  wire _11494_;
  wire _11495_;
  wire _11496_;
  wire _11497_;
  wire _11498_;
  wire _11499_;
  wire _11500_;
  wire _11501_;
  wire _11502_;
  wire _11503_;
  wire _11504_;
  wire _11505_;
  wire _11506_;
  wire _11507_;
  wire _11508_;
  wire _11509_;
  wire _11510_;
  wire _11511_;
  wire _11512_;
  wire _11513_;
  wire _11514_;
  wire _11515_;
  wire _11516_;
  wire _11517_;
  wire _11518_;
  wire _11519_;
  wire _11520_;
  wire _11521_;
  wire _11522_;
  wire _11523_;
  wire _11524_;
  wire _11525_;
  wire _11526_;
  wire _11527_;
  wire _11528_;
  wire _11529_;
  wire _11530_;
  wire _11531_;
  wire _11532_;
  wire _11533_;
  wire _11534_;
  wire _11535_;
  wire _11536_;
  wire _11537_;
  wire _11538_;
  wire _11539_;
  wire _11540_;
  wire _11541_;
  wire _11542_;
  wire _11543_;
  wire _11544_;
  wire _11545_;
  wire _11546_;
  wire _11547_;
  wire _11548_;
  wire _11549_;
  wire _11550_;
  wire _11551_;
  wire _11552_;
  wire _11553_;
  wire _11554_;
  wire _11555_;
  wire _11556_;
  wire _11557_;
  wire _11558_;
  wire _11559_;
  wire _11560_;
  wire _11561_;
  wire _11562_;
  wire _11563_;
  wire _11564_;
  wire _11565_;
  wire _11566_;
  wire _11567_;
  wire _11568_;
  wire _11569_;
  wire _11570_;
  wire _11571_;
  wire _11572_;
  wire _11573_;
  wire _11574_;
  wire _11575_;
  wire _11576_;
  wire _11577_;
  wire _11578_;
  wire _11579_;
  wire _11580_;
  wire _11581_;
  wire _11582_;
  wire _11583_;
  wire _11584_;
  wire _11585_;
  wire _11586_;
  wire _11587_;
  wire _11588_;
  wire _11589_;
  wire _11590_;
  wire _11591_;
  wire _11592_;
  wire _11593_;
  wire _11594_;
  wire _11595_;
  wire _11596_;
  wire _11597_;
  wire _11598_;
  wire _11599_;
  wire _11600_;
  wire _11601_;
  wire _11602_;
  wire _11603_;
  wire _11604_;
  wire _11605_;
  wire _11606_;
  wire _11607_;
  wire _11608_;
  wire _11609_;
  wire _11610_;
  wire _11611_;
  wire _11612_;
  wire _11613_;
  wire _11614_;
  wire _11615_;
  wire _11616_;
  wire _11617_;
  wire _11618_;
  wire _11619_;
  wire _11620_;
  wire _11621_;
  wire _11622_;
  wire _11623_;
  wire _11624_;
  wire _11625_;
  wire _11626_;
  wire _11627_;
  wire _11628_;
  wire _11629_;
  wire _11630_;
  wire _11631_;
  wire _11632_;
  wire _11633_;
  wire _11634_;
  wire _11635_;
  wire _11636_;
  wire _11637_;
  wire _11638_;
  wire _11639_;
  wire _11640_;
  wire _11641_;
  wire _11642_;
  wire _11643_;
  wire _11644_;
  wire _11645_;
  wire _11646_;
  wire _11647_;
  wire _11648_;
  wire _11649_;
  wire _11650_;
  wire _11651_;
  wire _11652_;
  wire _11653_;
  wire _11654_;
  wire _11655_;
  wire _11656_;
  wire _11657_;
  wire _11658_;
  wire _11659_;
  wire _11660_;
  wire _11661_;
  wire _11662_;
  wire _11663_;
  wire _11664_;
  wire _11665_;
  wire _11666_;
  wire _11667_;
  wire _11668_;
  wire _11669_;
  wire _11670_;
  wire _11671_;
  wire _11672_;
  wire _11673_;
  wire _11674_;
  wire _11675_;
  wire _11676_;
  wire _11677_;
  wire _11678_;
  wire _11679_;
  wire _11680_;
  wire _11681_;
  wire _11682_;
  wire _11683_;
  wire _11684_;
  wire _11685_;
  wire _11686_;
  wire _11687_;
  wire _11688_;
  wire _11689_;
  wire _11690_;
  wire _11691_;
  wire _11692_;
  wire _11693_;
  wire _11694_;
  wire _11695_;
  wire _11696_;
  wire _11697_;
  wire _11698_;
  wire _11699_;
  wire _11700_;
  wire _11701_;
  wire _11702_;
  wire _11703_;
  wire _11704_;
  wire _11705_;
  wire _11706_;
  wire _11707_;
  wire _11708_;
  wire _11709_;
  wire _11710_;
  wire _11711_;
  wire _11712_;
  wire _11713_;
  wire _11714_;
  wire _11715_;
  wire _11716_;
  wire _11717_;
  wire _11718_;
  wire _11719_;
  wire _11720_;
  wire _11721_;
  wire _11722_;
  wire _11723_;
  wire _11724_;
  wire _11725_;
  wire _11726_;
  wire _11727_;
  wire _11728_;
  wire _11729_;
  wire _11730_;
  wire _11731_;
  wire _11732_;
  wire _11733_;
  wire _11734_;
  wire _11735_;
  wire _11736_;
  wire _11737_;
  wire _11738_;
  wire _11739_;
  wire _11740_;
  wire _11741_;
  wire _11742_;
  wire _11743_;
  wire _11744_;
  wire _11745_;
  wire _11746_;
  wire _11747_;
  wire _11748_;
  wire _11749_;
  wire _11750_;
  wire _11751_;
  wire _11752_;
  wire _11753_;
  wire _11754_;
  wire _11755_;
  wire _11756_;
  wire _11757_;
  wire _11758_;
  wire _11759_;
  wire _11760_;
  wire _11761_;
  wire _11762_;
  wire _11763_;
  wire _11764_;
  wire _11765_;
  wire _11766_;
  wire _11767_;
  wire _11768_;
  wire _11769_;
  wire _11770_;
  wire _11771_;
  wire _11772_;
  wire _11773_;
  wire _11774_;
  wire _11775_;
  wire _11776_;
  wire _11777_;
  wire _11778_;
  wire _11779_;
  wire _11780_;
  wire _11781_;
  wire _11782_;
  wire _11783_;
  wire _11784_;
  wire _11785_;
  wire _11786_;
  wire _11787_;
  wire _11788_;
  wire _11789_;
  wire _11790_;
  wire _11791_;
  wire _11792_;
  wire _11793_;
  wire _11794_;
  wire _11795_;
  wire _11796_;
  wire _11797_;
  wire _11798_;
  wire _11799_;
  wire _11800_;
  wire _11801_;
  wire _11802_;
  wire _11803_;
  wire _11804_;
  wire _11805_;
  wire _11806_;
  wire _11807_;
  wire _11808_;
  wire _11809_;
  wire _11810_;
  wire _11811_;
  wire _11812_;
  wire _11813_;
  wire _11814_;
  wire _11815_;
  wire _11816_;
  wire _11817_;
  wire _11818_;
  wire _11819_;
  wire _11820_;
  wire _11821_;
  wire _11822_;
  wire _11823_;
  wire _11824_;
  wire _11825_;
  wire _11826_;
  wire _11827_;
  wire _11828_;
  wire _11829_;
  wire _11830_;
  wire _11831_;
  wire _11832_;
  wire _11833_;
  wire _11834_;
  wire _11835_;
  wire _11836_;
  wire _11837_;
  wire _11838_;
  wire _11839_;
  wire _11840_;
  wire _11841_;
  wire _11842_;
  wire _11843_;
  wire _11844_;
  wire _11845_;
  wire _11846_;
  wire _11847_;
  wire _11848_;
  wire _11849_;
  wire _11850_;
  wire _11851_;
  wire _11852_;
  wire _11853_;
  wire _11854_;
  wire _11855_;
  wire _11856_;
  wire _11857_;
  wire _11858_;
  wire _11859_;
  wire _11860_;
  wire _11861_;
  wire _11862_;
  wire _11863_;
  wire _11864_;
  wire _11865_;
  wire _11866_;
  wire _11867_;
  wire _11868_;
  wire _11869_;
  wire _11870_;
  wire _11871_;
  wire _11872_;
  wire _11873_;
  wire _11874_;
  wire _11875_;
  wire _11876_;
  wire _11877_;
  wire _11878_;
  wire _11879_;
  wire _11880_;
  wire _11881_;
  wire _11882_;
  wire _11883_;
  wire _11884_;
  wire _11885_;
  wire _11886_;
  wire _11887_;
  wire _11888_;
  wire _11889_;
  wire _11890_;
  wire _11891_;
  wire _11892_;
  wire _11893_;
  wire _11894_;
  wire _11895_;
  wire _11896_;
  wire _11897_;
  wire _11898_;
  wire _11899_;
  wire _11900_;
  wire _11901_;
  wire _11902_;
  wire _11903_;
  wire _11904_;
  wire _11905_;
  wire _11906_;
  wire _11907_;
  wire _11908_;
  wire _11909_;
  wire _11910_;
  wire _11911_;
  wire _11912_;
  wire _11913_;
  wire _11914_;
  wire _11915_;
  wire _11916_;
  wire _11917_;
  wire _11918_;
  wire _11919_;
  wire _11920_;
  wire _11921_;
  wire _11922_;
  wire _11923_;
  wire _11924_;
  wire _11925_;
  wire _11926_;
  wire _11927_;
  wire _11928_;
  wire _11929_;
  wire _11930_;
  wire _11931_;
  wire _11932_;
  wire _11933_;
  wire _11934_;
  wire _11935_;
  wire _11936_;
  wire _11937_;
  wire _11938_;
  wire _11939_;
  wire _11940_;
  wire _11941_;
  wire _11942_;
  wire _11943_;
  wire _11944_;
  wire _11945_;
  wire _11946_;
  wire _11947_;
  wire _11948_;
  wire _11949_;
  wire _11950_;
  wire _11951_;
  wire _11952_;
  wire _11953_;
  wire _11954_;
  wire _11955_;
  wire _11956_;
  wire _11957_;
  wire _11958_;
  wire _11959_;
  wire _11960_;
  wire _11961_;
  wire _11962_;
  wire _11963_;
  wire _11964_;
  wire _11965_;
  wire _11966_;
  wire _11967_;
  wire _11968_;
  wire _11969_;
  wire _11970_;
  wire _11971_;
  wire _11972_;
  wire _11973_;
  wire _11974_;
  wire _11975_;
  wire _11976_;
  wire _11977_;
  wire _11978_;
  wire _11979_;
  wire _11980_;
  wire _11981_;
  wire _11982_;
  wire _11983_;
  wire _11984_;
  wire _11985_;
  wire _11986_;
  wire _11987_;
  wire _11988_;
  wire _11989_;
  wire _11990_;
  wire _11991_;
  wire _11992_;
  wire _11993_;
  wire _11994_;
  wire _11995_;
  wire _11996_;
  wire _11997_;
  wire _11998_;
  wire _11999_;
  wire _12000_;
  wire _12001_;
  wire _12002_;
  wire _12003_;
  wire _12004_;
  wire _12005_;
  wire _12006_;
  wire _12007_;
  wire _12008_;
  wire _12009_;
  wire _12010_;
  wire _12011_;
  wire _12012_;
  wire _12013_;
  wire _12014_;
  wire _12015_;
  wire _12016_;
  wire _12017_;
  wire _12018_;
  wire _12019_;
  wire _12020_;
  wire _12021_;
  wire _12022_;
  wire _12023_;
  wire _12024_;
  wire _12025_;
  wire _12026_;
  wire _12027_;
  wire _12028_;
  wire _12029_;
  wire _12030_;
  wire _12031_;
  wire _12032_;
  wire _12033_;
  wire _12034_;
  wire _12035_;
  wire _12036_;
  wire _12037_;
  wire _12038_;
  wire _12039_;
  wire _12040_;
  wire _12041_;
  wire _12042_;
  wire _12043_;
  wire _12044_;
  wire _12045_;
  wire _12046_;
  wire _12047_;
  wire _12048_;
  wire _12049_;
  wire _12050_;
  wire _12051_;
  wire _12052_;
  wire _12053_;
  wire _12054_;
  wire _12055_;
  wire _12056_;
  wire _12057_;
  wire _12058_;
  wire _12059_;
  wire _12060_;
  wire _12061_;
  wire _12062_;
  wire _12063_;
  wire _12064_;
  wire _12065_;
  wire _12066_;
  wire _12067_;
  wire _12068_;
  wire _12069_;
  wire _12070_;
  wire _12071_;
  wire _12072_;
  wire _12073_;
  wire _12074_;
  wire _12075_;
  wire _12076_;
  wire _12077_;
  wire _12078_;
  wire _12079_;
  wire _12080_;
  wire _12081_;
  wire _12082_;
  wire _12083_;
  wire _12084_;
  wire _12085_;
  wire _12086_;
  wire _12087_;
  wire _12088_;
  wire _12089_;
  wire _12090_;
  wire _12091_;
  wire _12092_;
  wire _12093_;
  wire _12094_;
  wire _12095_;
  wire _12096_;
  wire _12097_;
  wire _12098_;
  wire _12099_;
  wire _12100_;
  wire _12101_;
  wire _12102_;
  wire _12103_;
  wire _12104_;
  wire _12105_;
  wire _12106_;
  wire _12107_;
  wire _12108_;
  wire _12109_;
  wire _12110_;
  wire _12111_;
  wire _12112_;
  wire _12113_;
  wire _12114_;
  wire _12115_;
  wire _12116_;
  wire _12117_;
  wire _12118_;
  wire _12119_;
  wire _12120_;
  wire _12121_;
  wire _12122_;
  wire _12123_;
  wire _12124_;
  wire _12125_;
  wire _12126_;
  wire _12127_;
  wire _12128_;
  wire _12129_;
  wire _12130_;
  wire _12131_;
  wire _12132_;
  wire _12133_;
  wire _12134_;
  wire _12135_;
  wire _12136_;
  wire _12137_;
  wire _12138_;
  wire _12139_;
  wire _12140_;
  wire _12141_;
  wire _12142_;
  wire _12143_;
  wire _12144_;
  wire _12145_;
  wire _12146_;
  wire _12147_;
  wire _12148_;
  wire _12149_;
  wire _12150_;
  wire _12151_;
  wire _12152_;
  wire _12153_;
  wire _12154_;
  wire _12155_;
  wire _12156_;
  wire _12157_;
  wire _12158_;
  wire _12159_;
  wire _12160_;
  wire _12161_;
  wire _12162_;
  wire _12163_;
  wire _12164_;
  wire _12165_;
  wire _12166_;
  wire _12167_;
  wire _12168_;
  wire _12169_;
  wire _12170_;
  wire _12171_;
  wire _12172_;
  wire _12173_;
  wire _12174_;
  wire _12175_;
  wire _12176_;
  wire _12177_;
  wire _12178_;
  wire _12179_;
  wire _12180_;
  wire _12181_;
  wire _12182_;
  wire _12183_;
  wire _12184_;
  wire _12185_;
  wire _12186_;
  wire _12187_;
  wire _12188_;
  wire _12189_;
  wire _12190_;
  wire _12191_;
  wire _12192_;
  wire _12193_;
  wire _12194_;
  wire _12195_;
  wire _12196_;
  wire _12197_;
  wire _12198_;
  wire _12199_;
  wire _12200_;
  wire _12201_;
  wire _12202_;
  wire _12203_;
  wire _12204_;
  wire _12205_;
  wire _12206_;
  wire _12207_;
  wire _12208_;
  wire _12209_;
  wire _12210_;
  wire _12211_;
  wire _12212_;
  wire _12213_;
  wire _12214_;
  wire _12215_;
  wire _12216_;
  wire _12217_;
  wire _12218_;
  wire _12219_;
  wire _12220_;
  wire _12221_;
  wire _12222_;
  wire _12223_;
  wire _12224_;
  wire _12225_;
  wire _12226_;
  wire _12227_;
  wire _12228_;
  wire _12229_;
  wire _12230_;
  wire _12231_;
  wire _12232_;
  wire _12233_;
  wire _12234_;
  wire _12235_;
  wire _12236_;
  wire _12237_;
  wire _12238_;
  wire _12239_;
  wire _12240_;
  wire _12241_;
  wire _12242_;
  wire _12243_;
  wire _12244_;
  wire _12245_;
  wire _12246_;
  wire _12247_;
  wire _12248_;
  wire _12249_;
  wire _12250_;
  wire _12251_;
  wire _12252_;
  wire _12253_;
  wire _12254_;
  wire _12255_;
  wire _12256_;
  wire _12257_;
  wire _12258_;
  wire _12259_;
  wire _12260_;
  wire _12261_;
  wire _12262_;
  wire _12263_;
  wire _12264_;
  wire _12265_;
  wire _12266_;
  wire _12267_;
  wire _12268_;
  wire _12269_;
  wire _12270_;
  wire _12271_;
  wire _12272_;
  wire _12273_;
  wire _12274_;
  wire _12275_;
  wire _12276_;
  wire _12277_;
  wire _12278_;
  wire _12279_;
  wire _12280_;
  wire _12281_;
  wire _12282_;
  wire _12283_;
  wire _12284_;
  wire _12285_;
  wire _12286_;
  wire _12287_;
  wire _12288_;
  wire _12289_;
  wire _12290_;
  wire _12291_;
  wire _12292_;
  wire _12293_;
  wire _12294_;
  wire _12295_;
  wire _12296_;
  wire _12297_;
  wire _12298_;
  wire _12299_;
  wire _12300_;
  wire _12301_;
  wire _12302_;
  wire _12303_;
  wire _12304_;
  wire _12305_;
  wire _12306_;
  wire _12307_;
  wire _12308_;
  wire _12309_;
  wire _12310_;
  wire _12311_;
  wire _12312_;
  wire _12313_;
  wire _12314_;
  wire _12315_;
  wire _12316_;
  wire _12317_;
  wire _12318_;
  wire _12319_;
  wire _12320_;
  wire _12321_;
  wire _12322_;
  wire _12323_;
  wire _12324_;
  wire _12325_;
  wire _12326_;
  wire _12327_;
  wire _12328_;
  wire _12329_;
  wire _12330_;
  wire _12331_;
  wire _12332_;
  wire _12333_;
  wire _12334_;
  wire _12335_;
  wire _12336_;
  wire _12337_;
  wire _12338_;
  wire _12339_;
  wire _12340_;
  wire _12341_;
  wire _12342_;
  wire _12343_;
  wire _12344_;
  wire _12345_;
  wire _12346_;
  wire _12347_;
  wire _12348_;
  wire _12349_;
  wire _12350_;
  wire _12351_;
  wire _12352_;
  wire _12353_;
  wire _12354_;
  wire _12355_;
  wire _12356_;
  wire _12357_;
  wire _12358_;
  wire _12359_;
  wire _12360_;
  wire _12361_;
  wire _12362_;
  wire _12363_;
  wire _12364_;
  wire _12365_;
  wire _12366_;
  wire _12367_;
  wire _12368_;
  wire _12369_;
  wire _12370_;
  wire _12371_;
  wire _12372_;
  wire _12373_;
  wire _12374_;
  wire _12375_;
  wire _12376_;
  wire _12377_;
  wire _12378_;
  wire _12379_;
  wire _12380_;
  wire _12381_;
  wire _12382_;
  wire _12383_;
  wire _12384_;
  wire _12385_;
  wire _12386_;
  wire _12387_;
  wire _12388_;
  wire _12389_;
  wire _12390_;
  wire _12391_;
  wire _12392_;
  wire _12393_;
  wire _12394_;
  wire _12395_;
  wire _12396_;
  wire _12397_;
  wire _12398_;
  wire _12399_;
  wire _12400_;
  wire _12401_;
  wire _12402_;
  wire _12403_;
  wire _12404_;
  wire _12405_;
  wire _12406_;
  wire _12407_;
  wire _12408_;
  wire _12409_;
  wire _12410_;
  wire _12411_;
  wire _12412_;
  wire _12413_;
  wire _12414_;
  wire _12415_;
  wire _12416_;
  wire _12417_;
  wire _12418_;
  wire _12419_;
  wire _12420_;
  wire _12421_;
  wire _12422_;
  wire _12423_;
  wire _12424_;
  wire _12425_;
  wire _12426_;
  wire _12427_;
  wire _12428_;
  wire _12429_;
  wire _12430_;
  wire _12431_;
  wire _12432_;
  wire _12433_;
  wire _12434_;
  wire _12435_;
  wire _12436_;
  wire _12437_;
  wire _12438_;
  wire _12439_;
  wire _12440_;
  wire _12441_;
  wire _12442_;
  wire _12443_;
  wire _12444_;
  wire _12445_;
  wire _12446_;
  wire _12447_;
  wire _12448_;
  wire _12449_;
  wire _12450_;
  wire _12451_;
  wire _12452_;
  wire _12453_;
  wire _12454_;
  wire _12455_;
  wire _12456_;
  wire _12457_;
  wire _12458_;
  wire _12459_;
  wire _12460_;
  wire _12461_;
  wire _12462_;
  wire _12463_;
  wire _12464_;
  wire _12465_;
  wire _12466_;
  wire _12467_;
  wire _12468_;
  wire _12469_;
  wire _12470_;
  wire _12471_;
  wire _12472_;
  wire _12473_;
  wire _12474_;
  wire _12475_;
  wire _12476_;
  wire _12477_;
  wire _12478_;
  wire _12479_;
  wire _12480_;
  wire _12481_;
  wire _12482_;
  wire _12483_;
  wire _12484_;
  wire _12485_;
  wire _12486_;
  wire _12487_;
  wire _12488_;
  wire _12489_;
  wire _12490_;
  wire _12491_;
  wire _12492_;
  wire _12493_;
  wire _12494_;
  wire _12495_;
  wire _12496_;
  wire _12497_;
  wire _12498_;
  wire _12499_;
  wire _12500_;
  wire _12501_;
  wire _12502_;
  wire _12503_;
  wire _12504_;
  wire _12505_;
  wire _12506_;
  wire _12507_;
  wire _12508_;
  wire _12509_;
  wire _12510_;
  wire _12511_;
  wire _12512_;
  wire _12513_;
  wire _12514_;
  wire _12515_;
  wire _12516_;
  wire _12517_;
  wire _12518_;
  wire _12519_;
  wire _12520_;
  wire _12521_;
  wire _12522_;
  wire _12523_;
  wire _12524_;
  wire _12525_;
  wire _12526_;
  wire _12527_;
  wire _12528_;
  wire _12529_;
  wire _12530_;
  wire _12531_;
  wire _12532_;
  wire _12533_;
  wire _12534_;
  wire _12535_;
  wire _12536_;
  wire _12537_;
  wire _12538_;
  wire _12539_;
  wire _12540_;
  wire _12541_;
  wire _12542_;
  wire _12543_;
  wire _12544_;
  wire _12545_;
  wire _12546_;
  wire _12547_;
  wire _12548_;
  wire _12549_;
  wire _12550_;
  wire _12551_;
  wire _12552_;
  wire _12553_;
  wire _12554_;
  wire _12555_;
  wire _12556_;
  wire _12557_;
  wire _12558_;
  wire _12559_;
  wire _12560_;
  wire _12561_;
  wire _12562_;
  wire _12563_;
  wire _12564_;
  wire _12565_;
  wire _12566_;
  wire _12567_;
  wire _12568_;
  wire _12569_;
  wire _12570_;
  wire _12571_;
  wire _12572_;
  wire _12573_;
  wire _12574_;
  wire _12575_;
  wire _12576_;
  wire _12577_;
  wire _12578_;
  wire _12579_;
  wire _12580_;
  wire _12581_;
  wire _12582_;
  wire _12583_;
  wire _12584_;
  wire _12585_;
  wire _12586_;
  wire _12587_;
  wire _12588_;
  wire _12589_;
  wire _12590_;
  wire _12591_;
  wire _12592_;
  wire _12593_;
  wire _12594_;
  wire _12595_;
  wire _12596_;
  wire _12597_;
  wire _12598_;
  wire _12599_;
  wire _12600_;
  wire _12601_;
  wire _12602_;
  wire _12603_;
  wire _12604_;
  wire _12605_;
  wire _12606_;
  wire _12607_;
  wire _12608_;
  wire _12609_;
  wire _12610_;
  wire _12611_;
  wire _12612_;
  wire _12613_;
  wire _12614_;
  wire _12615_;
  wire _12616_;
  wire _12617_;
  wire _12618_;
  wire _12619_;
  wire _12620_;
  wire _12621_;
  wire _12622_;
  wire _12623_;
  wire _12624_;
  wire _12625_;
  wire _12626_;
  wire _12627_;
  wire _12628_;
  wire _12629_;
  wire _12630_;
  wire _12631_;
  wire _12632_;
  wire _12633_;
  wire _12634_;
  wire _12635_;
  wire _12636_;
  wire _12637_;
  wire _12638_;
  wire _12639_;
  wire _12640_;
  wire _12641_;
  wire _12642_;
  wire _12643_;
  wire _12644_;
  wire _12645_;
  wire _12646_;
  wire _12647_;
  wire _12648_;
  wire _12649_;
  wire _12650_;
  wire _12651_;
  wire _12652_;
  wire _12653_;
  wire _12654_;
  wire _12655_;
  wire _12656_;
  wire _12657_;
  wire _12658_;
  wire _12659_;
  wire _12660_;
  wire _12661_;
  wire _12662_;
  wire _12663_;
  wire _12664_;
  wire _12665_;
  wire _12666_;
  wire _12667_;
  wire _12668_;
  wire _12669_;
  wire _12670_;
  wire _12671_;
  wire _12672_;
  wire _12673_;
  wire _12674_;
  wire _12675_;
  wire _12676_;
  wire _12677_;
  wire _12678_;
  wire _12679_;
  wire _12680_;
  wire _12681_;
  wire _12682_;
  wire _12683_;
  wire _12684_;
  wire _12685_;
  wire _12686_;
  wire _12687_;
  wire _12688_;
  wire _12689_;
  wire _12690_;
  wire _12691_;
  wire _12692_;
  wire _12693_;
  wire _12694_;
  wire _12695_;
  wire _12696_;
  wire _12697_;
  wire _12698_;
  wire _12699_;
  wire _12700_;
  wire _12701_;
  wire _12702_;
  wire _12703_;
  wire _12704_;
  wire _12705_;
  wire _12706_;
  wire _12707_;
  wire _12708_;
  wire _12709_;
  wire _12710_;
  wire _12711_;
  wire _12712_;
  wire _12713_;
  wire _12714_;
  wire _12715_;
  wire _12716_;
  wire _12717_;
  wire _12718_;
  wire _12719_;
  wire _12720_;
  wire _12721_;
  wire _12722_;
  wire _12723_;
  wire _12724_;
  wire _12725_;
  wire _12726_;
  wire _12727_;
  wire _12728_;
  wire _12729_;
  wire _12730_;
  wire _12731_;
  wire _12732_;
  wire _12733_;
  wire _12734_;
  wire _12735_;
  wire _12736_;
  wire _12737_;
  wire _12738_;
  wire _12739_;
  wire _12740_;
  wire _12741_;
  wire _12742_;
  wire _12743_;
  wire _12744_;
  wire _12745_;
  wire _12746_;
  wire _12747_;
  wire _12748_;
  wire _12749_;
  wire _12750_;
  wire _12751_;
  wire _12752_;
  wire _12753_;
  wire _12754_;
  wire _12755_;
  wire _12756_;
  wire _12757_;
  wire _12758_;
  wire _12759_;
  wire _12760_;
  wire _12761_;
  wire _12762_;
  wire _12763_;
  wire _12764_;
  wire _12765_;
  wire _12766_;
  wire _12767_;
  wire _12768_;
  wire _12769_;
  wire _12770_;
  wire _12771_;
  wire _12772_;
  wire _12773_;
  wire _12774_;
  wire _12775_;
  wire _12776_;
  wire _12777_;
  wire _12778_;
  wire _12779_;
  wire _12780_;
  wire _12781_;
  wire _12782_;
  wire _12783_;
  wire _12784_;
  wire _12785_;
  wire _12786_;
  wire _12787_;
  wire _12788_;
  wire _12789_;
  wire _12790_;
  wire _12791_;
  wire _12792_;
  wire _12793_;
  wire _12794_;
  wire _12795_;
  wire _12796_;
  wire _12797_;
  wire _12798_;
  wire _12799_;
  wire _12800_;
  wire _12801_;
  wire _12802_;
  wire _12803_;
  wire _12804_;
  wire _12805_;
  wire _12806_;
  wire _12807_;
  wire _12808_;
  wire _12809_;
  wire _12810_;
  wire _12811_;
  wire _12812_;
  wire _12813_;
  wire _12814_;
  wire _12815_;
  wire _12816_;
  wire _12817_;
  wire _12818_;
  wire _12819_;
  wire _12820_;
  wire _12821_;
  wire _12822_;
  wire _12823_;
  wire _12824_;
  wire _12825_;
  wire _12826_;
  wire _12827_;
  wire _12828_;
  wire _12829_;
  wire _12830_;
  wire _12831_;
  wire _12832_;
  wire _12833_;
  wire _12834_;
  wire _12835_;
  wire _12836_;
  wire _12837_;
  wire _12838_;
  wire _12839_;
  wire _12840_;
  wire _12841_;
  wire _12842_;
  wire _12843_;
  wire _12844_;
  wire _12845_;
  wire _12846_;
  wire _12847_;
  wire _12848_;
  wire _12849_;
  wire _12850_;
  wire _12851_;
  wire _12852_;
  wire _12853_;
  wire _12854_;
  wire _12855_;
  wire _12856_;
  wire _12857_;
  wire _12858_;
  wire _12859_;
  wire _12860_;
  wire _12861_;
  wire _12862_;
  wire _12863_;
  wire _12864_;
  wire _12865_;
  wire _12866_;
  wire _12867_;
  wire _12868_;
  wire _12869_;
  wire _12870_;
  wire _12871_;
  wire _12872_;
  wire _12873_;
  wire _12874_;
  wire _12875_;
  wire _12876_;
  wire _12877_;
  wire _12878_;
  wire _12879_;
  wire _12880_;
  wire _12881_;
  wire _12882_;
  wire _12883_;
  wire _12884_;
  wire _12885_;
  wire _12886_;
  wire _12887_;
  wire _12888_;
  wire _12889_;
  wire _12890_;
  wire _12891_;
  wire _12892_;
  wire _12893_;
  wire _12894_;
  wire _12895_;
  wire _12896_;
  wire _12897_;
  wire _12898_;
  wire _12899_;
  wire _12900_;
  wire _12901_;
  wire _12902_;
  wire _12903_;
  wire _12904_;
  wire _12905_;
  wire _12906_;
  wire _12907_;
  wire _12908_;
  wire _12909_;
  wire _12910_;
  wire _12911_;
  wire _12912_;
  wire _12913_;
  wire _12914_;
  wire _12915_;
  wire _12916_;
  wire _12917_;
  wire _12918_;
  wire _12919_;
  wire _12920_;
  wire _12921_;
  wire _12922_;
  wire _12923_;
  wire _12924_;
  wire _12925_;
  wire _12926_;
  wire _12927_;
  wire _12928_;
  wire _12929_;
  wire _12930_;
  wire _12931_;
  wire _12932_;
  wire _12933_;
  wire _12934_;
  wire _12935_;
  wire _12936_;
  wire _12937_;
  wire _12938_;
  wire _12939_;
  wire _12940_;
  wire _12941_;
  wire _12942_;
  wire _12943_;
  wire _12944_;
  wire _12945_;
  wire _12946_;
  wire _12947_;
  wire _12948_;
  wire _12949_;
  wire _12950_;
  wire _12951_;
  wire _12952_;
  wire _12953_;
  wire _12954_;
  wire _12955_;
  wire _12956_;
  wire _12957_;
  wire _12958_;
  wire _12959_;
  wire _12960_;
  wire _12961_;
  wire _12962_;
  wire _12963_;
  wire _12964_;
  wire _12965_;
  wire _12966_;
  wire _12967_;
  wire _12968_;
  wire _12969_;
  wire _12970_;
  wire _12971_;
  wire _12972_;
  wire _12973_;
  wire _12974_;
  wire _12975_;
  wire _12976_;
  wire _12977_;
  wire _12978_;
  wire _12979_;
  wire _12980_;
  wire _12981_;
  wire _12982_;
  wire _12983_;
  wire _12984_;
  wire _12985_;
  wire _12986_;
  wire _12987_;
  wire _12988_;
  wire _12989_;
  wire _12990_;
  wire _12991_;
  wire _12992_;
  wire _12993_;
  wire _12994_;
  wire _12995_;
  wire _12996_;
  wire _12997_;
  wire _12998_;
  wire _12999_;
  wire _13000_;
  wire _13001_;
  wire _13002_;
  wire _13003_;
  wire _13004_;
  wire _13005_;
  wire _13006_;
  wire _13007_;
  wire _13008_;
  wire _13009_;
  wire _13010_;
  wire _13011_;
  wire _13012_;
  wire _13013_;
  wire _13014_;
  wire _13015_;
  wire _13016_;
  wire _13017_;
  wire _13018_;
  wire _13019_;
  wire _13020_;
  wire _13021_;
  wire _13022_;
  wire _13023_;
  wire _13024_;
  wire _13025_;
  wire _13026_;
  wire _13027_;
  wire _13028_;
  wire _13029_;
  wire _13030_;
  wire _13031_;
  wire _13032_;
  wire _13033_;
  wire _13034_;
  wire _13035_;
  wire _13036_;
  wire _13037_;
  wire _13038_;
  wire _13039_;
  wire _13040_;
  wire _13041_;
  wire _13042_;
  wire _13043_;
  wire _13044_;
  wire _13045_;
  wire _13046_;
  wire _13047_;
  wire _13048_;
  wire _13049_;
  wire _13050_;
  wire _13051_;
  wire _13052_;
  wire _13053_;
  wire _13054_;
  wire _13055_;
  wire _13056_;
  wire _13057_;
  wire _13058_;
  wire _13059_;
  wire _13060_;
  wire _13061_;
  wire _13062_;
  wire _13063_;
  wire _13064_;
  wire _13065_;
  wire _13066_;
  wire _13067_;
  wire _13068_;
  wire _13069_;
  wire _13070_;
  wire _13071_;
  wire _13072_;
  wire _13073_;
  wire _13074_;
  wire _13075_;
  wire _13076_;
  wire _13077_;
  wire _13078_;
  wire _13079_;
  wire _13080_;
  wire _13081_;
  wire _13082_;
  wire _13083_;
  wire _13084_;
  wire _13085_;
  wire _13086_;
  wire _13087_;
  wire _13088_;
  wire _13089_;
  wire _13090_;
  wire _13091_;
  wire _13092_;
  wire _13093_;
  wire _13094_;
  wire _13095_;
  wire _13096_;
  wire _13097_;
  wire _13098_;
  wire _13099_;
  wire _13100_;
  wire _13101_;
  wire _13102_;
  wire _13103_;
  wire _13104_;
  wire _13105_;
  wire _13106_;
  wire _13107_;
  wire _13108_;
  wire _13109_;
  wire _13110_;
  wire _13111_;
  wire _13112_;
  wire _13113_;
  wire _13114_;
  wire _13115_;
  wire _13116_;
  wire _13117_;
  wire _13118_;
  wire _13119_;
  wire _13120_;
  wire _13121_;
  wire _13122_;
  wire _13123_;
  wire _13124_;
  wire _13125_;
  wire _13126_;
  wire _13127_;
  wire _13128_;
  wire _13129_;
  wire _13130_;
  wire _13131_;
  wire _13132_;
  wire _13133_;
  wire _13134_;
  wire _13135_;
  wire _13136_;
  wire _13137_;
  wire _13138_;
  wire _13139_;
  wire _13140_;
  wire _13141_;
  wire _13142_;
  wire _13143_;
  wire _13144_;
  wire _13145_;
  wire _13146_;
  wire _13147_;
  wire _13148_;
  wire _13149_;
  wire _13150_;
  wire _13151_;
  wire _13152_;
  wire _13153_;
  wire _13154_;
  wire _13155_;
  wire _13156_;
  wire _13157_;
  wire _13158_;
  wire _13159_;
  wire _13160_;
  wire _13161_;
  wire _13162_;
  wire _13163_;
  wire _13164_;
  wire _13165_;
  wire _13166_;
  wire _13167_;
  wire _13168_;
  wire _13169_;
  wire _13170_;
  wire _13171_;
  wire _13172_;
  wire _13173_;
  wire _13174_;
  wire _13175_;
  wire _13176_;
  wire _13177_;
  wire _13178_;
  wire _13179_;
  wire _13180_;
  wire _13181_;
  wire _13182_;
  wire _13183_;
  wire _13184_;
  wire _13185_;
  wire _13186_;
  wire _13187_;
  wire _13188_;
  wire _13189_;
  wire _13190_;
  wire _13191_;
  wire _13192_;
  wire _13193_;
  wire _13194_;
  wire _13195_;
  wire _13196_;
  wire _13197_;
  wire _13198_;
  wire _13199_;
  wire _13200_;
  wire _13201_;
  wire _13202_;
  wire _13203_;
  wire _13204_;
  wire _13205_;
  wire _13206_;
  wire _13207_;
  wire _13208_;
  wire _13209_;
  wire _13210_;
  wire _13211_;
  wire _13212_;
  wire _13213_;
  wire _13214_;
  wire _13215_;
  wire _13216_;
  wire _13217_;
  wire _13218_;
  wire _13219_;
  wire _13220_;
  wire _13221_;
  wire _13222_;
  wire _13223_;
  wire _13224_;
  wire _13225_;
  wire _13226_;
  wire _13227_;
  wire _13228_;
  wire _13229_;
  wire _13230_;
  wire _13231_;
  wire _13232_;
  wire _13233_;
  wire _13234_;
  wire _13235_;
  wire _13236_;
  wire _13237_;
  wire _13238_;
  wire _13239_;
  wire _13240_;
  wire _13241_;
  wire _13242_;
  wire _13243_;
  wire _13244_;
  wire _13245_;
  wire _13246_;
  wire _13247_;
  wire _13248_;
  wire _13249_;
  wire _13250_;
  wire _13251_;
  wire _13252_;
  wire _13253_;
  wire _13254_;
  wire _13255_;
  wire _13256_;
  wire _13257_;
  wire _13258_;
  wire _13259_;
  wire _13260_;
  wire _13261_;
  wire _13262_;
  wire _13263_;
  wire _13264_;
  wire _13265_;
  wire _13266_;
  wire _13267_;
  wire _13268_;
  wire _13269_;
  wire _13270_;
  wire _13271_;
  wire _13272_;
  wire _13273_;
  wire _13274_;
  wire _13275_;
  wire _13276_;
  wire _13277_;
  wire _13278_;
  wire _13279_;
  wire _13280_;
  wire _13281_;
  wire _13282_;
  wire _13283_;
  wire _13284_;
  wire _13285_;
  wire _13286_;
  wire _13287_;
  wire _13288_;
  wire _13289_;
  wire _13290_;
  wire _13291_;
  wire _13292_;
  wire _13293_;
  wire _13294_;
  wire _13295_;
  wire _13296_;
  wire _13297_;
  wire _13298_;
  wire _13299_;
  wire _13300_;
  wire _13301_;
  wire _13302_;
  wire _13303_;
  wire _13304_;
  wire _13305_;
  wire _13306_;
  wire _13307_;
  wire _13308_;
  wire _13309_;
  wire _13310_;
  wire _13311_;
  wire _13312_;
  wire _13313_;
  wire _13314_;
  wire _13315_;
  wire _13316_;
  wire _13317_;
  wire _13318_;
  wire _13319_;
  wire _13320_;
  wire _13321_;
  wire _13322_;
  wire _13323_;
  wire _13324_;
  wire _13325_;
  wire _13326_;
  wire _13327_;
  wire _13328_;
  wire _13329_;
  wire _13330_;
  wire _13331_;
  wire _13332_;
  wire _13333_;
  wire _13334_;
  wire _13335_;
  wire _13336_;
  wire _13337_;
  wire _13338_;
  wire _13339_;
  wire _13340_;
  wire _13341_;
  wire _13342_;
  wire _13343_;
  wire _13344_;
  wire _13345_;
  wire _13346_;
  wire _13347_;
  wire _13348_;
  wire _13349_;
  wire _13350_;
  wire _13351_;
  wire _13352_;
  wire _13353_;
  wire _13354_;
  wire _13355_;
  wire _13356_;
  wire _13357_;
  wire _13358_;
  wire _13359_;
  wire _13360_;
  wire _13361_;
  wire _13362_;
  wire _13363_;
  wire _13364_;
  wire _13365_;
  wire _13366_;
  wire _13367_;
  wire _13368_;
  wire _13369_;
  wire _13370_;
  wire _13371_;
  wire _13372_;
  wire _13373_;
  wire _13374_;
  wire _13375_;
  wire _13376_;
  wire _13377_;
  wire _13378_;
  wire _13379_;
  wire _13380_;
  wire _13381_;
  wire _13382_;
  wire _13383_;
  wire _13384_;
  wire _13385_;
  wire _13386_;
  wire _13387_;
  wire _13388_;
  wire _13389_;
  wire _13390_;
  wire _13391_;
  wire _13392_;
  wire _13393_;
  wire _13394_;
  wire _13395_;
  wire _13396_;
  wire _13397_;
  wire _13398_;
  wire _13399_;
  wire _13400_;
  wire _13401_;
  wire _13402_;
  wire _13403_;
  wire _13404_;
  wire _13405_;
  wire _13406_;
  wire _13407_;
  wire _13408_;
  wire _13409_;
  wire _13410_;
  wire _13411_;
  wire _13412_;
  wire _13413_;
  wire _13414_;
  wire _13415_;
  wire _13416_;
  wire _13417_;
  wire _13418_;
  wire _13419_;
  wire _13420_;
  wire _13421_;
  wire _13422_;
  wire _13423_;
  wire _13424_;
  wire _13425_;
  wire _13426_;
  wire _13427_;
  wire _13428_;
  wire _13429_;
  wire _13430_;
  wire _13431_;
  wire _13432_;
  wire _13433_;
  wire _13434_;
  wire _13435_;
  wire _13436_;
  wire _13437_;
  wire _13438_;
  wire _13439_;
  wire _13440_;
  wire _13441_;
  wire _13442_;
  wire _13443_;
  wire _13444_;
  wire _13445_;
  wire _13446_;
  wire _13447_;
  wire _13448_;
  wire _13449_;
  wire _13450_;
  wire _13451_;
  wire _13452_;
  wire _13453_;
  wire _13454_;
  wire _13455_;
  wire _13456_;
  wire _13457_;
  wire _13458_;
  wire _13459_;
  wire _13460_;
  wire _13461_;
  wire _13462_;
  wire _13463_;
  wire _13464_;
  wire _13465_;
  wire _13466_;
  wire _13467_;
  wire _13468_;
  wire _13469_;
  wire _13470_;
  wire _13471_;
  wire _13472_;
  wire _13473_;
  wire _13474_;
  wire _13475_;
  wire _13476_;
  wire _13477_;
  wire _13478_;
  wire _13479_;
  wire _13480_;
  wire _13481_;
  wire _13482_;
  wire _13483_;
  wire _13484_;
  wire _13485_;
  wire _13486_;
  wire _13487_;
  wire _13488_;
  wire _13489_;
  wire _13490_;
  wire _13491_;
  wire _13492_;
  wire _13493_;
  wire _13494_;
  wire _13495_;
  wire _13496_;
  wire _13497_;
  wire _13498_;
  wire _13499_;
  wire _13500_;
  wire _13501_;
  wire _13502_;
  wire _13503_;
  wire _13504_;
  wire _13505_;
  wire _13506_;
  wire _13507_;
  wire _13508_;
  wire _13509_;
  wire _13510_;
  wire _13511_;
  wire _13512_;
  wire _13513_;
  wire _13514_;
  wire _13515_;
  wire _13516_;
  wire _13517_;
  wire _13518_;
  wire _13519_;
  wire _13520_;
  wire _13521_;
  wire _13522_;
  wire _13523_;
  wire _13524_;
  wire _13525_;
  wire _13526_;
  wire _13527_;
  wire _13528_;
  wire _13529_;
  wire _13530_;
  wire _13531_;
  wire _13532_;
  wire _13533_;
  wire _13534_;
  wire _13535_;
  wire _13536_;
  wire _13537_;
  wire _13538_;
  wire _13539_;
  wire _13540_;
  wire _13541_;
  wire _13542_;
  wire _13543_;
  wire _13544_;
  wire _13545_;
  wire _13546_;
  wire _13547_;
  wire _13548_;
  wire _13549_;
  wire _13550_;
  wire _13551_;
  wire _13552_;
  wire _13553_;
  wire _13554_;
  wire _13555_;
  wire _13556_;
  wire _13557_;
  wire _13558_;
  wire _13559_;
  wire _13560_;
  wire _13561_;
  wire _13562_;
  wire _13563_;
  wire _13564_;
  wire _13565_;
  wire _13566_;
  wire _13567_;
  wire _13568_;
  wire _13569_;
  wire _13570_;
  wire _13571_;
  wire _13572_;
  wire _13573_;
  wire _13574_;
  wire _13575_;
  wire _13576_;
  wire _13577_;
  wire _13578_;
  wire _13579_;
  wire _13580_;
  wire _13581_;
  wire _13582_;
  wire _13583_;
  wire _13584_;
  wire _13585_;
  wire _13586_;
  wire _13587_;
  wire _13588_;
  wire _13589_;
  wire _13590_;
  wire _13591_;
  wire _13592_;
  wire _13593_;
  wire _13594_;
  wire _13595_;
  wire _13596_;
  wire _13597_;
  wire _13598_;
  wire _13599_;
  wire _13600_;
  wire _13601_;
  wire _13602_;
  wire _13603_;
  wire _13604_;
  wire _13605_;
  wire _13606_;
  wire _13607_;
  wire _13608_;
  wire _13609_;
  wire _13610_;
  wire _13611_;
  wire _13612_;
  wire _13613_;
  wire _13614_;
  wire _13615_;
  wire _13616_;
  wire _13617_;
  wire _13618_;
  wire _13619_;
  wire _13620_;
  wire _13621_;
  wire _13622_;
  wire _13623_;
  wire _13624_;
  wire _13625_;
  wire _13626_;
  wire _13627_;
  wire _13628_;
  wire _13629_;
  wire _13630_;
  wire _13631_;
  wire _13632_;
  wire _13633_;
  wire _13634_;
  wire _13635_;
  wire _13636_;
  wire _13637_;
  wire _13638_;
  wire _13639_;
  wire _13640_;
  wire _13641_;
  wire _13642_;
  wire _13643_;
  wire _13644_;
  wire _13645_;
  wire _13646_;
  wire _13647_;
  wire _13648_;
  wire _13649_;
  wire _13650_;
  wire _13651_;
  wire _13652_;
  wire _13653_;
  wire _13654_;
  wire _13655_;
  wire _13656_;
  wire _13657_;
  wire _13658_;
  wire _13659_;
  wire _13660_;
  wire _13661_;
  wire _13662_;
  wire _13663_;
  wire _13664_;
  wire _13665_;
  wire _13666_;
  wire _13667_;
  wire _13668_;
  wire _13669_;
  wire _13670_;
  wire _13671_;
  wire _13672_;
  wire _13673_;
  wire _13674_;
  wire _13675_;
  wire _13676_;
  wire _13677_;
  wire _13678_;
  wire _13679_;
  wire _13680_;
  wire _13681_;
  wire _13682_;
  wire _13683_;
  wire _13684_;
  wire _13685_;
  wire _13686_;
  wire _13687_;
  wire _13688_;
  wire _13689_;
  wire _13690_;
  wire _13691_;
  wire _13692_;
  wire _13693_;
  wire _13694_;
  wire _13695_;
  wire _13696_;
  wire _13697_;
  wire _13698_;
  wire _13699_;
  wire _13700_;
  wire _13701_;
  wire _13702_;
  wire _13703_;
  wire _13704_;
  wire _13705_;
  wire _13706_;
  wire _13707_;
  wire _13708_;
  wire _13709_;
  wire _13710_;
  wire _13711_;
  wire _13712_;
  wire _13713_;
  wire _13714_;
  wire _13715_;
  wire _13716_;
  wire _13717_;
  wire _13718_;
  wire _13719_;
  wire _13720_;
  wire _13721_;
  wire _13722_;
  wire _13723_;
  wire _13724_;
  wire _13725_;
  wire _13726_;
  wire _13727_;
  wire _13728_;
  wire _13729_;
  wire _13730_;
  wire _13731_;
  wire _13732_;
  wire _13733_;
  wire _13734_;
  wire _13735_;
  wire _13736_;
  wire _13737_;
  wire _13738_;
  wire _13739_;
  wire _13740_;
  wire _13741_;
  wire _13742_;
  wire _13743_;
  wire _13744_;
  wire _13745_;
  wire _13746_;
  wire _13747_;
  wire _13748_;
  wire _13749_;
  wire _13750_;
  wire _13751_;
  wire _13752_;
  wire _13753_;
  wire _13754_;
  wire _13755_;
  wire _13756_;
  wire _13757_;
  wire _13758_;
  wire _13759_;
  wire _13760_;
  wire _13761_;
  wire _13762_;
  wire _13763_;
  wire _13764_;
  wire _13765_;
  wire _13766_;
  wire _13767_;
  wire _13768_;
  wire _13769_;
  wire _13770_;
  wire _13771_;
  wire _13772_;
  wire _13773_;
  wire _13774_;
  wire _13775_;
  wire _13776_;
  wire _13777_;
  wire _13778_;
  wire _13779_;
  wire _13780_;
  wire _13781_;
  wire _13782_;
  wire _13783_;
  wire _13784_;
  wire _13785_;
  wire _13786_;
  wire _13787_;
  wire _13788_;
  wire _13789_;
  wire _13790_;
  wire _13791_;
  wire _13792_;
  wire _13793_;
  wire _13794_;
  wire _13795_;
  wire _13796_;
  wire _13797_;
  wire _13798_;
  wire _13799_;
  wire _13800_;
  wire _13801_;
  wire _13802_;
  wire _13803_;
  wire _13804_;
  wire _13805_;
  wire _13806_;
  wire _13807_;
  wire _13808_;
  wire _13809_;
  wire _13810_;
  wire _13811_;
  wire _13812_;
  wire _13813_;
  wire _13814_;
  wire _13815_;
  wire _13816_;
  wire _13817_;
  wire _13818_;
  wire _13819_;
  wire _13820_;
  wire _13821_;
  wire _13822_;
  wire _13823_;
  wire _13824_;
  wire _13825_;
  wire _13826_;
  wire _13827_;
  wire _13828_;
  wire _13829_;
  wire _13830_;
  wire _13831_;
  wire _13832_;
  wire _13833_;
  wire _13834_;
  wire _13835_;
  wire _13836_;
  wire _13837_;
  wire _13838_;
  wire _13839_;
  wire _13840_;
  wire _13841_;
  wire _13842_;
  wire _13843_;
  wire _13844_;
  wire _13845_;
  wire _13846_;
  wire _13847_;
  wire _13848_;
  wire _13849_;
  wire _13850_;
  wire _13851_;
  wire _13852_;
  wire _13853_;
  wire _13854_;
  wire _13855_;
  wire _13856_;
  wire _13857_;
  wire _13858_;
  wire _13859_;
  wire _13860_;
  wire _13861_;
  wire _13862_;
  wire _13863_;
  wire _13864_;
  wire _13865_;
  wire _13866_;
  wire _13867_;
  wire _13868_;
  wire _13869_;
  wire _13870_;
  wire _13871_;
  wire _13872_;
  wire _13873_;
  wire _13874_;
  wire _13875_;
  wire _13876_;
  wire _13877_;
  wire _13878_;
  wire _13879_;
  wire _13880_;
  wire _13881_;
  wire _13882_;
  wire _13883_;
  wire _13884_;
  wire _13885_;
  wire _13886_;
  wire _13887_;
  wire _13888_;
  wire _13889_;
  wire _13890_;
  wire _13891_;
  wire _13892_;
  wire _13893_;
  wire _13894_;
  wire _13895_;
  wire _13896_;
  wire _13897_;
  wire _13898_;
  wire _13899_;
  wire _13900_;
  wire _13901_;
  wire _13902_;
  wire _13903_;
  wire _13904_;
  wire _13905_;
  wire _13906_;
  wire _13907_;
  wire _13908_;
  wire _13909_;
  wire _13910_;
  wire _13911_;
  wire _13912_;
  wire _13913_;
  wire _13914_;
  wire _13915_;
  wire _13916_;
  wire _13917_;
  wire _13918_;
  wire _13919_;
  wire _13920_;
  wire _13921_;
  wire _13922_;
  wire _13923_;
  wire _13924_;
  wire _13925_;
  wire _13926_;
  wire _13927_;
  wire _13928_;
  wire _13929_;
  wire _13930_;
  wire _13931_;
  wire _13932_;
  wire _13933_;
  wire _13934_;
  wire _13935_;
  wire _13936_;
  wire _13937_;
  wire _13938_;
  wire _13939_;
  wire _13940_;
  wire _13941_;
  wire _13942_;
  wire _13943_;
  wire _13944_;
  wire _13945_;
  wire _13946_;
  wire _13947_;
  wire _13948_;
  wire _13949_;
  wire _13950_;
  wire _13951_;
  wire _13952_;
  wire _13953_;
  wire _13954_;
  wire _13955_;
  wire _13956_;
  wire _13957_;
  wire _13958_;
  wire _13959_;
  wire _13960_;
  wire _13961_;
  wire _13962_;
  wire _13963_;
  wire _13964_;
  wire _13965_;
  wire _13966_;
  wire _13967_;
  wire _13968_;
  wire _13969_;
  wire _13970_;
  wire _13971_;
  wire _13972_;
  wire _13973_;
  wire _13974_;
  wire _13975_;
  wire _13976_;
  wire _13977_;
  wire _13978_;
  wire _13979_;
  wire _13980_;
  wire _13981_;
  wire _13982_;
  wire _13983_;
  wire _13984_;
  wire _13985_;
  wire _13986_;
  wire _13987_;
  wire _13988_;
  wire _13989_;
  wire _13990_;
  wire _13991_;
  wire _13992_;
  wire _13993_;
  wire _13994_;
  wire _13995_;
  wire _13996_;
  wire _13997_;
  wire _13998_;
  wire _13999_;
  wire _14000_;
  wire _14001_;
  wire _14002_;
  wire _14003_;
  wire _14004_;
  wire _14005_;
  wire _14006_;
  wire _14007_;
  wire _14008_;
  wire _14009_;
  wire _14010_;
  wire _14011_;
  wire _14012_;
  wire _14013_;
  wire _14014_;
  wire _14015_;
  wire _14016_;
  wire _14017_;
  wire _14018_;
  wire _14019_;
  wire _14020_;
  wire _14021_;
  wire _14022_;
  wire _14023_;
  wire _14024_;
  wire _14025_;
  wire _14026_;
  wire _14027_;
  wire _14028_;
  wire _14029_;
  wire _14030_;
  wire _14031_;
  wire _14032_;
  wire _14033_;
  wire _14034_;
  wire _14035_;
  wire _14036_;
  wire _14037_;
  wire _14038_;
  wire _14039_;
  wire _14040_;
  wire _14041_;
  wire _14042_;
  wire _14043_;
  wire _14044_;
  wire _14045_;
  wire _14046_;
  wire _14047_;
  wire _14048_;
  wire _14049_;
  wire _14050_;
  wire _14051_;
  wire _14052_;
  wire _14053_;
  wire _14054_;
  wire _14055_;
  wire _14056_;
  wire _14057_;
  wire _14058_;
  wire _14059_;
  wire _14060_;
  wire _14061_;
  wire _14062_;
  wire _14063_;
  wire _14064_;
  wire _14065_;
  wire _14066_;
  wire _14067_;
  wire _14068_;
  wire _14069_;
  wire _14070_;
  wire _14071_;
  wire _14072_;
  wire _14073_;
  wire _14074_;
  wire _14075_;
  wire _14076_;
  wire _14077_;
  wire _14078_;
  wire _14079_;
  wire _14080_;
  wire _14081_;
  wire _14082_;
  wire _14083_;
  wire _14084_;
  wire _14085_;
  wire _14086_;
  wire _14087_;
  wire _14088_;
  wire _14089_;
  wire _14090_;
  wire _14091_;
  wire _14092_;
  wire _14093_;
  wire _14094_;
  wire _14095_;
  wire _14096_;
  wire _14097_;
  wire _14098_;
  wire _14099_;
  wire _14100_;
  wire _14101_;
  wire _14102_;
  wire _14103_;
  wire _14104_;
  wire _14105_;
  wire _14106_;
  wire _14107_;
  wire _14108_;
  wire _14109_;
  wire _14110_;
  wire _14111_;
  wire _14112_;
  wire _14113_;
  wire _14114_;
  wire _14115_;
  wire _14116_;
  wire _14117_;
  wire _14118_;
  wire _14119_;
  wire _14120_;
  wire _14121_;
  wire _14122_;
  wire _14123_;
  wire _14124_;
  wire _14125_;
  wire _14126_;
  wire _14127_;
  wire _14128_;
  wire _14129_;
  wire _14130_;
  wire _14131_;
  wire _14132_;
  wire _14133_;
  wire _14134_;
  wire _14135_;
  wire _14136_;
  wire _14137_;
  wire _14138_;
  wire _14139_;
  wire _14140_;
  wire _14141_;
  wire _14142_;
  wire _14143_;
  wire _14144_;
  wire _14145_;
  wire _14146_;
  wire _14147_;
  wire _14148_;
  wire _14149_;
  wire _14150_;
  wire _14151_;
  wire _14152_;
  wire _14153_;
  wire _14154_;
  wire _14155_;
  wire _14156_;
  wire _14157_;
  wire _14158_;
  wire _14159_;
  wire _14160_;
  wire _14161_;
  wire _14162_;
  wire _14163_;
  wire _14164_;
  wire _14165_;
  wire _14166_;
  wire _14167_;
  wire _14168_;
  wire _14169_;
  wire _14170_;
  wire _14171_;
  wire _14172_;
  wire _14173_;
  wire _14174_;
  wire _14175_;
  wire _14176_;
  wire _14177_;
  wire _14178_;
  wire _14179_;
  wire _14180_;
  wire _14181_;
  wire _14182_;
  wire _14183_;
  wire _14184_;
  wire _14185_;
  wire _14186_;
  wire _14187_;
  wire _14188_;
  wire _14189_;
  wire _14190_;
  wire _14191_;
  wire _14192_;
  wire _14193_;
  wire _14194_;
  wire _14195_;
  wire _14196_;
  wire _14197_;
  wire _14198_;
  wire _14199_;
  wire _14200_;
  wire _14201_;
  wire _14202_;
  wire _14203_;
  wire _14204_;
  wire _14205_;
  wire _14206_;
  wire _14207_;
  wire _14208_;
  wire _14209_;
  wire _14210_;
  wire _14211_;
  wire _14212_;
  wire _14213_;
  wire _14214_;
  wire _14215_;
  wire _14216_;
  wire _14217_;
  wire _14218_;
  wire _14219_;
  wire _14220_;
  wire _14221_;
  wire _14222_;
  wire _14223_;
  wire _14224_;
  wire _14225_;
  wire _14226_;
  wire _14227_;
  wire _14228_;
  wire _14229_;
  wire _14230_;
  wire _14231_;
  wire _14232_;
  wire _14233_;
  wire _14234_;
  wire _14235_;
  wire _14236_;
  wire _14237_;
  wire _14238_;
  wire _14239_;
  wire _14240_;
  wire _14241_;
  wire _14242_;
  wire _14243_;
  wire _14244_;
  wire _14245_;
  wire _14246_;
  wire _14247_;
  wire _14248_;
  wire _14249_;
  wire _14250_;
  wire _14251_;
  wire _14252_;
  wire _14253_;
  wire _14254_;
  wire _14255_;
  wire _14256_;
  wire _14257_;
  wire _14258_;
  wire _14259_;
  wire _14260_;
  wire _14261_;
  wire _14262_;
  wire _14263_;
  wire _14264_;
  wire _14265_;
  wire _14266_;
  wire _14267_;
  wire _14268_;
  wire _14269_;
  wire _14270_;
  wire _14271_;
  wire _14272_;
  wire _14273_;
  wire _14274_;
  wire _14275_;
  wire _14276_;
  wire _14277_;
  wire _14278_;
  wire _14279_;
  wire _14280_;
  wire _14281_;
  wire _14282_;
  wire _14283_;
  wire _14284_;
  wire _14285_;
  wire _14286_;
  wire _14287_;
  wire _14288_;
  wire _14289_;
  wire _14290_;
  wire _14291_;
  wire _14292_;
  wire _14293_;
  wire _14294_;
  wire _14295_;
  wire _14296_;
  wire _14297_;
  wire _14298_;
  wire _14299_;
  wire _14300_;
  wire _14301_;
  wire _14302_;
  wire _14303_;
  wire _14304_;
  wire _14305_;
  wire _14306_;
  wire _14307_;
  wire _14308_;
  wire _14309_;
  wire _14310_;
  wire _14311_;
  wire _14312_;
  wire _14313_;
  wire _14314_;
  wire _14315_;
  wire _14316_;
  wire _14317_;
  wire _14318_;
  wire _14319_;
  wire _14320_;
  wire _14321_;
  wire _14322_;
  wire _14323_;
  wire _14324_;
  wire _14325_;
  wire _14326_;
  wire _14327_;
  wire _14328_;
  wire _14329_;
  wire _14330_;
  wire _14331_;
  wire _14332_;
  wire _14333_;
  wire _14334_;
  wire _14335_;
  wire _14336_;
  wire _14337_;
  wire _14338_;
  wire _14339_;
  wire _14340_;
  wire _14341_;
  wire _14342_;
  wire _14343_;
  wire _14344_;
  wire _14345_;
  wire _14346_;
  wire _14347_;
  wire _14348_;
  wire _14349_;
  wire _14350_;
  wire _14351_;
  wire _14352_;
  wire _14353_;
  wire _14354_;
  wire _14355_;
  wire _14356_;
  wire _14357_;
  wire _14358_;
  wire _14359_;
  wire _14360_;
  wire _14361_;
  wire _14362_;
  wire _14363_;
  wire _14364_;
  wire _14365_;
  wire _14366_;
  wire _14367_;
  wire _14368_;
  wire _14369_;
  wire _14370_;
  wire _14371_;
  wire _14372_;
  wire _14373_;
  wire _14374_;
  wire _14375_;
  wire _14376_;
  wire _14377_;
  wire _14378_;
  wire _14379_;
  wire _14380_;
  wire _14381_;
  wire _14382_;
  wire _14383_;
  wire _14384_;
  wire _14385_;
  wire _14386_;
  wire _14387_;
  wire _14388_;
  wire _14389_;
  wire _14390_;
  wire _14391_;
  wire _14392_;
  wire _14393_;
  wire _14394_;
  wire _14395_;
  wire _14396_;
  wire _14397_;
  wire _14398_;
  wire _14399_;
  wire _14400_;
  wire _14401_;
  wire _14402_;
  wire _14403_;
  wire _14404_;
  wire _14405_;
  wire _14406_;
  wire _14407_;
  wire _14408_;
  wire _14409_;
  wire _14410_;
  wire _14411_;
  wire _14412_;
  wire _14413_;
  wire _14414_;
  wire _14415_;
  wire _14416_;
  wire _14417_;
  wire _14418_;
  wire _14419_;
  wire _14420_;
  wire _14421_;
  wire _14422_;
  wire _14423_;
  wire _14424_;
  wire _14425_;
  wire _14426_;
  wire _14427_;
  wire _14428_;
  wire _14429_;
  wire _14430_;
  wire _14431_;
  wire _14432_;
  wire _14433_;
  wire _14434_;
  wire _14435_;
  wire _14436_;
  wire _14437_;
  wire _14438_;
  wire _14439_;
  wire _14440_;
  wire _14441_;
  wire _14442_;
  wire _14443_;
  wire _14444_;
  wire _14445_;
  wire _14446_;
  wire _14447_;
  wire _14448_;
  wire _14449_;
  wire _14450_;
  wire _14451_;
  wire _14452_;
  wire _14453_;
  wire _14454_;
  wire _14455_;
  wire _14456_;
  wire _14457_;
  wire _14458_;
  wire _14459_;
  wire _14460_;
  wire _14461_;
  wire _14462_;
  wire _14463_;
  wire _14464_;
  wire _14465_;
  wire _14466_;
  wire _14467_;
  wire _14468_;
  wire _14469_;
  wire _14470_;
  wire _14471_;
  wire _14472_;
  wire _14473_;
  wire _14474_;
  wire _14475_;
  wire _14476_;
  wire _14477_;
  wire _14478_;
  wire _14479_;
  wire _14480_;
  wire _14481_;
  wire _14482_;
  wire _14483_;
  wire _14484_;
  wire _14485_;
  wire _14486_;
  wire _14487_;
  wire _14488_;
  wire _14489_;
  wire _14490_;
  wire _14491_;
  wire _14492_;
  wire _14493_;
  wire _14494_;
  wire _14495_;
  wire _14496_;
  wire _14497_;
  wire _14498_;
  wire _14499_;
  wire _14500_;
  wire _14501_;
  wire _14502_;
  wire _14503_;
  wire _14504_;
  wire _14505_;
  wire _14506_;
  wire _14507_;
  wire _14508_;
  wire _14509_;
  wire _14510_;
  wire _14511_;
  wire _14512_;
  wire _14513_;
  wire _14514_;
  wire _14515_;
  wire _14516_;
  wire _14517_;
  wire _14518_;
  wire _14519_;
  wire _14520_;
  wire _14521_;
  wire _14522_;
  wire _14523_;
  wire _14524_;
  wire _14525_;
  wire _14526_;
  wire _14527_;
  wire _14528_;
  wire _14529_;
  wire _14530_;
  wire _14531_;
  wire _14532_;
  wire _14533_;
  wire _14534_;
  wire _14535_;
  wire _14536_;
  wire _14537_;
  wire _14538_;
  wire _14539_;
  wire _14540_;
  wire _14541_;
  wire _14542_;
  wire _14543_;
  wire _14544_;
  wire _14545_;
  wire _14546_;
  wire _14547_;
  wire _14548_;
  wire _14549_;
  wire _14550_;
  wire _14551_;
  wire _14552_;
  wire _14553_;
  wire _14554_;
  wire _14555_;
  wire _14556_;
  wire _14557_;
  wire _14558_;
  wire _14559_;
  wire _14560_;
  wire _14561_;
  wire _14562_;
  wire _14563_;
  wire _14564_;
  wire _14565_;
  wire _14566_;
  wire _14567_;
  wire _14568_;
  wire _14569_;
  wire _14570_;
  wire _14571_;
  wire _14572_;
  wire _14573_;
  wire _14574_;
  wire _14575_;
  wire _14576_;
  wire _14577_;
  wire _14578_;
  wire _14579_;
  wire _14580_;
  wire _14581_;
  wire _14582_;
  wire _14583_;
  wire _14584_;
  wire _14585_;
  wire _14586_;
  wire _14587_;
  wire _14588_;
  wire _14589_;
  wire _14590_;
  wire _14591_;
  wire _14592_;
  wire _14593_;
  wire _14594_;
  wire _14595_;
  wire _14596_;
  wire _14597_;
  wire _14598_;
  wire _14599_;
  wire _14600_;
  wire _14601_;
  wire _14602_;
  wire _14603_;
  wire _14604_;
  wire _14605_;
  wire _14606_;
  wire _14607_;
  wire _14608_;
  wire _14609_;
  wire _14610_;
  wire _14611_;
  wire _14612_;
  wire _14613_;
  wire _14614_;
  wire _14615_;
  wire _14616_;
  wire _14617_;
  wire _14618_;
  wire _14619_;
  wire _14620_;
  wire _14621_;
  wire _14622_;
  wire _14623_;
  wire _14624_;
  wire _14625_;
  wire _14626_;
  wire _14627_;
  wire _14628_;
  wire _14629_;
  wire _14630_;
  wire _14631_;
  wire _14632_;
  wire _14633_;
  wire _14634_;
  wire _14635_;
  wire _14636_;
  wire _14637_;
  wire _14638_;
  wire _14639_;
  wire _14640_;
  wire _14641_;
  wire _14642_;
  wire _14643_;
  wire _14644_;
  wire _14645_;
  wire _14646_;
  wire _14647_;
  wire _14648_;
  wire _14649_;
  wire _14650_;
  wire _14651_;
  wire _14652_;
  wire _14653_;
  wire _14654_;
  wire _14655_;
  wire _14656_;
  wire _14657_;
  wire _14658_;
  wire _14659_;
  wire _14660_;
  wire _14661_;
  wire _14662_;
  wire _14663_;
  wire _14664_;
  wire _14665_;
  wire _14666_;
  wire _14667_;
  wire _14668_;
  wire _14669_;
  wire _14670_;
  wire _14671_;
  wire _14672_;
  wire _14673_;
  wire _14674_;
  wire _14675_;
  wire _14676_;
  wire _14677_;
  wire _14678_;
  wire _14679_;
  wire _14680_;
  wire _14681_;
  wire _14682_;
  wire _14683_;
  wire _14684_;
  wire _14685_;
  wire _14686_;
  wire _14687_;
  wire _14688_;
  wire _14689_;
  wire _14690_;
  wire _14691_;
  wire _14692_;
  wire _14693_;
  wire _14694_;
  wire _14695_;
  wire _14696_;
  wire _14697_;
  wire _14698_;
  wire _14699_;
  wire _14700_;
  wire _14701_;
  wire _14702_;
  wire _14703_;
  wire _14704_;
  wire _14705_;
  wire _14706_;
  wire _14707_;
  wire _14708_;
  wire _14709_;
  wire _14710_;
  wire _14711_;
  wire _14712_;
  wire _14713_;
  wire _14714_;
  wire _14715_;
  wire _14716_;
  wire _14717_;
  wire _14718_;
  wire _14719_;
  wire _14720_;
  wire _14721_;
  wire _14722_;
  wire _14723_;
  wire _14724_;
  wire _14725_;
  wire _14726_;
  wire _14727_;
  wire _14728_;
  wire _14729_;
  wire _14730_;
  wire _14731_;
  wire _14732_;
  wire _14733_;
  wire _14734_;
  wire _14735_;
  wire _14736_;
  wire _14737_;
  wire _14738_;
  wire _14739_;
  wire _14740_;
  wire _14741_;
  wire _14742_;
  wire _14743_;
  wire _14744_;
  wire _14745_;
  wire _14746_;
  wire _14747_;
  wire _14748_;
  wire _14749_;
  wire _14750_;
  wire _14751_;
  wire _14752_;
  wire _14753_;
  wire _14754_;
  wire _14755_;
  wire _14756_;
  wire _14757_;
  wire _14758_;
  wire _14759_;
  wire _14760_;
  wire _14761_;
  wire _14762_;
  wire _14763_;
  wire _14764_;
  wire _14765_;
  wire _14766_;
  wire _14767_;
  wire _14768_;
  wire _14769_;
  wire _14770_;
  wire _14771_;
  wire _14772_;
  wire _14773_;
  wire _14774_;
  wire _14775_;
  wire _14776_;
  wire _14777_;
  wire _14778_;
  wire _14779_;
  wire _14780_;
  wire _14781_;
  wire _14782_;
  wire _14783_;
  wire _14784_;
  wire _14785_;
  wire _14786_;
  wire _14787_;
  wire _14788_;
  wire _14789_;
  wire _14790_;
  wire _14791_;
  wire _14792_;
  wire _14793_;
  wire _14794_;
  wire _14795_;
  wire _14796_;
  wire _14797_;
  wire _14798_;
  wire _14799_;
  wire _14800_;
  wire _14801_;
  wire _14802_;
  wire _14803_;
  wire _14804_;
  wire _14805_;
  wire _14806_;
  wire _14807_;
  wire _14808_;
  wire _14809_;
  wire _14810_;
  wire _14811_;
  wire _14812_;
  wire _14813_;
  wire _14814_;
  wire _14815_;
  wire _14816_;
  wire _14817_;
  wire _14818_;
  wire _14819_;
  wire _14820_;
  wire _14821_;
  wire _14822_;
  wire _14823_;
  wire _14824_;
  wire _14825_;
  wire _14826_;
  wire _14827_;
  wire _14828_;
  wire _14829_;
  wire _14830_;
  wire _14831_;
  wire _14832_;
  wire _14833_;
  wire _14834_;
  wire _14835_;
  wire _14836_;
  wire _14837_;
  wire _14838_;
  wire _14839_;
  wire _14840_;
  wire _14841_;
  wire _14842_;
  wire _14843_;
  wire _14844_;
  wire _14845_;
  wire _14846_;
  wire _14847_;
  wire _14848_;
  wire _14849_;
  wire _14850_;
  wire _14851_;
  wire _14852_;
  wire _14853_;
  wire _14854_;
  wire _14855_;
  wire _14856_;
  wire _14857_;
  wire _14858_;
  wire _14859_;
  wire _14860_;
  wire _14861_;
  wire _14862_;
  wire _14863_;
  wire _14864_;
  wire _14865_;
  wire _14866_;
  wire _14867_;
  wire _14868_;
  wire _14869_;
  wire _14870_;
  wire _14871_;
  wire _14872_;
  wire _14873_;
  wire _14874_;
  wire _14875_;
  wire _14876_;
  wire _14877_;
  wire _14878_;
  wire _14879_;
  wire _14880_;
  wire _14881_;
  wire _14882_;
  wire _14883_;
  wire _14884_;
  wire _14885_;
  wire _14886_;
  wire _14887_;
  wire _14888_;
  wire _14889_;
  wire _14890_;
  wire _14891_;
  wire _14892_;
  wire _14893_;
  wire _14894_;
  wire _14895_;
  wire _14896_;
  wire _14897_;
  wire _14898_;
  wire _14899_;
  wire _14900_;
  wire _14901_;
  wire _14902_;
  wire _14903_;
  wire _14904_;
  wire _14905_;
  wire _14906_;
  wire _14907_;
  wire _14908_;
  wire _14909_;
  wire _14910_;
  wire _14911_;
  wire _14912_;
  wire _14913_;
  wire _14914_;
  wire _14915_;
  wire _14916_;
  wire _14917_;
  wire _14918_;
  wire _14919_;
  wire _14920_;
  wire _14921_;
  wire _14922_;
  wire _14923_;
  wire _14924_;
  wire _14925_;
  wire _14926_;
  wire _14927_;
  wire _14928_;
  wire _14929_;
  wire _14930_;
  wire _14931_;
  wire _14932_;
  wire _14933_;
  wire _14934_;
  wire _14935_;
  wire _14936_;
  wire _14937_;
  wire _14938_;
  wire _14939_;
  wire _14940_;
  wire _14941_;
  wire _14942_;
  wire _14943_;
  wire _14944_;
  wire _14945_;
  wire _14946_;
  wire _14947_;
  wire _14948_;
  wire _14949_;
  wire _14950_;
  wire _14951_;
  wire _14952_;
  wire _14953_;
  wire _14954_;
  wire _14955_;
  wire _14956_;
  wire _14957_;
  wire _14958_;
  wire _14959_;
  wire _14960_;
  wire _14961_;
  wire _14962_;
  wire _14963_;
  wire _14964_;
  wire _14965_;
  wire _14966_;
  wire _14967_;
  wire _14968_;
  wire _14969_;
  wire _14970_;
  wire _14971_;
  wire _14972_;
  wire _14973_;
  wire _14974_;
  wire _14975_;
  wire _14976_;
  wire _14977_;
  wire _14978_;
  wire _14979_;
  wire _14980_;
  wire _14981_;
  wire _14982_;
  wire _14983_;
  wire _14984_;
  wire _14985_;
  wire _14986_;
  wire _14987_;
  wire _14988_;
  wire _14989_;
  wire _14990_;
  wire _14991_;
  wire _14992_;
  wire _14993_;
  wire _14994_;
  wire _14995_;
  wire _14996_;
  wire _14997_;
  wire _14998_;
  wire _14999_;
  wire _15000_;
  wire _15001_;
  wire _15002_;
  wire _15003_;
  wire _15004_;
  wire _15005_;
  wire _15006_;
  wire _15007_;
  wire _15008_;
  wire _15009_;
  wire _15010_;
  wire _15011_;
  wire _15012_;
  wire _15013_;
  wire _15014_;
  wire _15015_;
  wire _15016_;
  wire _15017_;
  wire _15018_;
  wire _15019_;
  wire _15020_;
  wire _15021_;
  wire _15022_;
  wire _15023_;
  wire _15024_;
  wire _15025_;
  wire _15026_;
  wire _15027_;
  wire _15028_;
  wire _15029_;
  wire _15030_;
  wire _15031_;
  wire _15032_;
  wire _15033_;
  wire _15034_;
  wire _15035_;
  wire _15036_;
  wire _15037_;
  wire _15038_;
  wire _15039_;
  wire _15040_;
  wire _15041_;
  wire _15042_;
  wire _15043_;
  wire _15044_;
  wire _15045_;
  wire _15046_;
  wire _15047_;
  wire _15048_;
  wire _15049_;
  wire _15050_;
  wire _15051_;
  wire _15052_;
  wire _15053_;
  wire _15054_;
  wire _15055_;
  wire _15056_;
  wire _15057_;
  wire _15058_;
  wire _15059_;
  wire _15060_;
  wire _15061_;
  wire _15062_;
  wire _15063_;
  wire _15064_;
  wire _15065_;
  wire _15066_;
  wire _15067_;
  wire _15068_;
  wire _15069_;
  wire _15070_;
  wire _15071_;
  wire _15072_;
  wire _15073_;
  wire _15074_;
  wire _15075_;
  wire _15076_;
  wire _15077_;
  wire _15078_;
  wire _15079_;
  wire _15080_;
  wire _15081_;
  wire _15082_;
  wire _15083_;
  wire _15084_;
  wire _15085_;
  wire _15086_;
  wire _15087_;
  wire _15088_;
  wire _15089_;
  wire _15090_;
  wire _15091_;
  wire _15092_;
  wire _15093_;
  wire _15094_;
  wire _15095_;
  wire _15096_;
  wire _15097_;
  wire _15098_;
  wire _15099_;
  wire _15100_;
  wire _15101_;
  wire _15102_;
  wire _15103_;
  wire _15104_;
  wire _15105_;
  wire _15106_;
  wire _15107_;
  wire _15108_;
  wire _15109_;
  wire _15110_;
  wire _15111_;
  wire _15112_;
  wire _15113_;
  wire _15114_;
  wire _15115_;
  wire _15116_;
  wire _15117_;
  wire _15118_;
  wire _15119_;
  wire _15120_;
  wire _15121_;
  wire _15122_;
  wire _15123_;
  wire _15124_;
  wire _15125_;
  wire _15126_;
  wire _15127_;
  wire _15128_;
  wire _15129_;
  wire _15130_;
  wire _15131_;
  wire _15132_;
  wire _15133_;
  wire _15134_;
  wire _15135_;
  wire _15136_;
  wire _15137_;
  wire _15138_;
  wire _15139_;
  wire _15140_;
  wire _15141_;
  wire _15142_;
  wire _15143_;
  wire _15144_;
  wire _15145_;
  wire _15146_;
  wire _15147_;
  wire _15148_;
  wire _15149_;
  wire _15150_;
  wire _15151_;
  wire _15152_;
  wire _15153_;
  wire _15154_;
  wire _15155_;
  wire _15156_;
  wire _15157_;
  wire _15158_;
  wire _15159_;
  wire _15160_;
  wire _15161_;
  wire _15162_;
  wire _15163_;
  wire _15164_;
  wire _15165_;
  wire _15166_;
  wire _15167_;
  wire _15168_;
  wire _15169_;
  wire _15170_;
  wire _15171_;
  wire _15172_;
  wire _15173_;
  wire _15174_;
  wire _15175_;
  wire _15176_;
  wire _15177_;
  wire _15178_;
  wire _15179_;
  wire _15180_;
  wire _15181_;
  wire _15182_;
  wire _15183_;
  wire _15184_;
  wire _15185_;
  wire _15186_;
  wire _15187_;
  wire _15188_;
  wire _15189_;
  wire _15190_;
  wire _15191_;
  wire _15192_;
  wire _15193_;
  wire _15194_;
  wire _15195_;
  wire _15196_;
  wire _15197_;
  wire _15198_;
  wire _15199_;
  wire _15200_;
  wire _15201_;
  wire _15202_;
  wire _15203_;
  wire _15204_;
  wire _15205_;
  wire _15206_;
  wire _15207_;
  wire _15208_;
  wire _15209_;
  wire _15210_;
  wire _15211_;
  wire _15212_;
  wire _15213_;
  wire _15214_;
  wire _15215_;
  wire _15216_;
  wire _15217_;
  wire _15218_;
  wire _15219_;
  wire _15220_;
  wire _15221_;
  wire _15222_;
  wire _15223_;
  wire _15224_;
  wire _15225_;
  wire _15226_;
  wire _15227_;
  wire _15228_;
  wire _15229_;
  wire _15230_;
  wire _15231_;
  wire _15232_;
  wire _15233_;
  wire _15234_;
  wire _15235_;
  wire _15236_;
  wire _15237_;
  wire _15238_;
  wire _15239_;
  wire _15240_;
  wire _15241_;
  wire _15242_;
  wire _15243_;
  wire _15244_;
  wire _15245_;
  wire _15246_;
  wire _15247_;
  wire _15248_;
  wire _15249_;
  wire _15250_;
  wire _15251_;
  wire _15252_;
  wire _15253_;
  wire _15254_;
  wire _15255_;
  wire _15256_;
  wire _15257_;
  wire _15258_;
  wire _15259_;
  wire _15260_;
  wire _15261_;
  wire _15262_;
  wire _15263_;
  wire _15264_;
  wire _15265_;
  wire _15266_;
  wire _15267_;
  wire _15268_;
  wire _15269_;
  wire _15270_;
  wire _15271_;
  wire _15272_;
  wire _15273_;
  wire _15274_;
  wire _15275_;
  wire _15276_;
  wire _15277_;
  wire _15278_;
  wire _15279_;
  wire _15280_;
  wire _15281_;
  wire _15282_;
  wire _15283_;
  wire _15284_;
  wire _15285_;
  wire _15286_;
  wire _15287_;
  wire _15288_;
  wire _15289_;
  wire _15290_;
  wire _15291_;
  wire _15292_;
  wire _15293_;
  wire _15294_;
  wire _15295_;
  wire _15296_;
  wire _15297_;
  wire _15298_;
  wire _15299_;
  wire _15300_;
  wire _15301_;
  wire _15302_;
  wire _15303_;
  wire _15304_;
  wire _15305_;
  wire _15306_;
  wire _15307_;
  wire _15308_;
  wire _15309_;
  wire _15310_;
  wire _15311_;
  wire _15312_;
  wire _15313_;
  wire _15314_;
  wire _15315_;
  wire _15316_;
  wire _15317_;
  wire _15318_;
  wire _15319_;
  wire _15320_;
  wire _15321_;
  wire _15322_;
  wire _15323_;
  wire _15324_;
  wire _15325_;
  wire _15326_;
  wire _15327_;
  wire _15328_;
  wire _15329_;
  wire _15330_;
  wire _15331_;
  wire _15332_;
  wire _15333_;
  wire _15334_;
  wire _15335_;
  wire _15336_;
  wire _15337_;
  wire _15338_;
  wire _15339_;
  wire _15340_;
  wire _15341_;
  wire _15342_;
  wire _15343_;
  wire _15344_;
  wire _15345_;
  wire _15346_;
  wire _15347_;
  wire _15348_;
  wire _15349_;
  wire _15350_;
  wire _15351_;
  wire _15352_;
  wire _15353_;
  wire _15354_;
  wire _15355_;
  wire _15356_;
  wire _15357_;
  wire _15358_;
  wire _15359_;
  wire _15360_;
  wire _15361_;
  wire _15362_;
  wire _15363_;
  wire _15364_;
  wire _15365_;
  wire _15366_;
  wire _15367_;
  wire _15368_;
  wire _15369_;
  wire _15370_;
  wire _15371_;
  wire _15372_;
  wire _15373_;
  wire _15374_;
  wire _15375_;
  wire _15376_;
  wire _15377_;
  wire _15378_;
  wire _15379_;
  wire _15380_;
  wire _15381_;
  wire _15382_;
  wire _15383_;
  wire _15384_;
  wire _15385_;
  wire _15386_;
  wire _15387_;
  wire _15388_;
  wire _15389_;
  wire _15390_;
  wire _15391_;
  wire _15392_;
  wire _15393_;
  wire _15394_;
  wire _15395_;
  wire _15396_;
  wire _15397_;
  wire _15398_;
  wire _15399_;
  wire _15400_;
  wire _15401_;
  wire _15402_;
  wire _15403_;
  wire _15404_;
  wire _15405_;
  wire _15406_;
  wire _15407_;
  wire _15408_;
  wire _15409_;
  wire _15410_;
  wire _15411_;
  wire _15412_;
  wire _15413_;
  wire _15414_;
  wire _15415_;
  wire _15416_;
  wire _15417_;
  wire _15418_;
  wire _15419_;
  wire _15420_;
  wire _15421_;
  wire _15422_;
  wire _15423_;
  wire _15424_;
  wire _15425_;
  wire _15426_;
  wire _15427_;
  wire _15428_;
  wire _15429_;
  wire _15430_;
  wire _15431_;
  wire _15432_;
  wire _15433_;
  wire _15434_;
  wire _15435_;
  wire _15436_;
  wire _15437_;
  wire _15438_;
  wire _15439_;
  wire _15440_;
  wire _15441_;
  wire _15442_;
  wire _15443_;
  wire _15444_;
  wire _15445_;
  wire _15446_;
  wire _15447_;
  wire _15448_;
  wire _15449_;
  wire _15450_;
  wire _15451_;
  wire _15452_;
  wire _15453_;
  wire _15454_;
  wire _15455_;
  wire _15456_;
  wire _15457_;
  wire _15458_;
  wire _15459_;
  wire _15460_;
  wire _15461_;
  wire _15462_;
  wire _15463_;
  wire _15464_;
  wire _15465_;
  wire _15466_;
  wire _15467_;
  wire _15468_;
  wire _15469_;
  wire _15470_;
  wire _15471_;
  wire _15472_;
  wire _15473_;
  wire _15474_;
  wire _15475_;
  wire _15476_;
  wire _15477_;
  wire _15478_;
  wire _15479_;
  wire _15480_;
  wire _15481_;
  wire _15482_;
  wire _15483_;
  wire _15484_;
  wire _15485_;
  wire _15486_;
  wire _15487_;
  wire _15488_;
  wire _15489_;
  wire _15490_;
  wire _15491_;
  wire _15492_;
  wire _15493_;
  wire _15494_;
  wire _15495_;
  wire _15496_;
  wire _15497_;
  wire _15498_;
  wire _15499_;
  wire _15500_;
  wire _15501_;
  wire _15502_;
  wire _15503_;
  wire _15504_;
  wire _15505_;
  wire _15506_;
  wire _15507_;
  wire _15508_;
  wire _15509_;
  wire _15510_;
  wire _15511_;
  wire _15512_;
  wire _15513_;
  wire _15514_;
  wire _15515_;
  wire _15516_;
  wire _15517_;
  wire _15518_;
  wire _15519_;
  wire _15520_;
  wire _15521_;
  wire _15522_;
  wire _15523_;
  wire _15524_;
  wire _15525_;
  wire _15526_;
  wire _15527_;
  wire _15528_;
  wire _15529_;
  wire _15530_;
  wire _15531_;
  wire _15532_;
  wire _15533_;
  wire _15534_;
  wire _15535_;
  wire _15536_;
  wire _15537_;
  wire _15538_;
  wire _15539_;
  wire _15540_;
  wire _15541_;
  wire _15542_;
  wire _15543_;
  wire _15544_;
  wire _15545_;
  wire _15546_;
  wire _15547_;
  wire _15548_;
  wire _15549_;
  wire _15550_;
  wire _15551_;
  wire _15552_;
  wire _15553_;
  wire _15554_;
  wire _15555_;
  wire _15556_;
  wire _15557_;
  wire _15558_;
  wire _15559_;
  wire _15560_;
  wire _15561_;
  wire _15562_;
  wire _15563_;
  wire _15564_;
  wire _15565_;
  wire _15566_;
  wire _15567_;
  wire _15568_;
  wire _15569_;
  wire _15570_;
  wire _15571_;
  wire _15572_;
  wire _15573_;
  wire _15574_;
  wire _15575_;
  wire _15576_;
  wire _15577_;
  wire _15578_;
  wire _15579_;
  wire _15580_;
  wire _15581_;
  wire _15582_;
  wire _15583_;
  wire _15584_;
  wire _15585_;
  wire _15586_;
  wire _15587_;
  wire _15588_;
  wire _15589_;
  wire _15590_;
  wire _15591_;
  wire _15592_;
  wire _15593_;
  wire _15594_;
  wire _15595_;
  wire _15596_;
  wire _15597_;
  wire _15598_;
  wire _15599_;
  wire _15600_;
  wire _15601_;
  wire _15602_;
  wire _15603_;
  wire _15604_;
  wire _15605_;
  wire _15606_;
  wire _15607_;
  wire _15608_;
  wire _15609_;
  wire _15610_;
  wire _15611_;
  wire _15612_;
  wire _15613_;
  wire _15614_;
  wire _15615_;
  wire _15616_;
  wire _15617_;
  wire _15618_;
  wire _15619_;
  wire _15620_;
  wire _15621_;
  wire _15622_;
  wire _15623_;
  wire _15624_;
  wire _15625_;
  wire _15626_;
  wire _15627_;
  wire _15628_;
  wire _15629_;
  wire _15630_;
  wire _15631_;
  wire _15632_;
  wire _15633_;
  wire _15634_;
  wire _15635_;
  wire _15636_;
  wire _15637_;
  wire _15638_;
  wire _15639_;
  wire _15640_;
  wire _15641_;
  wire _15642_;
  wire _15643_;
  wire _15644_;
  wire _15645_;
  wire _15646_;
  wire _15647_;
  wire _15648_;
  wire _15649_;
  wire _15650_;
  wire _15651_;
  wire _15652_;
  wire _15653_;
  wire _15654_;
  wire _15655_;
  wire _15656_;
  wire _15657_;
  wire _15658_;
  wire _15659_;
  wire _15660_;
  wire _15661_;
  wire _15662_;
  wire _15663_;
  wire _15664_;
  wire _15665_;
  wire _15666_;
  wire _15667_;
  wire _15668_;
  wire _15669_;
  wire _15670_;
  wire _15671_;
  wire _15672_;
  wire _15673_;
  wire _15674_;
  wire _15675_;
  wire _15676_;
  wire _15677_;
  wire _15678_;
  wire _15679_;
  wire _15680_;
  wire _15681_;
  wire _15682_;
  wire _15683_;
  wire _15684_;
  wire _15685_;
  wire _15686_;
  wire _15687_;
  wire _15688_;
  wire _15689_;
  wire _15690_;
  wire _15691_;
  wire _15692_;
  wire _15693_;
  wire _15694_;
  wire _15695_;
  wire _15696_;
  wire _15697_;
  wire _15698_;
  wire _15699_;
  wire _15700_;
  wire _15701_;
  wire _15702_;
  wire _15703_;
  wire _15704_;
  wire _15705_;
  wire _15706_;
  wire _15707_;
  wire _15708_;
  wire _15709_;
  wire _15710_;
  wire _15711_;
  wire _15712_;
  wire _15713_;
  wire _15714_;
  wire _15715_;
  wire _15716_;
  wire _15717_;
  wire _15718_;
  wire _15719_;
  wire _15720_;
  wire _15721_;
  wire _15722_;
  wire _15723_;
  wire _15724_;
  wire _15725_;
  wire _15726_;
  wire _15727_;
  wire _15728_;
  wire _15729_;
  wire _15730_;
  wire _15731_;
  wire _15732_;
  wire _15733_;
  wire _15734_;
  wire _15735_;
  wire _15736_;
  wire _15737_;
  wire _15738_;
  wire _15739_;
  wire _15740_;
  wire _15741_;
  wire _15742_;
  wire _15743_;
  wire _15744_;
  wire _15745_;
  wire _15746_;
  wire _15747_;
  wire _15748_;
  wire _15749_;
  wire _15750_;
  wire _15751_;
  wire _15752_;
  wire _15753_;
  wire _15754_;
  wire _15755_;
  wire _15756_;
  wire _15757_;
  wire _15758_;
  wire _15759_;
  wire _15760_;
  wire _15761_;
  wire _15762_;
  wire _15763_;
  wire _15764_;
  wire _15765_;
  wire _15766_;
  wire _15767_;
  wire _15768_;
  wire _15769_;
  wire _15770_;
  wire _15771_;
  wire _15772_;
  wire _15773_;
  wire _15774_;
  wire _15775_;
  wire _15776_;
  wire _15777_;
  wire _15778_;
  wire _15779_;
  wire _15780_;
  wire _15781_;
  wire _15782_;
  wire _15783_;
  wire _15784_;
  wire _15785_;
  wire _15786_;
  wire _15787_;
  wire _15788_;
  wire _15789_;
  wire _15790_;
  wire _15791_;
  wire _15792_;
  wire _15793_;
  wire _15794_;
  wire _15795_;
  wire _15796_;
  wire _15797_;
  wire _15798_;
  wire _15799_;
  wire _15800_;
  wire _15801_;
  wire _15802_;
  wire _15803_;
  wire _15804_;
  wire _15805_;
  wire _15806_;
  wire _15807_;
  wire _15808_;
  wire _15809_;
  wire _15810_;
  wire _15811_;
  wire _15812_;
  wire _15813_;
  wire _15814_;
  wire _15815_;
  wire _15816_;
  wire _15817_;
  wire _15818_;
  wire _15819_;
  wire _15820_;
  wire _15821_;
  wire _15822_;
  wire _15823_;
  wire _15824_;
  wire _15825_;
  wire _15826_;
  wire _15827_;
  wire _15828_;
  wire _15829_;
  wire _15830_;
  wire _15831_;
  wire _15832_;
  wire _15833_;
  wire _15834_;
  wire _15835_;
  wire _15836_;
  wire _15837_;
  wire _15838_;
  wire _15839_;
  wire _15840_;
  wire _15841_;
  wire _15842_;
  wire _15843_;
  wire _15844_;
  wire _15845_;
  wire _15846_;
  wire _15847_;
  wire _15848_;
  wire _15849_;
  wire _15850_;
  wire _15851_;
  wire _15852_;
  wire _15853_;
  wire _15854_;
  wire _15855_;
  wire _15856_;
  wire _15857_;
  wire _15858_;
  wire _15859_;
  wire _15860_;
  wire _15861_;
  wire _15862_;
  wire _15863_;
  wire _15864_;
  wire _15865_;
  wire _15866_;
  wire _15867_;
  wire _15868_;
  wire _15869_;
  wire _15870_;
  wire _15871_;
  wire _15872_;
  wire _15873_;
  wire _15874_;
  wire _15875_;
  wire _15876_;
  wire _15877_;
  wire _15878_;
  wire _15879_;
  wire _15880_;
  wire _15881_;
  wire _15882_;
  wire _15883_;
  wire _15884_;
  wire _15885_;
  wire _15886_;
  wire _15887_;
  wire _15888_;
  wire _15889_;
  wire _15890_;
  wire _15891_;
  wire _15892_;
  wire _15893_;
  wire _15894_;
  wire _15895_;
  wire _15896_;
  wire _15897_;
  wire _15898_;
  wire _15899_;
  wire _15900_;
  wire _15901_;
  wire _15902_;
  wire _15903_;
  wire _15904_;
  wire _15905_;
  wire _15906_;
  wire _15907_;
  wire _15908_;
  wire _15909_;
  wire _15910_;
  wire _15911_;
  wire _15912_;
  wire _15913_;
  wire _15914_;
  wire _15915_;
  wire _15916_;
  wire _15917_;
  wire _15918_;
  wire _15919_;
  wire _15920_;
  wire _15921_;
  wire _15922_;
  wire _15923_;
  wire _15924_;
  wire _15925_;
  wire _15926_;
  wire _15927_;
  wire _15928_;
  wire _15929_;
  wire _15930_;
  wire _15931_;
  wire _15932_;
  wire _15933_;
  wire _15934_;
  wire _15935_;
  wire _15936_;
  wire _15937_;
  wire _15938_;
  wire _15939_;
  wire _15940_;
  wire _15941_;
  wire _15942_;
  wire _15943_;
  wire _15944_;
  wire _15945_;
  wire _15946_;
  wire _15947_;
  wire _15948_;
  wire _15949_;
  wire _15950_;
  wire _15951_;
  wire _15952_;
  wire _15953_;
  wire _15954_;
  wire _15955_;
  wire _15956_;
  wire _15957_;
  wire _15958_;
  wire _15959_;
  wire _15960_;
  wire _15961_;
  wire _15962_;
  wire _15963_;
  wire _15964_;
  wire _15965_;
  wire _15966_;
  wire _15967_;
  wire _15968_;
  wire _15969_;
  wire _15970_;
  wire _15971_;
  wire _15972_;
  wire _15973_;
  wire _15974_;
  wire _15975_;
  wire _15976_;
  wire _15977_;
  wire _15978_;
  wire _15979_;
  wire _15980_;
  wire _15981_;
  wire _15982_;
  wire _15983_;
  wire _15984_;
  wire _15985_;
  wire _15986_;
  wire _15987_;
  wire _15988_;
  wire _15989_;
  wire _15990_;
  wire _15991_;
  wire _15992_;
  wire _15993_;
  wire _15994_;
  wire _15995_;
  wire _15996_;
  wire _15997_;
  wire _15998_;
  wire _15999_;
  wire _16000_;
  wire _16001_;
  wire _16002_;
  wire _16003_;
  wire _16004_;
  wire _16005_;
  wire _16006_;
  wire _16007_;
  wire _16008_;
  wire _16009_;
  wire _16010_;
  wire _16011_;
  wire _16012_;
  wire _16013_;
  wire _16014_;
  wire _16015_;
  wire _16016_;
  wire _16017_;
  wire _16018_;
  wire _16019_;
  wire _16020_;
  wire _16021_;
  wire _16022_;
  wire _16023_;
  wire _16024_;
  wire _16025_;
  wire _16026_;
  wire _16027_;
  wire _16028_;
  wire _16029_;
  wire _16030_;
  wire _16031_;
  wire _16032_;
  wire _16033_;
  wire _16034_;
  wire _16035_;
  wire _16036_;
  wire _16037_;
  wire _16038_;
  wire _16039_;
  wire _16040_;
  wire _16041_;
  wire _16042_;
  wire _16043_;
  wire _16044_;
  wire _16045_;
  wire _16046_;
  wire _16047_;
  wire _16048_;
  wire _16049_;
  wire _16050_;
  wire _16051_;
  wire _16052_;
  wire _16053_;
  wire _16054_;
  wire _16055_;
  wire _16056_;
  wire _16057_;
  wire _16058_;
  wire _16059_;
  wire _16060_;
  wire _16061_;
  wire _16062_;
  wire _16063_;
  wire _16064_;
  wire _16065_;
  wire _16066_;
  wire _16067_;
  wire _16068_;
  wire _16069_;
  wire _16070_;
  wire _16071_;
  wire _16072_;
  wire _16073_;
  wire _16074_;
  wire _16075_;
  wire _16076_;
  wire _16077_;
  wire _16078_;
  wire _16079_;
  wire _16080_;
  wire _16081_;
  wire _16082_;
  wire _16083_;
  wire _16084_;
  wire _16085_;
  wire _16086_;
  wire _16087_;
  wire _16088_;
  wire _16089_;
  wire _16090_;
  wire _16091_;
  wire _16092_;
  wire _16093_;
  wire _16094_;
  wire _16095_;
  wire _16096_;
  wire _16097_;
  wire _16098_;
  wire _16099_;
  wire _16100_;
  wire _16101_;
  wire _16102_;
  wire _16103_;
  wire _16104_;
  wire _16105_;
  wire _16106_;
  wire _16107_;
  wire _16108_;
  wire _16109_;
  wire _16110_;
  wire _16111_;
  wire _16112_;
  wire _16113_;
  wire _16114_;
  wire _16115_;
  wire _16116_;
  wire _16117_;
  wire _16118_;
  wire _16119_;
  wire _16120_;
  wire _16121_;
  wire _16122_;
  wire _16123_;
  wire _16124_;
  wire _16125_;
  wire _16126_;
  wire _16127_;
  wire _16128_;
  wire _16129_;
  wire _16130_;
  wire _16131_;
  wire _16132_;
  wire _16133_;
  wire _16134_;
  wire _16135_;
  wire _16136_;
  wire _16137_;
  wire _16138_;
  wire _16139_;
  wire _16140_;
  wire _16141_;
  wire _16142_;
  wire _16143_;
  wire _16144_;
  wire _16145_;
  wire _16146_;
  wire _16147_;
  wire _16148_;
  wire _16149_;
  wire _16150_;
  wire _16151_;
  wire _16152_;
  wire _16153_;
  wire _16154_;
  wire _16155_;
  wire _16156_;
  wire _16157_;
  wire _16158_;
  wire _16159_;
  wire _16160_;
  wire _16161_;
  wire _16162_;
  wire _16163_;
  wire _16164_;
  wire _16165_;
  wire _16166_;
  wire _16167_;
  wire _16168_;
  wire _16169_;
  wire _16170_;
  wire _16171_;
  wire _16172_;
  wire _16173_;
  wire _16174_;
  wire _16175_;
  wire _16176_;
  wire _16177_;
  wire _16178_;
  wire _16179_;
  wire _16180_;
  wire _16181_;
  wire _16182_;
  wire _16183_;
  wire _16184_;
  wire _16185_;
  wire _16186_;
  wire _16187_;
  wire _16188_;
  wire _16189_;
  wire _16190_;
  wire _16191_;
  wire _16192_;
  wire _16193_;
  wire _16194_;
  wire _16195_;
  wire _16196_;
  wire _16197_;
  wire _16198_;
  wire _16199_;
  wire _16200_;
  wire _16201_;
  wire _16202_;
  wire _16203_;
  wire _16204_;
  wire _16205_;
  wire _16206_;
  wire _16207_;
  wire _16208_;
  wire _16209_;
  wire _16210_;
  wire _16211_;
  wire _16212_;
  wire _16213_;
  wire _16214_;
  wire _16215_;
  wire _16216_;
  wire _16217_;
  wire _16218_;
  wire _16219_;
  wire _16220_;
  wire _16221_;
  wire _16222_;
  wire _16223_;
  wire _16224_;
  wire _16225_;
  wire _16226_;
  wire _16227_;
  wire _16228_;
  wire _16229_;
  wire _16230_;
  wire _16231_;
  wire _16232_;
  wire _16233_;
  wire _16234_;
  wire _16235_;
  wire _16236_;
  wire _16237_;
  wire _16238_;
  wire _16239_;
  wire _16240_;
  wire _16241_;
  wire _16242_;
  wire _16243_;
  wire _16244_;
  wire _16245_;
  wire _16246_;
  wire _16247_;
  wire _16248_;
  wire _16249_;
  wire _16250_;
  wire _16251_;
  wire _16252_;
  wire _16253_;
  wire _16254_;
  wire _16255_;
  wire _16256_;
  wire _16257_;
  wire _16258_;
  wire _16259_;
  wire _16260_;
  wire _16261_;
  wire _16262_;
  wire _16263_;
  wire _16264_;
  wire _16265_;
  wire _16266_;
  wire _16267_;
  wire _16268_;
  wire _16269_;
  wire _16270_;
  wire _16271_;
  wire _16272_;
  wire _16273_;
  wire _16274_;
  wire _16275_;
  wire _16276_;
  wire _16277_;
  wire _16278_;
  wire _16279_;
  wire _16280_;
  wire _16281_;
  wire _16282_;
  wire _16283_;
  wire _16284_;
  wire _16285_;
  wire _16286_;
  wire _16287_;
  wire _16288_;
  wire _16289_;
  wire _16290_;
  wire _16291_;
  wire _16292_;
  wire _16293_;
  wire _16294_;
  wire _16295_;
  wire _16296_;
  wire _16297_;
  wire _16298_;
  wire _16299_;
  wire _16300_;
  wire _16301_;
  wire _16302_;
  wire _16303_;
  wire _16304_;
  wire _16305_;
  wire _16306_;
  wire _16307_;
  wire _16308_;
  wire _16309_;
  wire _16310_;
  wire _16311_;
  wire _16312_;
  wire _16313_;
  wire _16314_;
  wire _16315_;
  wire _16316_;
  wire _16317_;
  wire _16318_;
  wire _16319_;
  wire _16320_;
  wire _16321_;
  wire _16322_;
  wire _16323_;
  wire _16324_;
  wire _16325_;
  wire _16326_;
  wire _16327_;
  wire _16328_;
  wire _16329_;
  wire _16330_;
  wire _16331_;
  wire _16332_;
  wire _16333_;
  wire _16334_;
  wire _16335_;
  wire _16336_;
  wire _16337_;
  wire _16338_;
  wire _16339_;
  wire _16340_;
  wire _16341_;
  wire _16342_;
  wire _16343_;
  wire _16344_;
  wire _16345_;
  wire _16346_;
  wire _16347_;
  wire _16348_;
  wire _16349_;
  wire _16350_;
  wire _16351_;
  wire _16352_;
  wire _16353_;
  wire _16354_;
  wire _16355_;
  wire _16356_;
  wire _16357_;
  wire _16358_;
  wire _16359_;
  wire _16360_;
  wire _16361_;
  wire _16362_;
  wire _16363_;
  wire _16364_;
  wire _16365_;
  wire _16366_;
  wire _16367_;
  wire _16368_;
  wire _16369_;
  wire _16370_;
  wire _16371_;
  wire _16372_;
  wire _16373_;
  wire _16374_;
  wire _16375_;
  wire _16376_;
  wire _16377_;
  wire _16378_;
  wire _16379_;
  wire _16380_;
  wire _16381_;
  wire _16382_;
  wire _16383_;
  wire _16384_;
  wire _16385_;
  wire _16386_;
  wire _16387_;
  wire _16388_;
  wire _16389_;
  wire _16390_;
  wire _16391_;
  wire _16392_;
  wire _16393_;
  wire _16394_;
  wire _16395_;
  wire _16396_;
  wire _16397_;
  wire _16398_;
  wire _16399_;
  wire _16400_;
  wire _16401_;
  wire _16402_;
  wire _16403_;
  wire _16404_;
  wire _16405_;
  wire _16406_;
  wire _16407_;
  wire _16408_;
  wire _16409_;
  wire _16410_;
  wire _16411_;
  wire _16412_;
  wire _16413_;
  wire _16414_;
  wire _16415_;
  wire _16416_;
  wire _16417_;
  wire _16418_;
  wire _16419_;
  wire _16420_;
  wire _16421_;
  wire _16422_;
  wire _16423_;
  wire _16424_;
  wire _16425_;
  wire _16426_;
  wire _16427_;
  wire _16428_;
  wire _16429_;
  wire _16430_;
  wire _16431_;
  wire _16432_;
  wire _16433_;
  wire _16434_;
  wire _16435_;
  wire _16436_;
  wire _16437_;
  wire _16438_;
  wire _16439_;
  wire _16440_;
  wire _16441_;
  wire _16442_;
  wire _16443_;
  wire _16444_;
  wire _16445_;
  wire _16446_;
  wire _16447_;
  wire _16448_;
  wire _16449_;
  wire _16450_;
  wire _16451_;
  wire _16452_;
  wire _16453_;
  wire _16454_;
  wire _16455_;
  wire _16456_;
  wire _16457_;
  wire _16458_;
  wire _16459_;
  wire _16460_;
  wire _16461_;
  wire _16462_;
  wire _16463_;
  wire _16464_;
  wire _16465_;
  wire _16466_;
  wire _16467_;
  wire _16468_;
  wire _16469_;
  wire _16470_;
  wire _16471_;
  wire _16472_;
  wire _16473_;
  wire _16474_;
  wire _16475_;
  wire _16476_;
  wire _16477_;
  wire _16478_;
  wire _16479_;
  wire _16480_;
  wire _16481_;
  wire _16482_;
  wire _16483_;
  wire _16484_;
  wire _16485_;
  wire _16486_;
  wire _16487_;
  wire _16488_;
  wire _16489_;
  wire _16490_;
  wire _16491_;
  wire _16492_;
  wire _16493_;
  wire _16494_;
  wire _16495_;
  wire _16496_;
  wire _16497_;
  wire _16498_;
  wire _16499_;
  wire _16500_;
  wire _16501_;
  wire _16502_;
  wire _16503_;
  wire _16504_;
  wire _16505_;
  wire _16506_;
  wire _16507_;
  wire _16508_;
  wire _16509_;
  wire _16510_;
  wire _16511_;
  wire _16512_;
  wire _16513_;
  wire _16514_;
  wire _16515_;
  wire _16516_;
  wire _16517_;
  wire _16518_;
  wire _16519_;
  wire _16520_;
  wire _16521_;
  wire _16522_;
  wire _16523_;
  wire _16524_;
  wire _16525_;
  wire _16526_;
  wire _16527_;
  wire _16528_;
  wire _16529_;
  wire _16530_;
  wire _16531_;
  wire _16532_;
  wire _16533_;
  wire _16534_;
  wire _16535_;
  wire _16536_;
  wire _16537_;
  wire _16538_;
  wire _16539_;
  wire _16540_;
  wire _16541_;
  wire _16542_;
  wire _16543_;
  wire _16544_;
  wire _16545_;
  wire _16546_;
  wire _16547_;
  wire _16548_;
  wire _16549_;
  wire _16550_;
  wire _16551_;
  wire _16552_;
  wire _16553_;
  wire _16554_;
  wire _16555_;
  wire _16556_;
  wire _16557_;
  wire _16558_;
  wire _16559_;
  wire _16560_;
  wire _16561_;
  wire _16562_;
  wire _16563_;
  wire _16564_;
  wire _16565_;
  wire _16566_;
  wire _16567_;
  wire _16568_;
  wire _16569_;
  wire _16570_;
  wire _16571_;
  wire _16572_;
  wire _16573_;
  wire _16574_;
  wire _16575_;
  wire _16576_;
  wire _16577_;
  wire _16578_;
  wire _16579_;
  wire _16580_;
  wire _16581_;
  wire _16582_;
  wire _16583_;
  wire _16584_;
  wire _16585_;
  wire _16586_;
  wire _16587_;
  wire _16588_;
  wire _16589_;
  wire _16590_;
  wire _16591_;
  wire _16592_;
  wire _16593_;
  wire _16594_;
  wire _16595_;
  wire _16596_;
  wire _16597_;
  wire _16598_;
  wire _16599_;
  wire _16600_;
  wire _16601_;
  wire _16602_;
  wire _16603_;
  wire _16604_;
  wire _16605_;
  wire _16606_;
  wire _16607_;
  wire _16608_;
  wire _16609_;
  wire _16610_;
  wire _16611_;
  wire _16612_;
  wire _16613_;
  wire _16614_;
  wire _16615_;
  wire _16616_;
  wire _16617_;
  wire _16618_;
  wire _16619_;
  wire _16620_;
  wire _16621_;
  wire _16622_;
  wire _16623_;
  wire _16624_;
  wire _16625_;
  wire _16626_;
  wire _16627_;
  wire _16628_;
  wire _16629_;
  wire _16630_;
  wire _16631_;
  wire _16632_;
  wire _16633_;
  wire _16634_;
  wire _16635_;
  wire _16636_;
  wire _16637_;
  wire _16638_;
  wire _16639_;
  wire _16640_;
  wire _16641_;
  wire _16642_;
  wire _16643_;
  wire _16644_;
  wire _16645_;
  wire _16646_;
  wire _16647_;
  wire _16648_;
  wire _16649_;
  wire _16650_;
  wire _16651_;
  wire _16652_;
  wire _16653_;
  wire _16654_;
  wire _16655_;
  wire _16656_;
  wire _16657_;
  wire _16658_;
  wire _16659_;
  wire _16660_;
  wire _16661_;
  wire _16662_;
  wire _16663_;
  wire _16664_;
  wire _16665_;
  wire _16666_;
  wire _16667_;
  wire _16668_;
  wire _16669_;
  wire _16670_;
  wire _16671_;
  wire _16672_;
  wire _16673_;
  wire _16674_;
  wire _16675_;
  wire _16676_;
  wire _16677_;
  wire _16678_;
  wire _16679_;
  wire _16680_;
  wire _16681_;
  wire _16682_;
  wire _16683_;
  wire _16684_;
  wire _16685_;
  wire _16686_;
  wire _16687_;
  wire _16688_;
  wire _16689_;
  wire _16690_;
  wire _16691_;
  wire _16692_;
  wire _16693_;
  wire _16694_;
  wire _16695_;
  wire _16696_;
  wire _16697_;
  wire _16698_;
  wire _16699_;
  wire _16700_;
  wire _16701_;
  wire _16702_;
  wire _16703_;
  wire _16704_;
  wire _16705_;
  wire _16706_;
  wire _16707_;
  wire _16708_;
  wire _16709_;
  wire _16710_;
  wire _16711_;
  wire _16712_;
  wire _16713_;
  wire _16714_;
  wire _16715_;
  wire _16716_;
  wire _16717_;
  wire _16718_;
  wire _16719_;
  wire _16720_;
  wire _16721_;
  wire _16722_;
  wire _16723_;
  wire _16724_;
  wire _16725_;
  wire _16726_;
  wire _16727_;
  wire _16728_;
  wire _16729_;
  wire _16730_;
  wire _16731_;
  wire _16732_;
  wire _16733_;
  wire _16734_;
  wire _16735_;
  wire _16736_;
  wire _16737_;
  wire _16738_;
  wire _16739_;
  wire _16740_;
  wire _16741_;
  wire _16742_;
  wire _16743_;
  wire _16744_;
  wire _16745_;
  wire _16746_;
  wire _16747_;
  wire _16748_;
  wire _16749_;
  wire _16750_;
  wire _16751_;
  wire _16752_;
  wire _16753_;
  wire _16754_;
  wire _16755_;
  wire _16756_;
  wire _16757_;
  wire _16758_;
  wire _16759_;
  wire _16760_;
  wire _16761_;
  wire _16762_;
  wire _16763_;
  wire _16764_;
  wire _16765_;
  wire _16766_;
  wire _16767_;
  wire _16768_;
  wire _16769_;
  wire _16770_;
  wire _16771_;
  wire _16772_;
  wire _16773_;
  wire _16774_;
  wire _16775_;
  wire _16776_;
  wire _16777_;
  wire _16778_;
  wire _16779_;
  wire _16780_;
  wire _16781_;
  wire _16782_;
  wire _16783_;
  wire _16784_;
  wire _16785_;
  wire _16786_;
  wire _16787_;
  wire _16788_;
  wire _16789_;
  wire _16790_;
  wire _16791_;
  wire _16792_;
  wire _16793_;
  wire _16794_;
  wire _16795_;
  wire _16796_;
  wire _16797_;
  wire _16798_;
  wire _16799_;
  wire _16800_;
  wire _16801_;
  wire _16802_;
  wire _16803_;
  wire _16804_;
  wire _16805_;
  wire _16806_;
  wire _16807_;
  wire _16808_;
  wire _16809_;
  wire _16810_;
  wire _16811_;
  wire _16812_;
  wire _16813_;
  wire _16814_;
  wire _16815_;
  wire _16816_;
  wire _16817_;
  wire _16818_;
  wire _16819_;
  wire _16820_;
  wire _16821_;
  wire _16822_;
  wire _16823_;
  wire _16824_;
  wire _16825_;
  wire _16826_;
  wire _16827_;
  wire _16828_;
  wire _16829_;
  wire _16830_;
  wire _16831_;
  wire _16832_;
  wire _16833_;
  wire _16834_;
  wire _16835_;
  wire _16836_;
  wire _16837_;
  wire _16838_;
  wire _16839_;
  wire _16840_;
  wire _16841_;
  wire _16842_;
  wire _16843_;
  wire _16844_;
  wire _16845_;
  wire _16846_;
  wire _16847_;
  wire _16848_;
  wire _16849_;
  wire _16850_;
  wire _16851_;
  wire _16852_;
  wire _16853_;
  wire _16854_;
  wire _16855_;
  wire _16856_;
  wire _16857_;
  wire _16858_;
  wire _16859_;
  wire _16860_;
  wire _16861_;
  wire _16862_;
  wire _16863_;
  wire _16864_;
  wire _16865_;
  wire _16866_;
  wire _16867_;
  wire _16868_;
  wire _16869_;
  wire _16870_;
  wire _16871_;
  wire _16872_;
  wire _16873_;
  wire _16874_;
  wire _16875_;
  wire _16876_;
  wire _16877_;
  wire _16878_;
  wire _16879_;
  wire _16880_;
  wire _16881_;
  wire _16882_;
  wire _16883_;
  wire _16884_;
  wire _16885_;
  wire _16886_;
  wire _16887_;
  wire _16888_;
  wire _16889_;
  wire _16890_;
  wire _16891_;
  wire _16892_;
  wire _16893_;
  wire _16894_;
  wire _16895_;
  wire _16896_;
  wire _16897_;
  wire _16898_;
  wire _16899_;
  wire _16900_;
  wire _16901_;
  wire _16902_;
  wire _16903_;
  wire _16904_;
  wire _16905_;
  wire _16906_;
  wire _16907_;
  wire _16908_;
  wire _16909_;
  wire _16910_;
  wire _16911_;
  wire _16912_;
  wire _16913_;
  wire _16914_;
  wire _16915_;
  wire _16916_;
  wire _16917_;
  wire _16918_;
  wire _16919_;
  wire _16920_;
  wire _16921_;
  wire _16922_;
  wire _16923_;
  wire _16924_;
  wire _16925_;
  wire _16926_;
  wire _16927_;
  wire _16928_;
  wire _16929_;
  wire _16930_;
  wire _16931_;
  wire _16932_;
  wire _16933_;
  wire _16934_;
  wire _16935_;
  wire _16936_;
  wire _16937_;
  wire _16938_;
  wire _16939_;
  wire _16940_;
  wire _16941_;
  wire _16942_;
  wire _16943_;
  wire _16944_;
  wire _16945_;
  wire _16946_;
  wire _16947_;
  wire _16948_;
  wire _16949_;
  wire _16950_;
  wire _16951_;
  wire _16952_;
  wire _16953_;
  wire _16954_;
  wire _16955_;
  wire _16956_;
  wire _16957_;
  wire _16958_;
  wire _16959_;
  wire _16960_;
  wire _16961_;
  wire _16962_;
  wire _16963_;
  wire _16964_;
  wire _16965_;
  wire _16966_;
  wire _16967_;
  wire _16968_;
  wire _16969_;
  wire _16970_;
  wire _16971_;
  wire _16972_;
  wire _16973_;
  wire _16974_;
  wire _16975_;
  wire _16976_;
  wire _16977_;
  wire _16978_;
  wire _16979_;
  wire _16980_;
  wire _16981_;
  wire _16982_;
  wire _16983_;
  wire _16984_;
  wire _16985_;
  wire _16986_;
  wire _16987_;
  wire _16988_;
  wire _16989_;
  wire _16990_;
  wire _16991_;
  wire _16992_;
  wire _16993_;
  wire _16994_;
  wire _16995_;
  wire _16996_;
  wire _16997_;
  wire _16998_;
  wire _16999_;
  wire _17000_;
  wire _17001_;
  wire _17002_;
  wire _17003_;
  wire _17004_;
  wire _17005_;
  wire _17006_;
  wire _17007_;
  wire _17008_;
  wire _17009_;
  wire _17010_;
  wire _17011_;
  wire _17012_;
  wire _17013_;
  wire _17014_;
  wire _17015_;
  wire _17016_;
  wire _17017_;
  wire _17018_;
  wire _17019_;
  wire _17020_;
  wire _17021_;
  wire _17022_;
  wire _17023_;
  wire _17024_;
  wire _17025_;
  wire _17026_;
  wire _17027_;
  wire _17028_;
  wire _17029_;
  wire _17030_;
  wire _17031_;
  wire _17032_;
  wire _17033_;
  wire _17034_;
  wire _17035_;
  wire _17036_;
  wire _17037_;
  wire _17038_;
  wire _17039_;
  wire _17040_;
  wire _17041_;
  wire _17042_;
  wire _17043_;
  wire _17044_;
  wire _17045_;
  wire _17046_;
  wire _17047_;
  wire _17048_;
  wire _17049_;
  wire _17050_;
  wire _17051_;
  wire _17052_;
  wire _17053_;
  wire _17054_;
  wire _17055_;
  wire _17056_;
  wire _17057_;
  wire _17058_;
  wire _17059_;
  wire _17060_;
  wire _17061_;
  wire _17062_;
  wire _17063_;
  wire _17064_;
  wire _17065_;
  wire _17066_;
  wire _17067_;
  wire _17068_;
  wire _17069_;
  wire _17070_;
  wire _17071_;
  wire _17072_;
  wire _17073_;
  wire _17074_;
  wire _17075_;
  wire _17076_;
  wire _17077_;
  wire _17078_;
  wire _17079_;
  wire _17080_;
  wire _17081_;
  wire _17082_;
  wire _17083_;
  wire _17084_;
  wire _17085_;
  wire _17086_;
  wire _17087_;
  wire _17088_;
  wire _17089_;
  wire _17090_;
  wire _17091_;
  wire _17092_;
  wire _17093_;
  wire _17094_;
  wire _17095_;
  wire _17096_;
  wire _17097_;
  wire _17098_;
  wire _17099_;
  wire _17100_;
  wire _17101_;
  wire _17102_;
  wire _17103_;
  wire _17104_;
  wire _17105_;
  wire _17106_;
  wire _17107_;
  wire _17108_;
  wire _17109_;
  wire _17110_;
  wire _17111_;
  wire _17112_;
  wire _17113_;
  wire _17114_;
  wire _17115_;
  wire _17116_;
  wire _17117_;
  wire _17118_;
  wire _17119_;
  wire _17120_;
  wire _17121_;
  wire _17122_;
  wire _17123_;
  wire _17124_;
  wire _17125_;
  wire _17126_;
  wire _17127_;
  wire _17128_;
  wire _17129_;
  wire _17130_;
  wire _17131_;
  wire _17132_;
  wire _17133_;
  wire _17134_;
  wire _17135_;
  wire _17136_;
  wire _17137_;
  wire _17138_;
  wire _17139_;
  wire _17140_;
  wire _17141_;
  wire _17142_;
  wire _17143_;
  wire _17144_;
  wire _17145_;
  wire _17146_;
  wire _17147_;
  wire _17148_;
  wire _17149_;
  wire _17150_;
  wire _17151_;
  wire _17152_;
  wire _17153_;
  wire _17154_;
  wire _17155_;
  wire _17156_;
  wire _17157_;
  wire _17158_;
  wire _17159_;
  wire _17160_;
  wire _17161_;
  wire _17162_;
  wire _17163_;
  wire _17164_;
  wire _17165_;
  wire _17166_;
  wire _17167_;
  wire _17168_;
  wire _17169_;
  wire _17170_;
  wire _17171_;
  wire _17172_;
  wire _17173_;
  wire _17174_;
  wire _17175_;
  wire _17176_;
  wire _17177_;
  wire _17178_;
  wire _17179_;
  wire _17180_;
  wire _17181_;
  wire _17182_;
  wire _17183_;
  wire _17184_;
  wire _17185_;
  wire _17186_;
  wire _17187_;
  wire _17188_;
  wire _17189_;
  wire _17190_;
  wire _17191_;
  wire _17192_;
  wire _17193_;
  wire _17194_;
  wire _17195_;
  wire _17196_;
  wire _17197_;
  wire _17198_;
  wire _17199_;
  wire _17200_;
  wire _17201_;
  wire _17202_;
  wire _17203_;
  wire _17204_;
  wire _17205_;
  wire _17206_;
  wire _17207_;
  wire _17208_;
  wire _17209_;
  wire _17210_;
  wire _17211_;
  wire _17212_;
  wire _17213_;
  wire _17214_;
  wire _17215_;
  wire _17216_;
  wire _17217_;
  wire _17218_;
  wire _17219_;
  wire _17220_;
  wire _17221_;
  wire _17222_;
  wire _17223_;
  wire _17224_;
  wire _17225_;
  wire _17226_;
  wire _17227_;
  wire _17228_;
  wire _17229_;
  wire _17230_;
  wire _17231_;
  wire _17232_;
  wire _17233_;
  wire _17234_;
  wire _17235_;
  wire _17236_;
  wire _17237_;
  wire _17238_;
  wire _17239_;
  wire _17240_;
  wire _17241_;
  wire _17242_;
  wire _17243_;
  wire _17244_;
  wire _17245_;
  wire _17246_;
  wire _17247_;
  wire _17248_;
  wire _17249_;
  wire _17250_;
  wire _17251_;
  wire _17252_;
  wire _17253_;
  wire _17254_;
  wire _17255_;
  wire _17256_;
  wire _17257_;
  wire _17258_;
  wire _17259_;
  wire _17260_;
  wire _17261_;
  wire _17262_;
  wire _17263_;
  wire _17264_;
  wire _17265_;
  wire _17266_;
  wire _17267_;
  wire _17268_;
  wire _17269_;
  wire _17270_;
  wire _17271_;
  wire _17272_;
  wire _17273_;
  wire _17274_;
  wire _17275_;
  wire _17276_;
  wire _17277_;
  wire _17278_;
  wire _17279_;
  wire _17280_;
  wire _17281_;
  wire _17282_;
  wire _17283_;
  wire _17284_;
  wire _17285_;
  wire _17286_;
  wire _17287_;
  wire _17288_;
  wire _17289_;
  wire _17290_;
  wire _17291_;
  wire _17292_;
  wire _17293_;
  wire _17294_;
  wire _17295_;
  wire _17296_;
  wire _17297_;
  wire _17298_;
  wire _17299_;
  wire _17300_;
  wire _17301_;
  wire _17302_;
  wire _17303_;
  wire _17304_;
  wire _17305_;
  wire _17306_;
  wire _17307_;
  wire _17308_;
  wire _17309_;
  wire _17310_;
  wire _17311_;
  wire _17312_;
  wire _17313_;
  wire _17314_;
  wire _17315_;
  wire _17316_;
  wire _17317_;
  wire _17318_;
  wire _17319_;
  wire _17320_;
  wire _17321_;
  wire _17322_;
  wire _17323_;
  wire _17324_;
  wire _17325_;
  wire _17326_;
  wire _17327_;
  wire _17328_;
  wire _17329_;
  wire _17330_;
  wire _17331_;
  wire _17332_;
  wire _17333_;
  wire _17334_;
  wire _17335_;
  wire _17336_;
  wire _17337_;
  wire _17338_;
  wire _17339_;
  wire _17340_;
  wire _17341_;
  wire _17342_;
  wire _17343_;
  wire _17344_;
  wire _17345_;
  wire _17346_;
  wire _17347_;
  wire _17348_;
  wire _17349_;
  wire _17350_;
  wire _17351_;
  wire _17352_;
  wire _17353_;
  wire _17354_;
  wire _17355_;
  wire _17356_;
  wire _17357_;
  wire _17358_;
  wire _17359_;
  wire _17360_;
  wire _17361_;
  wire _17362_;
  wire _17363_;
  wire _17364_;
  wire _17365_;
  wire _17366_;
  wire _17367_;
  wire _17368_;
  wire _17369_;
  wire _17370_;
  wire _17371_;
  wire _17372_;
  wire _17373_;
  wire _17374_;
  wire _17375_;
  wire _17376_;
  wire _17377_;
  wire _17378_;
  wire _17379_;
  wire _17380_;
  wire _17381_;
  wire _17382_;
  wire _17383_;
  wire _17384_;
  wire _17385_;
  wire _17386_;
  wire _17387_;
  wire _17388_;
  wire _17389_;
  wire _17390_;
  wire _17391_;
  wire _17392_;
  wire _17393_;
  wire _17394_;
  wire _17395_;
  wire _17396_;
  wire _17397_;
  wire _17398_;
  wire _17399_;
  wire _17400_;
  wire _17401_;
  wire _17402_;
  wire _17403_;
  wire _17404_;
  wire _17405_;
  wire _17406_;
  wire _17407_;
  wire _17408_;
  wire _17409_;
  wire _17410_;
  wire _17411_;
  wire _17412_;
  wire _17413_;
  wire _17414_;
  wire _17415_;
  wire _17416_;
  wire _17417_;
  wire _17418_;
  wire _17419_;
  wire _17420_;
  wire _17421_;
  wire _17422_;
  wire _17423_;
  wire _17424_;
  wire _17425_;
  wire _17426_;
  wire _17427_;
  wire _17428_;
  wire _17429_;
  wire _17430_;
  wire _17431_;
  wire _17432_;
  wire _17433_;
  wire _17434_;
  wire _17435_;
  wire _17436_;
  wire _17437_;
  wire _17438_;
  wire _17439_;
  wire _17440_;
  wire _17441_;
  wire _17442_;
  wire _17443_;
  wire _17444_;
  wire _17445_;
  wire _17446_;
  wire _17447_;
  wire _17448_;
  wire _17449_;
  wire _17450_;
  wire _17451_;
  wire _17452_;
  wire _17453_;
  wire _17454_;
  wire _17455_;
  wire _17456_;
  wire _17457_;
  wire _17458_;
  wire _17459_;
  wire _17460_;
  wire _17461_;
  wire _17462_;
  wire _17463_;
  wire _17464_;
  wire _17465_;
  wire _17466_;
  wire _17467_;
  wire _17468_;
  wire _17469_;
  wire _17470_;
  wire _17471_;
  wire _17472_;
  wire _17473_;
  wire _17474_;
  wire _17475_;
  wire _17476_;
  wire _17477_;
  wire _17478_;
  wire _17479_;
  wire _17480_;
  wire _17481_;
  wire _17482_;
  wire _17483_;
  wire _17484_;
  wire _17485_;
  wire _17486_;
  wire _17487_;
  wire _17488_;
  wire _17489_;
  wire _17490_;
  wire _17491_;
  wire _17492_;
  wire _17493_;
  wire _17494_;
  wire _17495_;
  wire _17496_;
  wire _17497_;
  wire _17498_;
  wire _17499_;
  wire _17500_;
  wire _17501_;
  wire _17502_;
  wire _17503_;
  wire _17504_;
  wire _17505_;
  wire _17506_;
  wire _17507_;
  wire _17508_;
  wire _17509_;
  wire _17510_;
  wire _17511_;
  wire _17512_;
  wire _17513_;
  wire _17514_;
  wire _17515_;
  wire _17516_;
  wire _17517_;
  wire _17518_;
  wire _17519_;
  wire _17520_;
  wire _17521_;
  wire _17522_;
  wire _17523_;
  wire _17524_;
  wire _17525_;
  wire _17526_;
  wire _17527_;
  wire _17528_;
  wire _17529_;
  wire _17530_;
  wire _17531_;
  wire _17532_;
  wire _17533_;
  wire _17534_;
  wire _17535_;
  wire _17536_;
  wire _17537_;
  wire _17538_;
  wire _17539_;
  wire _17540_;
  wire _17541_;
  wire _17542_;
  wire _17543_;
  wire _17544_;
  wire _17545_;
  wire _17546_;
  wire _17547_;
  wire _17548_;
  wire _17549_;
  wire _17550_;
  wire _17551_;
  wire _17552_;
  wire _17553_;
  wire _17554_;
  wire _17555_;
  wire _17556_;
  wire _17557_;
  wire _17558_;
  wire _17559_;
  wire _17560_;
  wire _17561_;
  wire _17562_;
  wire _17563_;
  wire _17564_;
  wire _17565_;
  wire _17566_;
  wire _17567_;
  wire _17568_;
  wire _17569_;
  wire _17570_;
  wire _17571_;
  wire _17572_;
  wire _17573_;
  wire _17574_;
  wire _17575_;
  wire _17576_;
  wire _17577_;
  wire _17578_;
  wire _17579_;
  wire _17580_;
  wire _17581_;
  wire _17582_;
  wire _17583_;
  wire _17584_;
  wire _17585_;
  wire _17586_;
  wire _17587_;
  wire _17588_;
  wire _17589_;
  wire _17590_;
  wire _17591_;
  wire _17592_;
  wire _17593_;
  wire _17594_;
  wire _17595_;
  wire _17596_;
  wire _17597_;
  wire _17598_;
  wire _17599_;
  wire _17600_;
  wire _17601_;
  wire _17602_;
  wire _17603_;
  wire _17604_;
  wire _17605_;
  wire _17606_;
  wire _17607_;
  wire _17608_;
  wire _17609_;
  wire _17610_;
  wire _17611_;
  wire _17612_;
  wire _17613_;
  wire _17614_;
  wire _17615_;
  wire _17616_;
  wire _17617_;
  wire _17618_;
  wire _17619_;
  wire _17620_;
  wire _17621_;
  wire _17622_;
  wire _17623_;
  wire _17624_;
  wire _17625_;
  wire _17626_;
  wire _17627_;
  wire _17628_;
  wire _17629_;
  wire _17630_;
  wire _17631_;
  wire _17632_;
  wire _17633_;
  wire _17634_;
  wire _17635_;
  wire _17636_;
  wire _17637_;
  wire _17638_;
  wire _17639_;
  wire _17640_;
  wire _17641_;
  wire _17642_;
  wire _17643_;
  wire _17644_;
  wire _17645_;
  wire _17646_;
  wire _17647_;
  wire _17648_;
  wire _17649_;
  wire _17650_;
  wire _17651_;
  wire _17652_;
  wire _17653_;
  wire _17654_;
  wire _17655_;
  wire _17656_;
  wire _17657_;
  wire _17658_;
  wire _17659_;
  wire _17660_;
  wire _17661_;
  wire _17662_;
  wire _17663_;
  wire _17664_;
  wire _17665_;
  wire _17666_;
  wire _17667_;
  wire _17668_;
  wire _17669_;
  wire _17670_;
  wire _17671_;
  wire _17672_;
  wire _17673_;
  wire _17674_;
  wire _17675_;
  wire _17676_;
  wire _17677_;
  wire _17678_;
  wire _17679_;
  wire _17680_;
  wire _17681_;
  wire _17682_;
  wire _17683_;
  wire _17684_;
  wire _17685_;
  wire _17686_;
  wire _17687_;
  wire _17688_;
  wire _17689_;
  wire _17690_;
  wire _17691_;
  wire _17692_;
  wire _17693_;
  wire _17694_;
  wire _17695_;
  wire _17696_;
  wire _17697_;
  wire _17698_;
  wire _17699_;
  wire _17700_;
  wire _17701_;
  wire _17702_;
  wire _17703_;
  wire _17704_;
  wire _17705_;
  wire _17706_;
  wire _17707_;
  wire _17708_;
  wire _17709_;
  wire _17710_;
  wire _17711_;
  wire _17712_;
  wire _17713_;
  wire _17714_;
  wire _17715_;
  wire _17716_;
  wire _17717_;
  wire _17718_;
  wire _17719_;
  wire _17720_;
  wire _17721_;
  wire _17722_;
  wire _17723_;
  wire _17724_;
  wire _17725_;
  wire _17726_;
  wire _17727_;
  wire _17728_;
  wire _17729_;
  wire _17730_;
  wire _17731_;
  wire _17732_;
  wire _17733_;
  wire _17734_;
  wire _17735_;
  wire _17736_;
  wire _17737_;
  wire _17738_;
  wire _17739_;
  wire _17740_;
  wire _17741_;
  wire _17742_;
  wire _17743_;
  wire _17744_;
  wire _17745_;
  wire _17746_;
  wire _17747_;
  wire _17748_;
  wire _17749_;
  wire _17750_;
  wire _17751_;
  wire _17752_;
  wire _17753_;
  wire _17754_;
  wire _17755_;
  wire _17756_;
  wire _17757_;
  wire _17758_;
  wire _17759_;
  wire _17760_;
  wire _17761_;
  wire _17762_;
  wire _17763_;
  wire _17764_;
  wire _17765_;
  wire _17766_;
  wire _17767_;
  wire _17768_;
  wire _17769_;
  wire _17770_;
  wire _17771_;
  wire _17772_;
  wire _17773_;
  wire _17774_;
  wire _17775_;
  wire _17776_;
  wire _17777_;
  wire _17778_;
  wire _17779_;
  wire _17780_;
  wire _17781_;
  wire _17782_;
  wire _17783_;
  wire _17784_;
  wire _17785_;
  wire _17786_;
  wire _17787_;
  wire _17788_;
  wire _17789_;
  wire _17790_;
  wire _17791_;
  wire _17792_;
  wire _17793_;
  wire _17794_;
  wire _17795_;
  wire _17796_;
  wire _17797_;
  wire _17798_;
  wire _17799_;
  wire _17800_;
  wire _17801_;
  wire _17802_;
  wire _17803_;
  wire _17804_;
  wire _17805_;
  wire _17806_;
  wire _17807_;
  wire _17808_;
  wire _17809_;
  wire _17810_;
  wire _17811_;
  wire _17812_;
  wire _17813_;
  wire _17814_;
  wire _17815_;
  wire _17816_;
  wire _17817_;
  wire _17818_;
  wire _17819_;
  wire _17820_;
  wire _17821_;
  wire _17822_;
  wire _17823_;
  wire _17824_;
  wire _17825_;
  wire _17826_;
  wire _17827_;
  wire _17828_;
  wire _17829_;
  wire _17830_;
  wire _17831_;
  wire _17832_;
  wire _17833_;
  wire _17834_;
  wire _17835_;
  wire _17836_;
  wire _17837_;
  wire _17838_;
  wire _17839_;
  wire _17840_;
  wire _17841_;
  wire _17842_;
  wire _17843_;
  wire _17844_;
  wire _17845_;
  wire _17846_;
  wire _17847_;
  wire _17848_;
  wire _17849_;
  wire _17850_;
  wire _17851_;
  wire _17852_;
  wire _17853_;
  wire _17854_;
  wire _17855_;
  wire _17856_;
  wire _17857_;
  wire _17858_;
  wire _17859_;
  wire _17860_;
  wire _17861_;
  wire _17862_;
  wire _17863_;
  wire _17864_;
  wire _17865_;
  wire _17866_;
  wire _17867_;
  wire _17868_;
  wire _17869_;
  wire _17870_;
  wire _17871_;
  wire _17872_;
  wire _17873_;
  wire _17874_;
  wire _17875_;
  wire _17876_;
  wire _17877_;
  wire _17878_;
  wire _17879_;
  wire _17880_;
  wire _17881_;
  wire _17882_;
  wire _17883_;
  wire _17884_;
  wire _17885_;
  wire _17886_;
  wire _17887_;
  wire _17888_;
  wire _17889_;
  wire _17890_;
  wire _17891_;
  wire _17892_;
  wire _17893_;
  wire _17894_;
  wire _17895_;
  wire _17896_;
  wire _17897_;
  wire _17898_;
  wire _17899_;
  wire _17900_;
  wire _17901_;
  wire _17902_;
  wire _17903_;
  wire _17904_;
  wire _17905_;
  wire _17906_;
  wire _17907_;
  wire _17908_;
  wire _17909_;
  wire _17910_;
  wire _17911_;
  wire _17912_;
  wire _17913_;
  wire _17914_;
  wire _17915_;
  wire _17916_;
  wire _17917_;
  wire _17918_;
  wire _17919_;
  wire _17920_;
  wire _17921_;
  wire _17922_;
  wire _17923_;
  wire _17924_;
  wire _17925_;
  wire _17926_;
  wire _17927_;
  wire _17928_;
  wire _17929_;
  wire _17930_;
  wire _17931_;
  wire _17932_;
  wire _17933_;
  wire _17934_;
  wire _17935_;
  wire _17936_;
  wire _17937_;
  wire _17938_;
  wire _17939_;
  wire _17940_;
  wire _17941_;
  wire _17942_;
  wire _17943_;
  wire _17944_;
  wire _17945_;
  wire _17946_;
  wire _17947_;
  wire _17948_;
  wire _17949_;
  wire _17950_;
  wire _17951_;
  wire _17952_;
  wire _17953_;
  wire _17954_;
  wire _17955_;
  wire _17956_;
  wire _17957_;
  wire _17958_;
  wire _17959_;
  wire _17960_;
  wire _17961_;
  wire _17962_;
  wire _17963_;
  wire _17964_;
  wire _17965_;
  wire _17966_;
  wire _17967_;
  wire _17968_;
  wire _17969_;
  wire _17970_;
  wire _17971_;
  wire _17972_;
  wire _17973_;
  wire _17974_;
  wire _17975_;
  wire _17976_;
  wire _17977_;
  wire _17978_;
  wire _17979_;
  wire _17980_;
  wire _17981_;
  wire _17982_;
  wire _17983_;
  wire _17984_;
  wire _17985_;
  wire _17986_;
  wire _17987_;
  wire _17988_;
  wire _17989_;
  wire _17990_;
  wire _17991_;
  wire _17992_;
  wire _17993_;
  wire _17994_;
  wire _17995_;
  wire _17996_;
  wire _17997_;
  wire _17998_;
  wire _17999_;
  wire _18000_;
  wire _18001_;
  wire _18002_;
  wire _18003_;
  wire _18004_;
  wire _18005_;
  wire _18006_;
  wire _18007_;
  wire _18008_;
  wire _18009_;
  wire _18010_;
  wire _18011_;
  wire _18012_;
  wire _18013_;
  wire _18014_;
  wire _18015_;
  wire _18016_;
  wire _18017_;
  wire _18018_;
  wire _18019_;
  wire _18020_;
  wire _18021_;
  wire _18022_;
  wire _18023_;
  wire _18024_;
  wire _18025_;
  wire _18026_;
  wire _18027_;
  wire _18028_;
  wire _18029_;
  wire _18030_;
  wire _18031_;
  wire _18032_;
  wire _18033_;
  wire _18034_;
  wire _18035_;
  wire _18036_;
  wire _18037_;
  wire _18038_;
  wire _18039_;
  wire _18040_;
  wire _18041_;
  wire _18042_;
  wire _18043_;
  wire _18044_;
  wire _18045_;
  wire _18046_;
  wire _18047_;
  wire _18048_;
  wire _18049_;
  wire _18050_;
  wire _18051_;
  wire _18052_;
  wire _18053_;
  wire _18054_;
  wire _18055_;
  wire _18056_;
  wire _18057_;
  wire _18058_;
  wire _18059_;
  wire _18060_;
  wire _18061_;
  wire _18062_;
  wire _18063_;
  wire _18064_;
  wire _18065_;
  wire _18066_;
  wire _18067_;
  wire _18068_;
  wire _18069_;
  wire _18070_;
  wire _18071_;
  wire _18072_;
  wire _18073_;
  wire _18074_;
  wire _18075_;
  wire _18076_;
  wire _18077_;
  wire _18078_;
  wire _18079_;
  wire _18080_;
  wire _18081_;
  wire _18082_;
  wire _18083_;
  wire _18084_;
  wire _18085_;
  wire _18086_;
  wire _18087_;
  wire _18088_;
  wire _18089_;
  wire _18090_;
  wire _18091_;
  wire _18092_;
  wire _18093_;
  wire _18094_;
  wire _18095_;
  wire _18096_;
  wire _18097_;
  wire _18098_;
  wire _18099_;
  wire _18100_;
  wire _18101_;
  wire _18102_;
  wire _18103_;
  wire _18104_;
  wire _18105_;
  wire _18106_;
  wire _18107_;
  wire _18108_;
  wire _18109_;
  wire _18110_;
  wire _18111_;
  wire _18112_;
  wire _18113_;
  wire _18114_;
  wire _18115_;
  wire _18116_;
  wire _18117_;
  wire _18118_;
  wire _18119_;
  wire _18120_;
  wire _18121_;
  wire _18122_;
  wire _18123_;
  wire _18124_;
  wire _18125_;
  wire _18126_;
  wire _18127_;
  wire _18128_;
  wire _18129_;
  wire _18130_;
  wire _18131_;
  wire _18132_;
  wire _18133_;
  wire _18134_;
  wire _18135_;
  wire _18136_;
  wire _18137_;
  wire _18138_;
  wire _18139_;
  wire _18140_;
  wire _18141_;
  wire _18142_;
  wire _18143_;
  wire _18144_;
  wire _18145_;
  wire _18146_;
  wire _18147_;
  wire _18148_;
  wire _18149_;
  wire _18150_;
  wire _18151_;
  wire _18152_;
  wire _18153_;
  wire _18154_;
  wire _18155_;
  wire _18156_;
  wire _18157_;
  wire _18158_;
  wire _18159_;
  wire _18160_;
  wire _18161_;
  wire _18162_;
  wire _18163_;
  wire _18164_;
  wire _18165_;
  wire _18166_;
  wire _18167_;
  wire _18168_;
  wire _18169_;
  wire _18170_;
  wire _18171_;
  wire _18172_;
  wire _18173_;
  wire _18174_;
  wire _18175_;
  wire _18176_;
  wire _18177_;
  wire _18178_;
  wire _18179_;
  wire _18180_;
  wire _18181_;
  wire _18182_;
  wire _18183_;
  wire _18184_;
  wire _18185_;
  wire _18186_;
  wire _18187_;
  wire _18188_;
  wire _18189_;
  wire _18190_;
  wire _18191_;
  wire _18192_;
  wire _18193_;
  wire _18194_;
  wire _18195_;
  wire _18196_;
  wire _18197_;
  wire _18198_;
  wire _18199_;
  wire _18200_;
  wire _18201_;
  wire _18202_;
  wire _18203_;
  wire _18204_;
  wire _18205_;
  wire _18206_;
  wire _18207_;
  wire _18208_;
  wire _18209_;
  wire _18210_;
  wire _18211_;
  wire _18212_;
  wire _18213_;
  wire _18214_;
  wire _18215_;
  wire _18216_;
  wire _18217_;
  wire _18218_;
  wire _18219_;
  wire _18220_;
  wire _18221_;
  wire _18222_;
  wire _18223_;
  wire _18224_;
  wire _18225_;
  wire _18226_;
  wire _18227_;
  wire _18228_;
  wire _18229_;
  wire _18230_;
  wire _18231_;
  wire _18232_;
  wire _18233_;
  wire _18234_;
  wire _18235_;
  wire _18236_;
  wire _18237_;
  wire _18238_;
  wire _18239_;
  wire _18240_;
  wire _18241_;
  wire _18242_;
  wire _18243_;
  wire _18244_;
  wire _18245_;
  wire _18246_;
  wire _18247_;
  wire _18248_;
  wire _18249_;
  wire _18250_;
  wire _18251_;
  wire _18252_;
  wire _18253_;
  wire _18254_;
  wire _18255_;
  wire _18256_;
  wire _18257_;
  wire _18258_;
  wire _18259_;
  wire _18260_;
  wire _18261_;
  wire _18262_;
  wire _18263_;
  wire _18264_;
  wire _18265_;
  wire _18266_;
  wire _18267_;
  wire _18268_;
  wire _18269_;
  wire _18270_;
  wire _18271_;
  wire _18272_;
  wire _18273_;
  wire _18274_;
  wire _18275_;
  wire _18276_;
  wire _18277_;
  wire _18278_;
  wire _18279_;
  wire _18280_;
  wire _18281_;
  wire _18282_;
  wire _18283_;
  wire _18284_;
  wire _18285_;
  wire _18286_;
  wire _18287_;
  wire _18288_;
  wire _18289_;
  wire _18290_;
  wire _18291_;
  wire _18292_;
  wire _18293_;
  wire _18294_;
  wire _18295_;
  wire _18296_;
  wire _18297_;
  wire _18298_;
  wire _18299_;
  wire _18300_;
  wire _18301_;
  wire _18302_;
  wire _18303_;
  wire _18304_;
  wire _18305_;
  wire _18306_;
  wire _18307_;
  wire _18308_;
  wire _18309_;
  wire _18310_;
  wire _18311_;
  wire _18312_;
  wire _18313_;
  wire _18314_;
  wire _18315_;
  wire _18316_;
  wire _18317_;
  wire _18318_;
  wire _18319_;
  wire _18320_;
  wire _18321_;
  wire _18322_;
  wire _18323_;
  wire _18324_;
  wire _18325_;
  wire _18326_;
  wire _18327_;
  wire _18328_;
  wire _18329_;
  wire _18330_;
  wire _18331_;
  wire _18332_;
  wire _18333_;
  wire _18334_;
  wire _18335_;
  wire _18336_;
  wire _18337_;
  wire _18338_;
  wire _18339_;
  wire _18340_;
  wire _18341_;
  wire _18342_;
  wire _18343_;
  wire _18344_;
  wire _18345_;
  wire _18346_;
  wire _18347_;
  wire _18348_;
  wire _18349_;
  wire _18350_;
  wire _18351_;
  wire _18352_;
  wire _18353_;
  wire _18354_;
  wire _18355_;
  wire _18356_;
  wire _18357_;
  wire _18358_;
  wire _18359_;
  wire _18360_;
  wire _18361_;
  wire _18362_;
  wire _18363_;
  wire _18364_;
  wire _18365_;
  wire _18366_;
  wire _18367_;
  wire _18368_;
  wire _18369_;
  wire _18370_;
  wire _18371_;
  wire _18372_;
  wire _18373_;
  wire _18374_;
  wire _18375_;
  wire _18376_;
  wire _18377_;
  wire _18378_;
  wire _18379_;
  wire _18380_;
  wire _18381_;
  wire _18382_;
  wire _18383_;
  wire _18384_;
  wire _18385_;
  wire _18386_;
  wire _18387_;
  wire _18388_;
  wire _18389_;
  wire _18390_;
  wire _18391_;
  wire _18392_;
  wire _18393_;
  wire _18394_;
  wire _18395_;
  wire _18396_;
  wire _18397_;
  wire _18398_;
  wire _18399_;
  wire _18400_;
  wire _18401_;
  wire _18402_;
  wire _18403_;
  wire _18404_;
  wire _18405_;
  wire _18406_;
  wire _18407_;
  wire _18408_;
  wire _18409_;
  wire _18410_;
  wire _18411_;
  wire _18412_;
  wire _18413_;
  wire _18414_;
  wire _18415_;
  wire _18416_;
  wire _18417_;
  wire _18418_;
  wire _18419_;
  wire _18420_;
  wire _18421_;
  wire _18422_;
  wire _18423_;
  wire _18424_;
  wire _18425_;
  wire _18426_;
  wire _18427_;
  wire _18428_;
  wire _18429_;
  wire _18430_;
  wire _18431_;
  wire _18432_;
  wire _18433_;
  wire _18434_;
  wire _18435_;
  wire _18436_;
  wire _18437_;
  wire _18438_;
  wire _18439_;
  wire _18440_;
  wire _18441_;
  wire _18442_;
  wire _18443_;
  wire _18444_;
  wire _18445_;
  wire _18446_;
  wire _18447_;
  wire _18448_;
  wire _18449_;
  wire _18450_;
  wire _18451_;
  wire _18452_;
  wire _18453_;
  wire _18454_;
  wire _18455_;
  wire _18456_;
  wire _18457_;
  wire _18458_;
  wire _18459_;
  wire _18460_;
  wire _18461_;
  wire _18462_;
  wire _18463_;
  wire _18464_;
  wire _18465_;
  wire _18466_;
  wire _18467_;
  wire _18468_;
  wire _18469_;
  wire _18470_;
  wire _18471_;
  wire _18472_;
  wire _18473_;
  wire _18474_;
  wire _18475_;
  wire _18476_;
  wire _18477_;
  wire _18478_;
  wire _18479_;
  wire _18480_;
  wire _18481_;
  wire _18482_;
  wire _18483_;
  wire _18484_;
  wire _18485_;
  wire _18486_;
  wire _18487_;
  wire _18488_;
  wire _18489_;
  wire _18490_;
  wire _18491_;
  wire _18492_;
  wire _18493_;
  wire _18494_;
  wire _18495_;
  wire _18496_;
  wire _18497_;
  wire _18498_;
  wire _18499_;
  wire _18500_;
  wire _18501_;
  wire _18502_;
  wire _18503_;
  wire _18504_;
  wire _18505_;
  wire _18506_;
  wire _18507_;
  wire _18508_;
  wire _18509_;
  wire _18510_;
  wire _18511_;
  wire _18512_;
  wire _18513_;
  wire _18514_;
  wire _18515_;
  wire _18516_;
  wire _18517_;
  wire _18518_;
  wire _18519_;
  wire _18520_;
  wire _18521_;
  wire _18522_;
  wire _18523_;
  wire _18524_;
  wire _18525_;
  wire _18526_;
  wire _18527_;
  wire _18528_;
  wire _18529_;
  wire _18530_;
  wire _18531_;
  wire _18532_;
  wire _18533_;
  wire _18534_;
  wire _18535_;
  wire _18536_;
  wire _18537_;
  wire _18538_;
  wire _18539_;
  wire _18540_;
  wire _18541_;
  wire _18542_;
  wire _18543_;
  wire _18544_;
  wire _18545_;
  wire _18546_;
  wire _18547_;
  wire _18548_;
  wire _18549_;
  wire _18550_;
  wire _18551_;
  wire _18552_;
  wire _18553_;
  wire _18554_;
  wire _18555_;
  wire _18556_;
  wire _18557_;
  wire _18558_;
  wire _18559_;
  wire _18560_;
  wire _18561_;
  wire _18562_;
  wire _18563_;
  wire _18564_;
  wire _18565_;
  wire _18566_;
  wire _18567_;
  wire _18568_;
  wire _18569_;
  wire _18570_;
  wire _18571_;
  wire _18572_;
  wire _18573_;
  wire _18574_;
  wire _18575_;
  wire _18576_;
  wire _18577_;
  wire _18578_;
  wire _18579_;
  wire _18580_;
  wire _18581_;
  wire _18582_;
  wire _18583_;
  wire _18584_;
  wire _18585_;
  wire _18586_;
  wire _18587_;
  wire _18588_;
  wire _18589_;
  wire _18590_;
  wire _18591_;
  wire _18592_;
  wire _18593_;
  wire _18594_;
  wire _18595_;
  wire _18596_;
  wire _18597_;
  wire _18598_;
  wire _18599_;
  wire _18600_;
  wire _18601_;
  wire _18602_;
  wire _18603_;
  wire _18604_;
  wire _18605_;
  wire _18606_;
  wire _18607_;
  wire _18608_;
  wire _18609_;
  wire _18610_;
  wire _18611_;
  wire _18612_;
  wire _18613_;
  wire _18614_;
  wire _18615_;
  wire _18616_;
  wire _18617_;
  wire _18618_;
  wire _18619_;
  wire _18620_;
  wire _18621_;
  wire _18622_;
  wire _18623_;
  wire _18624_;
  wire _18625_;
  wire _18626_;
  wire _18627_;
  wire _18628_;
  wire _18629_;
  wire _18630_;
  wire _18631_;
  wire _18632_;
  wire _18633_;
  wire _18634_;
  wire _18635_;
  wire _18636_;
  wire _18637_;
  wire _18638_;
  wire _18639_;
  wire _18640_;
  wire _18641_;
  wire _18642_;
  wire _18643_;
  wire _18644_;
  wire _18645_;
  wire _18646_;
  wire _18647_;
  wire _18648_;
  wire _18649_;
  wire _18650_;
  wire _18651_;
  wire _18652_;
  wire _18653_;
  wire _18654_;
  wire _18655_;
  wire _18656_;
  wire _18657_;
  wire _18658_;
  wire _18659_;
  wire _18660_;
  wire _18661_;
  wire _18662_;
  wire _18663_;
  wire _18664_;
  wire _18665_;
  wire _18666_;
  wire _18667_;
  wire _18668_;
  wire _18669_;
  wire _18670_;
  wire _18671_;
  wire _18672_;
  wire _18673_;
  wire _18674_;
  wire _18675_;
  wire _18676_;
  wire _18677_;
  wire _18678_;
  wire _18679_;
  wire _18680_;
  wire _18681_;
  wire _18682_;
  wire _18683_;
  wire _18684_;
  wire _18685_;
  wire _18686_;
  wire _18687_;
  wire _18688_;
  wire _18689_;
  wire _18690_;
  wire _18691_;
  wire _18692_;
  wire _18693_;
  wire _18694_;
  wire _18695_;
  wire _18696_;
  wire _18697_;
  wire _18698_;
  wire _18699_;
  wire _18700_;
  wire _18701_;
  wire _18702_;
  wire _18703_;
  wire _18704_;
  wire _18705_;
  wire _18706_;
  wire _18707_;
  wire _18708_;
  wire _18709_;
  wire _18710_;
  wire _18711_;
  wire _18712_;
  wire _18713_;
  wire _18714_;
  wire _18715_;
  wire _18716_;
  wire _18717_;
  wire _18718_;
  wire _18719_;
  wire _18720_;
  wire _18721_;
  wire _18722_;
  wire _18723_;
  wire _18724_;
  wire _18725_;
  wire _18726_;
  wire _18727_;
  wire _18728_;
  wire _18729_;
  wire _18730_;
  wire _18731_;
  wire _18732_;
  wire _18733_;
  wire _18734_;
  wire _18735_;
  wire _18736_;
  wire _18737_;
  wire _18738_;
  wire _18739_;
  wire _18740_;
  wire _18741_;
  wire _18742_;
  wire _18743_;
  wire _18744_;
  wire _18745_;
  wire _18746_;
  wire _18747_;
  wire _18748_;
  wire _18749_;
  wire _18750_;
  wire _18751_;
  wire _18752_;
  wire _18753_;
  wire _18754_;
  wire _18755_;
  wire _18756_;
  wire _18757_;
  wire _18758_;
  wire _18759_;
  wire _18760_;
  wire _18761_;
  wire _18762_;
  wire _18763_;
  wire _18764_;
  wire _18765_;
  wire _18766_;
  wire _18767_;
  wire _18768_;
  wire _18769_;
  wire _18770_;
  wire _18771_;
  wire _18772_;
  wire _18773_;
  wire _18774_;
  wire _18775_;
  wire _18776_;
  wire _18777_;
  wire _18778_;
  wire _18779_;
  wire _18780_;
  wire _18781_;
  wire _18782_;
  wire _18783_;
  wire _18784_;
  wire _18785_;
  wire _18786_;
  wire _18787_;
  wire _18788_;
  wire _18789_;
  wire _18790_;
  wire _18791_;
  wire _18792_;
  wire _18793_;
  wire _18794_;
  wire _18795_;
  wire _18796_;
  wire _18797_;
  wire _18798_;
  wire _18799_;
  wire _18800_;
  wire _18801_;
  wire _18802_;
  wire _18803_;
  wire _18804_;
  wire _18805_;
  wire _18806_;
  wire _18807_;
  wire _18808_;
  wire _18809_;
  wire _18810_;
  wire _18811_;
  wire _18812_;
  wire _18813_;
  wire _18814_;
  wire _18815_;
  wire _18816_;
  wire _18817_;
  wire _18818_;
  wire _18819_;
  wire _18820_;
  wire _18821_;
  wire _18822_;
  wire _18823_;
  wire _18824_;
  wire _18825_;
  wire _18826_;
  wire _18827_;
  wire _18828_;
  wire _18829_;
  wire _18830_;
  wire _18831_;
  wire _18832_;
  wire _18833_;
  wire _18834_;
  wire _18835_;
  wire _18836_;
  wire _18837_;
  wire _18838_;
  wire _18839_;
  wire _18840_;
  wire _18841_;
  wire _18842_;
  wire _18843_;
  wire _18844_;
  wire _18845_;
  wire _18846_;
  wire _18847_;
  wire _18848_;
  wire _18849_;
  wire _18850_;
  wire _18851_;
  wire _18852_;
  wire _18853_;
  wire _18854_;
  wire _18855_;
  wire _18856_;
  wire _18857_;
  wire _18858_;
  wire _18859_;
  wire _18860_;
  wire _18861_;
  wire _18862_;
  wire _18863_;
  wire _18864_;
  wire _18865_;
  wire _18866_;
  wire _18867_;
  wire _18868_;
  wire _18869_;
  wire _18870_;
  wire _18871_;
  wire _18872_;
  wire _18873_;
  wire _18874_;
  wire _18875_;
  wire _18876_;
  wire _18877_;
  wire _18878_;
  wire _18879_;
  wire _18880_;
  wire _18881_;
  wire _18882_;
  wire _18883_;
  wire _18884_;
  wire _18885_;
  wire _18886_;
  wire _18887_;
  wire _18888_;
  wire _18889_;
  wire _18890_;
  wire _18891_;
  wire _18892_;
  wire _18893_;
  wire _18894_;
  wire _18895_;
  wire _18896_;
  wire _18897_;
  wire _18898_;
  wire _18899_;
  wire _18900_;
  wire _18901_;
  wire _18902_;
  wire _18903_;
  wire _18904_;
  wire _18905_;
  wire _18906_;
  wire _18907_;
  wire _18908_;
  wire _18909_;
  wire _18910_;
  wire _18911_;
  wire _18912_;
  wire _18913_;
  wire _18914_;
  wire _18915_;
  wire _18916_;
  wire _18917_;
  wire _18918_;
  wire _18919_;
  wire _18920_;
  wire _18921_;
  wire _18922_;
  wire _18923_;
  wire _18924_;
  wire _18925_;
  wire _18926_;
  wire _18927_;
  wire _18928_;
  wire _18929_;
  wire _18930_;
  wire _18931_;
  wire _18932_;
  wire _18933_;
  wire _18934_;
  wire _18935_;
  wire _18936_;
  wire _18937_;
  wire _18938_;
  wire _18939_;
  wire _18940_;
  wire _18941_;
  wire _18942_;
  wire _18943_;
  wire _18944_;
  wire _18945_;
  wire _18946_;
  wire _18947_;
  wire _18948_;
  wire _18949_;
  wire _18950_;
  wire _18951_;
  wire _18952_;
  wire _18953_;
  wire _18954_;
  wire _18955_;
  wire _18956_;
  wire _18957_;
  wire _18958_;
  wire _18959_;
  wire _18960_;
  wire _18961_;
  wire _18962_;
  wire _18963_;
  wire _18964_;
  wire _18965_;
  wire _18966_;
  wire _18967_;
  wire _18968_;
  wire _18969_;
  wire _18970_;
  wire _18971_;
  wire _18972_;
  wire _18973_;
  wire _18974_;
  wire _18975_;
  wire _18976_;
  wire _18977_;
  wire _18978_;
  wire _18979_;
  wire _18980_;
  wire _18981_;
  wire _18982_;
  wire _18983_;
  wire _18984_;
  wire _18985_;
  wire _18986_;
  wire _18987_;
  wire _18988_;
  wire _18989_;
  wire _18990_;
  wire _18991_;
  wire _18992_;
  wire _18993_;
  wire _18994_;
  wire _18995_;
  wire _18996_;
  wire _18997_;
  wire _18998_;
  wire _18999_;
  wire _19000_;
  wire _19001_;
  wire _19002_;
  wire _19003_;
  wire _19004_;
  wire _19005_;
  wire _19006_;
  wire _19007_;
  wire _19008_;
  wire _19009_;
  wire _19010_;
  wire _19011_;
  wire _19012_;
  wire _19013_;
  wire _19014_;
  wire _19015_;
  wire _19016_;
  wire _19017_;
  wire _19018_;
  wire _19019_;
  wire _19020_;
  wire _19021_;
  wire _19022_;
  wire _19023_;
  wire _19024_;
  wire _19025_;
  wire _19026_;
  wire _19027_;
  wire _19028_;
  wire _19029_;
  wire _19030_;
  wire _19031_;
  wire _19032_;
  wire _19033_;
  wire _19034_;
  wire _19035_;
  wire _19036_;
  wire _19037_;
  wire _19038_;
  wire _19039_;
  wire _19040_;
  wire _19041_;
  wire _19042_;
  wire _19043_;
  wire _19044_;
  wire _19045_;
  wire _19046_;
  wire _19047_;
  wire _19048_;
  wire _19049_;
  wire _19050_;
  wire _19051_;
  wire _19052_;
  wire _19053_;
  wire _19054_;
  wire _19055_;
  wire _19056_;
  wire _19057_;
  wire _19058_;
  wire _19059_;
  wire _19060_;
  wire _19061_;
  wire _19062_;
  wire _19063_;
  wire _19064_;
  wire _19065_;
  wire _19066_;
  wire _19067_;
  wire _19068_;
  wire _19069_;
  wire _19070_;
  wire _19071_;
  wire _19072_;
  wire _19073_;
  wire _19074_;
  wire _19075_;
  wire _19076_;
  wire _19077_;
  wire _19078_;
  wire _19079_;
  wire _19080_;
  wire _19081_;
  wire _19082_;
  wire _19083_;
  wire _19084_;
  wire _19085_;
  wire _19086_;
  wire _19087_;
  wire _19088_;
  wire _19089_;
  wire _19090_;
  wire _19091_;
  wire _19092_;
  wire _19093_;
  wire _19094_;
  wire _19095_;
  wire _19096_;
  wire _19097_;
  wire _19098_;
  wire _19099_;
  wire _19100_;
  wire _19101_;
  wire _19102_;
  wire _19103_;
  wire _19104_;
  wire _19105_;
  wire _19106_;
  wire _19107_;
  wire _19108_;
  wire _19109_;
  wire _19110_;
  wire _19111_;
  wire _19112_;
  wire _19113_;
  wire _19114_;
  wire _19115_;
  wire _19116_;
  wire _19117_;
  wire _19118_;
  wire _19119_;
  wire _19120_;
  wire _19121_;
  wire _19122_;
  wire _19123_;
  wire _19124_;
  wire _19125_;
  wire _19126_;
  wire _19127_;
  wire _19128_;
  wire _19129_;
  wire _19130_;
  wire _19131_;
  wire _19132_;
  wire _19133_;
  wire _19134_;
  wire _19135_;
  wire _19136_;
  wire _19137_;
  wire _19138_;
  wire _19139_;
  wire _19140_;
  wire _19141_;
  wire _19142_;
  wire _19143_;
  wire _19144_;
  wire _19145_;
  wire _19146_;
  wire _19147_;
  wire _19148_;
  wire _19149_;
  wire _19150_;
  wire _19151_;
  wire _19152_;
  wire _19153_;
  wire _19154_;
  wire _19155_;
  wire _19156_;
  wire _19157_;
  wire _19158_;
  wire _19159_;
  wire _19160_;
  wire _19161_;
  wire _19162_;
  wire _19163_;
  wire _19164_;
  wire _19165_;
  wire _19166_;
  wire _19167_;
  wire _19168_;
  wire _19169_;
  wire _19170_;
  wire _19171_;
  wire _19172_;
  wire _19173_;
  wire _19174_;
  wire _19175_;
  wire _19176_;
  wire _19177_;
  wire _19178_;
  wire _19179_;
  wire _19180_;
  wire _19181_;
  wire _19182_;
  wire _19183_;
  wire _19184_;
  wire _19185_;
  wire _19186_;
  wire _19187_;
  wire _19188_;
  wire _19189_;
  wire _19190_;
  wire _19191_;
  wire _19192_;
  wire _19193_;
  wire _19194_;
  wire _19195_;
  wire _19196_;
  wire _19197_;
  wire _19198_;
  wire _19199_;
  wire _19200_;
  wire _19201_;
  wire _19202_;
  wire _19203_;
  wire _19204_;
  wire _19205_;
  wire _19206_;
  wire _19207_;
  wire _19208_;
  wire _19209_;
  wire _19210_;
  wire _19211_;
  wire _19212_;
  wire _19213_;
  wire _19214_;
  wire _19215_;
  wire _19216_;
  wire _19217_;
  wire _19218_;
  wire _19219_;
  wire _19220_;
  wire _19221_;
  wire _19222_;
  wire _19223_;
  wire _19224_;
  wire _19225_;
  wire _19226_;
  wire _19227_;
  wire _19228_;
  wire _19229_;
  wire _19230_;
  wire _19231_;
  wire _19232_;
  wire _19233_;
  wire _19234_;
  wire _19235_;
  wire _19236_;
  wire _19237_;
  wire _19238_;
  wire _19239_;
  wire _19240_;
  wire _19241_;
  wire _19242_;
  wire _19243_;
  wire _19244_;
  wire _19245_;
  wire _19246_;
  wire _19247_;
  wire _19248_;
  wire _19249_;
  wire _19250_;
  wire _19251_;
  wire _19252_;
  wire _19253_;
  wire _19254_;
  wire _19255_;
  wire _19256_;
  wire _19257_;
  wire _19258_;
  wire _19259_;
  wire _19260_;
  wire _19261_;
  wire _19262_;
  wire _19263_;
  wire _19264_;
  wire _19265_;
  wire _19266_;
  wire _19267_;
  wire _19268_;
  wire _19269_;
  wire _19270_;
  wire _19271_;
  wire _19272_;
  wire _19273_;
  wire _19274_;
  wire _19275_;
  wire _19276_;
  wire _19277_;
  wire _19278_;
  wire _19279_;
  wire _19280_;
  wire _19281_;
  wire _19282_;
  wire _19283_;
  wire _19284_;
  wire _19285_;
  wire _19286_;
  wire _19287_;
  wire _19288_;
  wire _19289_;
  wire _19290_;
  wire _19291_;
  wire _19292_;
  wire _19293_;
  wire _19294_;
  wire _19295_;
  wire _19296_;
  wire _19297_;
  wire _19298_;
  wire _19299_;
  wire _19300_;
  wire _19301_;
  wire _19302_;
  wire _19303_;
  wire _19304_;
  wire _19305_;
  wire _19306_;
  wire _19307_;
  wire _19308_;
  wire _19309_;
  wire _19310_;
  wire _19311_;
  wire _19312_;
  wire _19313_;
  wire _19314_;
  wire _19315_;
  wire _19316_;
  wire _19317_;
  wire _19318_;
  wire _19319_;
  wire _19320_;
  wire _19321_;
  wire _19322_;
  wire _19323_;
  wire _19324_;
  wire _19325_;
  wire _19326_;
  wire _19327_;
  wire _19328_;
  wire _19329_;
  wire _19330_;
  wire _19331_;
  wire _19332_;
  wire _19333_;
  wire _19334_;
  wire _19335_;
  wire _19336_;
  wire _19337_;
  wire _19338_;
  wire _19339_;
  wire _19340_;
  wire _19341_;
  wire _19342_;
  wire _19343_;
  wire _19344_;
  wire _19345_;
  wire _19346_;
  wire _19347_;
  wire _19348_;
  wire _19349_;
  wire _19350_;
  wire _19351_;
  wire _19352_;
  wire _19353_;
  wire _19354_;
  wire _19355_;
  wire _19356_;
  wire _19357_;
  wire _19358_;
  wire _19359_;
  wire _19360_;
  wire _19361_;
  wire _19362_;
  wire _19363_;
  wire _19364_;
  wire _19365_;
  wire _19366_;
  wire _19367_;
  wire _19368_;
  wire _19369_;
  wire _19370_;
  wire _19371_;
  wire _19372_;
  wire _19373_;
  wire _19374_;
  wire _19375_;
  wire _19376_;
  wire _19377_;
  wire _19378_;
  wire _19379_;
  wire _19380_;
  wire _19381_;
  wire _19382_;
  wire _19383_;
  wire _19384_;
  wire _19385_;
  wire _19386_;
  wire _19387_;
  wire _19388_;
  wire _19389_;
  wire _19390_;
  wire _19391_;
  wire _19392_;
  wire _19393_;
  wire _19394_;
  wire _19395_;
  wire _19396_;
  wire _19397_;
  wire _19398_;
  wire _19399_;
  wire _19400_;
  wire _19401_;
  wire _19402_;
  wire _19403_;
  wire _19404_;
  wire _19405_;
  wire _19406_;
  wire _19407_;
  wire _19408_;
  wire _19409_;
  wire _19410_;
  wire _19411_;
  wire _19412_;
  wire _19413_;
  wire _19414_;
  wire _19415_;
  wire _19416_;
  wire _19417_;
  wire _19418_;
  wire _19419_;
  wire _19420_;
  wire _19421_;
  wire _19422_;
  wire _19423_;
  wire _19424_;
  wire _19425_;
  wire _19426_;
  wire _19427_;
  wire _19428_;
  wire _19429_;
  wire _19430_;
  wire _19431_;
  wire _19432_;
  wire _19433_;
  wire _19434_;
  wire _19435_;
  wire _19436_;
  wire _19437_;
  wire _19438_;
  wire _19439_;
  wire _19440_;
  wire _19441_;
  wire _19442_;
  wire _19443_;
  wire _19444_;
  wire _19445_;
  wire _19446_;
  wire _19447_;
  wire _19448_;
  wire _19449_;
  wire _19450_;
  wire _19451_;
  wire _19452_;
  wire _19453_;
  wire _19454_;
  wire _19455_;
  wire _19456_;
  wire _19457_;
  wire _19458_;
  wire _19459_;
  wire _19460_;
  wire _19461_;
  wire _19462_;
  wire _19463_;
  wire _19464_;
  wire _19465_;
  wire _19466_;
  wire _19467_;
  wire _19468_;
  wire _19469_;
  wire _19470_;
  wire _19471_;
  wire _19472_;
  wire _19473_;
  wire _19474_;
  wire _19475_;
  wire _19476_;
  wire _19477_;
  wire _19478_;
  wire _19479_;
  wire _19480_;
  wire _19481_;
  wire _19482_;
  wire _19483_;
  wire _19484_;
  wire _19485_;
  wire _19486_;
  wire _19487_;
  wire _19488_;
  wire _19489_;
  wire _19490_;
  wire _19491_;
  wire _19492_;
  wire _19493_;
  wire _19494_;
  wire _19495_;
  wire _19496_;
  wire _19497_;
  wire _19498_;
  wire _19499_;
  wire _19500_;
  wire _19501_;
  wire _19502_;
  wire _19503_;
  wire _19504_;
  wire _19505_;
  wire _19506_;
  wire _19507_;
  wire _19508_;
  wire _19509_;
  wire _19510_;
  wire _19511_;
  wire _19512_;
  wire _19513_;
  wire _19514_;
  wire _19515_;
  wire _19516_;
  wire _19517_;
  wire _19518_;
  wire _19519_;
  wire _19520_;
  wire _19521_;
  wire _19522_;
  wire _19523_;
  wire _19524_;
  wire _19525_;
  wire _19526_;
  wire _19527_;
  wire _19528_;
  wire _19529_;
  wire _19530_;
  wire _19531_;
  wire _19532_;
  wire _19533_;
  wire _19534_;
  wire _19535_;
  wire _19536_;
  wire _19537_;
  wire _19538_;
  wire _19539_;
  wire _19540_;
  wire _19541_;
  wire _19542_;
  wire _19543_;
  wire _19544_;
  wire _19545_;
  wire _19546_;
  wire _19547_;
  wire _19548_;
  wire _19549_;
  wire _19550_;
  wire _19551_;
  wire _19552_;
  wire _19553_;
  wire _19554_;
  wire _19555_;
  wire _19556_;
  wire _19557_;
  wire _19558_;
  wire _19559_;
  wire _19560_;
  wire _19561_;
  wire _19562_;
  wire _19563_;
  wire _19564_;
  wire _19565_;
  wire _19566_;
  wire _19567_;
  wire _19568_;
  wire _19569_;
  wire _19570_;
  wire _19571_;
  wire _19572_;
  wire _19573_;
  wire _19574_;
  wire _19575_;
  wire _19576_;
  wire _19577_;
  wire _19578_;
  wire _19579_;
  wire _19580_;
  wire _19581_;
  wire _19582_;
  wire _19583_;
  wire _19584_;
  wire _19585_;
  wire _19586_;
  wire _19587_;
  wire _19588_;
  wire _19589_;
  wire _19590_;
  wire _19591_;
  wire _19592_;
  wire _19593_;
  wire _19594_;
  wire _19595_;
  wire _19596_;
  wire _19597_;
  wire _19598_;
  wire _19599_;
  wire _19600_;
  wire _19601_;
  wire _19602_;
  wire _19603_;
  wire _19604_;
  wire _19605_;
  wire _19606_;
  wire _19607_;
  wire _19608_;
  wire _19609_;
  wire _19610_;
  wire _19611_;
  wire _19612_;
  wire _19613_;
  wire _19614_;
  wire _19615_;
  wire _19616_;
  wire _19617_;
  wire _19618_;
  wire _19619_;
  wire _19620_;
  wire _19621_;
  wire _19622_;
  wire _19623_;
  wire _19624_;
  wire _19625_;
  wire _19626_;
  wire _19627_;
  wire _19628_;
  wire _19629_;
  wire _19630_;
  wire _19631_;
  wire _19632_;
  wire _19633_;
  wire _19634_;
  wire _19635_;
  wire _19636_;
  wire _19637_;
  wire _19638_;
  wire _19639_;
  wire _19640_;
  wire _19641_;
  wire _19642_;
  wire _19643_;
  wire _19644_;
  wire _19645_;
  wire _19646_;
  wire _19647_;
  wire _19648_;
  wire _19649_;
  wire _19650_;
  wire _19651_;
  wire _19652_;
  wire _19653_;
  wire _19654_;
  wire _19655_;
  wire _19656_;
  wire _19657_;
  wire _19658_;
  wire _19659_;
  wire _19660_;
  wire _19661_;
  wire _19662_;
  wire _19663_;
  wire _19664_;
  wire _19665_;
  wire _19666_;
  wire _19667_;
  wire _19668_;
  wire _19669_;
  wire _19670_;
  wire _19671_;
  wire _19672_;
  wire _19673_;
  wire _19674_;
  wire _19675_;
  wire _19676_;
  wire _19677_;
  wire _19678_;
  wire _19679_;
  wire _19680_;
  wire _19681_;
  wire _19682_;
  wire _19683_;
  wire _19684_;
  wire _19685_;
  wire _19686_;
  wire _19687_;
  wire _19688_;
  wire _19689_;
  wire _19690_;
  wire _19691_;
  wire _19692_;
  wire _19693_;
  wire _19694_;
  wire _19695_;
  wire _19696_;
  wire _19697_;
  wire _19698_;
  wire _19699_;
  wire _19700_;
  wire _19701_;
  wire _19702_;
  wire _19703_;
  wire _19704_;
  wire _19705_;
  wire _19706_;
  wire _19707_;
  wire _19708_;
  wire _19709_;
  wire _19710_;
  wire _19711_;
  wire _19712_;
  wire _19713_;
  wire _19714_;
  wire _19715_;
  wire _19716_;
  wire _19717_;
  wire _19718_;
  wire _19719_;
  wire _19720_;
  wire _19721_;
  wire _19722_;
  wire _19723_;
  wire _19724_;
  wire _19725_;
  wire _19726_;
  wire _19727_;
  wire _19728_;
  wire _19729_;
  wire _19730_;
  wire _19731_;
  wire _19732_;
  wire _19733_;
  wire _19734_;
  wire _19735_;
  wire _19736_;
  wire _19737_;
  wire _19738_;
  wire _19739_;
  wire _19740_;
  wire _19741_;
  wire _19742_;
  wire _19743_;
  wire _19744_;
  wire _19745_;
  wire _19746_;
  wire _19747_;
  wire _19748_;
  wire _19749_;
  wire _19750_;
  wire _19751_;
  wire _19752_;
  wire _19753_;
  wire _19754_;
  wire _19755_;
  wire _19756_;
  wire _19757_;
  wire _19758_;
  wire _19759_;
  wire _19760_;
  wire _19761_;
  wire _19762_;
  wire _19763_;
  wire _19764_;
  wire _19765_;
  wire _19766_;
  wire _19767_;
  wire _19768_;
  wire _19769_;
  wire _19770_;
  wire _19771_;
  wire _19772_;
  wire _19773_;
  wire _19774_;
  wire _19775_;
  wire _19776_;
  wire _19777_;
  wire _19778_;
  wire _19779_;
  wire _19780_;
  wire _19781_;
  wire _19782_;
  wire _19783_;
  wire _19784_;
  wire _19785_;
  wire _19786_;
  wire _19787_;
  wire _19788_;
  wire _19789_;
  wire _19790_;
  wire _19791_;
  wire _19792_;
  wire _19793_;
  wire _19794_;
  wire _19795_;
  wire _19796_;
  wire _19797_;
  wire _19798_;
  wire _19799_;
  wire _19800_;
  wire _19801_;
  wire _19802_;
  wire _19803_;
  wire _19804_;
  wire _19805_;
  wire _19806_;
  wire _19807_;
  wire _19808_;
  wire _19809_;
  wire _19810_;
  wire _19811_;
  wire _19812_;
  wire _19813_;
  wire _19814_;
  wire _19815_;
  wire _19816_;
  wire _19817_;
  wire _19818_;
  wire _19819_;
  wire _19820_;
  wire _19821_;
  wire _19822_;
  wire _19823_;
  wire _19824_;
  wire _19825_;
  wire _19826_;
  wire _19827_;
  wire _19828_;
  wire _19829_;
  wire _19830_;
  wire _19831_;
  wire _19832_;
  wire _19833_;
  wire _19834_;
  wire _19835_;
  wire _19836_;
  wire _19837_;
  wire _19838_;
  wire _19839_;
  wire _19840_;
  wire _19841_;
  wire _19842_;
  wire _19843_;
  wire _19844_;
  wire _19845_;
  wire _19846_;
  wire _19847_;
  wire _19848_;
  wire _19849_;
  wire _19850_;
  wire _19851_;
  wire _19852_;
  wire _19853_;
  wire _19854_;
  wire _19855_;
  wire _19856_;
  wire _19857_;
  wire _19858_;
  wire _19859_;
  wire _19860_;
  wire _19861_;
  wire _19862_;
  wire _19863_;
  wire _19864_;
  wire _19865_;
  wire _19866_;
  wire _19867_;
  wire _19868_;
  wire _19869_;
  wire _19870_;
  wire _19871_;
  wire _19872_;
  wire _19873_;
  wire _19874_;
  wire _19875_;
  wire _19876_;
  wire _19877_;
  wire _19878_;
  wire _19879_;
  wire _19880_;
  wire _19881_;
  wire _19882_;
  wire _19883_;
  wire _19884_;
  wire _19885_;
  wire _19886_;
  wire _19887_;
  wire _19888_;
  wire _19889_;
  wire _19890_;
  wire _19891_;
  wire _19892_;
  wire _19893_;
  wire _19894_;
  wire _19895_;
  wire _19896_;
  wire _19897_;
  wire _19898_;
  wire _19899_;
  wire _19900_;
  wire _19901_;
  wire _19902_;
  wire _19903_;
  wire _19904_;
  wire _19905_;
  wire _19906_;
  wire _19907_;
  wire _19908_;
  wire _19909_;
  wire _19910_;
  wire _19911_;
  wire _19912_;
  wire _19913_;
  wire _19914_;
  wire _19915_;
  wire _19916_;
  wire _19917_;
  wire _19918_;
  wire _19919_;
  wire _19920_;
  wire _19921_;
  wire _19922_;
  wire _19923_;
  wire _19924_;
  wire _19925_;
  wire _19926_;
  wire _19927_;
  wire _19928_;
  wire _19929_;
  wire _19930_;
  wire _19931_;
  wire _19932_;
  wire _19933_;
  wire _19934_;
  wire _19935_;
  wire _19936_;
  wire _19937_;
  wire _19938_;
  wire _19939_;
  wire _19940_;
  wire _19941_;
  wire _19942_;
  wire _19943_;
  wire _19944_;
  wire _19945_;
  wire _19946_;
  wire _19947_;
  wire _19948_;
  wire _19949_;
  wire _19950_;
  wire _19951_;
  wire _19952_;
  wire _19953_;
  wire _19954_;
  wire _19955_;
  wire _19956_;
  wire _19957_;
  wire _19958_;
  wire _19959_;
  wire _19960_;
  wire _19961_;
  wire _19962_;
  wire _19963_;
  wire _19964_;
  wire _19965_;
  wire _19966_;
  wire _19967_;
  wire _19968_;
  wire _19969_;
  wire _19970_;
  wire _19971_;
  wire _19972_;
  wire _19973_;
  wire _19974_;
  wire _19975_;
  wire _19976_;
  wire _19977_;
  wire _19978_;
  wire _19979_;
  wire _19980_;
  wire _19981_;
  wire _19982_;
  wire _19983_;
  wire _19984_;
  wire _19985_;
  wire _19986_;
  wire _19987_;
  wire _19988_;
  wire _19989_;
  wire _19990_;
  wire _19991_;
  wire _19992_;
  wire _19993_;
  wire _19994_;
  wire _19995_;
  wire _19996_;
  wire _19997_;
  wire _19998_;
  wire _19999_;
  wire _20000_;
  wire _20001_;
  wire _20002_;
  wire _20003_;
  wire _20004_;
  wire _20005_;
  wire _20006_;
  wire _20007_;
  wire _20008_;
  wire _20009_;
  wire _20010_;
  wire _20011_;
  wire _20012_;
  wire _20013_;
  wire _20014_;
  wire _20015_;
  wire _20016_;
  wire _20017_;
  wire _20018_;
  wire _20019_;
  wire _20020_;
  wire _20021_;
  wire _20022_;
  wire _20023_;
  wire _20024_;
  wire _20025_;
  wire _20026_;
  wire _20027_;
  wire _20028_;
  wire _20029_;
  wire _20030_;
  wire _20031_;
  wire _20032_;
  wire _20033_;
  wire _20034_;
  wire _20035_;
  wire _20036_;
  wire _20037_;
  wire _20038_;
  wire _20039_;
  wire _20040_;
  wire _20041_;
  wire _20042_;
  wire _20043_;
  wire _20044_;
  wire _20045_;
  wire _20046_;
  wire _20047_;
  wire _20048_;
  wire _20049_;
  wire _20050_;
  wire _20051_;
  wire _20052_;
  wire _20053_;
  wire _20054_;
  wire _20055_;
  wire _20056_;
  wire _20057_;
  wire _20058_;
  wire _20059_;
  wire _20060_;
  wire _20061_;
  wire _20062_;
  wire _20063_;
  wire _20064_;
  wire _20065_;
  wire _20066_;
  wire _20067_;
  wire _20068_;
  wire _20069_;
  wire _20070_;
  wire _20071_;
  wire _20072_;
  wire _20073_;
  wire _20074_;
  wire _20075_;
  wire _20076_;
  wire _20077_;
  wire _20078_;
  wire _20079_;
  wire _20080_;
  wire _20081_;
  wire _20082_;
  wire _20083_;
  wire _20084_;
  wire _20085_;
  wire _20086_;
  wire _20087_;
  wire _20088_;
  wire _20089_;
  wire _20090_;
  wire _20091_;
  wire _20092_;
  wire _20093_;
  wire _20094_;
  wire _20095_;
  wire _20096_;
  wire _20097_;
  wire _20098_;
  wire _20099_;
  wire _20100_;
  wire _20101_;
  wire _20102_;
  wire _20103_;
  wire _20104_;
  wire _20105_;
  wire _20106_;
  wire _20107_;
  wire _20108_;
  wire _20109_;
  wire _20110_;
  wire _20111_;
  wire _20112_;
  wire _20113_;
  wire _20114_;
  wire _20115_;
  wire _20116_;
  wire _20117_;
  wire _20118_;
  wire _20119_;
  wire _20120_;
  wire _20121_;
  wire _20122_;
  wire _20123_;
  wire _20124_;
  wire _20125_;
  wire _20126_;
  wire _20127_;
  wire _20128_;
  wire _20129_;
  wire _20130_;
  wire _20131_;
  wire _20132_;
  wire _20133_;
  wire _20134_;
  wire _20135_;
  wire _20136_;
  wire _20137_;
  wire _20138_;
  wire _20139_;
  wire _20140_;
  wire _20141_;
  wire _20142_;
  wire _20143_;
  wire _20144_;
  wire _20145_;
  wire _20146_;
  wire _20147_;
  wire _20148_;
  wire _20149_;
  wire _20150_;
  wire _20151_;
  wire _20152_;
  wire _20153_;
  wire _20154_;
  wire _20155_;
  wire _20156_;
  wire _20157_;
  wire _20158_;
  wire _20159_;
  wire _20160_;
  wire _20161_;
  wire _20162_;
  wire _20163_;
  wire _20164_;
  wire _20165_;
  wire _20166_;
  wire _20167_;
  wire _20168_;
  wire _20169_;
  wire _20170_;
  wire _20171_;
  wire _20172_;
  wire _20173_;
  wire _20174_;
  wire _20175_;
  wire _20176_;
  wire _20177_;
  wire _20178_;
  wire _20179_;
  wire _20180_;
  wire _20181_;
  wire _20182_;
  wire _20183_;
  wire _20184_;
  wire _20185_;
  wire _20186_;
  wire _20187_;
  wire _20188_;
  wire _20189_;
  wire _20190_;
  wire _20191_;
  wire _20192_;
  wire _20193_;
  wire _20194_;
  wire _20195_;
  wire _20196_;
  wire _20197_;
  wire _20198_;
  wire _20199_;
  wire _20200_;
  wire _20201_;
  wire _20202_;
  wire _20203_;
  wire _20204_;
  wire _20205_;
  wire _20206_;
  wire _20207_;
  wire _20208_;
  wire _20209_;
  wire _20210_;
  wire _20211_;
  wire _20212_;
  wire _20213_;
  wire _20214_;
  wire _20215_;
  wire _20216_;
  wire _20217_;
  wire _20218_;
  wire _20219_;
  wire _20220_;
  wire _20221_;
  wire _20222_;
  wire _20223_;
  wire _20224_;
  wire _20225_;
  wire _20226_;
  wire _20227_;
  wire _20228_;
  wire _20229_;
  wire _20230_;
  wire _20231_;
  wire _20232_;
  wire _20233_;
  wire _20234_;
  wire _20235_;
  wire _20236_;
  wire _20237_;
  wire _20238_;
  wire _20239_;
  wire _20240_;
  wire _20241_;
  wire _20242_;
  wire _20243_;
  wire _20244_;
  wire _20245_;
  wire _20246_;
  wire _20247_;
  wire _20248_;
  wire _20249_;
  wire _20250_;
  wire _20251_;
  wire _20252_;
  wire _20253_;
  wire _20254_;
  wire _20255_;
  wire _20256_;
  wire _20257_;
  wire _20258_;
  wire _20259_;
  wire _20260_;
  wire _20261_;
  wire _20262_;
  wire _20263_;
  wire _20264_;
  wire _20265_;
  wire _20266_;
  wire _20267_;
  wire _20268_;
  wire _20269_;
  wire _20270_;
  wire _20271_;
  wire _20272_;
  wire _20273_;
  wire _20274_;
  wire _20275_;
  wire _20276_;
  wire _20277_;
  wire _20278_;
  wire _20279_;
  wire _20280_;
  wire _20281_;
  wire _20282_;
  wire _20283_;
  wire _20284_;
  wire _20285_;
  wire _20286_;
  wire _20287_;
  wire _20288_;
  wire _20289_;
  wire _20290_;
  wire _20291_;
  wire _20292_;
  wire _20293_;
  wire _20294_;
  wire _20295_;
  wire _20296_;
  wire _20297_;
  wire _20298_;
  wire _20299_;
  wire _20300_;
  wire _20301_;
  wire _20302_;
  wire _20303_;
  wire _20304_;
  wire _20305_;
  wire _20306_;
  wire _20307_;
  wire _20308_;
  wire _20309_;
  wire _20310_;
  wire _20311_;
  wire _20312_;
  wire _20313_;
  wire _20314_;
  wire _20315_;
  wire _20316_;
  wire _20317_;
  wire _20318_;
  wire _20319_;
  wire _20320_;
  wire _20321_;
  wire _20322_;
  wire _20323_;
  wire _20324_;
  wire _20325_;
  wire _20326_;
  wire _20327_;
  wire _20328_;
  wire _20329_;
  wire _20330_;
  wire _20331_;
  wire _20332_;
  wire _20333_;
  wire _20334_;
  wire _20335_;
  wire _20336_;
  wire _20337_;
  wire _20338_;
  wire _20339_;
  wire _20340_;
  wire _20341_;
  wire _20342_;
  wire _20343_;
  wire _20344_;
  wire _20345_;
  wire _20346_;
  wire _20347_;
  wire _20348_;
  wire _20349_;
  wire _20350_;
  wire _20351_;
  wire _20352_;
  wire _20353_;
  wire _20354_;
  wire _20355_;
  wire _20356_;
  wire _20357_;
  wire _20358_;
  wire _20359_;
  wire _20360_;
  wire _20361_;
  wire _20362_;
  wire _20363_;
  wire _20364_;
  wire _20365_;
  wire _20366_;
  wire _20367_;
  wire _20368_;
  wire _20369_;
  wire _20370_;
  wire _20371_;
  wire _20372_;
  wire _20373_;
  wire _20374_;
  wire _20375_;
  wire _20376_;
  wire _20377_;
  wire _20378_;
  wire _20379_;
  wire _20380_;
  wire _20381_;
  wire _20382_;
  wire _20383_;
  wire _20384_;
  wire _20385_;
  wire _20386_;
  wire _20387_;
  wire _20388_;
  wire _20389_;
  wire _20390_;
  wire _20391_;
  wire _20392_;
  wire _20393_;
  wire _20394_;
  wire _20395_;
  wire _20396_;
  wire _20397_;
  wire _20398_;
  wire _20399_;
  wire _20400_;
  wire _20401_;
  wire _20402_;
  wire _20403_;
  wire _20404_;
  wire _20405_;
  wire _20406_;
  wire _20407_;
  wire _20408_;
  wire _20409_;
  wire _20410_;
  wire _20411_;
  wire _20412_;
  wire _20413_;
  wire _20414_;
  wire _20415_;
  wire _20416_;
  wire _20417_;
  wire _20418_;
  wire _20419_;
  wire _20420_;
  wire _20421_;
  wire _20422_;
  wire _20423_;
  wire _20424_;
  wire _20425_;
  wire _20426_;
  wire _20427_;
  wire _20428_;
  wire _20429_;
  wire _20430_;
  wire _20431_;
  wire _20432_;
  wire _20433_;
  wire _20434_;
  wire _20435_;
  wire _20436_;
  wire _20437_;
  wire _20438_;
  wire _20439_;
  wire _20440_;
  wire _20441_;
  wire _20442_;
  wire _20443_;
  wire _20444_;
  wire _20445_;
  wire _20446_;
  wire _20447_;
  wire _20448_;
  wire _20449_;
  wire _20450_;
  wire _20451_;
  wire _20452_;
  wire _20453_;
  wire _20454_;
  wire _20455_;
  wire _20456_;
  wire _20457_;
  wire _20458_;
  wire _20459_;
  wire _20460_;
  wire _20461_;
  wire _20462_;
  wire _20463_;
  wire _20464_;
  wire _20465_;
  wire _20466_;
  wire _20467_;
  wire _20468_;
  wire _20469_;
  wire _20470_;
  wire _20471_;
  wire _20472_;
  wire _20473_;
  wire _20474_;
  wire _20475_;
  wire _20476_;
  wire _20477_;
  wire _20478_;
  wire _20479_;
  wire _20480_;
  wire _20481_;
  wire _20482_;
  wire _20483_;
  wire _20484_;
  wire _20485_;
  wire _20486_;
  wire _20487_;
  wire _20488_;
  wire _20489_;
  wire _20490_;
  wire _20491_;
  wire _20492_;
  wire _20493_;
  wire _20494_;
  wire _20495_;
  wire _20496_;
  wire _20497_;
  wire _20498_;
  wire _20499_;
  wire _20500_;
  wire _20501_;
  wire _20502_;
  wire _20503_;
  wire _20504_;
  wire _20505_;
  wire _20506_;
  wire _20507_;
  wire _20508_;
  wire _20509_;
  wire _20510_;
  wire _20511_;
  wire _20512_;
  wire _20513_;
  wire _20514_;
  wire _20515_;
  wire _20516_;
  wire _20517_;
  wire _20518_;
  wire _20519_;
  wire _20520_;
  wire _20521_;
  wire _20522_;
  wire _20523_;
  wire _20524_;
  wire _20525_;
  wire _20526_;
  wire _20527_;
  wire _20528_;
  wire _20529_;
  wire _20530_;
  wire _20531_;
  wire _20532_;
  wire _20533_;
  wire _20534_;
  wire _20535_;
  wire _20536_;
  wire _20537_;
  wire _20538_;
  wire _20539_;
  wire _20540_;
  wire _20541_;
  wire _20542_;
  wire _20543_;
  wire _20544_;
  wire _20545_;
  wire _20546_;
  wire _20547_;
  wire _20548_;
  wire _20549_;
  wire _20550_;
  wire _20551_;
  wire _20552_;
  wire _20553_;
  wire _20554_;
  wire _20555_;
  wire _20556_;
  wire _20557_;
  wire _20558_;
  wire _20559_;
  wire _20560_;
  wire _20561_;
  wire _20562_;
  wire _20563_;
  wire _20564_;
  wire _20565_;
  wire _20566_;
  wire _20567_;
  wire _20568_;
  wire _20569_;
  wire _20570_;
  wire _20571_;
  wire _20572_;
  wire _20573_;
  wire _20574_;
  wire _20575_;
  wire _20576_;
  wire _20577_;
  wire _20578_;
  wire _20579_;
  wire _20580_;
  wire _20581_;
  wire _20582_;
  wire _20583_;
  wire _20584_;
  wire _20585_;
  wire _20586_;
  wire _20587_;
  wire _20588_;
  wire _20589_;
  wire _20590_;
  wire _20591_;
  wire _20592_;
  wire _20593_;
  wire _20594_;
  wire _20595_;
  wire _20596_;
  wire _20597_;
  wire _20598_;
  wire _20599_;
  wire _20600_;
  wire _20601_;
  wire _20602_;
  wire _20603_;
  wire _20604_;
  wire _20605_;
  wire _20606_;
  wire _20607_;
  wire _20608_;
  wire _20609_;
  wire _20610_;
  wire _20611_;
  wire _20612_;
  wire _20613_;
  wire _20614_;
  wire _20615_;
  wire _20616_;
  wire _20617_;
  wire _20618_;
  wire _20619_;
  wire _20620_;
  wire _20621_;
  wire _20622_;
  wire _20623_;
  wire _20624_;
  wire _20625_;
  wire _20626_;
  wire _20627_;
  wire _20628_;
  wire _20629_;
  wire _20630_;
  wire _20631_;
  wire _20632_;
  wire _20633_;
  wire _20634_;
  wire _20635_;
  wire _20636_;
  wire _20637_;
  wire _20638_;
  wire _20639_;
  wire _20640_;
  wire _20641_;
  wire _20642_;
  wire _20643_;
  wire _20644_;
  wire _20645_;
  wire _20646_;
  wire _20647_;
  wire _20648_;
  wire _20649_;
  wire _20650_;
  wire _20651_;
  wire _20652_;
  wire _20653_;
  wire _20654_;
  wire _20655_;
  wire _20656_;
  wire _20657_;
  wire _20658_;
  wire _20659_;
  wire _20660_;
  wire _20661_;
  wire _20662_;
  wire _20663_;
  wire _20664_;
  wire _20665_;
  wire _20666_;
  wire _20667_;
  wire _20668_;
  wire _20669_;
  wire _20670_;
  wire _20671_;
  wire _20672_;
  wire _20673_;
  wire _20674_;
  wire _20675_;
  wire _20676_;
  wire _20677_;
  wire _20678_;
  wire _20679_;
  wire _20680_;
  wire _20681_;
  wire _20682_;
  wire _20683_;
  wire _20684_;
  wire _20685_;
  wire _20686_;
  wire _20687_;
  wire _20688_;
  wire _20689_;
  wire _20690_;
  wire _20691_;
  wire _20692_;
  wire _20693_;
  wire _20694_;
  wire _20695_;
  wire _20696_;
  wire _20697_;
  wire _20698_;
  wire _20699_;
  wire _20700_;
  wire _20701_;
  wire _20702_;
  wire _20703_;
  wire _20704_;
  wire _20705_;
  wire _20706_;
  wire _20707_;
  wire _20708_;
  wire _20709_;
  wire _20710_;
  wire _20711_;
  wire _20712_;
  wire _20713_;
  wire _20714_;
  wire _20715_;
  wire _20716_;
  wire _20717_;
  wire _20718_;
  wire _20719_;
  wire _20720_;
  wire _20721_;
  wire _20722_;
  wire _20723_;
  wire _20724_;
  wire _20725_;
  wire _20726_;
  wire _20727_;
  wire _20728_;
  wire _20729_;
  wire _20730_;
  wire _20731_;
  wire _20732_;
  wire _20733_;
  wire _20734_;
  wire _20735_;
  wire _20736_;
  wire _20737_;
  wire _20738_;
  wire _20739_;
  wire _20740_;
  wire _20741_;
  wire _20742_;
  wire _20743_;
  wire _20744_;
  wire _20745_;
  wire _20746_;
  wire _20747_;
  wire _20748_;
  wire _20749_;
  wire _20750_;
  wire _20751_;
  wire _20752_;
  wire _20753_;
  wire _20754_;
  wire _20755_;
  wire _20756_;
  wire _20757_;
  wire _20758_;
  wire _20759_;
  wire _20760_;
  wire _20761_;
  wire _20762_;
  wire _20763_;
  wire _20764_;
  wire _20765_;
  wire _20766_;
  wire _20767_;
  wire _20768_;
  wire _20769_;
  wire _20770_;
  wire _20771_;
  wire _20772_;
  wire _20773_;
  wire _20774_;
  wire _20775_;
  wire _20776_;
  wire _20777_;
  wire _20778_;
  wire _20779_;
  wire _20780_;
  wire _20781_;
  wire _20782_;
  wire _20783_;
  wire _20784_;
  wire _20785_;
  wire _20786_;
  wire _20787_;
  wire _20788_;
  wire _20789_;
  wire _20790_;
  wire _20791_;
  wire _20792_;
  wire _20793_;
  wire _20794_;
  wire _20795_;
  wire _20796_;
  wire _20797_;
  wire _20798_;
  wire _20799_;
  wire _20800_;
  wire _20801_;
  wire _20802_;
  wire _20803_;
  wire _20804_;
  wire _20805_;
  wire _20806_;
  wire _20807_;
  wire _20808_;
  wire _20809_;
  wire _20810_;
  wire _20811_;
  wire _20812_;
  wire _20813_;
  wire _20814_;
  wire _20815_;
  wire _20816_;
  wire _20817_;
  wire _20818_;
  wire _20819_;
  wire _20820_;
  wire _20821_;
  wire _20822_;
  wire _20823_;
  wire _20824_;
  wire _20825_;
  wire _20826_;
  wire _20827_;
  wire _20828_;
  wire _20829_;
  wire _20830_;
  wire _20831_;
  wire _20832_;
  wire _20833_;
  wire _20834_;
  wire _20835_;
  wire _20836_;
  wire _20837_;
  wire _20838_;
  wire _20839_;
  wire _20840_;
  wire _20841_;
  wire _20842_;
  wire _20843_;
  wire _20844_;
  wire _20845_;
  wire _20846_;
  wire _20847_;
  wire _20848_;
  wire _20849_;
  wire _20850_;
  wire _20851_;
  wire _20852_;
  wire _20853_;
  wire _20854_;
  wire _20855_;
  wire _20856_;
  wire _20857_;
  wire _20858_;
  wire _20859_;
  wire _20860_;
  wire _20861_;
  wire _20862_;
  wire _20863_;
  wire _20864_;
  wire _20865_;
  wire _20866_;
  wire _20867_;
  wire _20868_;
  wire _20869_;
  wire _20870_;
  wire _20871_;
  wire _20872_;
  wire _20873_;
  wire _20874_;
  wire _20875_;
  wire _20876_;
  wire _20877_;
  wire _20878_;
  wire _20879_;
  wire _20880_;
  wire _20881_;
  wire _20882_;
  wire _20883_;
  wire _20884_;
  wire _20885_;
  wire _20886_;
  wire _20887_;
  wire _20888_;
  wire _20889_;
  wire _20890_;
  wire _20891_;
  wire _20892_;
  wire _20893_;
  wire _20894_;
  wire _20895_;
  wire _20896_;
  wire _20897_;
  wire _20898_;
  wire _20899_;
  wire _20900_;
  wire _20901_;
  wire _20902_;
  wire _20903_;
  wire _20904_;
  wire _20905_;
  wire _20906_;
  wire _20907_;
  wire _20908_;
  wire _20909_;
  wire _20910_;
  wire _20911_;
  wire _20912_;
  wire _20913_;
  wire _20914_;
  wire _20915_;
  wire _20916_;
  wire _20917_;
  wire _20918_;
  wire _20919_;
  wire _20920_;
  wire _20921_;
  wire _20922_;
  wire _20923_;
  wire _20924_;
  wire _20925_;
  wire _20926_;
  wire _20927_;
  wire _20928_;
  wire _20929_;
  wire _20930_;
  wire _20931_;
  wire _20932_;
  wire _20933_;
  wire _20934_;
  wire _20935_;
  wire _20936_;
  wire _20937_;
  wire _20938_;
  wire _20939_;
  wire _20940_;
  wire _20941_;
  wire _20942_;
  wire _20943_;
  wire _20944_;
  wire _20945_;
  wire _20946_;
  wire _20947_;
  wire _20948_;
  wire _20949_;
  wire _20950_;
  wire _20951_;
  wire _20952_;
  wire _20953_;
  wire _20954_;
  wire _20955_;
  wire _20956_;
  wire _20957_;
  wire _20958_;
  wire _20959_;
  wire _20960_;
  wire _20961_;
  wire _20962_;
  wire _20963_;
  wire _20964_;
  wire _20965_;
  wire _20966_;
  wire _20967_;
  wire _20968_;
  wire _20969_;
  wire _20970_;
  wire _20971_;
  wire _20972_;
  wire _20973_;
  wire _20974_;
  wire _20975_;
  wire _20976_;
  wire _20977_;
  wire _20978_;
  wire _20979_;
  wire _20980_;
  wire _20981_;
  wire _20982_;
  wire _20983_;
  wire _20984_;
  wire _20985_;
  wire _20986_;
  wire _20987_;
  wire _20988_;
  wire _20989_;
  wire _20990_;
  wire _20991_;
  wire _20992_;
  wire _20993_;
  wire _20994_;
  wire _20995_;
  wire _20996_;
  wire _20997_;
  wire _20998_;
  wire _20999_;
  wire _21000_;
  wire _21001_;
  wire _21002_;
  wire _21003_;
  wire _21004_;
  wire _21005_;
  wire _21006_;
  wire _21007_;
  wire _21008_;
  wire _21009_;
  wire _21010_;
  wire _21011_;
  wire _21012_;
  wire _21013_;
  wire _21014_;
  wire _21015_;
  wire _21016_;
  wire _21017_;
  wire _21018_;
  wire _21019_;
  wire _21020_;
  wire _21021_;
  wire _21022_;
  wire _21023_;
  wire _21024_;
  wire _21025_;
  wire _21026_;
  wire _21027_;
  wire _21028_;
  wire _21029_;
  wire _21030_;
  wire _21031_;
  wire _21032_;
  wire _21033_;
  wire _21034_;
  wire _21035_;
  wire _21036_;
  wire _21037_;
  wire _21038_;
  wire _21039_;
  wire _21040_;
  wire _21041_;
  wire _21042_;
  wire _21043_;
  wire _21044_;
  wire _21045_;
  wire _21046_;
  wire _21047_;
  wire _21048_;
  wire _21049_;
  wire _21050_;
  wire _21051_;
  wire _21052_;
  wire _21053_;
  wire _21054_;
  wire _21055_;
  wire _21056_;
  wire _21057_;
  wire _21058_;
  wire _21059_;
  wire _21060_;
  wire _21061_;
  wire _21062_;
  wire _21063_;
  wire _21064_;
  wire _21065_;
  wire _21066_;
  wire _21067_;
  wire _21068_;
  wire _21069_;
  wire _21070_;
  wire _21071_;
  wire _21072_;
  wire _21073_;
  wire _21074_;
  wire _21075_;
  wire _21076_;
  wire _21077_;
  wire _21078_;
  wire _21079_;
  wire _21080_;
  wire _21081_;
  wire _21082_;
  wire _21083_;
  wire _21084_;
  wire _21085_;
  wire _21086_;
  wire _21087_;
  wire _21088_;
  wire _21089_;
  wire _21090_;
  wire _21091_;
  wire _21092_;
  wire _21093_;
  wire _21094_;
  wire _21095_;
  wire _21096_;
  wire _21097_;
  wire _21098_;
  wire _21099_;
  wire _21100_;
  wire _21101_;
  wire _21102_;
  wire _21103_;
  wire _21104_;
  wire _21105_;
  wire _21106_;
  wire _21107_;
  wire _21108_;
  wire _21109_;
  wire _21110_;
  wire _21111_;
  wire _21112_;
  wire _21113_;
  wire _21114_;
  wire _21115_;
  wire _21116_;
  wire _21117_;
  wire _21118_;
  wire _21119_;
  wire _21120_;
  wire _21121_;
  wire _21122_;
  wire _21123_;
  wire _21124_;
  wire _21125_;
  wire _21126_;
  wire _21127_;
  wire _21128_;
  wire _21129_;
  wire _21130_;
  wire _21131_;
  wire _21132_;
  wire _21133_;
  wire _21134_;
  wire _21135_;
  wire _21136_;
  wire _21137_;
  wire _21138_;
  wire _21139_;
  wire _21140_;
  wire _21141_;
  wire _21142_;
  wire _21143_;
  wire _21144_;
  wire _21145_;
  wire _21146_;
  wire _21147_;
  wire _21148_;
  wire _21149_;
  wire _21150_;
  wire _21151_;
  wire _21152_;
  wire _21153_;
  wire _21154_;
  wire _21155_;
  wire _21156_;
  wire _21157_;
  wire _21158_;
  wire _21159_;
  wire _21160_;
  wire _21161_;
  wire _21162_;
  wire _21163_;
  wire _21164_;
  wire _21165_;
  wire _21166_;
  wire _21167_;
  wire _21168_;
  wire _21169_;
  wire _21170_;
  wire _21171_;
  wire _21172_;
  wire _21173_;
  wire _21174_;
  wire _21175_;
  wire _21176_;
  wire _21177_;
  wire _21178_;
  wire _21179_;
  wire _21180_;
  wire _21181_;
  wire _21182_;
  wire _21183_;
  wire _21184_;
  wire _21185_;
  wire _21186_;
  wire _21187_;
  wire _21188_;
  wire _21189_;
  wire _21190_;
  wire _21191_;
  wire _21192_;
  wire _21193_;
  wire _21194_;
  wire _21195_;
  wire _21196_;
  wire _21197_;
  wire _21198_;
  wire _21199_;
  wire _21200_;
  wire _21201_;
  wire _21202_;
  wire _21203_;
  wire _21204_;
  wire _21205_;
  wire _21206_;
  wire _21207_;
  wire _21208_;
  wire _21209_;
  wire _21210_;
  wire _21211_;
  wire _21212_;
  wire _21213_;
  wire _21214_;
  wire _21215_;
  wire _21216_;
  wire _21217_;
  wire _21218_;
  wire _21219_;
  wire _21220_;
  wire _21221_;
  wire _21222_;
  wire _21223_;
  wire _21224_;
  wire _21225_;
  wire _21226_;
  wire _21227_;
  wire _21228_;
  wire _21229_;
  wire _21230_;
  wire _21231_;
  wire _21232_;
  wire _21233_;
  wire _21234_;
  wire _21235_;
  wire _21236_;
  wire _21237_;
  wire _21238_;
  wire _21239_;
  wire _21240_;
  wire _21241_;
  wire _21242_;
  wire _21243_;
  wire _21244_;
  wire _21245_;
  wire _21246_;
  wire _21247_;
  wire _21248_;
  wire _21249_;
  wire _21250_;
  wire _21251_;
  wire _21252_;
  wire _21253_;
  wire _21254_;
  wire _21255_;
  wire _21256_;
  wire _21257_;
  wire _21258_;
  wire _21259_;
  wire _21260_;
  wire _21261_;
  wire _21262_;
  wire _21263_;
  wire _21264_;
  wire _21265_;
  wire _21266_;
  wire _21267_;
  wire _21268_;
  wire _21269_;
  wire _21270_;
  wire _21271_;
  wire _21272_;
  wire _21273_;
  wire _21274_;
  wire _21275_;
  wire _21276_;
  wire _21277_;
  wire _21278_;
  wire _21279_;
  wire _21280_;
  wire _21281_;
  wire _21282_;
  wire _21283_;
  wire _21284_;
  wire _21285_;
  wire _21286_;
  wire _21287_;
  wire _21288_;
  wire _21289_;
  wire _21290_;
  wire _21291_;
  wire _21292_;
  wire _21293_;
  wire _21294_;
  wire _21295_;
  wire _21296_;
  wire _21297_;
  wire _21298_;
  wire _21299_;
  wire _21300_;
  wire _21301_;
  wire _21302_;
  wire _21303_;
  wire _21304_;
  wire _21305_;
  wire _21306_;
  wire _21307_;
  wire _21308_;
  wire _21309_;
  wire _21310_;
  wire _21311_;
  wire _21312_;
  wire _21313_;
  wire _21314_;
  wire _21315_;
  wire _21316_;
  wire _21317_;
  wire _21318_;
  wire _21319_;
  wire _21320_;
  wire _21321_;
  wire _21322_;
  wire _21323_;
  wire _21324_;
  wire _21325_;
  wire _21326_;
  wire _21327_;
  wire _21328_;
  wire _21329_;
  wire _21330_;
  wire _21331_;
  wire _21332_;
  wire _21333_;
  wire _21334_;
  wire _21335_;
  wire _21336_;
  wire _21337_;
  wire _21338_;
  wire _21339_;
  wire _21340_;
  wire _21341_;
  wire _21342_;
  wire _21343_;
  wire _21344_;
  wire _21345_;
  wire _21346_;
  wire _21347_;
  wire _21348_;
  wire _21349_;
  wire _21350_;
  wire _21351_;
  wire _21352_;
  wire _21353_;
  wire _21354_;
  wire _21355_;
  wire _21356_;
  wire _21357_;
  wire _21358_;
  wire _21359_;
  wire _21360_;
  wire _21361_;
  wire _21362_;
  wire _21363_;
  wire _21364_;
  wire _21365_;
  wire _21366_;
  wire _21367_;
  wire _21368_;
  wire _21369_;
  wire _21370_;
  wire _21371_;
  wire _21372_;
  wire _21373_;
  wire _21374_;
  wire _21375_;
  wire _21376_;
  wire _21377_;
  wire _21378_;
  wire _21379_;
  wire _21380_;
  wire _21381_;
  wire _21382_;
  wire _21383_;
  wire _21384_;
  wire _21385_;
  wire _21386_;
  wire _21387_;
  wire _21388_;
  wire _21389_;
  wire _21390_;
  wire _21391_;
  wire _21392_;
  wire _21393_;
  wire _21394_;
  wire _21395_;
  wire _21396_;
  wire _21397_;
  wire _21398_;
  wire _21399_;
  wire _21400_;
  wire _21401_;
  wire _21402_;
  wire _21403_;
  wire _21404_;
  wire _21405_;
  wire _21406_;
  wire _21407_;
  wire _21408_;
  wire _21409_;
  wire _21410_;
  wire _21411_;
  wire _21412_;
  wire _21413_;
  wire _21414_;
  wire _21415_;
  wire _21416_;
  wire _21417_;
  wire _21418_;
  wire _21419_;
  wire _21420_;
  wire _21421_;
  wire _21422_;
  wire _21423_;
  wire _21424_;
  wire _21425_;
  wire _21426_;
  wire _21427_;
  wire _21428_;
  wire _21429_;
  wire _21430_;
  wire _21431_;
  wire _21432_;
  wire _21433_;
  wire _21434_;
  wire _21435_;
  wire _21436_;
  wire _21437_;
  wire _21438_;
  wire _21439_;
  wire _21440_;
  wire _21441_;
  wire _21442_;
  wire _21443_;
  wire _21444_;
  wire _21445_;
  wire _21446_;
  wire _21447_;
  wire _21448_;
  wire _21449_;
  wire _21450_;
  wire _21451_;
  wire _21452_;
  wire _21453_;
  wire _21454_;
  wire _21455_;
  wire _21456_;
  wire _21457_;
  wire _21458_;
  wire _21459_;
  wire _21460_;
  wire _21461_;
  wire _21462_;
  wire _21463_;
  wire _21464_;
  wire _21465_;
  wire _21466_;
  wire _21467_;
  wire _21468_;
  wire _21469_;
  wire _21470_;
  wire _21471_;
  wire _21472_;
  wire _21473_;
  wire _21474_;
  wire _21475_;
  wire _21476_;
  wire _21477_;
  wire _21478_;
  wire _21479_;
  wire _21480_;
  wire _21481_;
  wire _21482_;
  wire _21483_;
  wire _21484_;
  wire _21485_;
  wire _21486_;
  wire _21487_;
  wire _21488_;
  wire _21489_;
  wire _21490_;
  wire _21491_;
  wire _21492_;
  wire _21493_;
  wire _21494_;
  wire _21495_;
  wire _21496_;
  wire _21497_;
  wire _21498_;
  wire _21499_;
  wire _21500_;
  wire _21501_;
  wire _21502_;
  wire _21503_;
  wire _21504_;
  wire _21505_;
  wire _21506_;
  wire _21507_;
  wire _21508_;
  wire _21509_;
  wire _21510_;
  wire _21511_;
  wire _21512_;
  wire _21513_;
  wire _21514_;
  wire _21515_;
  wire _21516_;
  wire _21517_;
  wire _21518_;
  wire _21519_;
  wire _21520_;
  wire _21521_;
  wire _21522_;
  wire _21523_;
  wire _21524_;
  wire _21525_;
  wire _21526_;
  wire _21527_;
  wire _21528_;
  wire _21529_;
  wire _21530_;
  wire _21531_;
  wire _21532_;
  wire _21533_;
  wire _21534_;
  wire _21535_;
  wire _21536_;
  wire _21537_;
  wire _21538_;
  wire _21539_;
  wire _21540_;
  wire _21541_;
  wire _21542_;
  wire _21543_;
  wire _21544_;
  wire _21545_;
  wire _21546_;
  wire _21547_;
  wire _21548_;
  wire _21549_;
  wire _21550_;
  wire _21551_;
  wire _21552_;
  wire _21553_;
  wire _21554_;
  wire _21555_;
  wire _21556_;
  wire _21557_;
  wire _21558_;
  wire _21559_;
  wire _21560_;
  wire _21561_;
  wire _21562_;
  wire _21563_;
  wire _21564_;
  wire _21565_;
  wire _21566_;
  wire _21567_;
  wire _21568_;
  wire _21569_;
  wire _21570_;
  wire _21571_;
  wire _21572_;
  wire _21573_;
  wire _21574_;
  wire _21575_;
  wire _21576_;
  wire _21577_;
  wire _21578_;
  wire _21579_;
  wire _21580_;
  wire _21581_;
  wire _21582_;
  wire _21583_;
  wire _21584_;
  wire _21585_;
  wire _21586_;
  wire _21587_;
  wire _21588_;
  wire _21589_;
  wire _21590_;
  wire _21591_;
  wire _21592_;
  wire _21593_;
  wire _21594_;
  wire _21595_;
  wire _21596_;
  wire _21597_;
  wire _21598_;
  wire _21599_;
  wire _21600_;
  wire _21601_;
  wire _21602_;
  wire _21603_;
  wire _21604_;
  wire _21605_;
  wire _21606_;
  wire _21607_;
  wire _21608_;
  wire _21609_;
  wire _21610_;
  wire _21611_;
  wire _21612_;
  wire _21613_;
  wire _21614_;
  wire _21615_;
  wire _21616_;
  wire _21617_;
  wire _21618_;
  wire _21619_;
  wire _21620_;
  wire _21621_;
  wire _21622_;
  wire _21623_;
  wire _21624_;
  wire _21625_;
  wire _21626_;
  wire _21627_;
  wire _21628_;
  wire _21629_;
  wire _21630_;
  wire _21631_;
  wire _21632_;
  wire _21633_;
  wire _21634_;
  wire _21635_;
  wire _21636_;
  wire _21637_;
  wire _21638_;
  wire _21639_;
  wire _21640_;
  wire _21641_;
  wire _21642_;
  wire _21643_;
  wire _21644_;
  wire _21645_;
  wire _21646_;
  wire _21647_;
  wire _21648_;
  wire _21649_;
  wire _21650_;
  wire _21651_;
  wire _21652_;
  wire _21653_;
  wire _21654_;
  wire _21655_;
  wire _21656_;
  wire _21657_;
  wire _21658_;
  wire _21659_;
  wire _21660_;
  wire _21661_;
  wire _21662_;
  wire _21663_;
  wire _21664_;
  wire _21665_;
  wire _21666_;
  wire _21667_;
  wire _21668_;
  wire _21669_;
  wire _21670_;
  wire _21671_;
  wire _21672_;
  wire _21673_;
  wire _21674_;
  wire _21675_;
  wire _21676_;
  wire _21677_;
  wire _21678_;
  wire _21679_;
  wire _21680_;
  wire _21681_;
  wire _21682_;
  wire _21683_;
  wire _21684_;
  wire _21685_;
  wire _21686_;
  wire _21687_;
  wire _21688_;
  wire _21689_;
  wire _21690_;
  wire _21691_;
  wire _21692_;
  wire _21693_;
  wire _21694_;
  wire _21695_;
  wire _21696_;
  wire _21697_;
  wire _21698_;
  wire _21699_;
  wire _21700_;
  wire _21701_;
  wire _21702_;
  wire _21703_;
  wire _21704_;
  wire _21705_;
  wire _21706_;
  wire _21707_;
  wire _21708_;
  wire _21709_;
  wire _21710_;
  wire _21711_;
  wire _21712_;
  wire _21713_;
  wire _21714_;
  wire _21715_;
  wire _21716_;
  wire _21717_;
  wire _21718_;
  wire _21719_;
  wire _21720_;
  wire _21721_;
  wire _21722_;
  wire _21723_;
  wire _21724_;
  wire _21725_;
  wire _21726_;
  wire _21727_;
  wire _21728_;
  wire _21729_;
  wire _21730_;
  wire _21731_;
  wire _21732_;
  wire _21733_;
  wire _21734_;
  wire _21735_;
  wire _21736_;
  wire _21737_;
  wire _21738_;
  wire _21739_;
  wire _21740_;
  wire _21741_;
  wire _21742_;
  wire _21743_;
  wire _21744_;
  wire _21745_;
  wire _21746_;
  wire _21747_;
  wire _21748_;
  wire _21749_;
  wire _21750_;
  wire _21751_;
  wire _21752_;
  wire _21753_;
  wire _21754_;
  wire _21755_;
  wire _21756_;
  wire _21757_;
  wire _21758_;
  wire _21759_;
  wire _21760_;
  wire _21761_;
  wire _21762_;
  wire _21763_;
  wire _21764_;
  wire _21765_;
  wire _21766_;
  wire _21767_;
  wire _21768_;
  wire _21769_;
  wire _21770_;
  wire _21771_;
  wire _21772_;
  wire _21773_;
  wire _21774_;
  wire _21775_;
  wire _21776_;
  wire _21777_;
  wire _21778_;
  wire _21779_;
  wire _21780_;
  wire _21781_;
  wire _21782_;
  wire _21783_;
  wire _21784_;
  wire _21785_;
  wire _21786_;
  wire _21787_;
  wire _21788_;
  wire _21789_;
  wire _21790_;
  wire _21791_;
  wire _21792_;
  wire _21793_;
  wire _21794_;
  wire _21795_;
  wire _21796_;
  wire _21797_;
  wire _21798_;
  wire _21799_;
  wire _21800_;
  wire _21801_;
  wire _21802_;
  wire _21803_;
  wire _21804_;
  wire _21805_;
  wire _21806_;
  wire _21807_;
  wire _21808_;
  wire _21809_;
  wire _21810_;
  wire _21811_;
  wire _21812_;
  wire _21813_;
  wire _21814_;
  wire _21815_;
  wire _21816_;
  wire _21817_;
  wire _21818_;
  wire _21819_;
  wire _21820_;
  wire _21821_;
  wire _21822_;
  wire _21823_;
  wire _21824_;
  wire _21825_;
  wire _21826_;
  wire _21827_;
  wire _21828_;
  wire _21829_;
  wire _21830_;
  wire _21831_;
  wire _21832_;
  wire _21833_;
  wire _21834_;
  wire _21835_;
  wire _21836_;
  wire _21837_;
  wire _21838_;
  wire _21839_;
  wire _21840_;
  wire _21841_;
  wire _21842_;
  wire _21843_;
  wire _21844_;
  wire _21845_;
  wire _21846_;
  wire _21847_;
  wire _21848_;
  wire _21849_;
  wire _21850_;
  wire _21851_;
  wire _21852_;
  wire _21853_;
  wire _21854_;
  wire _21855_;
  wire _21856_;
  wire _21857_;
  wire _21858_;
  wire _21859_;
  wire _21860_;
  wire _21861_;
  wire _21862_;
  wire _21863_;
  wire _21864_;
  wire _21865_;
  wire _21866_;
  wire _21867_;
  wire _21868_;
  wire _21869_;
  wire _21870_;
  wire _21871_;
  wire _21872_;
  wire _21873_;
  wire _21874_;
  wire _21875_;
  wire _21876_;
  wire _21877_;
  wire _21878_;
  wire _21879_;
  wire _21880_;
  wire _21881_;
  wire _21882_;
  wire _21883_;
  wire _21884_;
  wire _21885_;
  wire _21886_;
  wire _21887_;
  wire _21888_;
  wire _21889_;
  wire _21890_;
  wire _21891_;
  wire _21892_;
  wire _21893_;
  wire _21894_;
  wire _21895_;
  wire _21896_;
  wire _21897_;
  wire _21898_;
  wire _21899_;
  wire _21900_;
  wire _21901_;
  wire _21902_;
  wire _21903_;
  wire _21904_;
  wire _21905_;
  wire _21906_;
  wire _21907_;
  wire _21908_;
  wire _21909_;
  wire _21910_;
  wire _21911_;
  wire _21912_;
  wire _21913_;
  wire _21914_;
  wire _21915_;
  wire _21916_;
  wire _21917_;
  wire _21918_;
  wire _21919_;
  wire _21920_;
  wire _21921_;
  wire _21922_;
  wire _21923_;
  wire _21924_;
  wire _21925_;
  wire _21926_;
  wire _21927_;
  wire _21928_;
  wire _21929_;
  wire _21930_;
  wire _21931_;
  wire _21932_;
  wire _21933_;
  wire _21934_;
  wire _21935_;
  wire _21936_;
  wire _21937_;
  wire _21938_;
  wire _21939_;
  wire _21940_;
  wire _21941_;
  wire _21942_;
  wire _21943_;
  wire _21944_;
  wire _21945_;
  wire _21946_;
  wire _21947_;
  wire _21948_;
  wire _21949_;
  wire _21950_;
  wire _21951_;
  wire _21952_;
  wire _21953_;
  wire _21954_;
  wire _21955_;
  wire _21956_;
  wire _21957_;
  wire _21958_;
  wire _21959_;
  wire _21960_;
  wire _21961_;
  wire _21962_;
  wire _21963_;
  wire _21964_;
  wire _21965_;
  wire _21966_;
  wire _21967_;
  wire _21968_;
  wire _21969_;
  wire _21970_;
  wire _21971_;
  wire _21972_;
  wire _21973_;
  wire _21974_;
  wire _21975_;
  wire _21976_;
  wire _21977_;
  wire _21978_;
  wire _21979_;
  wire _21980_;
  wire _21981_;
  wire _21982_;
  wire _21983_;
  wire _21984_;
  wire _21985_;
  wire _21986_;
  wire _21987_;
  wire _21988_;
  wire _21989_;
  wire _21990_;
  wire _21991_;
  wire _21992_;
  wire _21993_;
  wire _21994_;
  wire _21995_;
  wire _21996_;
  wire _21997_;
  wire _21998_;
  wire _21999_;
  wire _22000_;
  wire _22001_;
  wire _22002_;
  wire _22003_;
  wire _22004_;
  wire _22005_;
  wire _22006_;
  wire _22007_;
  wire _22008_;
  wire _22009_;
  wire _22010_;
  wire _22011_;
  wire _22012_;
  wire _22013_;
  wire _22014_;
  wire _22015_;
  wire _22016_;
  wire _22017_;
  wire _22018_;
  wire _22019_;
  wire _22020_;
  wire _22021_;
  wire _22022_;
  wire _22023_;
  wire _22024_;
  wire _22025_;
  wire _22026_;
  wire _22027_;
  wire _22028_;
  wire _22029_;
  wire _22030_;
  wire _22031_;
  wire _22032_;
  wire _22033_;
  wire _22034_;
  wire _22035_;
  wire _22036_;
  wire _22037_;
  wire _22038_;
  wire _22039_;
  wire _22040_;
  wire _22041_;
  wire _22042_;
  wire _22043_;
  wire _22044_;
  wire _22045_;
  wire _22046_;
  wire _22047_;
  wire _22048_;
  wire _22049_;
  wire _22050_;
  wire _22051_;
  wire _22052_;
  wire _22053_;
  wire _22054_;
  wire _22055_;
  wire _22056_;
  wire _22057_;
  wire _22058_;
  wire _22059_;
  wire _22060_;
  wire _22061_;
  wire _22062_;
  wire _22063_;
  wire _22064_;
  wire _22065_;
  wire _22066_;
  wire _22067_;
  wire _22068_;
  wire _22069_;
  wire _22070_;
  wire _22071_;
  wire _22072_;
  wire _22073_;
  wire _22074_;
  wire _22075_;
  wire _22076_;
  wire _22077_;
  wire _22078_;
  wire _22079_;
  wire _22080_;
  wire _22081_;
  wire _22082_;
  wire _22083_;
  wire _22084_;
  wire _22085_;
  wire _22086_;
  wire _22087_;
  wire _22088_;
  wire _22089_;
  wire _22090_;
  wire _22091_;
  wire _22092_;
  wire _22093_;
  wire _22094_;
  wire _22095_;
  wire _22096_;
  wire _22097_;
  wire _22098_;
  wire _22099_;
  wire _22100_;
  wire _22101_;
  wire _22102_;
  wire _22103_;
  wire _22104_;
  wire _22105_;
  wire _22106_;
  wire _22107_;
  wire _22108_;
  wire _22109_;
  wire _22110_;
  wire _22111_;
  wire _22112_;
  wire _22113_;
  wire _22114_;
  wire _22115_;
  wire _22116_;
  wire _22117_;
  wire _22118_;
  wire _22119_;
  wire _22120_;
  wire _22121_;
  wire _22122_;
  wire _22123_;
  wire _22124_;
  wire _22125_;
  wire _22126_;
  wire _22127_;
  wire _22128_;
  wire _22129_;
  wire _22130_;
  wire _22131_;
  wire _22132_;
  wire _22133_;
  wire _22134_;
  wire _22135_;
  wire _22136_;
  wire _22137_;
  wire _22138_;
  wire _22139_;
  wire _22140_;
  wire _22141_;
  wire _22142_;
  wire _22143_;
  wire _22144_;
  wire _22145_;
  wire _22146_;
  wire _22147_;
  wire _22148_;
  wire _22149_;
  wire _22150_;
  wire _22151_;
  wire _22152_;
  wire _22153_;
  wire _22154_;
  wire _22155_;
  wire _22156_;
  wire _22157_;
  wire _22158_;
  wire _22159_;
  wire _22160_;
  wire _22161_;
  wire _22162_;
  wire _22163_;
  wire _22164_;
  wire _22165_;
  wire _22166_;
  wire _22167_;
  wire _22168_;
  wire _22169_;
  wire _22170_;
  wire _22171_;
  wire _22172_;
  wire _22173_;
  wire _22174_;
  wire _22175_;
  wire _22176_;
  wire _22177_;
  wire _22178_;
  wire _22179_;
  wire _22180_;
  wire _22181_;
  wire _22182_;
  wire _22183_;
  wire _22184_;
  wire _22185_;
  wire _22186_;
  wire _22187_;
  wire _22188_;
  wire _22189_;
  wire _22190_;
  wire _22191_;
  wire _22192_;
  wire _22193_;
  wire _22194_;
  wire _22195_;
  wire _22196_;
  wire _22197_;
  wire _22198_;
  wire _22199_;
  wire _22200_;
  wire _22201_;
  wire _22202_;
  wire _22203_;
  wire _22204_;
  wire _22205_;
  wire _22206_;
  wire _22207_;
  wire _22208_;
  wire _22209_;
  wire _22210_;
  wire _22211_;
  wire _22212_;
  wire _22213_;
  wire _22214_;
  wire _22215_;
  wire _22216_;
  wire _22217_;
  wire _22218_;
  wire _22219_;
  wire _22220_;
  wire _22221_;
  wire _22222_;
  wire _22223_;
  wire _22224_;
  wire _22225_;
  wire _22226_;
  wire _22227_;
  wire _22228_;
  wire _22229_;
  wire _22230_;
  wire _22231_;
  wire _22232_;
  wire _22233_;
  wire _22234_;
  wire _22235_;
  wire _22236_;
  wire _22237_;
  wire _22238_;
  wire _22239_;
  wire _22240_;
  wire _22241_;
  wire _22242_;
  wire _22243_;
  wire _22244_;
  wire _22245_;
  wire _22246_;
  wire _22247_;
  wire _22248_;
  wire _22249_;
  wire _22250_;
  wire _22251_;
  wire _22252_;
  wire _22253_;
  wire _22254_;
  wire _22255_;
  wire _22256_;
  wire _22257_;
  wire _22258_;
  wire _22259_;
  wire _22260_;
  wire _22261_;
  wire _22262_;
  wire _22263_;
  wire _22264_;
  wire _22265_;
  wire _22266_;
  wire _22267_;
  wire _22268_;
  wire _22269_;
  wire _22270_;
  wire _22271_;
  wire _22272_;
  wire _22273_;
  wire _22274_;
  wire _22275_;
  wire _22276_;
  wire _22277_;
  wire _22278_;
  wire _22279_;
  wire _22280_;
  wire _22281_;
  wire _22282_;
  wire _22283_;
  wire _22284_;
  wire _22285_;
  wire _22286_;
  wire _22287_;
  wire _22288_;
  wire _22289_;
  wire _22290_;
  wire _22291_;
  wire _22292_;
  wire _22293_;
  wire _22294_;
  wire _22295_;
  wire _22296_;
  wire _22297_;
  wire _22298_;
  wire _22299_;
  wire _22300_;
  wire _22301_;
  wire _22302_;
  wire _22303_;
  wire _22304_;
  wire _22305_;
  wire _22306_;
  wire _22307_;
  wire _22308_;
  wire _22309_;
  wire _22310_;
  wire _22311_;
  wire _22312_;
  wire _22313_;
  wire _22314_;
  wire _22315_;
  wire _22316_;
  wire _22317_;
  wire _22318_;
  wire _22319_;
  wire _22320_;
  wire _22321_;
  wire _22322_;
  wire _22323_;
  wire _22324_;
  wire _22325_;
  wire _22326_;
  wire _22327_;
  wire _22328_;
  wire _22329_;
  wire _22330_;
  wire _22331_;
  wire _22332_;
  wire _22333_;
  wire _22334_;
  wire _22335_;
  wire _22336_;
  wire _22337_;
  wire _22338_;
  wire _22339_;
  wire _22340_;
  wire _22341_;
  wire _22342_;
  wire _22343_;
  wire _22344_;
  wire _22345_;
  wire _22346_;
  wire _22347_;
  wire _22348_;
  wire _22349_;
  wire _22350_;
  wire _22351_;
  wire _22352_;
  wire _22353_;
  wire _22354_;
  wire _22355_;
  wire _22356_;
  wire _22357_;
  wire _22358_;
  wire _22359_;
  wire _22360_;
  wire _22361_;
  wire _22362_;
  wire _22363_;
  wire _22364_;
  wire _22365_;
  wire _22366_;
  wire _22367_;
  wire _22368_;
  wire _22369_;
  wire _22370_;
  wire _22371_;
  wire _22372_;
  wire _22373_;
  wire _22374_;
  wire _22375_;
  wire _22376_;
  wire _22377_;
  wire _22378_;
  wire _22379_;
  wire _22380_;
  wire _22381_;
  wire _22382_;
  wire _22383_;
  wire _22384_;
  wire _22385_;
  wire _22386_;
  wire _22387_;
  wire _22388_;
  wire _22389_;
  wire _22390_;
  wire _22391_;
  wire _22392_;
  wire _22393_;
  wire _22394_;
  wire _22395_;
  wire _22396_;
  wire _22397_;
  wire _22398_;
  wire _22399_;
  wire _22400_;
  wire _22401_;
  wire _22402_;
  wire _22403_;
  wire _22404_;
  wire _22405_;
  wire _22406_;
  wire _22407_;
  wire _22408_;
  wire _22409_;
  wire _22410_;
  wire _22411_;
  wire _22412_;
  wire _22413_;
  wire _22414_;
  wire _22415_;
  wire _22416_;
  wire _22417_;
  wire _22418_;
  wire _22419_;
  wire _22420_;
  wire _22421_;
  wire _22422_;
  wire _22423_;
  wire _22424_;
  wire _22425_;
  wire _22426_;
  wire _22427_;
  wire _22428_;
  wire _22429_;
  wire _22430_;
  wire _22431_;
  wire _22432_;
  wire _22433_;
  wire _22434_;
  wire _22435_;
  wire _22436_;
  wire _22437_;
  wire _22438_;
  wire _22439_;
  wire _22440_;
  wire _22441_;
  wire _22442_;
  wire _22443_;
  wire _22444_;
  wire _22445_;
  wire _22446_;
  wire _22447_;
  wire _22448_;
  wire _22449_;
  wire _22450_;
  wire _22451_;
  wire _22452_;
  wire _22453_;
  wire _22454_;
  wire _22455_;
  wire _22456_;
  wire _22457_;
  wire _22458_;
  wire _22459_;
  wire _22460_;
  wire _22461_;
  wire _22462_;
  wire _22463_;
  wire _22464_;
  wire _22465_;
  wire _22466_;
  wire _22467_;
  wire _22468_;
  wire _22469_;
  wire _22470_;
  wire _22471_;
  wire _22472_;
  wire _22473_;
  wire _22474_;
  wire _22475_;
  wire _22476_;
  wire _22477_;
  wire _22478_;
  wire _22479_;
  wire _22480_;
  wire _22481_;
  wire _22482_;
  wire _22483_;
  wire _22484_;
  wire _22485_;
  wire _22486_;
  wire _22487_;
  wire _22488_;
  wire _22489_;
  wire _22490_;
  wire _22491_;
  wire _22492_;
  wire _22493_;
  wire _22494_;
  wire _22495_;
  wire _22496_;
  wire _22497_;
  wire _22498_;
  wire _22499_;
  wire _22500_;
  wire _22501_;
  wire _22502_;
  wire _22503_;
  wire _22504_;
  wire _22505_;
  wire _22506_;
  wire _22507_;
  wire _22508_;
  wire _22509_;
  wire _22510_;
  wire _22511_;
  wire _22512_;
  wire _22513_;
  wire _22514_;
  wire _22515_;
  wire _22516_;
  wire _22517_;
  wire _22518_;
  wire _22519_;
  wire _22520_;
  wire _22521_;
  wire _22522_;
  wire _22523_;
  wire _22524_;
  wire _22525_;
  wire _22526_;
  wire _22527_;
  wire _22528_;
  wire _22529_;
  wire _22530_;
  wire _22531_;
  wire _22532_;
  wire _22533_;
  wire _22534_;
  wire _22535_;
  wire _22536_;
  wire _22537_;
  wire _22538_;
  wire _22539_;
  wire _22540_;
  wire _22541_;
  wire _22542_;
  wire _22543_;
  wire _22544_;
  wire _22545_;
  wire _22546_;
  wire _22547_;
  wire _22548_;
  wire _22549_;
  wire _22550_;
  wire _22551_;
  wire _22552_;
  wire _22553_;
  wire _22554_;
  wire _22555_;
  wire _22556_;
  wire _22557_;
  wire _22558_;
  wire _22559_;
  wire _22560_;
  wire _22561_;
  wire _22562_;
  wire _22563_;
  wire _22564_;
  wire _22565_;
  wire _22566_;
  wire _22567_;
  wire _22568_;
  wire _22569_;
  wire _22570_;
  wire _22571_;
  wire _22572_;
  wire _22573_;
  wire _22574_;
  wire _22575_;
  wire _22576_;
  wire _22577_;
  wire _22578_;
  wire _22579_;
  wire _22580_;
  wire _22581_;
  wire _22582_;
  wire _22583_;
  wire _22584_;
  wire _22585_;
  wire _22586_;
  wire _22587_;
  wire _22588_;
  wire _22589_;
  wire _22590_;
  wire _22591_;
  wire _22592_;
  wire _22593_;
  wire _22594_;
  wire _22595_;
  wire _22596_;
  wire _22597_;
  wire _22598_;
  wire _22599_;
  wire _22600_;
  wire _22601_;
  wire _22602_;
  wire _22603_;
  wire _22604_;
  wire _22605_;
  wire _22606_;
  wire _22607_;
  wire _22608_;
  wire _22609_;
  wire _22610_;
  wire _22611_;
  wire _22612_;
  wire _22613_;
  wire _22614_;
  wire _22615_;
  wire _22616_;
  wire _22617_;
  wire _22618_;
  wire _22619_;
  wire _22620_;
  wire _22621_;
  wire _22622_;
  wire _22623_;
  wire _22624_;
  wire _22625_;
  wire _22626_;
  wire _22627_;
  wire _22628_;
  wire _22629_;
  wire _22630_;
  wire _22631_;
  wire _22632_;
  wire _22633_;
  wire _22634_;
  wire _22635_;
  wire _22636_;
  wire _22637_;
  wire _22638_;
  wire _22639_;
  wire _22640_;
  wire _22641_;
  wire _22642_;
  wire _22643_;
  wire _22644_;
  wire _22645_;
  wire _22646_;
  wire _22647_;
  wire _22648_;
  wire _22649_;
  wire _22650_;
  wire _22651_;
  wire _22652_;
  wire _22653_;
  wire _22654_;
  wire _22655_;
  wire _22656_;
  wire _22657_;
  wire _22658_;
  wire _22659_;
  wire _22660_;
  wire _22661_;
  wire _22662_;
  wire _22663_;
  wire _22664_;
  wire _22665_;
  wire _22666_;
  wire _22667_;
  wire _22668_;
  wire _22669_;
  wire _22670_;
  wire _22671_;
  wire _22672_;
  wire _22673_;
  wire _22674_;
  wire _22675_;
  wire _22676_;
  wire _22677_;
  wire _22678_;
  wire _22679_;
  wire _22680_;
  wire _22681_;
  wire _22682_;
  wire _22683_;
  wire _22684_;
  wire _22685_;
  wire _22686_;
  wire _22687_;
  wire _22688_;
  wire _22689_;
  wire _22690_;
  wire _22691_;
  wire _22692_;
  wire _22693_;
  wire _22694_;
  wire _22695_;
  wire _22696_;
  wire _22697_;
  wire _22698_;
  wire _22699_;
  wire _22700_;
  wire _22701_;
  wire _22702_;
  wire _22703_;
  wire _22704_;
  wire _22705_;
  wire _22706_;
  wire _22707_;
  wire _22708_;
  wire _22709_;
  wire _22710_;
  wire _22711_;
  wire _22712_;
  wire _22713_;
  wire _22714_;
  wire _22715_;
  wire _22716_;
  wire _22717_;
  wire _22718_;
  wire _22719_;
  wire _22720_;
  wire _22721_;
  wire _22722_;
  wire _22723_;
  wire _22724_;
  wire _22725_;
  wire _22726_;
  wire _22727_;
  wire _22728_;
  wire _22729_;
  wire _22730_;
  wire _22731_;
  wire _22732_;
  wire _22733_;
  wire _22734_;
  wire _22735_;
  wire _22736_;
  wire _22737_;
  wire _22738_;
  wire _22739_;
  wire _22740_;
  wire _22741_;
  wire _22742_;
  wire _22743_;
  wire _22744_;
  wire _22745_;
  wire _22746_;
  wire _22747_;
  wire _22748_;
  wire _22749_;
  wire _22750_;
  wire _22751_;
  wire _22752_;
  wire _22753_;
  wire _22754_;
  wire _22755_;
  wire _22756_;
  wire _22757_;
  wire _22758_;
  wire _22759_;
  wire _22760_;
  wire _22761_;
  wire _22762_;
  wire _22763_;
  wire _22764_;
  wire _22765_;
  wire _22766_;
  wire _22767_;
  wire _22768_;
  wire _22769_;
  wire _22770_;
  wire _22771_;
  wire _22772_;
  wire _22773_;
  wire _22774_;
  wire _22775_;
  wire _22776_;
  wire _22777_;
  wire _22778_;
  wire _22779_;
  wire _22780_;
  wire _22781_;
  wire _22782_;
  wire _22783_;
  wire _22784_;
  wire _22785_;
  wire _22786_;
  wire _22787_;
  wire _22788_;
  wire _22789_;
  wire _22790_;
  wire _22791_;
  wire _22792_;
  wire _22793_;
  wire _22794_;
  wire _22795_;
  wire _22796_;
  wire _22797_;
  wire _22798_;
  wire _22799_;
  wire _22800_;
  wire _22801_;
  wire _22802_;
  wire _22803_;
  wire _22804_;
  wire _22805_;
  wire _22806_;
  wire _22807_;
  wire _22808_;
  wire _22809_;
  wire _22810_;
  wire _22811_;
  wire _22812_;
  wire _22813_;
  wire _22814_;
  wire _22815_;
  wire _22816_;
  wire _22817_;
  wire _22818_;
  wire _22819_;
  wire _22820_;
  wire _22821_;
  wire _22822_;
  wire _22823_;
  wire _22824_;
  wire _22825_;
  wire _22826_;
  wire _22827_;
  wire _22828_;
  wire _22829_;
  wire _22830_;
  wire _22831_;
  wire _22832_;
  wire _22833_;
  wire _22834_;
  wire _22835_;
  wire _22836_;
  wire _22837_;
  wire _22838_;
  wire _22839_;
  wire _22840_;
  wire _22841_;
  wire _22842_;
  wire _22843_;
  wire _22844_;
  wire _22845_;
  wire _22846_;
  wire _22847_;
  wire _22848_;
  wire _22849_;
  wire _22850_;
  wire _22851_;
  wire _22852_;
  wire _22853_;
  wire _22854_;
  wire _22855_;
  wire _22856_;
  wire _22857_;
  wire _22858_;
  wire _22859_;
  wire _22860_;
  wire _22861_;
  wire _22862_;
  wire _22863_;
  wire _22864_;
  wire _22865_;
  wire _22866_;
  wire _22867_;
  wire _22868_;
  wire _22869_;
  wire _22870_;
  wire _22871_;
  wire _22872_;
  wire _22873_;
  wire _22874_;
  wire _22875_;
  wire _22876_;
  wire _22877_;
  wire _22878_;
  wire _22879_;
  wire _22880_;
  wire _22881_;
  wire _22882_;
  wire _22883_;
  wire _22884_;
  wire _22885_;
  wire _22886_;
  wire _22887_;
  wire _22888_;
  wire _22889_;
  wire _22890_;
  wire _22891_;
  wire _22892_;
  wire _22893_;
  wire _22894_;
  wire _22895_;
  wire _22896_;
  wire _22897_;
  wire _22898_;
  wire _22899_;
  wire _22900_;
  wire _22901_;
  wire _22902_;
  wire _22903_;
  wire _22904_;
  wire _22905_;
  wire _22906_;
  wire _22907_;
  wire _22908_;
  wire _22909_;
  wire _22910_;
  wire _22911_;
  wire _22912_;
  wire _22913_;
  wire _22914_;
  wire _22915_;
  wire _22916_;
  wire _22917_;
  wire _22918_;
  wire _22919_;
  wire _22920_;
  wire _22921_;
  wire _22922_;
  wire _22923_;
  wire _22924_;
  wire _22925_;
  wire _22926_;
  wire _22927_;
  wire _22928_;
  wire _22929_;
  wire _22930_;
  wire _22931_;
  wire _22932_;
  wire _22933_;
  wire _22934_;
  wire _22935_;
  wire _22936_;
  wire _22937_;
  wire _22938_;
  wire _22939_;
  wire _22940_;
  wire _22941_;
  wire _22942_;
  wire _22943_;
  wire _22944_;
  wire _22945_;
  wire _22946_;
  wire _22947_;
  wire _22948_;
  wire _22949_;
  wire _22950_;
  wire _22951_;
  wire _22952_;
  wire _22953_;
  wire _22954_;
  wire _22955_;
  wire _22956_;
  wire _22957_;
  wire _22958_;
  wire _22959_;
  wire _22960_;
  wire _22961_;
  wire _22962_;
  wire _22963_;
  wire _22964_;
  wire _22965_;
  wire _22966_;
  wire _22967_;
  wire _22968_;
  wire _22969_;
  wire _22970_;
  wire _22971_;
  wire _22972_;
  wire _22973_;
  wire _22974_;
  wire _22975_;
  wire _22976_;
  wire _22977_;
  wire _22978_;
  wire _22979_;
  wire _22980_;
  wire _22981_;
  wire _22982_;
  wire _22983_;
  wire _22984_;
  wire _22985_;
  wire _22986_;
  wire _22987_;
  wire _22988_;
  wire _22989_;
  wire _22990_;
  wire _22991_;
  wire _22992_;
  wire _22993_;
  wire _22994_;
  wire _22995_;
  wire _22996_;
  wire _22997_;
  wire _22998_;
  wire _22999_;
  wire _23000_;
  wire _23001_;
  wire _23002_;
  wire _23003_;
  wire _23004_;
  wire _23005_;
  wire _23006_;
  wire _23007_;
  wire _23008_;
  wire _23009_;
  wire _23010_;
  wire _23011_;
  wire _23012_;
  wire _23013_;
  wire _23014_;
  wire _23015_;
  wire _23016_;
  wire _23017_;
  wire _23018_;
  wire _23019_;
  wire _23020_;
  wire _23021_;
  wire _23022_;
  wire _23023_;
  wire _23024_;
  wire _23025_;
  wire _23026_;
  wire _23027_;
  wire _23028_;
  wire _23029_;
  wire _23030_;
  wire _23031_;
  wire _23032_;
  wire _23033_;
  wire _23034_;
  wire _23035_;
  wire _23036_;
  wire _23037_;
  wire _23038_;
  wire _23039_;
  wire _23040_;
  wire _23041_;
  wire _23042_;
  wire _23043_;
  wire _23044_;
  wire _23045_;
  wire _23046_;
  wire _23047_;
  wire _23048_;
  wire _23049_;
  wire _23050_;
  wire _23051_;
  wire _23052_;
  wire _23053_;
  wire _23054_;
  wire _23055_;
  wire _23056_;
  wire _23057_;
  wire _23058_;
  wire _23059_;
  wire _23060_;
  wire _23061_;
  wire _23062_;
  wire _23063_;
  wire _23064_;
  wire _23065_;
  wire _23066_;
  wire _23067_;
  wire _23068_;
  wire _23069_;
  wire _23070_;
  wire _23071_;
  wire _23072_;
  wire _23073_;
  wire _23074_;
  wire _23075_;
  wire _23076_;
  wire _23077_;
  wire _23078_;
  wire _23079_;
  wire _23080_;
  wire _23081_;
  wire _23082_;
  wire _23083_;
  wire _23084_;
  wire _23085_;
  wire _23086_;
  wire _23087_;
  wire _23088_;
  wire _23089_;
  wire _23090_;
  wire _23091_;
  wire _23092_;
  wire _23093_;
  wire _23094_;
  wire _23095_;
  wire _23096_;
  wire _23097_;
  wire _23098_;
  wire _23099_;
  wire _23100_;
  wire _23101_;
  wire _23102_;
  wire _23103_;
  wire _23104_;
  wire _23105_;
  wire _23106_;
  wire _23107_;
  wire _23108_;
  wire _23109_;
  wire _23110_;
  wire _23111_;
  wire _23112_;
  wire _23113_;
  wire _23114_;
  wire _23115_;
  wire _23116_;
  wire _23117_;
  wire _23118_;
  wire _23119_;
  wire _23120_;
  wire _23121_;
  wire _23122_;
  wire _23123_;
  wire _23124_;
  wire _23125_;
  wire _23126_;
  wire _23127_;
  wire _23128_;
  wire _23129_;
  wire _23130_;
  wire _23131_;
  wire _23132_;
  wire _23133_;
  wire _23134_;
  wire _23135_;
  wire _23136_;
  wire _23137_;
  wire _23138_;
  wire _23139_;
  wire _23140_;
  wire _23141_;
  wire _23142_;
  wire _23143_;
  wire _23144_;
  wire _23145_;
  wire _23146_;
  wire _23147_;
  wire _23148_;
  wire _23149_;
  wire _23150_;
  wire _23151_;
  wire _23152_;
  wire _23153_;
  wire _23154_;
  wire _23155_;
  wire _23156_;
  wire _23157_;
  wire _23158_;
  wire _23159_;
  wire _23160_;
  wire _23161_;
  wire _23162_;
  wire _23163_;
  wire _23164_;
  wire _23165_;
  wire _23166_;
  wire _23167_;
  wire _23168_;
  wire _23169_;
  wire _23170_;
  wire _23171_;
  wire _23172_;
  wire _23173_;
  wire _23174_;
  wire _23175_;
  wire _23176_;
  wire _23177_;
  wire _23178_;
  wire _23179_;
  wire _23180_;
  wire _23181_;
  wire _23182_;
  wire _23183_;
  wire _23184_;
  wire _23185_;
  wire _23186_;
  wire _23187_;
  wire _23188_;
  wire _23189_;
  wire _23190_;
  wire _23191_;
  wire _23192_;
  wire _23193_;
  wire _23194_;
  wire _23195_;
  wire _23196_;
  wire _23197_;
  wire _23198_;
  wire _23199_;
  wire _23200_;
  wire _23201_;
  wire _23202_;
  wire _23203_;
  wire _23204_;
  wire _23205_;
  wire _23206_;
  wire _23207_;
  wire _23208_;
  wire _23209_;
  wire _23210_;
  wire _23211_;
  wire _23212_;
  wire _23213_;
  wire _23214_;
  wire _23215_;
  wire _23216_;
  wire _23217_;
  wire _23218_;
  wire _23219_;
  wire _23220_;
  wire _23221_;
  wire _23222_;
  wire _23223_;
  wire _23224_;
  wire _23225_;
  wire _23226_;
  wire _23227_;
  wire _23228_;
  wire _23229_;
  wire _23230_;
  wire _23231_;
  wire _23232_;
  wire _23233_;
  wire _23234_;
  wire _23235_;
  wire _23236_;
  wire _23237_;
  wire _23238_;
  wire _23239_;
  wire _23240_;
  wire _23241_;
  wire _23242_;
  wire _23243_;
  wire _23244_;
  wire _23245_;
  wire _23246_;
  wire _23247_;
  wire _23248_;
  wire _23249_;
  wire _23250_;
  wire _23251_;
  wire _23252_;
  wire _23253_;
  wire _23254_;
  wire _23255_;
  wire _23256_;
  wire _23257_;
  wire _23258_;
  wire _23259_;
  wire _23260_;
  wire _23261_;
  wire _23262_;
  wire _23263_;
  wire _23264_;
  wire _23265_;
  wire _23266_;
  wire _23267_;
  wire _23268_;
  wire _23269_;
  wire _23270_;
  wire _23271_;
  wire _23272_;
  wire _23273_;
  wire _23274_;
  wire _23275_;
  wire _23276_;
  wire _23277_;
  wire _23278_;
  wire _23279_;
  wire _23280_;
  wire _23281_;
  wire _23282_;
  wire _23283_;
  wire _23284_;
  wire _23285_;
  wire _23286_;
  wire _23287_;
  wire _23288_;
  wire _23289_;
  wire _23290_;
  wire _23291_;
  wire _23292_;
  wire _23293_;
  wire _23294_;
  wire _23295_;
  wire _23296_;
  wire _23297_;
  wire _23298_;
  wire _23299_;
  wire _23300_;
  wire _23301_;
  wire _23302_;
  wire _23303_;
  wire _23304_;
  wire _23305_;
  wire _23306_;
  wire _23307_;
  wire _23308_;
  wire _23309_;
  wire _23310_;
  wire _23311_;
  wire _23312_;
  wire _23313_;
  wire _23314_;
  wire _23315_;
  wire _23316_;
  wire _23317_;
  wire _23318_;
  wire _23319_;
  wire _23320_;
  wire _23321_;
  wire _23322_;
  wire _23323_;
  wire _23324_;
  wire _23325_;
  wire _23326_;
  wire _23327_;
  wire _23328_;
  wire _23329_;
  wire _23330_;
  wire _23331_;
  wire _23332_;
  wire _23333_;
  wire _23334_;
  wire _23335_;
  wire _23336_;
  wire _23337_;
  wire _23338_;
  wire _23339_;
  wire _23340_;
  wire _23341_;
  wire _23342_;
  wire _23343_;
  wire _23344_;
  wire _23345_;
  wire _23346_;
  wire _23347_;
  wire _23348_;
  wire _23349_;
  wire _23350_;
  wire _23351_;
  wire _23352_;
  wire _23353_;
  wire _23354_;
  wire _23355_;
  wire _23356_;
  wire _23357_;
  wire _23358_;
  wire _23359_;
  wire _23360_;
  wire _23361_;
  wire _23362_;
  wire _23363_;
  wire _23364_;
  wire _23365_;
  wire _23366_;
  wire _23367_;
  wire _23368_;
  wire _23369_;
  wire _23370_;
  wire _23371_;
  wire _23372_;
  wire _23373_;
  wire _23374_;
  wire _23375_;
  wire _23376_;
  wire _23377_;
  wire _23378_;
  wire _23379_;
  wire _23380_;
  wire _23381_;
  wire _23382_;
  wire _23383_;
  wire _23384_;
  wire _23385_;
  wire _23386_;
  wire _23387_;
  wire _23388_;
  wire _23389_;
  wire _23390_;
  wire _23391_;
  wire _23392_;
  wire _23393_;
  wire _23394_;
  wire _23395_;
  wire _23396_;
  wire _23397_;
  wire _23398_;
  wire _23399_;
  wire _23400_;
  wire _23401_;
  wire _23402_;
  wire _23403_;
  wire _23404_;
  wire _23405_;
  wire _23406_;
  wire _23407_;
  wire _23408_;
  wire _23409_;
  wire _23410_;
  wire _23411_;
  wire _23412_;
  wire _23413_;
  wire _23414_;
  wire _23415_;
  wire _23416_;
  wire _23417_;
  wire _23418_;
  wire _23419_;
  wire _23420_;
  wire _23421_;
  wire _23422_;
  wire _23423_;
  wire _23424_;
  wire _23425_;
  wire _23426_;
  wire _23427_;
  wire _23428_;
  wire _23429_;
  wire _23430_;
  wire _23431_;
  wire _23432_;
  wire _23433_;
  wire _23434_;
  wire _23435_;
  wire _23436_;
  wire _23437_;
  wire _23438_;
  wire _23439_;
  wire _23440_;
  wire _23441_;
  wire _23442_;
  wire _23443_;
  wire _23444_;
  wire _23445_;
  wire _23446_;
  wire _23447_;
  wire _23448_;
  wire _23449_;
  wire _23450_;
  wire _23451_;
  wire _23452_;
  wire _23453_;
  wire _23454_;
  wire _23455_;
  wire _23456_;
  wire _23457_;
  wire _23458_;
  wire _23459_;
  wire _23460_;
  wire _23461_;
  wire _23462_;
  wire _23463_;
  wire _23464_;
  wire _23465_;
  wire _23466_;
  wire _23467_;
  wire _23468_;
  wire _23469_;
  wire _23470_;
  wire _23471_;
  wire _23472_;
  wire _23473_;
  wire _23474_;
  wire _23475_;
  wire _23476_;
  wire _23477_;
  wire _23478_;
  wire _23479_;
  wire _23480_;
  wire _23481_;
  wire _23482_;
  wire _23483_;
  wire _23484_;
  wire _23485_;
  wire _23486_;
  wire _23487_;
  wire _23488_;
  wire _23489_;
  wire _23490_;
  wire _23491_;
  wire _23492_;
  wire _23493_;
  wire _23494_;
  wire _23495_;
  wire _23496_;
  wire _23497_;
  wire _23498_;
  wire _23499_;
  wire _23500_;
  wire _23501_;
  wire _23502_;
  wire _23503_;
  wire _23504_;
  wire _23505_;
  wire _23506_;
  wire _23507_;
  wire _23508_;
  wire _23509_;
  wire _23510_;
  wire _23511_;
  wire _23512_;
  wire _23513_;
  wire _23514_;
  wire _23515_;
  wire _23516_;
  wire _23517_;
  wire _23518_;
  wire _23519_;
  wire _23520_;
  wire _23521_;
  wire _23522_;
  wire _23523_;
  wire _23524_;
  wire _23525_;
  wire _23526_;
  wire _23527_;
  wire _23528_;
  wire _23529_;
  wire _23530_;
  wire _23531_;
  wire _23532_;
  wire _23533_;
  wire _23534_;
  wire _23535_;
  wire _23536_;
  wire _23537_;
  wire _23538_;
  wire _23539_;
  wire _23540_;
  wire _23541_;
  wire _23542_;
  wire _23543_;
  wire _23544_;
  wire _23545_;
  wire _23546_;
  wire _23547_;
  wire _23548_;
  wire _23549_;
  wire _23550_;
  wire _23551_;
  wire _23552_;
  wire _23553_;
  wire _23554_;
  wire _23555_;
  wire _23556_;
  wire _23557_;
  wire _23558_;
  wire _23559_;
  wire _23560_;
  wire _23561_;
  wire _23562_;
  wire _23563_;
  wire _23564_;
  wire _23565_;
  wire _23566_;
  wire _23567_;
  wire _23568_;
  wire _23569_;
  wire _23570_;
  wire _23571_;
  wire _23572_;
  wire _23573_;
  wire _23574_;
  wire _23575_;
  wire _23576_;
  wire _23577_;
  wire _23578_;
  wire _23579_;
  wire _23580_;
  wire _23581_;
  wire _23582_;
  wire _23583_;
  wire _23584_;
  wire _23585_;
  wire _23586_;
  wire _23587_;
  wire _23588_;
  wire _23589_;
  wire _23590_;
  wire _23591_;
  wire _23592_;
  wire _23593_;
  wire _23594_;
  wire _23595_;
  wire _23596_;
  wire _23597_;
  wire _23598_;
  wire _23599_;
  wire _23600_;
  wire _23601_;
  wire _23602_;
  wire _23603_;
  wire _23604_;
  wire _23605_;
  wire _23606_;
  wire _23607_;
  wire _23608_;
  wire _23609_;
  wire _23610_;
  wire _23611_;
  wire _23612_;
  wire _23613_;
  wire _23614_;
  wire _23615_;
  wire _23616_;
  wire _23617_;
  wire _23618_;
  wire _23619_;
  wire _23620_;
  wire _23621_;
  wire _23622_;
  wire _23623_;
  wire _23624_;
  wire _23625_;
  wire _23626_;
  wire _23627_;
  wire _23628_;
  wire _23629_;
  wire _23630_;
  wire _23631_;
  wire _23632_;
  wire _23633_;
  wire _23634_;
  wire _23635_;
  wire _23636_;
  wire _23637_;
  wire _23638_;
  wire _23639_;
  wire _23640_;
  wire _23641_;
  wire _23642_;
  wire _23643_;
  wire _23644_;
  wire _23645_;
  wire _23646_;
  wire _23647_;
  wire _23648_;
  wire _23649_;
  wire _23650_;
  wire _23651_;
  wire _23652_;
  wire _23653_;
  wire _23654_;
  wire _23655_;
  wire _23656_;
  wire _23657_;
  wire _23658_;
  wire _23659_;
  wire _23660_;
  wire _23661_;
  wire _23662_;
  wire _23663_;
  wire _23664_;
  wire _23665_;
  wire _23666_;
  wire _23667_;
  wire _23668_;
  wire _23669_;
  wire _23670_;
  wire _23671_;
  wire _23672_;
  wire _23673_;
  wire _23674_;
  wire _23675_;
  wire _23676_;
  wire _23677_;
  wire _23678_;
  wire _23679_;
  wire _23680_;
  wire _23681_;
  wire _23682_;
  wire _23683_;
  wire _23684_;
  wire _23685_;
  wire _23686_;
  wire _23687_;
  wire _23688_;
  wire _23689_;
  wire _23690_;
  wire _23691_;
  wire _23692_;
  wire _23693_;
  wire _23694_;
  wire _23695_;
  wire _23696_;
  wire _23697_;
  wire _23698_;
  wire _23699_;
  wire _23700_;
  wire _23701_;
  wire _23702_;
  wire _23703_;
  wire _23704_;
  wire _23705_;
  wire _23706_;
  wire _23707_;
  wire _23708_;
  wire _23709_;
  wire _23710_;
  wire _23711_;
  wire _23712_;
  wire _23713_;
  wire _23714_;
  wire _23715_;
  wire _23716_;
  wire _23717_;
  wire _23718_;
  wire _23719_;
  wire _23720_;
  wire _23721_;
  wire _23722_;
  wire _23723_;
  wire _23724_;
  wire _23725_;
  wire _23726_;
  wire _23727_;
  wire _23728_;
  wire _23729_;
  wire _23730_;
  wire _23731_;
  wire _23732_;
  wire _23733_;
  wire _23734_;
  wire _23735_;
  wire _23736_;
  wire _23737_;
  wire _23738_;
  wire _23739_;
  wire _23740_;
  wire _23741_;
  wire _23742_;
  wire _23743_;
  wire _23744_;
  wire _23745_;
  wire _23746_;
  wire _23747_;
  wire _23748_;
  wire _23749_;
  wire _23750_;
  wire _23751_;
  wire _23752_;
  wire _23753_;
  wire _23754_;
  wire _23755_;
  wire _23756_;
  wire _23757_;
  wire _23758_;
  wire _23759_;
  wire _23760_;
  wire _23761_;
  wire _23762_;
  wire _23763_;
  wire _23764_;
  wire _23765_;
  wire _23766_;
  wire _23767_;
  wire _23768_;
  wire _23769_;
  wire _23770_;
  wire _23771_;
  wire _23772_;
  wire _23773_;
  wire _23774_;
  wire _23775_;
  wire _23776_;
  wire _23777_;
  wire _23778_;
  wire _23779_;
  wire _23780_;
  wire _23781_;
  wire _23782_;
  wire _23783_;
  wire _23784_;
  wire _23785_;
  wire _23786_;
  wire _23787_;
  wire _23788_;
  wire _23789_;
  wire _23790_;
  wire _23791_;
  wire _23792_;
  wire _23793_;
  wire _23794_;
  wire _23795_;
  wire _23796_;
  wire _23797_;
  wire _23798_;
  wire _23799_;
  wire _23800_;
  wire _23801_;
  wire _23802_;
  wire _23803_;
  wire _23804_;
  wire _23805_;
  wire _23806_;
  wire _23807_;
  wire _23808_;
  wire _23809_;
  wire _23810_;
  wire _23811_;
  wire _23812_;
  wire _23813_;
  wire _23814_;
  wire _23815_;
  wire _23816_;
  wire _23817_;
  wire _23818_;
  wire _23819_;
  wire _23820_;
  wire _23821_;
  wire _23822_;
  wire _23823_;
  wire _23824_;
  wire _23825_;
  wire _23826_;
  wire _23827_;
  wire _23828_;
  wire _23829_;
  wire _23830_;
  wire _23831_;
  wire _23832_;
  wire _23833_;
  wire _23834_;
  wire _23835_;
  wire _23836_;
  wire _23837_;
  wire _23838_;
  wire _23839_;
  wire _23840_;
  wire _23841_;
  wire _23842_;
  wire _23843_;
  wire _23844_;
  wire _23845_;
  wire _23846_;
  wire _23847_;
  wire _23848_;
  wire _23849_;
  wire _23850_;
  wire _23851_;
  wire _23852_;
  wire _23853_;
  wire _23854_;
  wire _23855_;
  wire _23856_;
  wire _23857_;
  wire _23858_;
  wire _23859_;
  wire _23860_;
  wire _23861_;
  wire _23862_;
  wire _23863_;
  wire _23864_;
  wire _23865_;
  wire _23866_;
  wire _23867_;
  wire _23868_;
  wire _23869_;
  wire _23870_;
  wire _23871_;
  wire _23872_;
  wire _23873_;
  wire _23874_;
  wire _23875_;
  wire _23876_;
  wire _23877_;
  wire _23878_;
  wire _23879_;
  wire _23880_;
  wire _23881_;
  wire _23882_;
  wire _23883_;
  wire _23884_;
  wire _23885_;
  wire _23886_;
  wire _23887_;
  wire _23888_;
  wire _23889_;
  wire _23890_;
  wire _23891_;
  wire _23892_;
  wire _23893_;
  wire _23894_;
  wire _23895_;
  wire _23896_;
  wire _23897_;
  wire _23898_;
  wire _23899_;
  wire _23900_;
  wire _23901_;
  wire _23902_;
  wire _23903_;
  wire _23904_;
  wire _23905_;
  wire _23906_;
  wire _23907_;
  wire _23908_;
  wire _23909_;
  wire _23910_;
  wire _23911_;
  wire _23912_;
  wire _23913_;
  wire _23914_;
  wire _23915_;
  wire _23916_;
  wire _23917_;
  wire _23918_;
  wire _23919_;
  wire _23920_;
  wire _23921_;
  wire _23922_;
  wire _23923_;
  wire _23924_;
  wire _23925_;
  wire _23926_;
  wire _23927_;
  wire _23928_;
  wire _23929_;
  wire _23930_;
  wire _23931_;
  wire _23932_;
  wire _23933_;
  wire _23934_;
  wire _23935_;
  wire _23936_;
  wire _23937_;
  wire _23938_;
  wire _23939_;
  wire _23940_;
  wire _23941_;
  wire _23942_;
  wire _23943_;
  wire _23944_;
  wire _23945_;
  wire _23946_;
  wire _23947_;
  wire _23948_;
  wire _23949_;
  wire _23950_;
  wire _23951_;
  wire _23952_;
  wire _23953_;
  wire _23954_;
  wire _23955_;
  wire _23956_;
  wire _23957_;
  wire _23958_;
  wire _23959_;
  wire _23960_;
  wire _23961_;
  wire _23962_;
  wire _23963_;
  wire _23964_;
  wire _23965_;
  wire _23966_;
  wire _23967_;
  wire _23968_;
  wire _23969_;
  wire _23970_;
  wire _23971_;
  wire _23972_;
  wire _23973_;
  wire _23974_;
  wire _23975_;
  wire _23976_;
  wire _23977_;
  wire _23978_;
  wire _23979_;
  wire _23980_;
  wire _23981_;
  wire _23982_;
  wire _23983_;
  wire _23984_;
  wire _23985_;
  wire _23986_;
  wire _23987_;
  wire _23988_;
  wire _23989_;
  wire _23990_;
  wire _23991_;
  wire _23992_;
  wire _23993_;
  wire _23994_;
  wire _23995_;
  wire _23996_;
  wire _23997_;
  wire _23998_;
  wire _23999_;
  wire _24000_;
  wire _24001_;
  wire _24002_;
  wire _24003_;
  wire _24004_;
  wire _24005_;
  wire _24006_;
  wire _24007_;
  wire _24008_;
  wire _24009_;
  wire _24010_;
  wire _24011_;
  wire _24012_;
  wire _24013_;
  wire _24014_;
  wire _24015_;
  wire _24016_;
  wire _24017_;
  wire _24018_;
  wire _24019_;
  wire _24020_;
  wire _24021_;
  wire _24022_;
  wire _24023_;
  wire _24024_;
  wire _24025_;
  wire _24026_;
  wire _24027_;
  wire _24028_;
  wire _24029_;
  wire _24030_;
  wire _24031_;
  wire _24032_;
  wire _24033_;
  wire _24034_;
  wire _24035_;
  wire _24036_;
  wire _24037_;
  wire _24038_;
  wire _24039_;
  wire _24040_;
  wire _24041_;
  wire _24042_;
  wire _24043_;
  wire _24044_;
  wire _24045_;
  wire _24046_;
  wire _24047_;
  wire _24048_;
  wire _24049_;
  wire _24050_;
  wire _24051_;
  wire _24052_;
  wire _24053_;
  wire _24054_;
  wire _24055_;
  wire _24056_;
  wire _24057_;
  wire _24058_;
  wire _24059_;
  wire _24060_;
  wire _24061_;
  wire _24062_;
  wire _24063_;
  wire _24064_;
  wire _24065_;
  wire _24066_;
  wire _24067_;
  wire _24068_;
  wire _24069_;
  wire _24070_;
  wire _24071_;
  wire _24072_;
  wire _24073_;
  wire _24074_;
  wire _24075_;
  wire _24076_;
  wire _24077_;
  wire _24078_;
  wire _24079_;
  wire _24080_;
  wire _24081_;
  wire _24082_;
  wire _24083_;
  wire _24084_;
  wire _24085_;
  wire _24086_;
  wire _24087_;
  wire _24088_;
  wire _24089_;
  wire _24090_;
  wire _24091_;
  wire _24092_;
  wire _24093_;
  wire _24094_;
  wire _24095_;
  wire _24096_;
  wire _24097_;
  wire _24098_;
  wire _24099_;
  wire _24100_;
  wire _24101_;
  wire _24102_;
  wire _24103_;
  wire _24104_;
  wire _24105_;
  wire _24106_;
  wire _24107_;
  wire _24108_;
  wire _24109_;
  wire _24110_;
  wire _24111_;
  wire _24112_;
  wire _24113_;
  wire _24114_;
  wire _24115_;
  wire _24116_;
  wire _24117_;
  wire _24118_;
  wire _24119_;
  wire _24120_;
  wire _24121_;
  wire _24122_;
  wire _24123_;
  wire _24124_;
  wire _24125_;
  wire _24126_;
  wire _24127_;
  wire _24128_;
  wire _24129_;
  wire _24130_;
  wire _24131_;
  wire _24132_;
  wire _24133_;
  wire _24134_;
  wire _24135_;
  wire _24136_;
  wire _24137_;
  wire _24138_;
  wire _24139_;
  wire _24140_;
  wire _24141_;
  wire _24142_;
  wire _24143_;
  wire _24144_;
  wire _24145_;
  wire _24146_;
  wire _24147_;
  wire _24148_;
  wire _24149_;
  wire _24150_;
  wire _24151_;
  wire _24152_;
  wire _24153_;
  wire _24154_;
  wire _24155_;
  wire _24156_;
  wire _24157_;
  wire _24158_;
  wire _24159_;
  wire _24160_;
  wire _24161_;
  wire _24162_;
  wire _24163_;
  wire _24164_;
  wire _24165_;
  wire _24166_;
  wire _24167_;
  wire _24168_;
  wire _24169_;
  wire _24170_;
  wire _24171_;
  wire _24172_;
  wire _24173_;
  wire _24174_;
  wire _24175_;
  wire _24176_;
  wire _24177_;
  wire _24178_;
  wire _24179_;
  wire _24180_;
  wire _24181_;
  wire _24182_;
  wire _24183_;
  wire _24184_;
  wire _24185_;
  wire _24186_;
  wire _24187_;
  wire _24188_;
  wire _24189_;
  wire _24190_;
  wire _24191_;
  wire _24192_;
  wire _24193_;
  wire _24194_;
  wire _24195_;
  wire _24196_;
  wire _24197_;
  wire _24198_;
  wire _24199_;
  wire _24200_;
  wire _24201_;
  wire _24202_;
  wire _24203_;
  wire _24204_;
  wire _24205_;
  wire _24206_;
  wire _24207_;
  wire _24208_;
  wire _24209_;
  wire _24210_;
  wire _24211_;
  wire _24212_;
  wire _24213_;
  wire _24214_;
  wire _24215_;
  wire _24216_;
  wire _24217_;
  wire _24218_;
  wire _24219_;
  wire _24220_;
  wire _24221_;
  wire _24222_;
  wire _24223_;
  wire _24224_;
  wire _24225_;
  wire _24226_;
  wire _24227_;
  wire _24228_;
  wire _24229_;
  wire _24230_;
  wire _24231_;
  wire _24232_;
  wire _24233_;
  wire _24234_;
  wire _24235_;
  wire _24236_;
  wire _24237_;
  wire _24238_;
  wire _24239_;
  wire _24240_;
  wire _24241_;
  wire _24242_;
  wire _24243_;
  wire _24244_;
  wire _24245_;
  wire _24246_;
  wire _24247_;
  wire _24248_;
  wire _24249_;
  wire _24250_;
  wire _24251_;
  wire _24252_;
  wire _24253_;
  wire _24254_;
  wire _24255_;
  wire _24256_;
  wire _24257_;
  wire _24258_;
  wire _24259_;
  wire _24260_;
  wire _24261_;
  wire _24262_;
  wire _24263_;
  wire _24264_;
  wire _24265_;
  wire _24266_;
  wire _24267_;
  wire _24268_;
  wire _24269_;
  wire _24270_;
  wire _24271_;
  wire _24272_;
  wire _24273_;
  wire _24274_;
  wire _24275_;
  wire _24276_;
  wire _24277_;
  wire _24278_;
  wire _24279_;
  wire _24280_;
  wire _24281_;
  wire _24282_;
  wire _24283_;
  wire _24284_;
  wire _24285_;
  wire _24286_;
  wire _24287_;
  wire _24288_;
  wire _24289_;
  wire _24290_;
  wire _24291_;
  wire _24292_;
  wire _24293_;
  wire _24294_;
  wire _24295_;
  wire _24296_;
  wire _24297_;
  wire _24298_;
  wire _24299_;
  wire _24300_;
  wire _24301_;
  wire _24302_;
  wire _24303_;
  wire _24304_;
  wire _24305_;
  wire _24306_;
  wire _24307_;
  wire _24308_;
  wire _24309_;
  wire _24310_;
  wire _24311_;
  wire _24312_;
  wire _24313_;
  wire _24314_;
  wire _24315_;
  wire _24316_;
  wire _24317_;
  wire _24318_;
  wire _24319_;
  wire _24320_;
  wire _24321_;
  wire _24322_;
  wire _24323_;
  wire _24324_;
  wire _24325_;
  wire _24326_;
  wire _24327_;
  wire _24328_;
  wire _24329_;
  wire _24330_;
  wire _24331_;
  wire _24332_;
  wire _24333_;
  wire _24334_;
  wire _24335_;
  wire _24336_;
  wire _24337_;
  wire _24338_;
  wire _24339_;
  wire _24340_;
  wire _24341_;
  wire _24342_;
  wire _24343_;
  wire _24344_;
  wire _24345_;
  wire _24346_;
  wire _24347_;
  wire _24348_;
  wire _24349_;
  wire _24350_;
  wire _24351_;
  wire _24352_;
  wire _24353_;
  wire _24354_;
  wire _24355_;
  wire _24356_;
  wire _24357_;
  wire _24358_;
  wire _24359_;
  wire _24360_;
  wire _24361_;
  wire _24362_;
  wire _24363_;
  wire _24364_;
  wire _24365_;
  wire _24366_;
  wire _24367_;
  wire _24368_;
  wire _24369_;
  wire _24370_;
  wire _24371_;
  wire _24372_;
  wire _24373_;
  wire _24374_;
  wire _24375_;
  wire _24376_;
  wire _24377_;
  wire _24378_;
  wire _24379_;
  wire _24380_;
  wire _24381_;
  wire _24382_;
  wire _24383_;
  wire _24384_;
  wire _24385_;
  wire _24386_;
  wire _24387_;
  wire _24388_;
  wire _24389_;
  wire _24390_;
  wire _24391_;
  wire _24392_;
  wire _24393_;
  wire _24394_;
  wire _24395_;
  wire _24396_;
  wire _24397_;
  wire _24398_;
  wire _24399_;
  wire _24400_;
  wire _24401_;
  wire _24402_;
  wire _24403_;
  wire _24404_;
  wire _24405_;
  wire _24406_;
  wire _24407_;
  wire _24408_;
  wire _24409_;
  wire _24410_;
  wire _24411_;
  wire _24412_;
  wire _24413_;
  wire _24414_;
  wire _24415_;
  wire _24416_;
  wire _24417_;
  wire _24418_;
  wire _24419_;
  wire _24420_;
  wire _24421_;
  wire _24422_;
  wire _24423_;
  wire _24424_;
  wire _24425_;
  wire _24426_;
  wire _24427_;
  wire _24428_;
  wire _24429_;
  wire _24430_;
  wire _24431_;
  wire _24432_;
  wire _24433_;
  wire _24434_;
  wire _24435_;
  wire _24436_;
  wire _24437_;
  wire _24438_;
  wire _24439_;
  wire _24440_;
  wire _24441_;
  wire _24442_;
  wire _24443_;
  wire _24444_;
  wire _24445_;
  wire _24446_;
  wire _24447_;
  wire _24448_;
  wire _24449_;
  wire _24450_;
  wire _24451_;
  wire _24452_;
  wire _24453_;
  wire _24454_;
  wire _24455_;
  wire _24456_;
  wire _24457_;
  wire _24458_;
  wire _24459_;
  wire _24460_;
  wire _24461_;
  wire _24462_;
  wire _24463_;
  wire _24464_;
  wire _24465_;
  wire _24466_;
  wire _24467_;
  wire _24468_;
  wire _24469_;
  wire _24470_;
  wire _24471_;
  wire _24472_;
  wire _24473_;
  wire _24474_;
  wire _24475_;
  wire _24476_;
  wire _24477_;
  wire _24478_;
  wire _24479_;
  wire _24480_;
  wire _24481_;
  wire _24482_;
  wire _24483_;
  wire _24484_;
  wire _24485_;
  wire _24486_;
  wire _24487_;
  wire _24488_;
  wire _24489_;
  wire _24490_;
  wire _24491_;
  wire _24492_;
  wire _24493_;
  wire _24494_;
  wire _24495_;
  wire _24496_;
  wire _24497_;
  wire _24498_;
  wire _24499_;
  wire _24500_;
  wire _24501_;
  wire _24502_;
  wire _24503_;
  wire _24504_;
  wire _24505_;
  wire _24506_;
  wire _24507_;
  wire _24508_;
  wire _24509_;
  wire _24510_;
  wire _24511_;
  wire _24512_;
  wire _24513_;
  wire _24514_;
  wire _24515_;
  wire _24516_;
  wire _24517_;
  wire _24518_;
  wire _24519_;
  wire _24520_;
  wire _24521_;
  wire _24522_;
  wire _24523_;
  wire _24524_;
  wire _24525_;
  wire _24526_;
  wire _24527_;
  wire _24528_;
  wire _24529_;
  wire _24530_;
  wire _24531_;
  wire _24532_;
  wire _24533_;
  wire _24534_;
  wire _24535_;
  wire _24536_;
  wire _24537_;
  wire _24538_;
  wire _24539_;
  wire _24540_;
  wire _24541_;
  wire _24542_;
  wire _24543_;
  wire _24544_;
  wire _24545_;
  wire _24546_;
  wire _24547_;
  wire _24548_;
  wire _24549_;
  wire _24550_;
  wire _24551_;
  wire _24552_;
  wire _24553_;
  wire _24554_;
  wire _24555_;
  wire _24556_;
  wire _24557_;
  wire _24558_;
  wire _24559_;
  wire _24560_;
  wire _24561_;
  wire _24562_;
  wire _24563_;
  wire _24564_;
  wire _24565_;
  wire _24566_;
  wire _24567_;
  wire _24568_;
  wire _24569_;
  wire _24570_;
  wire _24571_;
  wire _24572_;
  wire _24573_;
  wire _24574_;
  wire _24575_;
  wire _24576_;
  wire _24577_;
  wire _24578_;
  wire _24579_;
  wire _24580_;
  wire _24581_;
  wire _24582_;
  wire _24583_;
  wire _24584_;
  wire _24585_;
  wire _24586_;
  wire _24587_;
  wire _24588_;
  wire _24589_;
  wire _24590_;
  wire _24591_;
  wire _24592_;
  wire _24593_;
  wire _24594_;
  wire _24595_;
  wire _24596_;
  wire _24597_;
  wire _24598_;
  wire _24599_;
  wire _24600_;
  wire _24601_;
  wire _24602_;
  wire _24603_;
  wire _24604_;
  wire _24605_;
  wire _24606_;
  wire _24607_;
  wire _24608_;
  wire _24609_;
  wire _24610_;
  wire _24611_;
  wire _24612_;
  wire _24613_;
  wire _24614_;
  wire _24615_;
  wire _24616_;
  wire _24617_;
  wire _24618_;
  wire _24619_;
  wire _24620_;
  wire _24621_;
  wire _24622_;
  wire _24623_;
  wire _24624_;
  wire _24625_;
  wire _24626_;
  wire _24627_;
  wire _24628_;
  wire _24629_;
  wire _24630_;
  wire _24631_;
  wire _24632_;
  wire _24633_;
  wire _24634_;
  wire _24635_;
  wire _24636_;
  wire _24637_;
  wire _24638_;
  wire _24639_;
  wire _24640_;
  wire _24641_;
  wire _24642_;
  wire _24643_;
  wire _24644_;
  wire _24645_;
  wire _24646_;
  wire _24647_;
  wire _24648_;
  wire _24649_;
  wire _24650_;
  wire _24651_;
  wire _24652_;
  wire _24653_;
  wire _24654_;
  wire _24655_;
  wire _24656_;
  wire _24657_;
  wire _24658_;
  wire _24659_;
  wire _24660_;
  wire _24661_;
  wire _24662_;
  wire _24663_;
  wire _24664_;
  wire _24665_;
  wire _24666_;
  wire _24667_;
  wire _24668_;
  wire _24669_;
  wire _24670_;
  wire _24671_;
  wire _24672_;
  wire _24673_;
  wire _24674_;
  wire _24675_;
  wire _24676_;
  wire _24677_;
  wire _24678_;
  wire _24679_;
  wire _24680_;
  wire _24681_;
  wire _24682_;
  wire _24683_;
  wire _24684_;
  wire _24685_;
  wire _24686_;
  wire _24687_;
  wire _24688_;
  wire _24689_;
  wire _24690_;
  wire _24691_;
  wire _24692_;
  wire _24693_;
  wire _24694_;
  wire _24695_;
  wire _24696_;
  wire _24697_;
  wire _24698_;
  wire _24699_;
  wire _24700_;
  wire _24701_;
  wire _24702_;
  wire _24703_;
  wire _24704_;
  wire _24705_;
  wire _24706_;
  wire _24707_;
  wire _24708_;
  wire _24709_;
  wire _24710_;
  wire _24711_;
  wire _24712_;
  wire _24713_;
  wire _24714_;
  wire _24715_;
  wire _24716_;
  wire _24717_;
  wire _24718_;
  wire _24719_;
  wire _24720_;
  wire _24721_;
  wire _24722_;
  wire _24723_;
  wire _24724_;
  wire _24725_;
  wire _24726_;
  wire _24727_;
  wire _24728_;
  wire _24729_;
  wire _24730_;
  wire _24731_;
  wire _24732_;
  wire _24733_;
  wire _24734_;
  wire _24735_;
  wire _24736_;
  wire _24737_;
  wire _24738_;
  wire _24739_;
  wire _24740_;
  wire _24741_;
  wire _24742_;
  wire _24743_;
  wire _24744_;
  wire _24745_;
  wire _24746_;
  wire _24747_;
  wire _24748_;
  wire _24749_;
  wire _24750_;
  wire _24751_;
  wire _24752_;
  wire _24753_;
  wire _24754_;
  wire _24755_;
  wire _24756_;
  wire _24757_;
  wire _24758_;
  wire _24759_;
  wire _24760_;
  wire _24761_;
  wire _24762_;
  wire _24763_;
  wire _24764_;
  wire _24765_;
  wire _24766_;
  wire _24767_;
  wire _24768_;
  wire _24769_;
  wire _24770_;
  wire _24771_;
  wire _24772_;
  wire _24773_;
  wire _24774_;
  wire _24775_;
  wire _24776_;
  wire _24777_;
  wire _24778_;
  wire _24779_;
  wire _24780_;
  wire _24781_;
  wire _24782_;
  wire _24783_;
  wire _24784_;
  wire _24785_;
  wire _24786_;
  wire _24787_;
  wire _24788_;
  wire _24789_;
  wire _24790_;
  wire _24791_;
  wire _24792_;
  wire _24793_;
  wire _24794_;
  wire _24795_;
  wire _24796_;
  wire _24797_;
  wire _24798_;
  wire _24799_;
  wire _24800_;
  wire _24801_;
  wire _24802_;
  wire _24803_;
  wire _24804_;
  wire _24805_;
  wire _24806_;
  wire _24807_;
  wire _24808_;
  wire _24809_;
  wire _24810_;
  wire _24811_;
  wire _24812_;
  wire _24813_;
  wire _24814_;
  wire _24815_;
  wire _24816_;
  wire _24817_;
  wire _24818_;
  wire _24819_;
  wire _24820_;
  wire _24821_;
  wire _24822_;
  wire _24823_;
  wire _24824_;
  wire _24825_;
  wire _24826_;
  wire _24827_;
  wire _24828_;
  wire _24829_;
  wire _24830_;
  wire _24831_;
  wire _24832_;
  wire _24833_;
  wire _24834_;
  wire _24835_;
  wire _24836_;
  wire _24837_;
  wire _24838_;
  wire _24839_;
  wire _24840_;
  wire _24841_;
  wire _24842_;
  wire _24843_;
  wire _24844_;
  wire _24845_;
  wire _24846_;
  wire _24847_;
  wire _24848_;
  wire _24849_;
  wire _24850_;
  wire _24851_;
  wire _24852_;
  wire _24853_;
  wire _24854_;
  wire _24855_;
  wire _24856_;
  wire _24857_;
  wire _24858_;
  wire _24859_;
  wire _24860_;
  wire _24861_;
  wire _24862_;
  wire _24863_;
  wire _24864_;
  wire _24865_;
  wire _24866_;
  wire _24867_;
  wire _24868_;
  wire _24869_;
  wire _24870_;
  wire _24871_;
  wire _24872_;
  wire _24873_;
  wire _24874_;
  wire _24875_;
  wire _24876_;
  wire _24877_;
  wire _24878_;
  wire _24879_;
  wire _24880_;
  wire _24881_;
  wire _24882_;
  wire _24883_;
  wire _24884_;
  wire _24885_;
  wire _24886_;
  wire _24887_;
  wire _24888_;
  wire _24889_;
  wire _24890_;
  wire _24891_;
  wire _24892_;
  wire _24893_;
  wire _24894_;
  wire _24895_;
  wire _24896_;
  wire _24897_;
  wire _24898_;
  wire _24899_;
  wire _24900_;
  wire _24901_;
  wire _24902_;
  wire _24903_;
  wire _24904_;
  wire _24905_;
  wire _24906_;
  wire _24907_;
  wire _24908_;
  wire _24909_;
  wire _24910_;
  wire _24911_;
  wire _24912_;
  wire _24913_;
  wire _24914_;
  wire _24915_;
  wire _24916_;
  wire _24917_;
  wire _24918_;
  wire _24919_;
  wire _24920_;
  wire _24921_;
  wire _24922_;
  wire _24923_;
  wire _24924_;
  wire _24925_;
  wire _24926_;
  wire _24927_;
  wire _24928_;
  wire _24929_;
  wire _24930_;
  wire _24931_;
  wire _24932_;
  wire _24933_;
  wire _24934_;
  wire _24935_;
  wire _24936_;
  wire _24937_;
  wire _24938_;
  wire _24939_;
  wire _24940_;
  wire _24941_;
  wire _24942_;
  wire _24943_;
  wire _24944_;
  wire _24945_;
  wire _24946_;
  wire _24947_;
  wire _24948_;
  wire _24949_;
  wire _24950_;
  wire _24951_;
  wire _24952_;
  wire _24953_;
  wire _24954_;
  wire _24955_;
  wire _24956_;
  wire _24957_;
  wire _24958_;
  wire _24959_;
  wire _24960_;
  wire _24961_;
  wire _24962_;
  wire _24963_;
  wire _24964_;
  wire _24965_;
  wire _24966_;
  wire _24967_;
  wire _24968_;
  wire _24969_;
  wire _24970_;
  wire _24971_;
  wire _24972_;
  wire _24973_;
  wire _24974_;
  wire _24975_;
  wire _24976_;
  wire _24977_;
  wire _24978_;
  wire _24979_;
  wire _24980_;
  wire _24981_;
  wire _24982_;
  wire _24983_;
  wire _24984_;
  wire _24985_;
  wire _24986_;
  wire _24987_;
  wire _24988_;
  wire _24989_;
  wire _24990_;
  wire _24991_;
  wire _24992_;
  wire _24993_;
  wire _24994_;
  wire _24995_;
  wire _24996_;
  wire _24997_;
  wire _24998_;
  wire _24999_;
  wire _25000_;
  wire _25001_;
  wire _25002_;
  wire _25003_;
  wire _25004_;
  wire _25005_;
  wire _25006_;
  wire _25007_;
  wire _25008_;
  wire _25009_;
  wire _25010_;
  wire _25011_;
  wire _25012_;
  wire _25013_;
  wire _25014_;
  wire _25015_;
  wire _25016_;
  wire _25017_;
  wire _25018_;
  wire _25019_;
  wire _25020_;
  wire _25021_;
  wire _25022_;
  wire _25023_;
  wire _25024_;
  wire _25025_;
  wire _25026_;
  wire _25027_;
  wire _25028_;
  wire _25029_;
  wire _25030_;
  wire _25031_;
  wire _25032_;
  wire _25033_;
  wire _25034_;
  wire _25035_;
  wire _25036_;
  wire _25037_;
  wire _25038_;
  wire _25039_;
  wire _25040_;
  wire _25041_;
  wire _25042_;
  wire _25043_;
  wire _25044_;
  wire _25045_;
  wire _25046_;
  wire _25047_;
  wire _25048_;
  wire _25049_;
  wire _25050_;
  wire _25051_;
  wire _25052_;
  wire _25053_;
  wire _25054_;
  wire _25055_;
  wire _25056_;
  wire _25057_;
  wire _25058_;
  wire _25059_;
  wire _25060_;
  wire _25061_;
  wire _25062_;
  wire _25063_;
  wire _25064_;
  wire _25065_;
  wire _25066_;
  wire _25067_;
  wire _25068_;
  wire _25069_;
  wire _25070_;
  wire _25071_;
  wire _25072_;
  wire _25073_;
  wire _25074_;
  wire _25075_;
  wire _25076_;
  wire _25077_;
  wire _25078_;
  wire _25079_;
  wire _25080_;
  wire _25081_;
  wire _25082_;
  wire _25083_;
  wire _25084_;
  wire _25085_;
  wire _25086_;
  wire _25087_;
  wire _25088_;
  wire _25089_;
  wire _25090_;
  wire _25091_;
  wire _25092_;
  wire _25093_;
  wire _25094_;
  wire _25095_;
  wire _25096_;
  wire _25097_;
  wire _25098_;
  wire _25099_;
  wire _25100_;
  wire _25101_;
  wire _25102_;
  wire _25103_;
  wire _25104_;
  wire _25105_;
  wire _25106_;
  wire _25107_;
  wire _25108_;
  wire _25109_;
  wire _25110_;
  wire _25111_;
  wire _25112_;
  wire _25113_;
  wire _25114_;
  wire _25115_;
  wire _25116_;
  wire _25117_;
  wire _25118_;
  wire _25119_;
  wire _25120_;
  wire _25121_;
  wire _25122_;
  wire _25123_;
  wire _25124_;
  wire _25125_;
  wire _25126_;
  wire _25127_;
  wire _25128_;
  wire _25129_;
  wire _25130_;
  wire _25131_;
  wire _25132_;
  wire _25133_;
  wire _25134_;
  wire _25135_;
  wire _25136_;
  wire _25137_;
  wire _25138_;
  wire _25139_;
  wire _25140_;
  wire _25141_;
  wire _25142_;
  wire _25143_;
  wire _25144_;
  wire _25145_;
  wire _25146_;
  wire _25147_;
  wire _25148_;
  wire _25149_;
  wire _25150_;
  wire _25151_;
  wire _25152_;
  wire _25153_;
  wire _25154_;
  wire _25155_;
  wire _25156_;
  wire _25157_;
  wire _25158_;
  wire _25159_;
  wire _25160_;
  wire _25161_;
  wire _25162_;
  wire _25163_;
  wire _25164_;
  wire _25165_;
  wire _25166_;
  wire _25167_;
  wire _25168_;
  wire _25169_;
  wire _25170_;
  wire _25171_;
  wire _25172_;
  wire _25173_;
  wire _25174_;
  wire _25175_;
  wire _25176_;
  wire _25177_;
  wire _25178_;
  wire _25179_;
  wire _25180_;
  wire _25181_;
  wire _25182_;
  wire _25183_;
  wire _25184_;
  wire _25185_;
  wire _25186_;
  wire _25187_;
  wire _25188_;
  wire _25189_;
  wire _25190_;
  wire _25191_;
  wire _25192_;
  wire _25193_;
  wire _25194_;
  wire _25195_;
  wire _25196_;
  wire _25197_;
  wire _25198_;
  wire _25199_;
  wire _25200_;
  wire _25201_;
  wire _25202_;
  wire _25203_;
  wire _25204_;
  wire _25205_;
  wire _25206_;
  wire _25207_;
  wire _25208_;
  wire _25209_;
  wire _25210_;
  wire _25211_;
  wire _25212_;
  wire _25213_;
  wire _25214_;
  wire _25215_;
  wire _25216_;
  wire _25217_;
  wire _25218_;
  wire _25219_;
  wire _25220_;
  wire _25221_;
  wire _25222_;
  wire _25223_;
  wire _25224_;
  wire _25225_;
  wire _25226_;
  wire _25227_;
  wire _25228_;
  wire _25229_;
  wire _25230_;
  wire _25231_;
  wire _25232_;
  wire _25233_;
  wire _25234_;
  wire _25235_;
  wire _25236_;
  wire _25237_;
  wire _25238_;
  wire _25239_;
  wire _25240_;
  wire _25241_;
  wire _25242_;
  wire _25243_;
  wire _25244_;
  wire _25245_;
  wire _25246_;
  wire _25247_;
  wire _25248_;
  wire _25249_;
  wire _25250_;
  wire _25251_;
  wire _25252_;
  wire _25253_;
  wire _25254_;
  wire _25255_;
  wire _25256_;
  wire _25257_;
  wire _25258_;
  wire _25259_;
  wire _25260_;
  wire _25261_;
  wire _25262_;
  wire _25263_;
  wire _25264_;
  wire _25265_;
  wire _25266_;
  wire _25267_;
  wire _25268_;
  wire _25269_;
  wire _25270_;
  wire _25271_;
  wire _25272_;
  wire _25273_;
  wire _25274_;
  wire _25275_;
  wire _25276_;
  wire _25277_;
  wire _25278_;
  wire _25279_;
  wire _25280_;
  wire _25281_;
  wire _25282_;
  wire _25283_;
  wire _25284_;
  wire _25285_;
  wire _25286_;
  wire _25287_;
  wire _25288_;
  wire _25289_;
  wire _25290_;
  wire _25291_;
  wire _25292_;
  wire _25293_;
  wire _25294_;
  wire _25295_;
  wire _25296_;
  wire _25297_;
  wire _25298_;
  wire _25299_;
  wire _25300_;
  wire _25301_;
  wire _25302_;
  wire _25303_;
  wire _25304_;
  wire _25305_;
  wire _25306_;
  wire _25307_;
  wire _25308_;
  wire _25309_;
  wire _25310_;
  wire _25311_;
  wire _25312_;
  wire _25313_;
  wire _25314_;
  wire _25315_;
  wire _25316_;
  wire _25317_;
  wire _25318_;
  wire _25319_;
  wire _25320_;
  wire _25321_;
  wire _25322_;
  wire _25323_;
  wire _25324_;
  wire _25325_;
  wire _25326_;
  wire _25327_;
  wire _25328_;
  wire _25329_;
  wire _25330_;
  wire _25331_;
  wire _25332_;
  wire _25333_;
  wire _25334_;
  wire _25335_;
  wire _25336_;
  wire _25337_;
  wire _25338_;
  wire _25339_;
  wire _25340_;
  wire _25341_;
  wire _25342_;
  wire _25343_;
  wire _25344_;
  wire _25345_;
  wire _25346_;
  wire _25347_;
  wire _25348_;
  wire _25349_;
  wire _25350_;
  wire _25351_;
  wire _25352_;
  wire _25353_;
  wire _25354_;
  wire _25355_;
  wire _25356_;
  wire _25357_;
  wire _25358_;
  wire _25359_;
  wire _25360_;
  wire _25361_;
  wire _25362_;
  wire _25363_;
  wire _25364_;
  wire _25365_;
  wire _25366_;
  wire _25367_;
  wire _25368_;
  wire _25369_;
  wire _25370_;
  wire _25371_;
  wire _25372_;
  wire _25373_;
  wire _25374_;
  wire _25375_;
  wire _25376_;
  wire _25377_;
  wire _25378_;
  wire _25379_;
  wire _25380_;
  wire _25381_;
  wire _25382_;
  wire _25383_;
  wire _25384_;
  wire _25385_;
  wire _25386_;
  wire _25387_;
  wire _25388_;
  wire _25389_;
  wire _25390_;
  wire _25391_;
  wire _25392_;
  wire _25393_;
  wire _25394_;
  wire _25395_;
  wire _25396_;
  wire _25397_;
  wire _25398_;
  wire _25399_;
  wire _25400_;
  wire _25401_;
  wire _25402_;
  wire _25403_;
  wire _25404_;
  wire _25405_;
  wire _25406_;
  wire _25407_;
  wire _25408_;
  wire _25409_;
  wire _25410_;
  wire _25411_;
  wire _25412_;
  wire _25413_;
  wire _25414_;
  wire _25415_;
  wire _25416_;
  wire _25417_;
  wire _25418_;
  wire _25419_;
  wire _25420_;
  wire _25421_;
  wire _25422_;
  wire _25423_;
  wire _25424_;
  wire _25425_;
  wire _25426_;
  wire _25427_;
  wire _25428_;
  wire _25429_;
  wire _25430_;
  wire _25431_;
  wire _25432_;
  wire _25433_;
  wire _25434_;
  wire _25435_;
  wire _25436_;
  wire _25437_;
  wire _25438_;
  wire _25439_;
  wire _25440_;
  wire _25441_;
  wire _25442_;
  wire _25443_;
  wire _25444_;
  wire _25445_;
  wire _25446_;
  wire _25447_;
  wire _25448_;
  wire _25449_;
  wire _25450_;
  wire _25451_;
  wire _25452_;
  wire _25453_;
  wire _25454_;
  wire _25455_;
  wire _25456_;
  wire _25457_;
  wire _25458_;
  wire _25459_;
  wire _25460_;
  wire _25461_;
  wire _25462_;
  wire _25463_;
  wire _25464_;
  wire _25465_;
  wire _25466_;
  wire _25467_;
  wire _25468_;
  wire _25469_;
  wire _25470_;
  wire _25471_;
  wire _25472_;
  wire _25473_;
  wire _25474_;
  wire _25475_;
  wire _25476_;
  wire _25477_;
  wire _25478_;
  wire _25479_;
  wire _25480_;
  wire _25481_;
  wire _25482_;
  wire _25483_;
  wire _25484_;
  wire _25485_;
  wire _25486_;
  wire _25487_;
  wire _25488_;
  wire _25489_;
  wire _25490_;
  wire _25491_;
  wire _25492_;
  wire _25493_;
  wire _25494_;
  wire _25495_;
  wire _25496_;
  wire _25497_;
  wire _25498_;
  wire _25499_;
  wire _25500_;
  wire _25501_;
  wire _25502_;
  wire _25503_;
  wire _25504_;
  wire _25505_;
  wire _25506_;
  wire _25507_;
  wire _25508_;
  wire _25509_;
  wire _25510_;
  wire _25511_;
  wire _25512_;
  wire _25513_;
  wire _25514_;
  wire _25515_;
  wire _25516_;
  wire _25517_;
  wire _25518_;
  wire _25519_;
  wire _25520_;
  wire _25521_;
  wire _25522_;
  wire _25523_;
  wire _25524_;
  wire _25525_;
  wire _25526_;
  wire _25527_;
  wire _25528_;
  wire _25529_;
  wire _25530_;
  wire _25531_;
  wire _25532_;
  wire _25533_;
  wire _25534_;
  wire _25535_;
  wire _25536_;
  wire _25537_;
  wire _25538_;
  wire _25539_;
  wire _25540_;
  wire _25541_;
  wire _25542_;
  wire _25543_;
  wire _25544_;
  wire _25545_;
  wire _25546_;
  wire _25547_;
  wire _25548_;
  wire _25549_;
  wire _25550_;
  wire _25551_;
  wire _25552_;
  wire _25553_;
  wire _25554_;
  wire _25555_;
  wire _25556_;
  wire _25557_;
  wire _25558_;
  wire _25559_;
  wire _25560_;
  wire _25561_;
  wire _25562_;
  wire _25563_;
  wire _25564_;
  wire _25565_;
  wire _25566_;
  wire _25567_;
  wire _25568_;
  wire _25569_;
  wire _25570_;
  wire _25571_;
  wire _25572_;
  wire _25573_;
  wire _25574_;
  wire _25575_;
  wire _25576_;
  wire _25577_;
  wire _25578_;
  wire _25579_;
  wire _25580_;
  wire _25581_;
  wire _25582_;
  wire _25583_;
  wire _25584_;
  wire _25585_;
  wire _25586_;
  wire _25587_;
  wire _25588_;
  wire _25589_;
  wire _25590_;
  wire _25591_;
  wire _25592_;
  wire _25593_;
  wire _25594_;
  wire _25595_;
  wire _25596_;
  wire _25597_;
  wire _25598_;
  wire _25599_;
  wire _25600_;
  wire _25601_;
  wire _25602_;
  wire _25603_;
  wire _25604_;
  wire _25605_;
  wire _25606_;
  wire _25607_;
  wire _25608_;
  wire _25609_;
  wire _25610_;
  wire _25611_;
  wire _25612_;
  wire _25613_;
  wire _25614_;
  wire _25615_;
  wire _25616_;
  wire _25617_;
  wire _25618_;
  wire _25619_;
  wire _25620_;
  wire _25621_;
  wire _25622_;
  wire _25623_;
  wire _25624_;
  wire _25625_;
  wire _25626_;
  wire _25627_;
  wire _25628_;
  wire _25629_;
  wire _25630_;
  wire _25631_;
  wire _25632_;
  wire _25633_;
  wire _25634_;
  wire _25635_;
  wire _25636_;
  wire _25637_;
  wire _25638_;
  wire _25639_;
  wire _25640_;
  wire _25641_;
  wire _25642_;
  wire _25643_;
  wire _25644_;
  wire _25645_;
  wire _25646_;
  wire _25647_;
  wire _25648_;
  wire _25649_;
  wire _25650_;
  wire _25651_;
  wire _25652_;
  wire _25653_;
  wire _25654_;
  wire _25655_;
  wire _25656_;
  wire _25657_;
  wire _25658_;
  wire _25659_;
  wire _25660_;
  wire _25661_;
  wire _25662_;
  wire _25663_;
  wire _25664_;
  wire _25665_;
  wire _25666_;
  wire _25667_;
  wire _25668_;
  wire _25669_;
  wire _25670_;
  wire _25671_;
  wire _25672_;
  wire _25673_;
  wire _25674_;
  wire _25675_;
  wire _25676_;
  wire _25677_;
  wire _25678_;
  wire _25679_;
  wire _25680_;
  wire _25681_;
  wire _25682_;
  wire _25683_;
  wire _25684_;
  wire _25685_;
  wire _25686_;
  wire _25687_;
  wire _25688_;
  wire _25689_;
  wire _25690_;
  wire _25691_;
  wire _25692_;
  wire _25693_;
  wire _25694_;
  wire _25695_;
  wire _25696_;
  wire _25697_;
  wire _25698_;
  wire _25699_;
  wire _25700_;
  wire _25701_;
  wire _25702_;
  wire _25703_;
  wire _25704_;
  wire _25705_;
  wire _25706_;
  wire _25707_;
  wire _25708_;
  wire _25709_;
  wire _25710_;
  wire _25711_;
  wire _25712_;
  wire _25713_;
  wire _25714_;
  wire _25715_;
  wire _25716_;
  wire _25717_;
  wire _25718_;
  wire _25719_;
  wire _25720_;
  wire _25721_;
  wire _25722_;
  wire _25723_;
  wire _25724_;
  wire _25725_;
  wire _25726_;
  wire _25727_;
  wire _25728_;
  wire _25729_;
  wire _25730_;
  wire _25731_;
  wire _25732_;
  wire _25733_;
  wire _25734_;
  wire _25735_;
  wire _25736_;
  wire _25737_;
  wire _25738_;
  wire _25739_;
  wire _25740_;
  wire _25741_;
  wire _25742_;
  wire _25743_;
  wire _25744_;
  wire _25745_;
  wire _25746_;
  wire _25747_;
  wire _25748_;
  wire _25749_;
  wire _25750_;
  wire _25751_;
  wire _25752_;
  wire _25753_;
  wire _25754_;
  wire _25755_;
  wire _25756_;
  wire _25757_;
  wire _25758_;
  wire _25759_;
  wire _25760_;
  wire _25761_;
  wire _25762_;
  wire _25763_;
  wire _25764_;
  wire _25765_;
  wire _25766_;
  wire _25767_;
  wire _25768_;
  wire _25769_;
  wire _25770_;
  wire _25771_;
  wire _25772_;
  wire _25773_;
  wire _25774_;
  wire _25775_;
  wire _25776_;
  wire _25777_;
  wire _25778_;
  wire _25779_;
  wire _25780_;
  wire _25781_;
  wire _25782_;
  wire _25783_;
  wire _25784_;
  wire _25785_;
  wire _25786_;
  wire _25787_;
  wire _25788_;
  wire _25789_;
  wire _25790_;
  wire _25791_;
  wire _25792_;
  wire _25793_;
  wire _25794_;
  wire _25795_;
  wire _25796_;
  wire _25797_;
  wire _25798_;
  wire _25799_;
  wire _25800_;
  wire _25801_;
  wire _25802_;
  wire _25803_;
  wire _25804_;
  wire _25805_;
  wire _25806_;
  wire _25807_;
  wire _25808_;
  wire _25809_;
  wire _25810_;
  wire _25811_;
  wire _25812_;
  wire _25813_;
  wire _25814_;
  wire _25815_;
  wire _25816_;
  wire _25817_;
  wire _25818_;
  wire _25819_;
  wire _25820_;
  wire _25821_;
  wire _25822_;
  wire _25823_;
  wire _25824_;
  wire _25825_;
  wire _25826_;
  wire _25827_;
  wire _25828_;
  wire _25829_;
  wire _25830_;
  wire _25831_;
  wire _25832_;
  wire _25833_;
  wire _25834_;
  wire _25835_;
  wire _25836_;
  wire _25837_;
  wire _25838_;
  wire _25839_;
  wire _25840_;
  wire _25841_;
  wire _25842_;
  wire _25843_;
  wire _25844_;
  wire _25845_;
  wire _25846_;
  wire _25847_;
  wire _25848_;
  wire _25849_;
  wire _25850_;
  wire _25851_;
  wire _25852_;
  wire _25853_;
  wire _25854_;
  wire _25855_;
  wire _25856_;
  wire _25857_;
  wire _25858_;
  wire _25859_;
  wire _25860_;
  wire _25861_;
  wire _25862_;
  wire _25863_;
  wire _25864_;
  wire _25865_;
  wire _25866_;
  wire _25867_;
  wire _25868_;
  wire _25869_;
  wire _25870_;
  wire _25871_;
  wire _25872_;
  wire _25873_;
  wire _25874_;
  wire _25875_;
  wire _25876_;
  wire _25877_;
  wire _25878_;
  wire _25879_;
  wire _25880_;
  wire _25881_;
  wire _25882_;
  wire _25883_;
  wire _25884_;
  wire _25885_;
  wire _25886_;
  wire _25887_;
  wire _25888_;
  wire _25889_;
  wire _25890_;
  wire _25891_;
  wire _25892_;
  wire _25893_;
  wire _25894_;
  wire _25895_;
  wire _25896_;
  wire _25897_;
  wire _25898_;
  wire _25899_;
  wire _25900_;
  wire _25901_;
  wire _25902_;
  wire _25903_;
  wire _25904_;
  wire _25905_;
  wire _25906_;
  wire _25907_;
  wire _25908_;
  wire _25909_;
  wire _25910_;
  wire _25911_;
  wire _25912_;
  wire _25913_;
  wire _25914_;
  wire _25915_;
  wire _25916_;
  wire _25917_;
  wire _25918_;
  wire _25919_;
  wire _25920_;
  wire _25921_;
  wire _25922_;
  wire _25923_;
  wire _25924_;
  wire _25925_;
  wire _25926_;
  wire _25927_;
  wire _25928_;
  wire _25929_;
  wire _25930_;
  wire _25931_;
  wire _25932_;
  wire _25933_;
  wire _25934_;
  wire _25935_;
  wire _25936_;
  wire _25937_;
  wire _25938_;
  wire _25939_;
  wire _25940_;
  wire _25941_;
  wire _25942_;
  wire _25943_;
  wire _25944_;
  wire _25945_;
  wire _25946_;
  wire _25947_;
  wire _25948_;
  wire _25949_;
  wire _25950_;
  wire _25951_;
  wire _25952_;
  wire _25953_;
  wire _25954_;
  wire _25955_;
  wire _25956_;
  wire _25957_;
  wire _25958_;
  wire _25959_;
  wire _25960_;
  wire _25961_;
  wire _25962_;
  wire _25963_;
  wire _25964_;
  wire _25965_;
  wire _25966_;
  wire _25967_;
  wire _25968_;
  wire _25969_;
  wire _25970_;
  wire _25971_;
  wire _25972_;
  wire _25973_;
  wire _25974_;
  wire _25975_;
  wire _25976_;
  wire _25977_;
  wire _25978_;
  wire _25979_;
  wire _25980_;
  wire _25981_;
  wire _25982_;
  wire _25983_;
  wire _25984_;
  wire _25985_;
  wire _25986_;
  wire _25987_;
  wire _25988_;
  wire _25989_;
  wire _25990_;
  wire _25991_;
  wire _25992_;
  wire _25993_;
  wire _25994_;
  wire _25995_;
  wire _25996_;
  wire _25997_;
  wire _25998_;
  wire _25999_;
  wire _26000_;
  wire _26001_;
  wire _26002_;
  wire _26003_;
  wire _26004_;
  wire _26005_;
  wire _26006_;
  wire _26007_;
  wire _26008_;
  wire _26009_;
  wire _26010_;
  wire _26011_;
  wire _26012_;
  wire _26013_;
  wire _26014_;
  wire _26015_;
  wire _26016_;
  wire _26017_;
  wire _26018_;
  wire _26019_;
  wire _26020_;
  wire _26021_;
  wire _26022_;
  wire _26023_;
  wire _26024_;
  wire _26025_;
  wire _26026_;
  wire _26027_;
  wire _26028_;
  wire _26029_;
  wire _26030_;
  wire _26031_;
  wire _26032_;
  wire _26033_;
  wire _26034_;
  wire _26035_;
  wire _26036_;
  wire _26037_;
  wire _26038_;
  wire _26039_;
  wire _26040_;
  wire _26041_;
  wire _26042_;
  wire _26043_;
  wire _26044_;
  wire _26045_;
  wire _26046_;
  wire _26047_;
  wire _26048_;
  wire _26049_;
  wire _26050_;
  wire _26051_;
  wire _26052_;
  wire _26053_;
  wire _26054_;
  wire _26055_;
  wire _26056_;
  wire _26057_;
  wire _26058_;
  wire _26059_;
  wire _26060_;
  wire _26061_;
  wire _26062_;
  wire _26063_;
  wire _26064_;
  wire _26065_;
  wire _26066_;
  wire _26067_;
  wire _26068_;
  wire _26069_;
  wire _26070_;
  wire _26071_;
  wire _26072_;
  wire _26073_;
  wire _26074_;
  wire _26075_;
  wire _26076_;
  wire _26077_;
  wire _26078_;
  wire _26079_;
  wire _26080_;
  wire _26081_;
  wire _26082_;
  wire _26083_;
  wire _26084_;
  wire _26085_;
  wire _26086_;
  wire _26087_;
  wire _26088_;
  wire _26089_;
  wire _26090_;
  wire _26091_;
  wire _26092_;
  wire _26093_;
  wire _26094_;
  wire _26095_;
  wire _26096_;
  wire _26097_;
  wire _26098_;
  wire _26099_;
  wire _26100_;
  wire _26101_;
  wire _26102_;
  wire _26103_;
  wire _26104_;
  wire _26105_;
  wire _26106_;
  wire _26107_;
  wire _26108_;
  wire _26109_;
  wire _26110_;
  wire _26111_;
  wire _26112_;
  wire _26113_;
  wire _26114_;
  wire _26115_;
  wire _26116_;
  wire _26117_;
  wire _26118_;
  wire _26119_;
  wire _26120_;
  wire _26121_;
  wire _26122_;
  wire _26123_;
  wire _26124_;
  wire _26125_;
  wire _26126_;
  wire _26127_;
  wire _26128_;
  wire _26129_;
  wire _26130_;
  wire _26131_;
  wire _26132_;
  wire _26133_;
  wire _26134_;
  wire _26135_;
  wire _26136_;
  wire _26137_;
  wire _26138_;
  wire _26139_;
  wire _26140_;
  wire _26141_;
  wire _26142_;
  wire _26143_;
  wire _26144_;
  wire _26145_;
  wire _26146_;
  wire _26147_;
  wire _26148_;
  wire _26149_;
  wire _26150_;
  wire _26151_;
  wire _26152_;
  wire _26153_;
  wire _26154_;
  wire _26155_;
  wire _26156_;
  wire _26157_;
  wire _26158_;
  wire _26159_;
  wire _26160_;
  wire _26161_;
  wire _26162_;
  wire _26163_;
  wire _26164_;
  wire _26165_;
  wire _26166_;
  wire _26167_;
  wire _26168_;
  wire _26169_;
  wire _26170_;
  wire _26171_;
  wire _26172_;
  wire _26173_;
  wire _26174_;
  wire _26175_;
  wire _26176_;
  wire _26177_;
  wire _26178_;
  wire _26179_;
  wire _26180_;
  wire _26181_;
  wire _26182_;
  wire _26183_;
  wire _26184_;
  wire _26185_;
  wire _26186_;
  wire _26187_;
  wire _26188_;
  wire _26189_;
  wire _26190_;
  wire _26191_;
  wire _26192_;
  wire _26193_;
  wire _26194_;
  wire _26195_;
  wire _26196_;
  wire _26197_;
  wire _26198_;
  wire _26199_;
  wire _26200_;
  wire _26201_;
  wire _26202_;
  wire _26203_;
  wire _26204_;
  wire _26205_;
  wire _26206_;
  wire _26207_;
  wire _26208_;
  wire _26209_;
  wire _26210_;
  wire _26211_;
  wire _26212_;
  wire _26213_;
  wire _26214_;
  wire _26215_;
  wire _26216_;
  wire _26217_;
  wire _26218_;
  wire _26219_;
  wire _26220_;
  wire _26221_;
  wire _26222_;
  wire _26223_;
  wire _26224_;
  wire _26225_;
  wire _26226_;
  wire _26227_;
  wire _26228_;
  wire _26229_;
  wire _26230_;
  wire _26231_;
  wire _26232_;
  wire _26233_;
  wire _26234_;
  wire _26235_;
  wire _26236_;
  wire _26237_;
  wire _26238_;
  wire _26239_;
  wire _26240_;
  wire _26241_;
  wire _26242_;
  wire _26243_;
  wire _26244_;
  wire _26245_;
  wire _26246_;
  wire _26247_;
  wire _26248_;
  wire _26249_;
  wire _26250_;
  wire _26251_;
  wire _26252_;
  wire _26253_;
  wire _26254_;
  wire _26255_;
  wire _26256_;
  wire _26257_;
  wire _26258_;
  wire _26259_;
  wire _26260_;
  wire _26261_;
  wire _26262_;
  wire _26263_;
  wire _26264_;
  wire _26265_;
  wire _26266_;
  wire _26267_;
  wire _26268_;
  wire _26269_;
  wire _26270_;
  wire _26271_;
  wire _26272_;
  wire _26273_;
  wire _26274_;
  wire _26275_;
  wire _26276_;
  wire _26277_;
  wire _26278_;
  wire _26279_;
  wire _26280_;
  wire _26281_;
  wire _26282_;
  wire _26283_;
  wire _26284_;
  wire _26285_;
  wire _26286_;
  wire _26287_;
  wire _26288_;
  wire _26289_;
  wire _26290_;
  wire _26291_;
  wire _26292_;
  wire _26293_;
  wire _26294_;
  wire _26295_;
  wire _26296_;
  wire _26297_;
  wire _26298_;
  wire _26299_;
  wire _26300_;
  wire _26301_;
  wire _26302_;
  wire _26303_;
  wire _26304_;
  wire _26305_;
  wire _26306_;
  wire _26307_;
  wire _26308_;
  wire _26309_;
  wire _26310_;
  wire _26311_;
  wire _26312_;
  wire _26313_;
  wire _26314_;
  wire _26315_;
  wire _26316_;
  wire _26317_;
  wire _26318_;
  wire _26319_;
  wire _26320_;
  wire _26321_;
  wire _26322_;
  wire _26323_;
  wire _26324_;
  wire _26325_;
  wire _26326_;
  wire _26327_;
  wire _26328_;
  wire _26329_;
  wire _26330_;
  wire _26331_;
  wire _26332_;
  wire _26333_;
  wire _26334_;
  wire _26335_;
  wire _26336_;
  wire _26337_;
  wire _26338_;
  wire _26339_;
  wire _26340_;
  wire _26341_;
  wire _26342_;
  wire _26343_;
  wire _26344_;
  wire _26345_;
  wire _26346_;
  wire _26347_;
  wire _26348_;
  wire _26349_;
  wire _26350_;
  wire _26351_;
  wire _26352_;
  wire _26353_;
  wire _26354_;
  wire _26355_;
  wire _26356_;
  wire _26357_;
  wire _26358_;
  wire _26359_;
  wire _26360_;
  wire _26361_;
  wire _26362_;
  wire _26363_;
  wire _26364_;
  wire _26365_;
  wire _26366_;
  wire _26367_;
  wire _26368_;
  wire _26369_;
  wire _26370_;
  wire _26371_;
  wire _26372_;
  wire _26373_;
  wire _26374_;
  wire _26375_;
  wire _26376_;
  wire _26377_;
  wire _26378_;
  wire _26379_;
  wire _26380_;
  wire _26381_;
  wire _26382_;
  wire _26383_;
  wire _26384_;
  wire _26385_;
  wire _26386_;
  wire _26387_;
  wire _26388_;
  wire _26389_;
  wire _26390_;
  wire _26391_;
  wire _26392_;
  wire _26393_;
  wire _26394_;
  wire _26395_;
  wire _26396_;
  wire _26397_;
  wire _26398_;
  wire _26399_;
  wire _26400_;
  wire _26401_;
  wire _26402_;
  wire _26403_;
  wire _26404_;
  wire _26405_;
  wire _26406_;
  wire _26407_;
  wire _26408_;
  wire _26409_;
  wire _26410_;
  wire _26411_;
  wire _26412_;
  wire _26413_;
  wire _26414_;
  wire _26415_;
  wire _26416_;
  wire _26417_;
  wire _26418_;
  wire _26419_;
  wire _26420_;
  wire _26421_;
  wire _26422_;
  wire _26423_;
  wire _26424_;
  wire _26425_;
  wire _26426_;
  wire _26427_;
  wire _26428_;
  wire _26429_;
  wire _26430_;
  wire _26431_;
  wire _26432_;
  wire _26433_;
  wire _26434_;
  wire _26435_;
  wire _26436_;
  wire _26437_;
  wire _26438_;
  wire _26439_;
  wire _26440_;
  wire _26441_;
  wire _26442_;
  wire _26443_;
  wire _26444_;
  wire _26445_;
  wire _26446_;
  wire _26447_;
  wire _26448_;
  wire _26449_;
  wire _26450_;
  wire _26451_;
  wire _26452_;
  wire _26453_;
  wire _26454_;
  wire _26455_;
  wire _26456_;
  wire _26457_;
  wire _26458_;
  wire _26459_;
  wire _26460_;
  wire _26461_;
  wire _26462_;
  wire _26463_;
  wire _26464_;
  wire _26465_;
  wire _26466_;
  wire _26467_;
  wire _26468_;
  wire _26469_;
  wire _26470_;
  wire _26471_;
  wire _26472_;
  wire _26473_;
  wire _26474_;
  wire _26475_;
  wire _26476_;
  wire _26477_;
  wire _26478_;
  wire _26479_;
  wire _26480_;
  wire _26481_;
  wire _26482_;
  wire _26483_;
  wire _26484_;
  wire _26485_;
  wire _26486_;
  wire _26487_;
  wire _26488_;
  wire _26489_;
  wire _26490_;
  wire _26491_;
  wire _26492_;
  wire _26493_;
  wire _26494_;
  wire _26495_;
  wire _26496_;
  wire _26497_;
  wire _26498_;
  wire _26499_;
  wire _26500_;
  wire _26501_;
  wire _26502_;
  wire _26503_;
  wire _26504_;
  wire _26505_;
  wire _26506_;
  wire _26507_;
  wire _26508_;
  wire _26509_;
  wire _26510_;
  wire _26511_;
  wire _26512_;
  wire _26513_;
  wire _26514_;
  wire _26515_;
  wire _26516_;
  wire _26517_;
  wire _26518_;
  wire _26519_;
  wire _26520_;
  wire _26521_;
  wire _26522_;
  wire _26523_;
  wire _26524_;
  wire _26525_;
  wire _26526_;
  wire _26527_;
  wire _26528_;
  wire _26529_;
  wire _26530_;
  wire _26531_;
  wire _26532_;
  wire _26533_;
  wire _26534_;
  wire _26535_;
  wire _26536_;
  wire _26537_;
  wire _26538_;
  wire _26539_;
  wire _26540_;
  wire _26541_;
  wire _26542_;
  wire _26543_;
  wire _26544_;
  wire _26545_;
  wire _26546_;
  wire _26547_;
  wire _26548_;
  wire _26549_;
  wire _26550_;
  wire _26551_;
  wire _26552_;
  wire _26553_;
  wire _26554_;
  wire _26555_;
  wire _26556_;
  wire _26557_;
  wire _26558_;
  wire _26559_;
  wire _26560_;
  wire _26561_;
  wire _26562_;
  wire _26563_;
  wire _26564_;
  wire _26565_;
  wire _26566_;
  wire _26567_;
  wire _26568_;
  wire _26569_;
  wire _26570_;
  wire _26571_;
  wire _26572_;
  wire _26573_;
  wire _26574_;
  wire _26575_;
  wire _26576_;
  wire _26577_;
  wire _26578_;
  wire _26579_;
  wire _26580_;
  wire _26581_;
  wire _26582_;
  wire _26583_;
  wire _26584_;
  wire _26585_;
  wire _26586_;
  wire _26587_;
  wire _26588_;
  wire _26589_;
  wire _26590_;
  wire _26591_;
  wire _26592_;
  wire _26593_;
  wire _26594_;
  wire _26595_;
  wire _26596_;
  wire _26597_;
  wire _26598_;
  wire _26599_;
  wire _26600_;
  wire _26601_;
  wire _26602_;
  wire _26603_;
  wire _26604_;
  wire _26605_;
  wire _26606_;
  wire _26607_;
  wire _26608_;
  wire _26609_;
  wire _26610_;
  wire _26611_;
  wire _26612_;
  wire _26613_;
  wire _26614_;
  wire _26615_;
  wire _26616_;
  wire _26617_;
  wire _26618_;
  wire _26619_;
  wire _26620_;
  wire _26621_;
  wire _26622_;
  wire _26623_;
  wire _26624_;
  wire _26625_;
  wire _26626_;
  wire _26627_;
  wire _26628_;
  wire _26629_;
  wire _26630_;
  wire _26631_;
  wire _26632_;
  wire _26633_;
  wire _26634_;
  wire _26635_;
  wire _26636_;
  wire _26637_;
  wire _26638_;
  wire _26639_;
  wire _26640_;
  wire _26641_;
  wire _26642_;
  wire _26643_;
  wire _26644_;
  wire _26645_;
  wire _26646_;
  wire _26647_;
  wire _26648_;
  wire _26649_;
  wire _26650_;
  wire _26651_;
  wire _26652_;
  wire _26653_;
  wire _26654_;
  wire _26655_;
  wire _26656_;
  wire _26657_;
  wire _26658_;
  wire _26659_;
  wire _26660_;
  wire _26661_;
  wire _26662_;
  wire _26663_;
  wire _26664_;
  wire _26665_;
  wire _26666_;
  wire _26667_;
  wire _26668_;
  wire _26669_;
  wire _26670_;
  wire _26671_;
  wire _26672_;
  wire _26673_;
  wire _26674_;
  wire _26675_;
  wire _26676_;
  wire _26677_;
  wire _26678_;
  wire _26679_;
  wire _26680_;
  wire _26681_;
  wire _26682_;
  wire _26683_;
  wire _26684_;
  wire _26685_;
  wire _26686_;
  wire _26687_;
  wire _26688_;
  wire _26689_;
  wire _26690_;
  wire _26691_;
  wire _26692_;
  wire _26693_;
  wire _26694_;
  wire _26695_;
  wire _26696_;
  wire _26697_;
  wire _26698_;
  wire _26699_;
  wire _26700_;
  wire _26701_;
  wire _26702_;
  wire _26703_;
  wire _26704_;
  wire _26705_;
  wire _26706_;
  wire _26707_;
  wire _26708_;
  wire _26709_;
  wire _26710_;
  wire _26711_;
  wire _26712_;
  wire _26713_;
  wire _26714_;
  wire _26715_;
  wire _26716_;
  wire _26717_;
  wire _26718_;
  wire _26719_;
  wire _26720_;
  wire _26721_;
  wire _26722_;
  wire _26723_;
  wire _26724_;
  wire _26725_;
  wire _26726_;
  wire _26727_;
  wire _26728_;
  wire _26729_;
  wire _26730_;
  wire _26731_;
  wire _26732_;
  wire _26733_;
  wire _26734_;
  wire _26735_;
  wire _26736_;
  wire _26737_;
  wire _26738_;
  wire _26739_;
  wire _26740_;
  wire _26741_;
  wire _26742_;
  wire _26743_;
  wire _26744_;
  wire _26745_;
  wire _26746_;
  wire _26747_;
  wire _26748_;
  wire _26749_;
  wire _26750_;
  wire _26751_;
  wire _26752_;
  wire _26753_;
  wire _26754_;
  wire _26755_;
  wire _26756_;
  wire _26757_;
  wire _26758_;
  wire _26759_;
  wire _26760_;
  wire _26761_;
  wire _26762_;
  wire _26763_;
  wire _26764_;
  wire _26765_;
  wire _26766_;
  wire _26767_;
  wire _26768_;
  wire _26769_;
  wire _26770_;
  wire _26771_;
  wire _26772_;
  wire _26773_;
  wire _26774_;
  wire _26775_;
  wire _26776_;
  wire _26777_;
  wire _26778_;
  wire _26779_;
  wire _26780_;
  wire _26781_;
  wire _26782_;
  wire _26783_;
  wire _26784_;
  wire _26785_;
  wire _26786_;
  wire _26787_;
  wire _26788_;
  wire _26789_;
  wire _26790_;
  wire _26791_;
  wire _26792_;
  wire _26793_;
  wire _26794_;
  wire _26795_;
  wire _26796_;
  wire _26797_;
  wire _26798_;
  wire _26799_;
  wire _26800_;
  wire _26801_;
  wire _26802_;
  wire _26803_;
  wire _26804_;
  wire _26805_;
  wire _26806_;
  wire _26807_;
  wire _26808_;
  wire _26809_;
  wire _26810_;
  wire _26811_;
  wire _26812_;
  wire _26813_;
  wire _26814_;
  wire _26815_;
  wire _26816_;
  wire _26817_;
  wire _26818_;
  wire _26819_;
  wire _26820_;
  wire _26821_;
  wire _26822_;
  wire _26823_;
  wire _26824_;
  wire _26825_;
  wire _26826_;
  wire _26827_;
  wire _26828_;
  wire _26829_;
  wire _26830_;
  wire _26831_;
  wire _26832_;
  wire _26833_;
  wire _26834_;
  wire _26835_;
  wire _26836_;
  wire _26837_;
  wire _26838_;
  wire _26839_;
  wire _26840_;
  wire _26841_;
  wire _26842_;
  wire _26843_;
  wire _26844_;
  wire _26845_;
  wire _26846_;
  wire _26847_;
  wire _26848_;
  wire _26849_;
  wire _26850_;
  wire _26851_;
  wire _26852_;
  wire _26853_;
  wire _26854_;
  wire _26855_;
  wire _26856_;
  wire _26857_;
  wire _26858_;
  wire _26859_;
  wire _26860_;
  wire _26861_;
  wire _26862_;
  wire _26863_;
  wire _26864_;
  wire _26865_;
  wire _26866_;
  wire _26867_;
  wire _26868_;
  wire _26869_;
  wire _26870_;
  wire _26871_;
  wire _26872_;
  wire _26873_;
  wire _26874_;
  wire _26875_;
  wire _26876_;
  wire _26877_;
  wire _26878_;
  wire _26879_;
  wire _26880_;
  wire _26881_;
  wire _26882_;
  wire _26883_;
  wire _26884_;
  wire _26885_;
  wire _26886_;
  wire _26887_;
  wire _26888_;
  wire _26889_;
  wire _26890_;
  wire _26891_;
  wire _26892_;
  wire _26893_;
  wire _26894_;
  wire _26895_;
  wire _26896_;
  wire _26897_;
  wire _26898_;
  wire _26899_;
  wire _26900_;
  wire _26901_;
  wire _26902_;
  wire _26903_;
  wire _26904_;
  wire _26905_;
  wire _26906_;
  wire _26907_;
  wire _26908_;
  wire _26909_;
  wire _26910_;
  wire _26911_;
  wire _26912_;
  wire _26913_;
  wire _26914_;
  wire _26915_;
  wire _26916_;
  wire _26917_;
  wire _26918_;
  wire _26919_;
  wire _26920_;
  wire _26921_;
  wire _26922_;
  wire _26923_;
  wire _26924_;
  wire _26925_;
  wire _26926_;
  wire _26927_;
  wire _26928_;
  wire _26929_;
  wire _26930_;
  wire _26931_;
  wire _26932_;
  wire _26933_;
  wire _26934_;
  wire _26935_;
  wire _26936_;
  wire _26937_;
  wire _26938_;
  wire _26939_;
  wire _26940_;
  wire _26941_;
  wire _26942_;
  wire _26943_;
  wire _26944_;
  wire _26945_;
  wire _26946_;
  wire _26947_;
  wire _26948_;
  wire _26949_;
  wire _26950_;
  wire _26951_;
  wire _26952_;
  wire _26953_;
  wire _26954_;
  wire _26955_;
  wire _26956_;
  wire _26957_;
  wire _26958_;
  wire _26959_;
  wire _26960_;
  wire _26961_;
  wire _26962_;
  wire _26963_;
  wire _26964_;
  wire _26965_;
  wire _26966_;
  wire _26967_;
  wire _26968_;
  wire _26969_;
  wire _26970_;
  wire _26971_;
  wire _26972_;
  wire _26973_;
  wire _26974_;
  wire _26975_;
  wire _26976_;
  wire _26977_;
  wire _26978_;
  wire _26979_;
  wire _26980_;
  wire _26981_;
  wire _26982_;
  wire _26983_;
  wire _26984_;
  wire _26985_;
  wire _26986_;
  wire _26987_;
  wire _26988_;
  wire _26989_;
  wire _26990_;
  wire _26991_;
  wire _26992_;
  wire _26993_;
  wire _26994_;
  wire _26995_;
  wire _26996_;
  wire _26997_;
  wire _26998_;
  wire _26999_;
  wire _27000_;
  wire _27001_;
  wire _27002_;
  wire _27003_;
  wire _27004_;
  wire _27005_;
  wire _27006_;
  wire _27007_;
  wire _27008_;
  wire _27009_;
  wire _27010_;
  wire _27011_;
  wire _27012_;
  wire _27013_;
  wire _27014_;
  wire _27015_;
  wire _27016_;
  wire _27017_;
  wire _27018_;
  wire _27019_;
  wire _27020_;
  wire _27021_;
  wire _27022_;
  wire _27023_;
  wire _27024_;
  wire _27025_;
  wire _27026_;
  wire _27027_;
  wire _27028_;
  wire _27029_;
  wire _27030_;
  wire _27031_;
  wire _27032_;
  wire _27033_;
  wire _27034_;
  wire _27035_;
  wire _27036_;
  wire _27037_;
  wire _27038_;
  wire _27039_;
  wire _27040_;
  wire _27041_;
  wire _27042_;
  wire _27043_;
  wire _27044_;
  wire _27045_;
  wire _27046_;
  wire _27047_;
  wire _27048_;
  wire _27049_;
  wire _27050_;
  wire _27051_;
  wire _27052_;
  wire _27053_;
  wire _27054_;
  wire _27055_;
  wire _27056_;
  wire _27057_;
  wire _27058_;
  wire _27059_;
  wire _27060_;
  wire _27061_;
  wire _27062_;
  wire _27063_;
  wire _27064_;
  wire _27065_;
  wire _27066_;
  wire _27067_;
  wire _27068_;
  wire _27069_;
  wire _27070_;
  wire _27071_;
  wire _27072_;
  wire _27073_;
  wire _27074_;
  wire _27075_;
  wire _27076_;
  wire _27077_;
  wire _27078_;
  wire _27079_;
  wire _27080_;
  wire _27081_;
  wire _27082_;
  wire _27083_;
  wire _27084_;
  wire _27085_;
  wire _27086_;
  wire _27087_;
  wire _27088_;
  wire _27089_;
  wire _27090_;
  wire _27091_;
  wire _27092_;
  wire _27093_;
  wire _27094_;
  wire _27095_;
  wire _27096_;
  wire _27097_;
  wire _27098_;
  wire _27099_;
  wire _27100_;
  wire _27101_;
  wire _27102_;
  wire _27103_;
  wire _27104_;
  wire _27105_;
  wire _27106_;
  wire _27107_;
  wire _27108_;
  wire _27109_;
  wire _27110_;
  wire _27111_;
  wire _27112_;
  wire _27113_;
  wire _27114_;
  wire _27115_;
  wire _27116_;
  wire _27117_;
  wire _27118_;
  wire _27119_;
  wire _27120_;
  wire _27121_;
  wire _27122_;
  wire _27123_;
  wire _27124_;
  wire _27125_;
  wire _27126_;
  wire _27127_;
  wire _27128_;
  wire _27129_;
  wire _27130_;
  wire _27131_;
  wire _27132_;
  wire _27133_;
  wire _27134_;
  wire _27135_;
  wire _27136_;
  wire _27137_;
  wire _27138_;
  wire _27139_;
  wire _27140_;
  wire _27141_;
  wire _27142_;
  wire _27143_;
  wire _27144_;
  wire _27145_;
  wire _27146_;
  wire _27147_;
  wire _27148_;
  wire _27149_;
  wire _27150_;
  wire _27151_;
  wire _27152_;
  wire _27153_;
  wire _27154_;
  wire _27155_;
  wire _27156_;
  wire _27157_;
  wire _27158_;
  wire _27159_;
  wire _27160_;
  wire _27161_;
  wire _27162_;
  wire _27163_;
  wire _27164_;
  wire _27165_;
  wire _27166_;
  wire _27167_;
  wire _27168_;
  wire _27169_;
  wire _27170_;
  wire _27171_;
  wire _27172_;
  wire _27173_;
  wire _27174_;
  wire _27175_;
  wire _27176_;
  wire _27177_;
  wire _27178_;
  wire _27179_;
  wire _27180_;
  wire _27181_;
  wire _27182_;
  wire _27183_;
  wire _27184_;
  wire _27185_;
  wire _27186_;
  wire _27187_;
  wire _27188_;
  wire _27189_;
  wire _27190_;
  wire _27191_;
  wire _27192_;
  wire _27193_;
  wire _27194_;
  wire _27195_;
  wire _27196_;
  wire _27197_;
  wire _27198_;
  wire _27199_;
  wire _27200_;
  wire _27201_;
  wire _27202_;
  wire _27203_;
  wire _27204_;
  wire _27205_;
  wire _27206_;
  wire _27207_;
  wire _27208_;
  wire _27209_;
  wire _27210_;
  wire _27211_;
  wire _27212_;
  wire _27213_;
  wire _27214_;
  wire _27215_;
  wire _27216_;
  wire _27217_;
  wire _27218_;
  wire _27219_;
  wire _27220_;
  wire _27221_;
  wire _27222_;
  wire _27223_;
  wire _27224_;
  wire _27225_;
  wire _27226_;
  wire _27227_;
  wire _27228_;
  wire _27229_;
  wire _27230_;
  wire _27231_;
  wire _27232_;
  wire _27233_;
  wire _27234_;
  wire _27235_;
  wire _27236_;
  wire _27237_;
  wire _27238_;
  wire _27239_;
  wire _27240_;
  wire _27241_;
  wire _27242_;
  wire _27243_;
  wire _27244_;
  wire _27245_;
  wire _27246_;
  wire _27247_;
  wire _27248_;
  wire _27249_;
  wire _27250_;
  wire _27251_;
  wire _27252_;
  wire _27253_;
  wire _27254_;
  wire _27255_;
  wire _27256_;
  wire _27257_;
  wire _27258_;
  wire _27259_;
  wire _27260_;
  wire _27261_;
  wire _27262_;
  wire _27263_;
  wire _27264_;
  wire _27265_;
  wire _27266_;
  wire _27267_;
  wire _27268_;
  wire _27269_;
  wire _27270_;
  wire _27271_;
  wire _27272_;
  wire _27273_;
  wire _27274_;
  wire _27275_;
  wire _27276_;
  wire _27277_;
  wire _27278_;
  wire _27279_;
  wire _27280_;
  wire _27281_;
  wire _27282_;
  wire _27283_;
  wire _27284_;
  wire _27285_;
  wire _27286_;
  wire _27287_;
  wire _27288_;
  wire _27289_;
  wire _27290_;
  wire _27291_;
  wire _27292_;
  wire _27293_;
  wire _27294_;
  wire _27295_;
  wire _27296_;
  wire _27297_;
  wire _27298_;
  wire _27299_;
  wire _27300_;
  wire _27301_;
  wire _27302_;
  wire _27303_;
  wire _27304_;
  wire _27305_;
  wire _27306_;
  wire _27307_;
  wire _27308_;
  wire _27309_;
  wire _27310_;
  wire _27311_;
  wire _27312_;
  wire _27313_;
  wire _27314_;
  wire _27315_;
  wire _27316_;
  wire _27317_;
  wire _27318_;
  wire _27319_;
  wire _27320_;
  wire _27321_;
  wire _27322_;
  wire _27323_;
  wire _27324_;
  wire _27325_;
  wire _27326_;
  wire _27327_;
  wire _27328_;
  wire _27329_;
  wire _27330_;
  wire _27331_;
  wire _27332_;
  wire _27333_;
  wire _27334_;
  wire _27335_;
  wire _27336_;
  wire _27337_;
  wire _27338_;
  wire _27339_;
  wire _27340_;
  wire _27341_;
  wire _27342_;
  wire _27343_;
  wire _27344_;
  wire _27345_;
  wire _27346_;
  wire _27347_;
  wire _27348_;
  wire _27349_;
  wire _27350_;
  wire _27351_;
  wire _27352_;
  wire _27353_;
  wire _27354_;
  wire _27355_;
  wire _27356_;
  wire _27357_;
  wire _27358_;
  wire _27359_;
  wire _27360_;
  wire _27361_;
  wire _27362_;
  wire _27363_;
  wire _27364_;
  wire _27365_;
  wire _27366_;
  wire _27367_;
  wire _27368_;
  wire _27369_;
  wire _27370_;
  wire _27371_;
  wire _27372_;
  wire _27373_;
  wire _27374_;
  wire _27375_;
  wire _27376_;
  wire _27377_;
  wire _27378_;
  wire _27379_;
  wire _27380_;
  wire _27381_;
  wire _27382_;
  wire _27383_;
  wire _27384_;
  wire _27385_;
  wire _27386_;
  wire _27387_;
  wire _27388_;
  wire _27389_;
  wire _27390_;
  wire _27391_;
  wire _27392_;
  wire _27393_;
  wire _27394_;
  wire _27395_;
  wire _27396_;
  wire _27397_;
  wire _27398_;
  wire _27399_;
  wire _27400_;
  wire _27401_;
  wire _27402_;
  wire _27403_;
  wire _27404_;
  wire _27405_;
  wire _27406_;
  wire _27407_;
  wire _27408_;
  wire _27409_;
  wire _27410_;
  wire _27411_;
  wire _27412_;
  wire _27413_;
  wire _27414_;
  wire _27415_;
  wire _27416_;
  wire _27417_;
  wire _27418_;
  wire _27419_;
  wire _27420_;
  wire _27421_;
  wire _27422_;
  wire _27423_;
  wire _27424_;
  wire _27425_;
  wire _27426_;
  wire _27427_;
  wire _27428_;
  wire _27429_;
  wire _27430_;
  wire _27431_;
  wire _27432_;
  wire _27433_;
  wire _27434_;
  wire _27435_;
  wire _27436_;
  wire _27437_;
  wire _27438_;
  wire _27439_;
  wire _27440_;
  wire _27441_;
  wire _27442_;
  wire _27443_;
  wire _27444_;
  wire _27445_;
  wire _27446_;
  wire _27447_;
  wire _27448_;
  wire _27449_;
  wire _27450_;
  wire _27451_;
  wire _27452_;
  wire _27453_;
  wire _27454_;
  wire _27455_;
  wire _27456_;
  wire _27457_;
  wire _27458_;
  wire _27459_;
  wire _27460_;
  wire _27461_;
  wire _27462_;
  wire _27463_;
  wire _27464_;
  wire _27465_;
  wire _27466_;
  wire _27467_;
  wire _27468_;
  wire _27469_;
  wire _27470_;
  wire _27471_;
  wire _27472_;
  wire _27473_;
  wire _27474_;
  wire _27475_;
  wire _27476_;
  wire _27477_;
  wire _27478_;
  wire _27479_;
  wire _27480_;
  wire _27481_;
  wire _27482_;
  wire _27483_;
  wire _27484_;
  wire _27485_;
  wire _27486_;
  wire _27487_;
  wire _27488_;
  wire _27489_;
  wire _27490_;
  wire _27491_;
  wire _27492_;
  wire _27493_;
  wire _27494_;
  wire _27495_;
  wire _27496_;
  wire _27497_;
  wire _27498_;
  wire _27499_;
  wire _27500_;
  wire _27501_;
  wire _27502_;
  wire _27503_;
  wire _27504_;
  wire _27505_;
  wire _27506_;
  wire _27507_;
  wire _27508_;
  wire _27509_;
  wire _27510_;
  wire _27511_;
  wire _27512_;
  wire _27513_;
  wire _27514_;
  wire _27515_;
  wire _27516_;
  wire _27517_;
  wire _27518_;
  wire _27519_;
  wire _27520_;
  wire _27521_;
  wire _27522_;
  wire _27523_;
  wire _27524_;
  wire _27525_;
  wire _27526_;
  wire _27527_;
  wire _27528_;
  wire _27529_;
  wire _27530_;
  wire _27531_;
  wire _27532_;
  wire _27533_;
  wire _27534_;
  wire _27535_;
  wire _27536_;
  wire _27537_;
  wire _27538_;
  wire _27539_;
  wire _27540_;
  wire _27541_;
  wire _27542_;
  wire _27543_;
  wire _27544_;
  wire _27545_;
  wire _27546_;
  wire _27547_;
  wire _27548_;
  wire _27549_;
  wire _27550_;
  wire _27551_;
  wire _27552_;
  wire _27553_;
  wire _27554_;
  wire _27555_;
  wire _27556_;
  wire _27557_;
  wire _27558_;
  wire _27559_;
  wire _27560_;
  wire _27561_;
  wire _27562_;
  wire _27563_;
  wire _27564_;
  wire _27565_;
  wire _27566_;
  wire _27567_;
  wire _27568_;
  wire _27569_;
  wire _27570_;
  wire _27571_;
  wire _27572_;
  wire _27573_;
  wire _27574_;
  wire _27575_;
  wire _27576_;
  wire _27577_;
  wire _27578_;
  wire _27579_;
  wire _27580_;
  wire _27581_;
  wire _27582_;
  wire _27583_;
  wire _27584_;
  wire _27585_;
  wire _27586_;
  wire _27587_;
  wire _27588_;
  wire _27589_;
  wire _27590_;
  wire _27591_;
  wire _27592_;
  wire _27593_;
  wire _27594_;
  wire _27595_;
  wire _27596_;
  wire _27597_;
  wire _27598_;
  wire _27599_;
  wire _27600_;
  wire _27601_;
  wire _27602_;
  wire _27603_;
  wire _27604_;
  wire _27605_;
  wire _27606_;
  wire _27607_;
  wire _27608_;
  wire _27609_;
  wire _27610_;
  wire _27611_;
  wire _27612_;
  wire _27613_;
  wire _27614_;
  wire _27615_;
  wire _27616_;
  wire _27617_;
  wire _27618_;
  wire _27619_;
  wire _27620_;
  wire _27621_;
  wire _27622_;
  wire _27623_;
  wire _27624_;
  wire _27625_;
  wire _27626_;
  wire _27627_;
  wire _27628_;
  wire _27629_;
  wire _27630_;
  wire _27631_;
  wire _27632_;
  wire _27633_;
  wire _27634_;
  wire _27635_;
  wire _27636_;
  wire _27637_;
  wire _27638_;
  wire _27639_;
  wire _27640_;
  wire _27641_;
  wire _27642_;
  wire _27643_;
  wire _27644_;
  wire _27645_;
  wire _27646_;
  wire _27647_;
  wire _27648_;
  wire _27649_;
  wire _27650_;
  wire _27651_;
  wire _27652_;
  wire _27653_;
  wire _27654_;
  wire _27655_;
  wire _27656_;
  wire _27657_;
  wire _27658_;
  wire _27659_;
  wire _27660_;
  wire _27661_;
  wire _27662_;
  wire _27663_;
  wire _27664_;
  wire _27665_;
  wire _27666_;
  wire _27667_;
  wire _27668_;
  wire _27669_;
  wire _27670_;
  wire _27671_;
  wire _27672_;
  wire _27673_;
  wire _27674_;
  wire _27675_;
  wire _27676_;
  wire _27677_;
  wire _27678_;
  wire _27679_;
  wire _27680_;
  wire _27681_;
  wire _27682_;
  wire _27683_;
  wire _27684_;
  wire _27685_;
  wire _27686_;
  wire _27687_;
  wire _27688_;
  wire _27689_;
  wire _27690_;
  wire _27691_;
  wire _27692_;
  wire _27693_;
  wire _27694_;
  wire _27695_;
  wire _27696_;
  wire _27697_;
  wire _27698_;
  wire _27699_;
  wire _27700_;
  wire _27701_;
  wire _27702_;
  wire _27703_;
  wire _27704_;
  wire _27705_;
  wire _27706_;
  wire _27707_;
  wire _27708_;
  wire _27709_;
  wire _27710_;
  wire _27711_;
  wire _27712_;
  wire _27713_;
  wire _27714_;
  wire _27715_;
  wire _27716_;
  wire _27717_;
  wire _27718_;
  wire _27719_;
  wire _27720_;
  wire _27721_;
  wire _27722_;
  wire _27723_;
  wire _27724_;
  wire _27725_;
  wire _27726_;
  wire _27727_;
  wire _27728_;
  wire _27729_;
  wire _27730_;
  wire _27731_;
  wire _27732_;
  wire _27733_;
  wire _27734_;
  wire _27735_;
  wire _27736_;
  wire _27737_;
  wire _27738_;
  wire _27739_;
  wire _27740_;
  wire _27741_;
  wire _27742_;
  wire _27743_;
  wire _27744_;
  wire _27745_;
  wire _27746_;
  wire _27747_;
  wire _27748_;
  wire _27749_;
  wire _27750_;
  wire _27751_;
  wire _27752_;
  wire _27753_;
  wire _27754_;
  wire _27755_;
  wire _27756_;
  wire _27757_;
  wire _27758_;
  wire _27759_;
  wire _27760_;
  wire _27761_;
  wire _27762_;
  wire _27763_;
  wire _27764_;
  wire _27765_;
  wire _27766_;
  wire _27767_;
  wire _27768_;
  wire _27769_;
  wire _27770_;
  wire _27771_;
  wire _27772_;
  wire _27773_;
  wire _27774_;
  wire _27775_;
  wire _27776_;
  wire _27777_;
  wire _27778_;
  wire _27779_;
  wire _27780_;
  wire _27781_;
  wire _27782_;
  wire _27783_;
  wire _27784_;
  wire _27785_;
  wire _27786_;
  wire _27787_;
  wire _27788_;
  wire _27789_;
  wire _27790_;
  wire _27791_;
  wire _27792_;
  wire _27793_;
  wire _27794_;
  wire _27795_;
  wire _27796_;
  wire _27797_;
  wire _27798_;
  wire _27799_;
  wire _27800_;
  wire _27801_;
  wire _27802_;
  wire _27803_;
  wire _27804_;
  wire _27805_;
  wire _27806_;
  wire _27807_;
  wire _27808_;
  wire _27809_;
  wire _27810_;
  wire _27811_;
  wire _27812_;
  wire _27813_;
  wire _27814_;
  wire _27815_;
  wire _27816_;
  wire _27817_;
  wire _27818_;
  wire _27819_;
  wire _27820_;
  wire _27821_;
  wire _27822_;
  wire _27823_;
  wire _27824_;
  wire _27825_;
  wire _27826_;
  wire _27827_;
  wire _27828_;
  wire _27829_;
  wire _27830_;
  wire _27831_;
  wire _27832_;
  wire _27833_;
  wire _27834_;
  wire _27835_;
  wire _27836_;
  wire _27837_;
  wire _27838_;
  wire _27839_;
  wire _27840_;
  wire _27841_;
  wire _27842_;
  wire _27843_;
  wire _27844_;
  wire _27845_;
  wire _27846_;
  wire _27847_;
  wire _27848_;
  wire _27849_;
  wire _27850_;
  wire _27851_;
  wire _27852_;
  wire _27853_;
  wire _27854_;
  wire _27855_;
  wire _27856_;
  wire _27857_;
  wire _27858_;
  wire _27859_;
  wire _27860_;
  wire _27861_;
  wire _27862_;
  wire _27863_;
  wire _27864_;
  wire _27865_;
  wire _27866_;
  wire _27867_;
  wire _27868_;
  wire _27869_;
  wire _27870_;
  wire _27871_;
  wire _27872_;
  wire _27873_;
  wire _27874_;
  wire _27875_;
  wire _27876_;
  wire _27877_;
  wire _27878_;
  wire _27879_;
  wire _27880_;
  wire _27881_;
  wire _27882_;
  wire _27883_;
  wire _27884_;
  wire _27885_;
  wire _27886_;
  wire _27887_;
  wire _27888_;
  wire _27889_;
  wire _27890_;
  wire _27891_;
  wire _27892_;
  wire _27893_;
  wire _27894_;
  wire _27895_;
  wire _27896_;
  wire _27897_;
  wire _27898_;
  wire _27899_;
  wire _27900_;
  wire _27901_;
  wire _27902_;
  wire _27903_;
  wire _27904_;
  wire _27905_;
  wire _27906_;
  wire _27907_;
  wire _27908_;
  wire _27909_;
  wire _27910_;
  wire _27911_;
  wire _27912_;
  wire _27913_;
  wire _27914_;
  wire _27915_;
  wire _27916_;
  wire _27917_;
  wire _27918_;
  wire _27919_;
  wire _27920_;
  wire _27921_;
  wire _27922_;
  wire _27923_;
  wire _27924_;
  wire _27925_;
  wire _27926_;
  wire _27927_;
  wire _27928_;
  wire _27929_;
  wire _27930_;
  wire _27931_;
  wire _27932_;
  wire _27933_;
  wire _27934_;
  wire _27935_;
  wire _27936_;
  wire _27937_;
  wire _27938_;
  wire _27939_;
  wire _27940_;
  wire _27941_;
  wire _27942_;
  wire _27943_;
  wire _27944_;
  wire _27945_;
  wire _27946_;
  wire _27947_;
  wire _27948_;
  wire _27949_;
  wire _27950_;
  wire _27951_;
  wire _27952_;
  wire _27953_;
  wire _27954_;
  wire _27955_;
  wire _27956_;
  wire _27957_;
  wire _27958_;
  wire _27959_;
  wire _27960_;
  wire _27961_;
  wire _27962_;
  wire _27963_;
  wire _27964_;
  wire _27965_;
  wire _27966_;
  wire _27967_;
  wire _27968_;
  wire _27969_;
  wire _27970_;
  wire _27971_;
  wire _27972_;
  wire _27973_;
  wire _27974_;
  wire _27975_;
  wire _27976_;
  wire _27977_;
  wire _27978_;
  wire _27979_;
  wire _27980_;
  wire _27981_;
  wire _27982_;
  wire _27983_;
  wire _27984_;
  wire _27985_;
  wire _27986_;
  wire _27987_;
  wire _27988_;
  wire _27989_;
  wire _27990_;
  wire _27991_;
  wire _27992_;
  wire _27993_;
  wire _27994_;
  wire _27995_;
  wire _27996_;
  wire _27997_;
  wire _27998_;
  wire _27999_;
  wire _28000_;
  wire _28001_;
  wire _28002_;
  wire _28003_;
  wire _28004_;
  wire _28005_;
  wire _28006_;
  wire _28007_;
  wire _28008_;
  wire _28009_;
  wire _28010_;
  wire _28011_;
  wire _28012_;
  wire _28013_;
  wire _28014_;
  wire _28015_;
  wire _28016_;
  wire _28017_;
  wire _28018_;
  wire _28019_;
  wire _28020_;
  wire _28021_;
  wire _28022_;
  wire _28023_;
  wire _28024_;
  wire _28025_;
  wire _28026_;
  wire _28027_;
  wire _28028_;
  wire _28029_;
  wire _28030_;
  wire _28031_;
  wire _28032_;
  wire _28033_;
  wire _28034_;
  wire _28035_;
  wire _28036_;
  wire _28037_;
  wire _28038_;
  wire _28039_;
  wire _28040_;
  wire _28041_;
  wire _28042_;
  wire _28043_;
  wire _28044_;
  wire _28045_;
  wire _28046_;
  wire _28047_;
  wire _28048_;
  wire _28049_;
  wire _28050_;
  wire _28051_;
  wire _28052_;
  wire _28053_;
  wire _28054_;
  wire _28055_;
  wire _28056_;
  wire _28057_;
  wire _28058_;
  wire _28059_;
  wire _28060_;
  wire _28061_;
  wire _28062_;
  wire _28063_;
  wire _28064_;
  wire _28065_;
  wire _28066_;
  wire _28067_;
  wire _28068_;
  wire _28069_;
  wire _28070_;
  wire _28071_;
  wire _28072_;
  wire _28073_;
  wire _28074_;
  wire _28075_;
  wire _28076_;
  wire _28077_;
  wire _28078_;
  wire _28079_;
  wire _28080_;
  wire _28081_;
  wire _28082_;
  wire _28083_;
  wire _28084_;
  wire _28085_;
  wire _28086_;
  wire _28087_;
  wire _28088_;
  wire _28089_;
  wire _28090_;
  wire _28091_;
  wire _28092_;
  wire _28093_;
  wire _28094_;
  wire _28095_;
  wire _28096_;
  wire _28097_;
  wire _28098_;
  wire _28099_;
  wire _28100_;
  wire _28101_;
  wire _28102_;
  wire _28103_;
  wire _28104_;
  wire _28105_;
  wire _28106_;
  wire _28107_;
  wire _28108_;
  wire _28109_;
  wire _28110_;
  wire _28111_;
  wire _28112_;
  wire _28113_;
  wire _28114_;
  wire _28115_;
  wire _28116_;
  wire _28117_;
  wire _28118_;
  wire _28119_;
  wire _28120_;
  wire _28121_;
  wire _28122_;
  wire _28123_;
  wire _28124_;
  wire _28125_;
  wire _28126_;
  wire _28127_;
  wire _28128_;
  wire _28129_;
  wire _28130_;
  wire _28131_;
  wire _28132_;
  wire _28133_;
  wire _28134_;
  wire _28135_;
  wire _28136_;
  wire _28137_;
  wire _28138_;
  wire _28139_;
  wire _28140_;
  wire _28141_;
  wire _28142_;
  wire _28143_;
  wire _28144_;
  wire _28145_;
  wire _28146_;
  wire _28147_;
  wire _28148_;
  wire _28149_;
  wire _28150_;
  wire _28151_;
  wire _28152_;
  wire _28153_;
  wire _28154_;
  wire _28155_;
  wire _28156_;
  wire _28157_;
  wire _28158_;
  wire _28159_;
  wire _28160_;
  wire _28161_;
  wire _28162_;
  wire _28163_;
  wire _28164_;
  wire _28165_;
  wire _28166_;
  wire _28167_;
  wire _28168_;
  wire _28169_;
  wire _28170_;
  wire _28171_;
  wire _28172_;
  wire _28173_;
  wire _28174_;
  wire _28175_;
  wire _28176_;
  wire _28177_;
  wire _28178_;
  wire _28179_;
  wire _28180_;
  wire _28181_;
  wire _28182_;
  wire _28183_;
  wire _28184_;
  wire _28185_;
  wire _28186_;
  wire _28187_;
  wire _28188_;
  wire _28189_;
  wire _28190_;
  wire _28191_;
  wire _28192_;
  wire _28193_;
  wire _28194_;
  wire _28195_;
  wire _28196_;
  wire _28197_;
  wire _28198_;
  wire _28199_;
  wire _28200_;
  wire _28201_;
  wire _28202_;
  wire _28203_;
  wire _28204_;
  wire _28205_;
  wire _28206_;
  wire _28207_;
  wire _28208_;
  wire _28209_;
  wire _28210_;
  wire _28211_;
  wire _28212_;
  wire _28213_;
  wire _28214_;
  wire _28215_;
  wire _28216_;
  wire _28217_;
  wire _28218_;
  wire _28219_;
  wire _28220_;
  wire _28221_;
  wire _28222_;
  wire _28223_;
  wire _28224_;
  wire _28225_;
  wire _28226_;
  wire _28227_;
  wire _28228_;
  wire _28229_;
  wire _28230_;
  wire _28231_;
  wire _28232_;
  wire _28233_;
  wire _28234_;
  wire _28235_;
  wire _28236_;
  wire _28237_;
  wire _28238_;
  wire _28239_;
  wire _28240_;
  wire _28241_;
  wire _28242_;
  wire _28243_;
  wire _28244_;
  wire _28245_;
  wire _28246_;
  wire _28247_;
  wire _28248_;
  wire _28249_;
  wire _28250_;
  wire _28251_;
  wire _28252_;
  wire _28253_;
  wire _28254_;
  wire _28255_;
  wire _28256_;
  wire _28257_;
  wire _28258_;
  wire _28259_;
  wire _28260_;
  wire _28261_;
  wire _28262_;
  wire _28263_;
  wire _28264_;
  wire _28265_;
  wire _28266_;
  wire _28267_;
  wire _28268_;
  wire _28269_;
  wire _28270_;
  wire _28271_;
  wire _28272_;
  wire _28273_;
  wire _28274_;
  wire _28275_;
  wire _28276_;
  wire _28277_;
  wire _28278_;
  wire _28279_;
  wire _28280_;
  wire _28281_;
  wire _28282_;
  wire _28283_;
  wire _28284_;
  wire _28285_;
  wire _28286_;
  wire _28287_;
  wire _28288_;
  wire _28289_;
  wire _28290_;
  wire _28291_;
  wire _28292_;
  wire _28293_;
  wire _28294_;
  wire _28295_;
  wire _28296_;
  wire _28297_;
  wire _28298_;
  wire _28299_;
  wire _28300_;
  wire _28301_;
  wire _28302_;
  wire _28303_;
  wire _28304_;
  wire _28305_;
  wire _28306_;
  wire _28307_;
  wire _28308_;
  wire _28309_;
  wire _28310_;
  wire _28311_;
  wire _28312_;
  wire _28313_;
  wire _28314_;
  wire _28315_;
  wire _28316_;
  wire _28317_;
  wire _28318_;
  wire _28319_;
  wire _28320_;
  wire _28321_;
  wire _28322_;
  wire _28323_;
  wire _28324_;
  wire _28325_;
  wire _28326_;
  wire _28327_;
  wire _28328_;
  wire _28329_;
  wire _28330_;
  wire _28331_;
  wire _28332_;
  wire _28333_;
  wire _28334_;
  wire _28335_;
  wire _28336_;
  wire _28337_;
  wire _28338_;
  wire _28339_;
  wire _28340_;
  wire _28341_;
  wire _28342_;
  wire _28343_;
  wire _28344_;
  wire _28345_;
  wire _28346_;
  wire _28347_;
  wire _28348_;
  wire _28349_;
  wire _28350_;
  wire _28351_;
  wire _28352_;
  wire _28353_;
  wire _28354_;
  wire _28355_;
  wire _28356_;
  wire _28357_;
  wire _28358_;
  wire _28359_;
  wire _28360_;
  wire _28361_;
  wire _28362_;
  wire _28363_;
  wire _28364_;
  wire _28365_;
  wire _28366_;
  wire _28367_;
  wire _28368_;
  wire _28369_;
  wire _28370_;
  wire _28371_;
  wire _28372_;
  wire _28373_;
  wire _28374_;
  wire _28375_;
  wire _28376_;
  wire _28377_;
  wire _28378_;
  wire _28379_;
  wire _28380_;
  wire _28381_;
  wire _28382_;
  wire _28383_;
  wire _28384_;
  wire _28385_;
  wire _28386_;
  wire _28387_;
  wire _28388_;
  wire _28389_;
  wire _28390_;
  wire _28391_;
  wire _28392_;
  wire _28393_;
  wire _28394_;
  wire _28395_;
  wire _28396_;
  wire _28397_;
  wire _28398_;
  wire _28399_;
  wire _28400_;
  wire _28401_;
  wire _28402_;
  wire _28403_;
  wire _28404_;
  wire _28405_;
  wire _28406_;
  wire _28407_;
  wire _28408_;
  wire _28409_;
  wire _28410_;
  wire _28411_;
  wire _28412_;
  wire _28413_;
  wire _28414_;
  wire _28415_;
  wire _28416_;
  wire _28417_;
  wire _28418_;
  wire _28419_;
  wire _28420_;
  wire _28421_;
  wire _28422_;
  wire _28423_;
  wire _28424_;
  wire _28425_;
  wire _28426_;
  wire _28427_;
  wire _28428_;
  wire _28429_;
  wire _28430_;
  wire _28431_;
  wire _28432_;
  wire _28433_;
  wire _28434_;
  wire _28435_;
  wire _28436_;
  wire _28437_;
  wire _28438_;
  wire _28439_;
  wire _28440_;
  wire _28441_;
  wire _28442_;
  wire _28443_;
  wire _28444_;
  wire _28445_;
  wire _28446_;
  wire _28447_;
  wire _28448_;
  wire _28449_;
  wire _28450_;
  wire _28451_;
  wire _28452_;
  wire _28453_;
  wire _28454_;
  wire _28455_;
  wire _28456_;
  wire _28457_;
  wire _28458_;
  wire _28459_;
  wire _28460_;
  wire _28461_;
  wire _28462_;
  wire _28463_;
  wire _28464_;
  wire _28465_;
  wire _28466_;
  wire _28467_;
  wire _28468_;
  wire _28469_;
  wire _28470_;
  wire _28471_;
  wire _28472_;
  wire _28473_;
  wire _28474_;
  wire _28475_;
  wire _28476_;
  wire _28477_;
  wire _28478_;
  wire _28479_;
  wire _28480_;
  wire _28481_;
  wire _28482_;
  wire _28483_;
  wire _28484_;
  wire _28485_;
  wire _28486_;
  wire _28487_;
  wire _28488_;
  wire _28489_;
  wire _28490_;
  wire _28491_;
  wire _28492_;
  wire _28493_;
  wire _28494_;
  wire _28495_;
  wire _28496_;
  wire _28497_;
  wire _28498_;
  wire _28499_;
  wire _28500_;
  wire _28501_;
  wire _28502_;
  wire _28503_;
  wire _28504_;
  wire _28505_;
  wire _28506_;
  wire _28507_;
  wire _28508_;
  wire _28509_;
  wire _28510_;
  wire _28511_;
  wire _28512_;
  wire _28513_;
  wire _28514_;
  wire _28515_;
  wire _28516_;
  wire _28517_;
  wire _28518_;
  wire _28519_;
  wire _28520_;
  wire _28521_;
  wire _28522_;
  wire _28523_;
  wire _28524_;
  wire _28525_;
  wire _28526_;
  wire _28527_;
  wire _28528_;
  wire _28529_;
  wire _28530_;
  wire _28531_;
  wire _28532_;
  wire _28533_;
  wire _28534_;
  wire _28535_;
  wire _28536_;
  wire _28537_;
  wire _28538_;
  wire _28539_;
  wire _28540_;
  wire _28541_;
  wire _28542_;
  wire _28543_;
  wire _28544_;
  wire _28545_;
  wire _28546_;
  wire _28547_;
  wire _28548_;
  wire _28549_;
  wire _28550_;
  wire _28551_;
  wire _28552_;
  wire _28553_;
  wire _28554_;
  wire _28555_;
  wire _28556_;
  wire _28557_;
  wire _28558_;
  wire _28559_;
  wire _28560_;
  wire _28561_;
  wire _28562_;
  wire _28563_;
  wire _28564_;
  wire _28565_;
  wire _28566_;
  wire _28567_;
  wire _28568_;
  wire _28569_;
  wire _28570_;
  wire _28571_;
  wire _28572_;
  wire _28573_;
  wire _28574_;
  wire _28575_;
  wire _28576_;
  wire _28577_;
  wire _28578_;
  wire _28579_;
  wire _28580_;
  wire _28581_;
  wire _28582_;
  wire _28583_;
  wire _28584_;
  wire _28585_;
  wire _28586_;
  wire _28587_;
  wire _28588_;
  wire _28589_;
  wire _28590_;
  wire _28591_;
  wire _28592_;
  wire _28593_;
  wire _28594_;
  wire _28595_;
  wire _28596_;
  wire _28597_;
  wire _28598_;
  wire _28599_;
  wire _28600_;
  wire _28601_;
  wire _28602_;
  wire _28603_;
  wire _28604_;
  wire _28605_;
  wire _28606_;
  wire _28607_;
  wire _28608_;
  wire _28609_;
  wire _28610_;
  wire _28611_;
  wire _28612_;
  wire _28613_;
  wire _28614_;
  wire _28615_;
  wire _28616_;
  wire _28617_;
  wire _28618_;
  wire _28619_;
  wire _28620_;
  wire _28621_;
  wire _28622_;
  wire _28623_;
  wire _28624_;
  wire _28625_;
  wire _28626_;
  wire _28627_;
  wire _28628_;
  wire _28629_;
  wire _28630_;
  wire _28631_;
  wire _28632_;
  wire _28633_;
  wire _28634_;
  wire _28635_;
  wire _28636_;
  wire _28637_;
  wire _28638_;
  wire _28639_;
  wire _28640_;
  wire _28641_;
  wire _28642_;
  wire _28643_;
  wire _28644_;
  wire _28645_;
  wire _28646_;
  wire _28647_;
  wire _28648_;
  wire _28649_;
  wire _28650_;
  wire _28651_;
  wire _28652_;
  wire _28653_;
  wire _28654_;
  wire _28655_;
  wire _28656_;
  wire _28657_;
  wire _28658_;
  wire _28659_;
  wire _28660_;
  wire _28661_;
  wire _28662_;
  wire _28663_;
  wire _28664_;
  wire _28665_;
  wire _28666_;
  wire _28667_;
  wire _28668_;
  wire _28669_;
  wire _28670_;
  wire _28671_;
  wire _28672_;
  wire _28673_;
  wire _28674_;
  wire _28675_;
  wire _28676_;
  wire _28677_;
  wire _28678_;
  wire _28679_;
  wire _28680_;
  wire _28681_;
  wire _28682_;
  wire _28683_;
  wire _28684_;
  wire _28685_;
  wire _28686_;
  wire _28687_;
  wire _28688_;
  wire _28689_;
  wire _28690_;
  wire _28691_;
  wire _28692_;
  wire _28693_;
  wire _28694_;
  wire _28695_;
  wire _28696_;
  wire _28697_;
  wire _28698_;
  wire _28699_;
  wire _28700_;
  wire _28701_;
  wire _28702_;
  wire _28703_;
  wire _28704_;
  wire _28705_;
  wire _28706_;
  wire _28707_;
  wire _28708_;
  wire _28709_;
  wire _28710_;
  wire _28711_;
  wire _28712_;
  wire _28713_;
  wire _28714_;
  wire _28715_;
  wire _28716_;
  wire _28717_;
  wire _28718_;
  wire _28719_;
  wire _28720_;
  wire _28721_;
  wire _28722_;
  wire _28723_;
  wire _28724_;
  wire _28725_;
  wire _28726_;
  wire _28727_;
  wire _28728_;
  wire _28729_;
  wire _28730_;
  wire _28731_;
  wire _28732_;
  wire _28733_;
  wire _28734_;
  wire _28735_;
  wire _28736_;
  wire _28737_;
  wire _28738_;
  wire _28739_;
  wire _28740_;
  wire _28741_;
  wire _28742_;
  wire _28743_;
  wire _28744_;
  wire _28745_;
  wire _28746_;
  wire _28747_;
  wire _28748_;
  wire _28749_;
  wire _28750_;
  wire _28751_;
  wire _28752_;
  wire _28753_;
  wire _28754_;
  wire _28755_;
  wire _28756_;
  wire _28757_;
  wire _28758_;
  wire _28759_;
  wire _28760_;
  wire _28761_;
  wire _28762_;
  wire _28763_;
  wire _28764_;
  wire _28765_;
  wire _28766_;
  wire _28767_;
  wire _28768_;
  wire _28769_;
  wire _28770_;
  wire _28771_;
  wire _28772_;
  wire _28773_;
  wire _28774_;
  wire _28775_;
  wire _28776_;
  wire _28777_;
  wire _28778_;
  wire _28779_;
  wire _28780_;
  wire _28781_;
  wire _28782_;
  wire _28783_;
  wire _28784_;
  wire _28785_;
  wire _28786_;
  wire _28787_;
  wire _28788_;
  wire _28789_;
  wire _28790_;
  wire _28791_;
  wire _28792_;
  wire _28793_;
  wire _28794_;
  wire _28795_;
  wire _28796_;
  wire _28797_;
  wire _28798_;
  wire _28799_;
  wire _28800_;
  wire _28801_;
  wire _28802_;
  wire _28803_;
  wire _28804_;
  wire _28805_;
  wire _28806_;
  wire _28807_;
  wire _28808_;
  wire _28809_;
  wire _28810_;
  wire _28811_;
  wire _28812_;
  wire _28813_;
  wire _28814_;
  wire _28815_;
  wire _28816_;
  wire _28817_;
  wire _28818_;
  wire _28819_;
  wire _28820_;
  wire _28821_;
  wire _28822_;
  wire _28823_;
  wire _28824_;
  wire _28825_;
  wire _28826_;
  wire _28827_;
  wire _28828_;
  wire _28829_;
  wire _28830_;
  wire _28831_;
  wire _28832_;
  wire _28833_;
  wire _28834_;
  wire _28835_;
  wire _28836_;
  wire _28837_;
  wire _28838_;
  wire _28839_;
  wire _28840_;
  wire _28841_;
  wire _28842_;
  wire _28843_;
  wire _28844_;
  wire _28845_;
  wire _28846_;
  wire _28847_;
  wire _28848_;
  wire _28849_;
  wire _28850_;
  wire _28851_;
  wire _28852_;
  wire _28853_;
  wire _28854_;
  wire _28855_;
  wire _28856_;
  wire _28857_;
  wire _28858_;
  wire _28859_;
  wire _28860_;
  wire _28861_;
  wire _28862_;
  wire _28863_;
  wire _28864_;
  wire _28865_;
  wire _28866_;
  wire _28867_;
  wire _28868_;
  wire _28869_;
  wire _28870_;
  wire _28871_;
  wire _28872_;
  wire _28873_;
  wire _28874_;
  wire _28875_;
  wire _28876_;
  wire _28877_;
  wire _28878_;
  wire _28879_;
  wire _28880_;
  wire _28881_;
  wire _28882_;
  wire _28883_;
  wire _28884_;
  wire _28885_;
  wire _28886_;
  wire _28887_;
  wire _28888_;
  wire _28889_;
  wire _28890_;
  wire _28891_;
  wire _28892_;
  wire _28893_;
  wire _28894_;
  wire _28895_;
  wire _28896_;
  wire _28897_;
  wire _28898_;
  wire _28899_;
  wire _28900_;
  wire _28901_;
  wire _28902_;
  wire _28903_;
  wire _28904_;
  wire _28905_;
  wire _28906_;
  wire _28907_;
  wire _28908_;
  wire _28909_;
  wire _28910_;
  wire _28911_;
  wire _28912_;
  wire _28913_;
  wire _28914_;
  wire _28915_;
  wire _28916_;
  wire _28917_;
  wire _28918_;
  wire _28919_;
  wire _28920_;
  wire _28921_;
  wire _28922_;
  wire _28923_;
  wire _28924_;
  wire _28925_;
  wire _28926_;
  wire _28927_;
  wire _28928_;
  wire _28929_;
  wire _28930_;
  wire _28931_;
  wire _28932_;
  wire _28933_;
  wire _28934_;
  wire _28935_;
  wire _28936_;
  wire _28937_;
  wire _28938_;
  wire _28939_;
  wire _28940_;
  wire _28941_;
  wire _28942_;
  wire _28943_;
  wire _28944_;
  wire _28945_;
  wire _28946_;
  wire _28947_;
  wire _28948_;
  wire _28949_;
  wire _28950_;
  wire _28951_;
  wire _28952_;
  wire _28953_;
  wire _28954_;
  wire _28955_;
  wire _28956_;
  wire _28957_;
  wire _28958_;
  wire _28959_;
  wire _28960_;
  wire _28961_;
  wire _28962_;
  wire _28963_;
  wire _28964_;
  wire _28965_;
  wire _28966_;
  wire _28967_;
  wire _28968_;
  wire _28969_;
  wire _28970_;
  wire _28971_;
  wire _28972_;
  wire _28973_;
  wire _28974_;
  wire _28975_;
  wire _28976_;
  wire _28977_;
  wire _28978_;
  wire _28979_;
  wire _28980_;
  wire _28981_;
  wire _28982_;
  wire _28983_;
  wire _28984_;
  wire _28985_;
  wire _28986_;
  wire _28987_;
  wire _28988_;
  wire _28989_;
  wire _28990_;
  wire _28991_;
  wire _28992_;
  wire _28993_;
  wire _28994_;
  wire _28995_;
  wire _28996_;
  wire _28997_;
  wire _28998_;
  wire _28999_;
  wire _29000_;
  wire _29001_;
  wire _29002_;
  wire _29003_;
  wire _29004_;
  wire _29005_;
  wire _29006_;
  wire _29007_;
  wire _29008_;
  wire _29009_;
  wire _29010_;
  wire _29011_;
  wire _29012_;
  wire _29013_;
  wire _29014_;
  wire _29015_;
  wire _29016_;
  wire _29017_;
  wire _29018_;
  wire _29019_;
  wire _29020_;
  wire _29021_;
  wire _29022_;
  wire _29023_;
  wire _29024_;
  wire _29025_;
  wire _29026_;
  wire _29027_;
  wire _29028_;
  wire _29029_;
  wire _29030_;
  wire _29031_;
  wire _29032_;
  wire _29033_;
  wire _29034_;
  wire _29035_;
  wire _29036_;
  wire _29037_;
  wire _29038_;
  wire _29039_;
  wire _29040_;
  wire _29041_;
  wire _29042_;
  wire _29043_;
  wire _29044_;
  wire _29045_;
  wire _29046_;
  wire _29047_;
  wire _29048_;
  wire _29049_;
  wire _29050_;
  wire _29051_;
  wire _29052_;
  wire _29053_;
  wire _29054_;
  wire _29055_;
  wire _29056_;
  wire _29057_;
  wire _29058_;
  wire _29059_;
  wire _29060_;
  wire _29061_;
  wire _29062_;
  wire _29063_;
  wire _29064_;
  wire _29065_;
  wire _29066_;
  wire _29067_;
  wire _29068_;
  wire _29069_;
  wire _29070_;
  wire _29071_;
  wire _29072_;
  wire _29073_;
  wire _29074_;
  wire _29075_;
  wire _29076_;
  wire _29077_;
  wire _29078_;
  wire _29079_;
  wire _29080_;
  wire _29081_;
  wire _29082_;
  wire _29083_;
  wire _29084_;
  wire _29085_;
  wire _29086_;
  wire _29087_;
  wire _29088_;
  wire _29089_;
  wire _29090_;
  wire _29091_;
  wire _29092_;
  wire _29093_;
  wire _29094_;
  wire _29095_;
  wire _29096_;
  wire _29097_;
  wire _29098_;
  wire _29099_;
  wire _29100_;
  wire _29101_;
  wire _29102_;
  wire _29103_;
  wire _29104_;
  wire _29105_;
  wire _29106_;
  wire _29107_;
  wire _29108_;
  wire _29109_;
  wire _29110_;
  wire _29111_;
  wire _29112_;
  wire _29113_;
  wire _29114_;
  wire _29115_;
  wire _29116_;
  wire _29117_;
  wire _29118_;
  wire _29119_;
  wire _29120_;
  wire _29121_;
  wire _29122_;
  wire _29123_;
  wire _29124_;
  wire _29125_;
  wire _29126_;
  wire _29127_;
  wire _29128_;
  wire _29129_;
  wire _29130_;
  wire _29131_;
  wire _29132_;
  wire _29133_;
  wire _29134_;
  wire _29135_;
  wire _29136_;
  wire _29137_;
  wire _29138_;
  wire _29139_;
  wire _29140_;
  wire _29141_;
  wire _29142_;
  wire _29143_;
  wire _29144_;
  wire _29145_;
  wire _29146_;
  wire _29147_;
  wire _29148_;
  wire _29149_;
  wire _29150_;
  wire _29151_;
  wire _29152_;
  wire _29153_;
  wire _29154_;
  wire _29155_;
  wire _29156_;
  wire _29157_;
  wire _29158_;
  wire _29159_;
  wire _29160_;
  wire _29161_;
  wire _29162_;
  wire _29163_;
  wire _29164_;
  wire _29165_;
  wire _29166_;
  wire _29167_;
  wire _29168_;
  wire _29169_;
  wire _29170_;
  wire _29171_;
  wire _29172_;
  wire _29173_;
  wire _29174_;
  wire _29175_;
  wire _29176_;
  wire _29177_;
  wire _29178_;
  wire _29179_;
  wire _29180_;
  wire _29181_;
  wire _29182_;
  wire _29183_;
  wire _29184_;
  wire _29185_;
  wire _29186_;
  wire _29187_;
  wire _29188_;
  wire _29189_;
  wire _29190_;
  wire _29191_;
  wire _29192_;
  wire _29193_;
  wire _29194_;
  wire _29195_;
  wire _29196_;
  wire _29197_;
  wire _29198_;
  wire _29199_;
  wire _29200_;
  wire _29201_;
  wire _29202_;
  wire _29203_;
  wire _29204_;
  wire _29205_;
  wire _29206_;
  wire _29207_;
  wire _29208_;
  wire _29209_;
  wire _29210_;
  wire _29211_;
  wire _29212_;
  wire _29213_;
  wire _29214_;
  wire _29215_;
  wire _29216_;
  wire _29217_;
  wire _29218_;
  wire _29219_;
  wire _29220_;
  wire _29221_;
  wire _29222_;
  wire _29223_;
  wire _29224_;
  wire _29225_;
  wire _29226_;
  wire _29227_;
  wire _29228_;
  wire _29229_;
  wire _29230_;
  wire _29231_;
  wire _29232_;
  wire _29233_;
  wire _29234_;
  wire _29235_;
  wire _29236_;
  wire _29237_;
  wire _29238_;
  wire _29239_;
  wire _29240_;
  wire _29241_;
  wire _29242_;
  wire _29243_;
  wire _29244_;
  wire _29245_;
  wire _29246_;
  wire _29247_;
  wire _29248_;
  wire _29249_;
  wire _29250_;
  wire _29251_;
  wire _29252_;
  wire _29253_;
  wire _29254_;
  wire _29255_;
  wire _29256_;
  wire _29257_;
  wire _29258_;
  wire _29259_;
  wire _29260_;
  wire _29261_;
  wire _29262_;
  wire _29263_;
  wire _29264_;
  wire _29265_;
  wire _29266_;
  wire _29267_;
  wire _29268_;
  wire _29269_;
  wire _29270_;
  wire _29271_;
  wire _29272_;
  wire _29273_;
  wire _29274_;
  wire _29275_;
  wire _29276_;
  wire _29277_;
  wire _29278_;
  wire _29279_;
  wire _29280_;
  wire _29281_;
  wire _29282_;
  wire _29283_;
  wire _29284_;
  wire _29285_;
  wire _29286_;
  wire _29287_;
  wire _29288_;
  wire _29289_;
  wire _29290_;
  wire _29291_;
  wire _29292_;
  wire _29293_;
  wire _29294_;
  wire _29295_;
  wire _29296_;
  wire _29297_;
  wire _29298_;
  wire _29299_;
  wire _29300_;
  wire _29301_;
  wire _29302_;
  wire _29303_;
  wire _29304_;
  wire _29305_;
  wire _29306_;
  wire _29307_;
  wire _29308_;
  wire _29309_;
  wire _29310_;
  wire _29311_;
  wire _29312_;
  wire _29313_;
  wire _29314_;
  wire _29315_;
  wire _29316_;
  wire _29317_;
  wire _29318_;
  wire _29319_;
  wire _29320_;
  wire _29321_;
  wire _29322_;
  wire _29323_;
  wire _29324_;
  wire _29325_;
  wire _29326_;
  wire _29327_;
  wire _29328_;
  wire _29329_;
  wire _29330_;
  wire _29331_;
  wire _29332_;
  wire _29333_;
  wire _29334_;
  wire _29335_;
  wire _29336_;
  wire _29337_;
  wire _29338_;
  wire _29339_;
  wire _29340_;
  wire _29341_;
  wire _29342_;
  wire _29343_;
  wire _29344_;
  wire _29345_;
  wire _29346_;
  wire _29347_;
  wire _29348_;
  wire _29349_;
  wire _29350_;
  wire _29351_;
  wire _29352_;
  wire _29353_;
  wire _29354_;
  wire _29355_;
  wire _29356_;
  wire _29357_;
  wire _29358_;
  wire _29359_;
  wire _29360_;
  wire _29361_;
  wire _29362_;
  wire _29363_;
  wire _29364_;
  wire _29365_;
  wire _29366_;
  wire _29367_;
  wire _29368_;
  wire _29369_;
  wire _29370_;
  wire _29371_;
  wire _29372_;
  wire _29373_;
  wire _29374_;
  wire _29375_;
  wire _29376_;
  wire _29377_;
  wire _29378_;
  wire _29379_;
  wire _29380_;
  wire _29381_;
  wire _29382_;
  wire _29383_;
  wire _29384_;
  wire _29385_;
  wire _29386_;
  wire _29387_;
  wire _29388_;
  wire _29389_;
  wire _29390_;
  wire _29391_;
  wire _29392_;
  wire _29393_;
  wire _29394_;
  wire _29395_;
  wire _29396_;
  wire _29397_;
  wire _29398_;
  wire _29399_;
  wire _29400_;
  wire _29401_;
  wire _29402_;
  wire _29403_;
  wire _29404_;
  wire _29405_;
  wire _29406_;
  wire _29407_;
  wire _29408_;
  wire _29409_;
  wire _29410_;
  wire _29411_;
  wire _29412_;
  wire _29413_;
  wire _29414_;
  wire _29415_;
  wire _29416_;
  wire _29417_;
  wire _29418_;
  wire _29419_;
  wire _29420_;
  wire _29421_;
  wire _29422_;
  wire _29423_;
  wire _29424_;
  wire _29425_;
  wire _29426_;
  wire _29427_;
  wire _29428_;
  wire _29429_;
  wire _29430_;
  wire _29431_;
  wire _29432_;
  wire _29433_;
  wire _29434_;
  wire _29435_;
  wire _29436_;
  wire _29437_;
  wire _29438_;
  wire _29439_;
  wire _29440_;
  wire _29441_;
  wire _29442_;
  wire _29443_;
  wire _29444_;
  wire _29445_;
  wire _29446_;
  wire _29447_;
  wire _29448_;
  wire _29449_;
  wire _29450_;
  wire _29451_;
  wire _29452_;
  wire _29453_;
  wire _29454_;
  wire _29455_;
  wire _29456_;
  wire _29457_;
  wire _29458_;
  wire _29459_;
  wire _29460_;
  wire _29461_;
  wire _29462_;
  wire _29463_;
  wire _29464_;
  wire _29465_;
  wire _29466_;
  wire _29467_;
  wire _29468_;
  wire _29469_;
  wire _29470_;
  wire _29471_;
  wire _29472_;
  wire _29473_;
  wire _29474_;
  wire _29475_;
  wire _29476_;
  wire _29477_;
  wire _29478_;
  wire _29479_;
  wire _29480_;
  wire _29481_;
  wire _29482_;
  wire _29483_;
  wire _29484_;
  wire _29485_;
  wire _29486_;
  wire _29487_;
  wire _29488_;
  wire _29489_;
  wire _29490_;
  wire _29491_;
  wire _29492_;
  wire _29493_;
  wire _29494_;
  wire _29495_;
  wire _29496_;
  wire _29497_;
  wire _29498_;
  wire _29499_;
  wire _29500_;
  wire _29501_;
  wire _29502_;
  wire _29503_;
  wire _29504_;
  wire _29505_;
  wire _29506_;
  wire _29507_;
  wire _29508_;
  wire _29509_;
  wire _29510_;
  wire _29511_;
  wire _29512_;
  wire _29513_;
  wire _29514_;
  wire _29515_;
  wire _29516_;
  wire _29517_;
  wire _29518_;
  wire _29519_;
  wire _29520_;
  wire _29521_;
  wire _29522_;
  wire _29523_;
  wire _29524_;
  wire _29525_;
  wire _29526_;
  wire _29527_;
  wire _29528_;
  wire _29529_;
  wire _29530_;
  wire _29531_;
  wire _29532_;
  wire _29533_;
  wire _29534_;
  wire _29535_;
  wire _29536_;
  wire _29537_;
  wire _29538_;
  wire _29539_;
  wire _29540_;
  wire _29541_;
  wire _29542_;
  wire _29543_;
  wire _29544_;
  wire _29545_;
  wire _29546_;
  wire _29547_;
  wire _29548_;
  wire _29549_;
  wire _29550_;
  wire _29551_;
  wire _29552_;
  wire _29553_;
  wire _29554_;
  wire _29555_;
  wire _29556_;
  wire _29557_;
  wire _29558_;
  wire _29559_;
  wire _29560_;
  wire _29561_;
  wire _29562_;
  wire _29563_;
  wire _29564_;
  wire _29565_;
  wire _29566_;
  wire _29567_;
  wire _29568_;
  wire _29569_;
  wire _29570_;
  wire _29571_;
  wire _29572_;
  wire _29573_;
  wire _29574_;
  wire _29575_;
  wire _29576_;
  wire _29577_;
  wire _29578_;
  wire _29579_;
  wire _29580_;
  wire _29581_;
  wire _29582_;
  wire _29583_;
  wire _29584_;
  wire _29585_;
  wire _29586_;
  wire _29587_;
  wire _29588_;
  wire _29589_;
  wire _29590_;
  wire _29591_;
  wire _29592_;
  wire _29593_;
  wire _29594_;
  wire _29595_;
  wire _29596_;
  wire _29597_;
  wire _29598_;
  wire _29599_;
  wire _29600_;
  wire _29601_;
  wire _29602_;
  wire _29603_;
  wire _29604_;
  wire _29605_;
  wire _29606_;
  wire _29607_;
  wire _29608_;
  wire _29609_;
  wire _29610_;
  wire _29611_;
  wire _29612_;
  wire _29613_;
  wire _29614_;
  wire _29615_;
  wire _29616_;
  wire _29617_;
  wire _29618_;
  wire _29619_;
  wire _29620_;
  wire _29621_;
  wire _29622_;
  wire _29623_;
  wire _29624_;
  wire _29625_;
  wire _29626_;
  wire _29627_;
  wire _29628_;
  wire _29629_;
  wire _29630_;
  wire _29631_;
  wire _29632_;
  wire _29633_;
  wire _29634_;
  wire _29635_;
  wire _29636_;
  wire _29637_;
  wire _29638_;
  wire _29639_;
  wire _29640_;
  wire _29641_;
  wire _29642_;
  wire _29643_;
  wire _29644_;
  wire _29645_;
  wire _29646_;
  wire _29647_;
  wire _29648_;
  wire _29649_;
  wire _29650_;
  wire _29651_;
  wire _29652_;
  wire _29653_;
  wire _29654_;
  wire _29655_;
  wire _29656_;
  wire _29657_;
  wire _29658_;
  wire _29659_;
  wire _29660_;
  wire _29661_;
  wire _29662_;
  wire _29663_;
  wire _29664_;
  wire _29665_;
  wire _29666_;
  wire _29667_;
  wire _29668_;
  wire _29669_;
  wire _29670_;
  wire _29671_;
  wire _29672_;
  wire _29673_;
  wire _29674_;
  wire _29675_;
  wire _29676_;
  wire _29677_;
  wire _29678_;
  wire _29679_;
  wire _29680_;
  wire _29681_;
  wire _29682_;
  wire _29683_;
  wire _29684_;
  wire _29685_;
  wire _29686_;
  wire _29687_;
  wire _29688_;
  wire _29689_;
  wire _29690_;
  wire _29691_;
  wire _29692_;
  wire _29693_;
  wire _29694_;
  wire _29695_;
  wire _29696_;
  wire _29697_;
  wire _29698_;
  wire _29699_;
  wire _29700_;
  wire _29701_;
  wire _29702_;
  wire _29703_;
  wire _29704_;
  wire _29705_;
  wire _29706_;
  wire _29707_;
  wire _29708_;
  wire _29709_;
  wire _29710_;
  wire _29711_;
  wire _29712_;
  wire _29713_;
  wire _29714_;
  wire _29715_;
  wire _29716_;
  wire _29717_;
  wire _29718_;
  wire _29719_;
  wire _29720_;
  wire _29721_;
  wire _29722_;
  wire _29723_;
  wire _29724_;
  wire _29725_;
  wire _29726_;
  wire _29727_;
  wire _29728_;
  wire _29729_;
  wire _29730_;
  wire _29731_;
  wire _29732_;
  wire _29733_;
  wire _29734_;
  wire _29735_;
  wire _29736_;
  wire _29737_;
  wire _29738_;
  wire _29739_;
  wire _29740_;
  wire _29741_;
  wire _29742_;
  wire _29743_;
  wire _29744_;
  wire _29745_;
  wire _29746_;
  wire _29747_;
  wire _29748_;
  wire _29749_;
  wire _29750_;
  wire _29751_;
  wire _29752_;
  wire _29753_;
  wire _29754_;
  wire _29755_;
  wire _29756_;
  wire _29757_;
  wire _29758_;
  wire _29759_;
  wire _29760_;
  wire _29761_;
  wire _29762_;
  wire _29763_;
  wire _29764_;
  wire _29765_;
  wire _29766_;
  wire _29767_;
  wire _29768_;
  wire _29769_;
  wire _29770_;
  wire _29771_;
  wire _29772_;
  wire _29773_;
  wire _29774_;
  wire _29775_;
  wire _29776_;
  wire _29777_;
  wire _29778_;
  wire _29779_;
  wire _29780_;
  wire _29781_;
  wire _29782_;
  wire _29783_;
  wire _29784_;
  wire _29785_;
  wire _29786_;
  wire _29787_;
  wire _29788_;
  wire _29789_;
  wire _29790_;
  wire _29791_;
  wire _29792_;
  wire _29793_;
  wire _29794_;
  wire _29795_;
  wire _29796_;
  wire _29797_;
  wire _29798_;
  wire _29799_;
  wire _29800_;
  wire _29801_;
  wire _29802_;
  wire _29803_;
  wire _29804_;
  wire _29805_;
  wire _29806_;
  wire _29807_;
  wire _29808_;
  wire _29809_;
  wire _29810_;
  wire _29811_;
  wire _29812_;
  wire _29813_;
  wire _29814_;
  wire _29815_;
  wire _29816_;
  wire _29817_;
  wire _29818_;
  wire _29819_;
  wire _29820_;
  wire _29821_;
  wire _29822_;
  wire _29823_;
  wire _29824_;
  wire _29825_;
  wire _29826_;
  wire _29827_;
  wire _29828_;
  wire _29829_;
  wire _29830_;
  wire _29831_;
  wire _29832_;
  wire _29833_;
  wire _29834_;
  wire _29835_;
  wire _29836_;
  wire _29837_;
  wire _29838_;
  wire _29839_;
  wire _29840_;
  wire _29841_;
  wire _29842_;
  wire _29843_;
  wire _29844_;
  wire _29845_;
  wire _29846_;
  wire _29847_;
  wire _29848_;
  wire _29849_;
  wire _29850_;
  wire _29851_;
  wire _29852_;
  wire _29853_;
  wire _29854_;
  wire _29855_;
  wire _29856_;
  wire _29857_;
  wire _29858_;
  wire _29859_;
  wire _29860_;
  wire _29861_;
  wire _29862_;
  wire _29863_;
  wire _29864_;
  wire _29865_;
  wire _29866_;
  wire _29867_;
  wire _29868_;
  wire _29869_;
  wire _29870_;
  wire _29871_;
  wire _29872_;
  wire _29873_;
  wire _29874_;
  wire _29875_;
  wire _29876_;
  wire _29877_;
  wire _29878_;
  wire _29879_;
  wire _29880_;
  wire _29881_;
  wire _29882_;
  wire _29883_;
  wire _29884_;
  wire _29885_;
  wire _29886_;
  wire _29887_;
  wire _29888_;
  wire _29889_;
  wire _29890_;
  wire _29891_;
  wire _29892_;
  wire _29893_;
  wire _29894_;
  wire _29895_;
  wire _29896_;
  wire _29897_;
  wire _29898_;
  wire _29899_;
  wire _29900_;
  wire _29901_;
  wire _29902_;
  wire _29903_;
  wire _29904_;
  wire _29905_;
  wire _29906_;
  wire _29907_;
  wire _29908_;
  wire _29909_;
  wire _29910_;
  wire _29911_;
  wire _29912_;
  wire _29913_;
  wire _29914_;
  wire _29915_;
  wire _29916_;
  wire _29917_;
  wire _29918_;
  wire _29919_;
  wire _29920_;
  wire _29921_;
  wire _29922_;
  wire _29923_;
  wire _29924_;
  wire _29925_;
  wire _29926_;
  wire _29927_;
  wire _29928_;
  wire _29929_;
  wire _29930_;
  wire _29931_;
  wire _29932_;
  wire _29933_;
  wire _29934_;
  wire _29935_;
  wire _29936_;
  wire _29937_;
  wire _29938_;
  wire _29939_;
  wire _29940_;
  wire _29941_;
  wire _29942_;
  wire _29943_;
  wire _29944_;
  wire _29945_;
  wire _29946_;
  wire _29947_;
  wire _29948_;
  wire _29949_;
  wire _29950_;
  wire _29951_;
  wire _29952_;
  wire _29953_;
  wire _29954_;
  wire _29955_;
  wire _29956_;
  wire _29957_;
  wire _29958_;
  wire _29959_;
  wire _29960_;
  wire _29961_;
  wire _29962_;
  wire _29963_;
  wire _29964_;
  wire _29965_;
  wire _29966_;
  wire _29967_;
  wire _29968_;
  wire _29969_;
  wire _29970_;
  wire _29971_;
  wire _29972_;
  wire _29973_;
  wire _29974_;
  wire _29975_;
  wire _29976_;
  wire _29977_;
  wire _29978_;
  wire _29979_;
  wire _29980_;
  wire _29981_;
  wire _29982_;
  wire _29983_;
  wire _29984_;
  wire _29985_;
  wire _29986_;
  wire _29987_;
  wire _29988_;
  wire _29989_;
  wire _29990_;
  wire _29991_;
  wire _29992_;
  wire _29993_;
  wire _29994_;
  wire _29995_;
  wire _29996_;
  wire _29997_;
  wire _29998_;
  wire _29999_;
  wire _30000_;
  wire _30001_;
  wire _30002_;
  wire _30003_;
  wire _30004_;
  wire _30005_;
  wire _30006_;
  wire _30007_;
  wire _30008_;
  wire _30009_;
  wire _30010_;
  wire _30011_;
  wire _30012_;
  wire _30013_;
  wire _30014_;
  wire _30015_;
  wire _30016_;
  wire _30017_;
  wire _30018_;
  wire _30019_;
  wire _30020_;
  wire _30021_;
  wire _30022_;
  wire _30023_;
  wire _30024_;
  wire _30025_;
  wire _30026_;
  wire _30027_;
  wire _30028_;
  wire _30029_;
  wire _30030_;
  wire _30031_;
  wire _30032_;
  wire _30033_;
  wire _30034_;
  wire _30035_;
  wire _30036_;
  wire _30037_;
  wire _30038_;
  wire _30039_;
  wire _30040_;
  wire _30041_;
  wire _30042_;
  wire _30043_;
  wire _30044_;
  wire _30045_;
  wire _30046_;
  wire _30047_;
  wire _30048_;
  wire _30049_;
  wire _30050_;
  wire _30051_;
  wire _30052_;
  wire _30053_;
  wire _30054_;
  wire _30055_;
  wire _30056_;
  wire _30057_;
  wire _30058_;
  wire _30059_;
  wire _30060_;
  wire _30061_;
  wire _30062_;
  wire _30063_;
  wire _30064_;
  wire _30065_;
  wire _30066_;
  wire _30067_;
  wire _30068_;
  wire _30069_;
  wire _30070_;
  wire _30071_;
  wire _30072_;
  wire _30073_;
  wire _30074_;
  wire _30075_;
  wire _30076_;
  wire _30077_;
  wire _30078_;
  wire _30079_;
  wire _30080_;
  wire _30081_;
  wire _30082_;
  wire _30083_;
  wire _30084_;
  wire _30085_;
  wire _30086_;
  wire _30087_;
  wire _30088_;
  wire _30089_;
  wire _30090_;
  wire _30091_;
  wire _30092_;
  wire _30093_;
  wire _30094_;
  wire _30095_;
  wire _30096_;
  wire _30097_;
  wire _30098_;
  wire _30099_;
  wire _30100_;
  wire _30101_;
  wire _30102_;
  wire _30103_;
  wire _30104_;
  wire _30105_;
  wire _30106_;
  wire _30107_;
  wire _30108_;
  wire _30109_;
  wire _30110_;
  wire _30111_;
  wire _30112_;
  wire _30113_;
  wire _30114_;
  wire _30115_;
  wire _30116_;
  wire _30117_;
  wire _30118_;
  wire _30119_;
  wire _30120_;
  wire _30121_;
  wire _30122_;
  wire _30123_;
  wire _30124_;
  wire _30125_;
  wire _30126_;
  wire _30127_;
  wire _30128_;
  wire _30129_;
  wire _30130_;
  wire _30131_;
  wire _30132_;
  wire _30133_;
  wire _30134_;
  wire _30135_;
  wire _30136_;
  wire _30137_;
  wire _30138_;
  wire _30139_;
  wire _30140_;
  wire _30141_;
  wire _30142_;
  wire _30143_;
  wire _30144_;
  wire _30145_;
  wire _30146_;
  wire _30147_;
  wire _30148_;
  wire _30149_;
  wire _30150_;
  wire _30151_;
  wire _30152_;
  wire _30153_;
  wire _30154_;
  wire _30155_;
  wire _30156_;
  wire _30157_;
  wire _30158_;
  wire _30159_;
  wire _30160_;
  wire _30161_;
  wire _30162_;
  wire _30163_;
  wire _30164_;
  wire _30165_;
  wire _30166_;
  wire _30167_;
  wire _30168_;
  wire _30169_;
  wire _30170_;
  wire _30171_;
  wire _30172_;
  wire _30173_;
  wire _30174_;
  wire _30175_;
  wire _30176_;
  wire _30177_;
  wire _30178_;
  wire _30179_;
  wire _30180_;
  wire _30181_;
  wire _30182_;
  wire _30183_;
  wire _30184_;
  wire _30185_;
  wire _30186_;
  wire _30187_;
  wire _30188_;
  wire _30189_;
  wire _30190_;
  wire _30191_;
  wire _30192_;
  wire _30193_;
  wire _30194_;
  wire _30195_;
  wire _30196_;
  wire _30197_;
  wire _30198_;
  wire _30199_;
  wire _30200_;
  wire _30201_;
  wire _30202_;
  wire _30203_;
  wire _30204_;
  wire _30205_;
  wire _30206_;
  wire _30207_;
  wire _30208_;
  wire _30209_;
  wire _30210_;
  wire _30211_;
  wire _30212_;
  wire _30213_;
  wire _30214_;
  wire _30215_;
  wire _30216_;
  wire _30217_;
  wire _30218_;
  wire _30219_;
  wire _30220_;
  wire _30221_;
  wire _30222_;
  wire _30223_;
  wire _30224_;
  wire _30225_;
  wire _30226_;
  wire _30227_;
  wire _30228_;
  wire _30229_;
  wire _30230_;
  wire _30231_;
  wire _30232_;
  wire _30233_;
  wire _30234_;
  wire _30235_;
  wire _30236_;
  wire _30237_;
  wire _30238_;
  wire _30239_;
  wire _30240_;
  wire _30241_;
  wire _30242_;
  wire _30243_;
  wire _30244_;
  wire _30245_;
  wire _30246_;
  wire _30247_;
  wire _30248_;
  wire _30249_;
  wire _30250_;
  wire _30251_;
  wire _30252_;
  wire _30253_;
  wire _30254_;
  wire _30255_;
  wire _30256_;
  wire _30257_;
  wire _30258_;
  wire _30259_;
  wire _30260_;
  wire _30261_;
  wire _30262_;
  wire _30263_;
  wire _30264_;
  wire _30265_;
  wire _30266_;
  wire _30267_;
  wire _30268_;
  wire _30269_;
  wire _30270_;
  wire _30271_;
  wire _30272_;
  wire _30273_;
  wire _30274_;
  wire _30275_;
  wire _30276_;
  wire _30277_;
  wire _30278_;
  wire _30279_;
  wire _30280_;
  wire _30281_;
  wire _30282_;
  wire _30283_;
  wire _30284_;
  wire _30285_;
  wire _30286_;
  wire _30287_;
  wire _30288_;
  wire _30289_;
  wire _30290_;
  wire _30291_;
  wire _30292_;
  wire _30293_;
  wire _30294_;
  wire _30295_;
  wire _30296_;
  wire _30297_;
  wire _30298_;
  wire _30299_;
  wire _30300_;
  wire _30301_;
  wire _30302_;
  wire _30303_;
  wire _30304_;
  wire _30305_;
  wire _30306_;
  wire _30307_;
  wire _30308_;
  wire _30309_;
  wire _30310_;
  wire _30311_;
  wire _30312_;
  wire _30313_;
  wire _30314_;
  wire _30315_;
  wire _30316_;
  wire _30317_;
  wire _30318_;
  wire _30319_;
  wire _30320_;
  wire _30321_;
  wire _30322_;
  wire _30323_;
  wire _30324_;
  wire _30325_;
  wire _30326_;
  wire _30327_;
  wire _30328_;
  wire _30329_;
  wire _30330_;
  wire _30331_;
  wire _30332_;
  wire _30333_;
  wire _30334_;
  wire _30335_;
  wire _30336_;
  wire _30337_;
  wire _30338_;
  wire _30339_;
  wire _30340_;
  wire _30341_;
  wire _30342_;
  wire _30343_;
  wire _30344_;
  wire _30345_;
  wire _30346_;
  wire _30347_;
  wire _30348_;
  wire _30349_;
  wire _30350_;
  wire _30351_;
  wire _30352_;
  wire _30353_;
  wire _30354_;
  wire _30355_;
  wire _30356_;
  wire _30357_;
  wire _30358_;
  wire _30359_;
  wire _30360_;
  wire _30361_;
  wire _30362_;
  wire _30363_;
  wire _30364_;
  wire _30365_;
  wire _30366_;
  wire _30367_;
  wire _30368_;
  wire _30369_;
  wire _30370_;
  wire _30371_;
  wire _30372_;
  wire _30373_;
  wire _30374_;
  wire _30375_;
  wire _30376_;
  wire _30377_;
  wire _30378_;
  wire _30379_;
  wire _30380_;
  wire _30381_;
  wire _30382_;
  wire _30383_;
  wire _30384_;
  wire _30385_;
  wire _30386_;
  wire _30387_;
  wire _30388_;
  wire _30389_;
  wire _30390_;
  wire _30391_;
  wire _30392_;
  wire _30393_;
  wire _30394_;
  wire _30395_;
  wire _30396_;
  wire _30397_;
  wire _30398_;
  wire _30399_;
  wire _30400_;
  wire _30401_;
  wire _30402_;
  wire _30403_;
  wire _30404_;
  wire _30405_;
  wire _30406_;
  wire _30407_;
  wire _30408_;
  wire _30409_;
  wire _30410_;
  wire _30411_;
  wire _30412_;
  wire _30413_;
  wire _30414_;
  wire _30415_;
  wire _30416_;
  wire _30417_;
  wire _30418_;
  wire _30419_;
  wire _30420_;
  wire _30421_;
  wire _30422_;
  wire _30423_;
  wire _30424_;
  wire _30425_;
  wire _30426_;
  wire _30427_;
  wire _30428_;
  wire _30429_;
  wire _30430_;
  wire _30431_;
  wire _30432_;
  wire _30433_;
  wire _30434_;
  wire _30435_;
  wire _30436_;
  wire _30437_;
  wire _30438_;
  wire _30439_;
  wire _30440_;
  wire _30441_;
  wire _30442_;
  wire _30443_;
  wire _30444_;
  wire _30445_;
  wire _30446_;
  wire _30447_;
  wire _30448_;
  wire _30449_;
  wire _30450_;
  wire _30451_;
  wire _30452_;
  wire _30453_;
  wire _30454_;
  wire _30455_;
  wire _30456_;
  wire _30457_;
  wire _30458_;
  wire _30459_;
  wire _30460_;
  wire _30461_;
  wire _30462_;
  wire _30463_;
  wire _30464_;
  wire _30465_;
  wire _30466_;
  wire _30467_;
  wire _30468_;
  wire _30469_;
  wire _30470_;
  wire _30471_;
  wire _30472_;
  wire _30473_;
  wire _30474_;
  wire _30475_;
  wire _30476_;
  wire _30477_;
  wire _30478_;
  wire _30479_;
  wire _30480_;
  wire _30481_;
  wire _30482_;
  wire _30483_;
  wire _30484_;
  wire _30485_;
  wire _30486_;
  wire _30487_;
  wire _30488_;
  wire _30489_;
  wire _30490_;
  wire _30491_;
  wire _30492_;
  wire _30493_;
  wire _30494_;
  wire _30495_;
  wire _30496_;
  wire _30497_;
  wire _30498_;
  wire _30499_;
  wire _30500_;
  wire _30501_;
  wire _30502_;
  wire _30503_;
  wire _30504_;
  wire _30505_;
  wire _30506_;
  wire _30507_;
  wire _30508_;
  wire _30509_;
  wire _30510_;
  wire _30511_;
  wire _30512_;
  wire _30513_;
  wire _30514_;
  wire _30515_;
  wire _30516_;
  wire _30517_;
  wire _30518_;
  wire _30519_;
  wire _30520_;
  wire _30521_;
  wire _30522_;
  wire _30523_;
  wire _30524_;
  wire _30525_;
  wire _30526_;
  wire _30527_;
  wire _30528_;
  wire _30529_;
  wire _30530_;
  wire _30531_;
  wire _30532_;
  wire _30533_;
  wire _30534_;
  wire _30535_;
  wire _30536_;
  wire _30537_;
  wire _30538_;
  wire _30539_;
  wire _30540_;
  wire _30541_;
  wire _30542_;
  wire _30543_;
  wire _30544_;
  wire _30545_;
  wire _30546_;
  wire _30547_;
  wire _30548_;
  wire _30549_;
  wire _30550_;
  wire _30551_;
  wire _30552_;
  wire _30553_;
  wire _30554_;
  wire _30555_;
  wire _30556_;
  wire _30557_;
  wire _30558_;
  wire _30559_;
  wire _30560_;
  wire _30561_;
  wire _30562_;
  wire _30563_;
  wire _30564_;
  wire _30565_;
  wire _30566_;
  wire _30567_;
  wire _30568_;
  wire _30569_;
  wire _30570_;
  wire _30571_;
  wire _30572_;
  wire _30573_;
  wire _30574_;
  wire _30575_;
  wire _30576_;
  wire _30577_;
  wire _30578_;
  wire _30579_;
  wire _30580_;
  wire _30581_;
  wire _30582_;
  wire _30583_;
  wire _30584_;
  wire _30585_;
  wire _30586_;
  wire _30587_;
  wire _30588_;
  wire _30589_;
  wire _30590_;
  wire _30591_;
  wire _30592_;
  wire _30593_;
  wire _30594_;
  wire _30595_;
  wire _30596_;
  wire _30597_;
  wire _30598_;
  wire _30599_;
  wire _30600_;
  wire _30601_;
  wire _30602_;
  wire _30603_;
  wire _30604_;
  wire _30605_;
  wire _30606_;
  wire _30607_;
  wire _30608_;
  wire _30609_;
  wire _30610_;
  wire _30611_;
  wire _30612_;
  wire _30613_;
  wire _30614_;
  wire _30615_;
  wire _30616_;
  wire _30617_;
  wire _30618_;
  wire _30619_;
  wire _30620_;
  wire _30621_;
  wire _30622_;
  wire _30623_;
  wire _30624_;
  wire _30625_;
  wire _30626_;
  wire _30627_;
  wire _30628_;
  wire _30629_;
  wire _30630_;
  wire _30631_;
  wire _30632_;
  wire _30633_;
  wire _30634_;
  wire _30635_;
  wire _30636_;
  wire _30637_;
  wire _30638_;
  wire _30639_;
  wire _30640_;
  wire _30641_;
  wire _30642_;
  wire _30643_;
  wire _30644_;
  wire _30645_;
  wire _30646_;
  wire _30647_;
  wire _30648_;
  wire _30649_;
  wire _30650_;
  wire _30651_;
  wire _30652_;
  wire _30653_;
  wire _30654_;
  wire _30655_;
  wire _30656_;
  wire _30657_;
  wire _30658_;
  wire _30659_;
  wire _30660_;
  wire _30661_;
  wire _30662_;
  wire _30663_;
  wire _30664_;
  wire _30665_;
  wire _30666_;
  wire _30667_;
  wire _30668_;
  wire _30669_;
  wire _30670_;
  wire _30671_;
  wire _30672_;
  wire _30673_;
  wire _30674_;
  wire _30675_;
  wire _30676_;
  wire _30677_;
  wire _30678_;
  wire _30679_;
  wire _30680_;
  wire _30681_;
  wire _30682_;
  wire _30683_;
  wire _30684_;
  wire _30685_;
  wire _30686_;
  wire _30687_;
  wire _30688_;
  wire _30689_;
  wire _30690_;
  wire _30691_;
  wire _30692_;
  wire _30693_;
  wire _30694_;
  wire _30695_;
  wire _30696_;
  wire _30697_;
  wire _30698_;
  wire _30699_;
  wire _30700_;
  wire _30701_;
  wire _30702_;
  wire _30703_;
  wire _30704_;
  wire _30705_;
  wire _30706_;
  wire _30707_;
  wire _30708_;
  wire _30709_;
  wire _30710_;
  wire _30711_;
  wire _30712_;
  wire _30713_;
  wire _30714_;
  wire _30715_;
  wire _30716_;
  wire _30717_;
  wire _30718_;
  wire _30719_;
  wire _30720_;
  wire _30721_;
  wire _30722_;
  wire _30723_;
  wire _30724_;
  wire _30725_;
  wire _30726_;
  wire _30727_;
  wire _30728_;
  wire _30729_;
  wire _30730_;
  wire _30731_;
  wire _30732_;
  wire _30733_;
  wire _30734_;
  wire _30735_;
  wire _30736_;
  wire _30737_;
  wire _30738_;
  wire _30739_;
  wire _30740_;
  wire _30741_;
  wire _30742_;
  wire _30743_;
  wire _30744_;
  wire _30745_;
  wire _30746_;
  wire _30747_;
  wire _30748_;
  wire _30749_;
  wire _30750_;
  wire _30751_;
  wire _30752_;
  wire _30753_;
  wire _30754_;
  wire _30755_;
  wire _30756_;
  wire _30757_;
  wire _30758_;
  wire _30759_;
  wire _30760_;
  wire _30761_;
  wire _30762_;
  wire _30763_;
  wire _30764_;
  wire _30765_;
  wire _30766_;
  wire _30767_;
  wire _30768_;
  wire _30769_;
  wire _30770_;
  wire _30771_;
  wire _30772_;
  wire _30773_;
  wire _30774_;
  wire _30775_;
  wire _30776_;
  wire _30777_;
  wire _30778_;
  wire _30779_;
  wire _30780_;
  wire _30781_;
  wire _30782_;
  wire _30783_;
  wire _30784_;
  wire _30785_;
  wire _30786_;
  wire _30787_;
  wire _30788_;
  wire _30789_;
  wire _30790_;
  wire _30791_;
  wire _30792_;
  wire _30793_;
  wire _30794_;
  wire _30795_;
  wire _30796_;
  wire _30797_;
  wire _30798_;
  wire _30799_;
  wire _30800_;
  wire _30801_;
  wire _30802_;
  wire _30803_;
  wire _30804_;
  wire _30805_;
  wire _30806_;
  wire _30807_;
  wire _30808_;
  wire _30809_;
  wire _30810_;
  wire _30811_;
  wire _30812_;
  wire _30813_;
  wire _30814_;
  wire _30815_;
  wire _30816_;
  wire _30817_;
  wire _30818_;
  wire _30819_;
  wire _30820_;
  wire _30821_;
  wire _30822_;
  wire _30823_;
  wire _30824_;
  wire _30825_;
  wire _30826_;
  wire _30827_;
  wire _30828_;
  wire _30829_;
  wire _30830_;
  wire _30831_;
  wire _30832_;
  wire _30833_;
  wire _30834_;
  wire _30835_;
  wire _30836_;
  wire _30837_;
  wire _30838_;
  wire _30839_;
  wire _30840_;
  wire _30841_;
  wire _30842_;
  wire _30843_;
  wire _30844_;
  wire _30845_;
  wire _30846_;
  wire _30847_;
  wire _30848_;
  wire _30849_;
  wire _30850_;
  wire _30851_;
  wire _30852_;
  wire _30853_;
  wire _30854_;
  wire _30855_;
  wire _30856_;
  wire _30857_;
  wire _30858_;
  wire _30859_;
  wire _30860_;
  wire _30861_;
  wire _30862_;
  wire _30863_;
  wire _30864_;
  wire _30865_;
  wire _30866_;
  wire _30867_;
  wire _30868_;
  wire _30869_;
  wire _30870_;
  wire _30871_;
  wire _30872_;
  wire _30873_;
  wire _30874_;
  wire _30875_;
  wire _30876_;
  wire _30877_;
  wire _30878_;
  wire _30879_;
  wire _30880_;
  wire _30881_;
  wire _30882_;
  wire _30883_;
  wire _30884_;
  wire _30885_;
  wire _30886_;
  wire _30887_;
  wire _30888_;
  wire _30889_;
  wire _30890_;
  wire _30891_;
  wire _30892_;
  wire _30893_;
  wire _30894_;
  wire _30895_;
  wire _30896_;
  wire _30897_;
  wire _30898_;
  wire _30899_;
  wire _30900_;
  wire _30901_;
  wire _30902_;
  wire _30903_;
  wire _30904_;
  wire _30905_;
  wire _30906_;
  wire _30907_;
  wire _30908_;
  wire _30909_;
  wire _30910_;
  wire _30911_;
  wire _30912_;
  wire _30913_;
  wire _30914_;
  wire _30915_;
  wire _30916_;
  wire _30917_;
  wire _30918_;
  wire _30919_;
  wire _30920_;
  wire _30921_;
  wire _30922_;
  wire _30923_;
  wire _30924_;
  wire _30925_;
  wire _30926_;
  wire _30927_;
  wire _30928_;
  wire _30929_;
  wire _30930_;
  wire _30931_;
  wire _30932_;
  wire _30933_;
  wire _30934_;
  wire _30935_;
  wire _30936_;
  wire _30937_;
  wire _30938_;
  wire _30939_;
  wire _30940_;
  wire _30941_;
  wire _30942_;
  wire _30943_;
  wire _30944_;
  wire _30945_;
  wire _30946_;
  wire _30947_;
  wire _30948_;
  wire _30949_;
  wire _30950_;
  wire _30951_;
  wire _30952_;
  wire _30953_;
  wire _30954_;
  wire _30955_;
  wire _30956_;
  wire _30957_;
  wire _30958_;
  wire _30959_;
  wire _30960_;
  wire _30961_;
  wire _30962_;
  wire _30963_;
  wire _30964_;
  wire _30965_;
  wire _30966_;
  wire _30967_;
  wire _30968_;
  wire _30969_;
  wire _30970_;
  wire _30971_;
  wire _30972_;
  wire _30973_;
  wire _30974_;
  wire _30975_;
  wire _30976_;
  wire _30977_;
  wire _30978_;
  wire _30979_;
  wire _30980_;
  wire _30981_;
  wire _30982_;
  wire _30983_;
  wire _30984_;
  wire _30985_;
  wire _30986_;
  wire _30987_;
  wire _30988_;
  wire _30989_;
  wire _30990_;
  wire _30991_;
  wire _30992_;
  wire _30993_;
  wire _30994_;
  wire _30995_;
  wire _30996_;
  wire _30997_;
  wire _30998_;
  wire _30999_;
  wire _31000_;
  wire _31001_;
  wire _31002_;
  wire _31003_;
  wire _31004_;
  wire _31005_;
  wire _31006_;
  wire _31007_;
  wire _31008_;
  wire _31009_;
  wire _31010_;
  wire _31011_;
  wire _31012_;
  wire _31013_;
  wire _31014_;
  wire _31015_;
  wire _31016_;
  wire _31017_;
  wire _31018_;
  wire _31019_;
  wire _31020_;
  wire _31021_;
  wire _31022_;
  wire _31023_;
  wire _31024_;
  wire _31025_;
  wire _31026_;
  wire _31027_;
  wire _31028_;
  wire _31029_;
  wire _31030_;
  wire _31031_;
  wire _31032_;
  wire _31033_;
  wire _31034_;
  wire _31035_;
  wire _31036_;
  wire _31037_;
  wire _31038_;
  wire _31039_;
  wire _31040_;
  wire _31041_;
  wire _31042_;
  wire _31043_;
  wire _31044_;
  wire _31045_;
  wire _31046_;
  wire _31047_;
  wire _31048_;
  wire _31049_;
  wire _31050_;
  wire _31051_;
  wire _31052_;
  wire _31053_;
  wire _31054_;
  wire _31055_;
  wire _31056_;
  wire _31057_;
  wire _31058_;
  wire _31059_;
  wire _31060_;
  wire _31061_;
  wire _31062_;
  wire _31063_;
  wire _31064_;
  wire _31065_;
  wire _31066_;
  wire _31067_;
  wire _31068_;
  wire _31069_;
  wire _31070_;
  wire _31071_;
  wire _31072_;
  wire _31073_;
  wire _31074_;
  wire _31075_;
  wire _31076_;
  wire _31077_;
  wire _31078_;
  wire _31079_;
  wire _31080_;
  wire _31081_;
  wire _31082_;
  wire _31083_;
  wire _31084_;
  wire _31085_;
  wire _31086_;
  wire _31087_;
  wire _31088_;
  wire _31089_;
  wire _31090_;
  wire _31091_;
  wire _31092_;
  wire _31093_;
  wire _31094_;
  wire _31095_;
  wire _31096_;
  wire _31097_;
  wire _31098_;
  wire _31099_;
  wire _31100_;
  wire _31101_;
  wire _31102_;
  wire _31103_;
  wire _31104_;
  wire _31105_;
  wire _31106_;
  wire _31107_;
  wire _31108_;
  wire _31109_;
  wire _31110_;
  wire _31111_;
  wire _31112_;
  wire _31113_;
  wire _31114_;
  wire _31115_;
  wire _31116_;
  wire _31117_;
  wire _31118_;
  wire _31119_;
  wire _31120_;
  wire _31121_;
  wire _31122_;
  wire _31123_;
  wire _31124_;
  wire _31125_;
  wire _31126_;
  wire _31127_;
  wire _31128_;
  wire _31129_;
  wire _31130_;
  wire _31131_;
  wire _31132_;
  wire _31133_;
  wire _31134_;
  wire _31135_;
  wire _31136_;
  wire _31137_;
  wire _31138_;
  wire _31139_;
  wire _31140_;
  wire _31141_;
  wire _31142_;
  wire _31143_;
  wire _31144_;
  wire _31145_;
  wire _31146_;
  wire _31147_;
  wire _31148_;
  wire _31149_;
  wire _31150_;
  wire _31151_;
  wire _31152_;
  wire _31153_;
  wire _31154_;
  wire _31155_;
  wire _31156_;
  wire _31157_;
  wire _31158_;
  wire _31159_;
  wire _31160_;
  wire _31161_;
  wire _31162_;
  wire _31163_;
  wire _31164_;
  wire _31165_;
  wire _31166_;
  wire _31167_;
  wire _31168_;
  wire _31169_;
  wire _31170_;
  wire _31171_;
  wire _31172_;
  wire _31173_;
  wire _31174_;
  wire _31175_;
  wire _31176_;
  wire _31177_;
  wire _31178_;
  wire _31179_;
  wire _31180_;
  wire _31181_;
  wire _31182_;
  wire _31183_;
  wire _31184_;
  wire _31185_;
  wire _31186_;
  wire _31187_;
  wire _31188_;
  wire _31189_;
  wire _31190_;
  wire _31191_;
  wire _31192_;
  wire _31193_;
  wire _31194_;
  wire _31195_;
  wire _31196_;
  wire _31197_;
  wire _31198_;
  wire _31199_;
  wire _31200_;
  wire _31201_;
  wire _31202_;
  wire _31203_;
  wire _31204_;
  wire _31205_;
  wire _31206_;
  wire _31207_;
  wire _31208_;
  wire _31209_;
  wire _31210_;
  wire _31211_;
  wire _31212_;
  wire _31213_;
  wire _31214_;
  wire _31215_;
  wire _31216_;
  wire _31217_;
  wire _31218_;
  wire _31219_;
  wire _31220_;
  wire _31221_;
  wire _31222_;
  wire _31223_;
  wire _31224_;
  wire _31225_;
  wire _31226_;
  wire _31227_;
  wire _31228_;
  wire _31229_;
  wire _31230_;
  wire _31231_;
  wire _31232_;
  wire _31233_;
  wire _31234_;
  wire _31235_;
  wire _31236_;
  wire _31237_;
  wire _31238_;
  wire _31239_;
  wire _31240_;
  wire _31241_;
  wire _31242_;
  wire _31243_;
  wire _31244_;
  wire _31245_;
  wire _31246_;
  wire _31247_;
  wire _31248_;
  wire _31249_;
  wire _31250_;
  wire _31251_;
  wire _31252_;
  wire _31253_;
  wire _31254_;
  wire _31255_;
  wire _31256_;
  wire _31257_;
  wire _31258_;
  wire _31259_;
  wire _31260_;
  wire _31261_;
  wire _31262_;
  wire _31263_;
  wire _31264_;
  wire _31265_;
  wire _31266_;
  wire _31267_;
  wire _31268_;
  wire _31269_;
  wire _31270_;
  wire _31271_;
  wire _31272_;
  wire _31273_;
  wire _31274_;
  wire _31275_;
  wire _31276_;
  wire _31277_;
  wire _31278_;
  wire _31279_;
  wire _31280_;
  wire _31281_;
  wire _31282_;
  wire _31283_;
  wire _31284_;
  wire _31285_;
  wire _31286_;
  wire _31287_;
  wire _31288_;
  wire _31289_;
  wire _31290_;
  wire _31291_;
  wire _31292_;
  wire _31293_;
  wire _31294_;
  wire _31295_;
  wire _31296_;
  wire _31297_;
  wire _31298_;
  wire _31299_;
  wire _31300_;
  wire _31301_;
  wire _31302_;
  wire _31303_;
  wire _31304_;
  wire _31305_;
  wire _31306_;
  wire _31307_;
  wire _31308_;
  wire _31309_;
  wire _31310_;
  wire _31311_;
  wire _31312_;
  wire _31313_;
  wire _31314_;
  wire _31315_;
  wire _31316_;
  wire _31317_;
  wire _31318_;
  wire _31319_;
  wire _31320_;
  wire _31321_;
  wire _31322_;
  wire _31323_;
  wire _31324_;
  wire _31325_;
  wire _31326_;
  wire _31327_;
  wire _31328_;
  wire _31329_;
  wire _31330_;
  wire _31331_;
  wire _31332_;
  wire _31333_;
  wire _31334_;
  wire _31335_;
  wire _31336_;
  wire _31337_;
  wire _31338_;
  wire _31339_;
  wire _31340_;
  wire _31341_;
  wire _31342_;
  wire _31343_;
  wire _31344_;
  wire _31345_;
  wire _31346_;
  wire _31347_;
  wire _31348_;
  wire _31349_;
  wire _31350_;
  wire _31351_;
  wire _31352_;
  wire _31353_;
  wire _31354_;
  wire _31355_;
  wire _31356_;
  wire _31357_;
  wire _31358_;
  wire _31359_;
  wire _31360_;
  wire _31361_;
  wire _31362_;
  wire _31363_;
  wire _31364_;
  wire _31365_;
  wire _31366_;
  wire _31367_;
  wire _31368_;
  wire _31369_;
  wire _31370_;
  wire _31371_;
  wire _31372_;
  wire _31373_;
  wire _31374_;
  wire _31375_;
  wire _31376_;
  wire _31377_;
  wire _31378_;
  wire _31379_;
  wire _31380_;
  wire _31381_;
  wire _31382_;
  wire _31383_;
  wire _31384_;
  wire _31385_;
  wire _31386_;
  wire _31387_;
  wire _31388_;
  wire _31389_;
  wire _31390_;
  wire _31391_;
  wire _31392_;
  wire _31393_;
  wire _31394_;
  wire _31395_;
  wire _31396_;
  wire _31397_;
  wire _31398_;
  wire _31399_;
  wire _31400_;
  wire _31401_;
  wire _31402_;
  wire _31403_;
  wire _31404_;
  wire _31405_;
  wire _31406_;
  wire _31407_;
  wire _31408_;
  wire _31409_;
  wire _31410_;
  wire _31411_;
  wire _31412_;
  wire _31413_;
  wire _31414_;
  wire _31415_;
  wire _31416_;
  wire _31417_;
  wire _31418_;
  wire _31419_;
  wire _31420_;
  wire _31421_;
  wire _31422_;
  wire _31423_;
  wire _31424_;
  wire _31425_;
  wire _31426_;
  wire _31427_;
  wire _31428_;
  wire _31429_;
  wire _31430_;
  wire _31431_;
  wire _31432_;
  wire _31433_;
  wire _31434_;
  wire _31435_;
  wire _31436_;
  wire _31437_;
  wire _31438_;
  wire _31439_;
  wire _31440_;
  wire _31441_;
  wire _31442_;
  wire _31443_;
  wire _31444_;
  wire _31445_;
  wire _31446_;
  wire _31447_;
  wire _31448_;
  wire _31449_;
  wire _31450_;
  wire _31451_;
  wire _31452_;
  wire _31453_;
  wire _31454_;
  wire _31455_;
  wire _31456_;
  wire _31457_;
  wire _31458_;
  wire _31459_;
  wire _31460_;
  wire _31461_;
  wire _31462_;
  wire _31463_;
  wire _31464_;
  wire _31465_;
  wire _31466_;
  wire _31467_;
  wire _31468_;
  wire _31469_;
  wire _31470_;
  wire _31471_;
  wire _31472_;
  wire _31473_;
  wire _31474_;
  wire _31475_;
  wire _31476_;
  wire _31477_;
  wire _31478_;
  wire _31479_;
  wire _31480_;
  wire _31481_;
  wire _31482_;
  wire _31483_;
  wire _31484_;
  wire _31485_;
  wire _31486_;
  wire _31487_;
  wire _31488_;
  wire _31489_;
  wire _31490_;
  wire _31491_;
  wire _31492_;
  wire _31493_;
  wire _31494_;
  wire _31495_;
  wire _31496_;
  wire _31497_;
  wire _31498_;
  wire _31499_;
  wire _31500_;
  wire _31501_;
  wire _31502_;
  wire _31503_;
  wire _31504_;
  wire _31505_;
  wire _31506_;
  wire _31507_;
  wire _31508_;
  wire _31509_;
  wire _31510_;
  wire _31511_;
  wire _31512_;
  wire _31513_;
  wire _31514_;
  wire _31515_;
  wire _31516_;
  wire _31517_;
  wire _31518_;
  wire _31519_;
  wire _31520_;
  wire _31521_;
  wire _31522_;
  wire _31523_;
  wire _31524_;
  wire _31525_;
  wire _31526_;
  wire _31527_;
  wire _31528_;
  wire _31529_;
  wire _31530_;
  wire _31531_;
  wire _31532_;
  wire _31533_;
  wire _31534_;
  wire _31535_;
  wire _31536_;
  wire _31537_;
  wire _31538_;
  wire _31539_;
  wire _31540_;
  wire _31541_;
  wire _31542_;
  wire _31543_;
  wire _31544_;
  wire _31545_;
  wire _31546_;
  wire _31547_;
  wire _31548_;
  wire _31549_;
  wire _31550_;
  wire _31551_;
  wire _31552_;
  wire _31553_;
  wire _31554_;
  wire _31555_;
  wire _31556_;
  wire _31557_;
  wire _31558_;
  wire _31559_;
  wire _31560_;
  wire _31561_;
  wire _31562_;
  wire _31563_;
  wire _31564_;
  wire _31565_;
  wire _31566_;
  wire _31567_;
  wire _31568_;
  wire _31569_;
  wire _31570_;
  wire _31571_;
  wire _31572_;
  wire _31573_;
  wire _31574_;
  wire _31575_;
  wire _31576_;
  wire _31577_;
  wire _31578_;
  wire _31579_;
  wire _31580_;
  wire _31581_;
  wire _31582_;
  wire _31583_;
  wire _31584_;
  wire _31585_;
  wire _31586_;
  wire _31587_;
  wire _31588_;
  wire _31589_;
  wire _31590_;
  wire _31591_;
  wire _31592_;
  wire _31593_;
  wire _31594_;
  wire _31595_;
  wire _31596_;
  wire _31597_;
  wire _31598_;
  wire _31599_;
  wire _31600_;
  wire _31601_;
  wire _31602_;
  wire _31603_;
  wire _31604_;
  wire _31605_;
  wire _31606_;
  wire _31607_;
  wire _31608_;
  wire _31609_;
  wire _31610_;
  wire _31611_;
  wire _31612_;
  wire _31613_;
  wire _31614_;
  wire _31615_;
  wire _31616_;
  wire _31617_;
  wire _31618_;
  wire _31619_;
  wire _31620_;
  wire _31621_;
  wire _31622_;
  wire _31623_;
  wire _31624_;
  wire _31625_;
  wire _31626_;
  wire _31627_;
  wire _31628_;
  wire _31629_;
  wire _31630_;
  wire _31631_;
  wire _31632_;
  wire _31633_;
  wire _31634_;
  wire _31635_;
  wire _31636_;
  wire _31637_;
  wire _31638_;
  wire _31639_;
  wire _31640_;
  wire _31641_;
  wire _31642_;
  wire _31643_;
  wire _31644_;
  wire _31645_;
  wire _31646_;
  wire _31647_;
  wire _31648_;
  wire _31649_;
  wire _31650_;
  wire _31651_;
  wire _31652_;
  wire _31653_;
  wire _31654_;
  wire _31655_;
  wire _31656_;
  wire _31657_;
  wire _31658_;
  wire _31659_;
  wire _31660_;
  wire _31661_;
  wire _31662_;
  wire _31663_;
  wire _31664_;
  wire _31665_;
  wire _31666_;
  wire _31667_;
  wire _31668_;
  wire _31669_;
  wire _31670_;
  wire _31671_;
  wire _31672_;
  wire _31673_;
  wire _31674_;
  wire _31675_;
  wire _31676_;
  wire _31677_;
  wire _31678_;
  wire _31679_;
  wire _31680_;
  wire _31681_;
  wire _31682_;
  wire _31683_;
  wire _31684_;
  wire _31685_;
  wire _31686_;
  wire _31687_;
  wire _31688_;
  wire _31689_;
  wire _31690_;
  wire _31691_;
  wire _31692_;
  wire _31693_;
  wire _31694_;
  wire _31695_;
  wire _31696_;
  wire _31697_;
  wire _31698_;
  wire _31699_;
  wire _31700_;
  wire _31701_;
  wire _31702_;
  wire _31703_;
  wire _31704_;
  wire _31705_;
  wire _31706_;
  wire _31707_;
  wire _31708_;
  wire _31709_;
  wire _31710_;
  wire _31711_;
  wire _31712_;
  wire _31713_;
  wire _31714_;
  wire _31715_;
  wire _31716_;
  wire _31717_;
  wire _31718_;
  wire _31719_;
  wire _31720_;
  wire _31721_;
  wire _31722_;
  wire _31723_;
  wire _31724_;
  wire _31725_;
  wire _31726_;
  wire _31727_;
  wire _31728_;
  wire _31729_;
  wire _31730_;
  wire _31731_;
  wire _31732_;
  wire _31733_;
  wire _31734_;
  wire _31735_;
  wire _31736_;
  wire _31737_;
  wire _31738_;
  wire _31739_;
  wire _31740_;
  wire _31741_;
  wire _31742_;
  wire _31743_;
  wire _31744_;
  wire _31745_;
  wire _31746_;
  wire _31747_;
  wire _31748_;
  wire _31749_;
  wire _31750_;
  wire _31751_;
  wire _31752_;
  wire _31753_;
  wire _31754_;
  wire _31755_;
  wire _31756_;
  wire _31757_;
  wire _31758_;
  wire _31759_;
  wire _31760_;
  wire _31761_;
  wire _31762_;
  wire _31763_;
  wire _31764_;
  wire _31765_;
  wire _31766_;
  wire _31767_;
  wire _31768_;
  wire _31769_;
  wire _31770_;
  wire _31771_;
  wire _31772_;
  wire _31773_;
  wire _31774_;
  wire _31775_;
  wire _31776_;
  wire _31777_;
  wire _31778_;
  wire _31779_;
  wire _31780_;
  wire _31781_;
  wire _31782_;
  wire _31783_;
  wire _31784_;
  wire _31785_;
  wire _31786_;
  wire _31787_;
  wire _31788_;
  wire _31789_;
  wire _31790_;
  wire _31791_;
  wire _31792_;
  wire _31793_;
  wire _31794_;
  wire _31795_;
  wire _31796_;
  wire _31797_;
  wire _31798_;
  wire _31799_;
  wire _31800_;
  wire _31801_;
  wire _31802_;
  wire _31803_;
  wire _31804_;
  wire _31805_;
  wire _31806_;
  wire _31807_;
  wire _31808_;
  wire _31809_;
  wire _31810_;
  wire _31811_;
  wire _31812_;
  wire _31813_;
  wire _31814_;
  wire _31815_;
  wire _31816_;
  wire _31817_;
  wire _31818_;
  wire _31819_;
  wire _31820_;
  wire _31821_;
  wire _31822_;
  wire _31823_;
  wire _31824_;
  wire _31825_;
  wire _31826_;
  wire _31827_;
  wire _31828_;
  wire _31829_;
  wire _31830_;
  wire _31831_;
  wire _31832_;
  wire _31833_;
  wire _31834_;
  wire _31835_;
  wire _31836_;
  wire _31837_;
  wire _31838_;
  wire _31839_;
  wire _31840_;
  wire _31841_;
  wire _31842_;
  wire _31843_;
  wire _31844_;
  wire _31845_;
  wire _31846_;
  wire _31847_;
  wire _31848_;
  wire _31849_;
  wire _31850_;
  wire _31851_;
  wire _31852_;
  wire _31853_;
  wire _31854_;
  wire _31855_;
  wire _31856_;
  wire _31857_;
  wire _31858_;
  wire _31859_;
  wire _31860_;
  wire _31861_;
  wire _31862_;
  wire _31863_;
  wire _31864_;
  wire _31865_;
  wire _31866_;
  wire _31867_;
  wire _31868_;
  wire _31869_;
  wire _31870_;
  wire _31871_;
  wire _31872_;
  wire _31873_;
  wire _31874_;
  wire _31875_;
  wire _31876_;
  wire _31877_;
  wire _31878_;
  wire _31879_;
  wire _31880_;
  wire _31881_;
  wire _31882_;
  wire _31883_;
  wire _31884_;
  wire _31885_;
  wire _31886_;
  wire _31887_;
  wire _31888_;
  wire _31889_;
  wire _31890_;
  wire _31891_;
  wire _31892_;
  wire _31893_;
  wire _31894_;
  wire _31895_;
  wire _31896_;
  wire _31897_;
  wire _31898_;
  wire _31899_;
  wire _31900_;
  wire _31901_;
  wire _31902_;
  wire _31903_;
  wire _31904_;
  wire _31905_;
  wire _31906_;
  wire _31907_;
  wire _31908_;
  wire _31909_;
  wire _31910_;
  wire _31911_;
  wire _31912_;
  wire _31913_;
  wire _31914_;
  wire _31915_;
  wire _31916_;
  wire _31917_;
  wire _31918_;
  wire _31919_;
  wire _31920_;
  wire _31921_;
  wire _31922_;
  wire _31923_;
  wire _31924_;
  wire _31925_;
  wire _31926_;
  wire _31927_;
  wire _31928_;
  wire _31929_;
  wire _31930_;
  wire _31931_;
  wire _31932_;
  wire _31933_;
  wire _31934_;
  wire _31935_;
  wire _31936_;
  wire _31937_;
  wire _31938_;
  wire _31939_;
  wire _31940_;
  wire _31941_;
  wire _31942_;
  wire _31943_;
  wire _31944_;
  wire _31945_;
  wire _31946_;
  wire _31947_;
  wire _31948_;
  wire _31949_;
  wire _31950_;
  wire _31951_;
  wire _31952_;
  wire _31953_;
  wire _31954_;
  wire _31955_;
  wire _31956_;
  wire _31957_;
  wire _31958_;
  wire _31959_;
  wire _31960_;
  wire _31961_;
  wire _31962_;
  wire _31963_;
  wire _31964_;
  wire _31965_;
  wire _31966_;
  wire _31967_;
  wire _31968_;
  wire _31969_;
  wire _31970_;
  wire _31971_;
  wire _31972_;
  wire _31973_;
  wire _31974_;
  wire _31975_;
  wire _31976_;
  wire _31977_;
  wire _31978_;
  wire _31979_;
  wire _31980_;
  wire _31981_;
  wire _31982_;
  wire _31983_;
  wire _31984_;
  wire _31985_;
  wire _31986_;
  wire _31987_;
  wire _31988_;
  wire _31989_;
  wire _31990_;
  wire _31991_;
  wire _31992_;
  wire _31993_;
  wire _31994_;
  wire _31995_;
  wire _31996_;
  wire _31997_;
  wire _31998_;
  wire _31999_;
  wire _32000_;
  wire _32001_;
  wire _32002_;
  wire _32003_;
  wire _32004_;
  wire _32005_;
  wire _32006_;
  wire _32007_;
  wire _32008_;
  wire _32009_;
  wire _32010_;
  wire _32011_;
  wire _32012_;
  wire _32013_;
  wire _32014_;
  wire _32015_;
  wire _32016_;
  wire _32017_;
  wire _32018_;
  wire _32019_;
  wire _32020_;
  wire _32021_;
  wire _32022_;
  wire _32023_;
  wire _32024_;
  wire _32025_;
  wire _32026_;
  wire _32027_;
  wire _32028_;
  wire _32029_;
  wire _32030_;
  wire _32031_;
  wire _32032_;
  wire _32033_;
  wire _32034_;
  wire _32035_;
  wire _32036_;
  wire _32037_;
  wire _32038_;
  wire _32039_;
  wire _32040_;
  wire _32041_;
  wire _32042_;
  wire _32043_;
  wire _32044_;
  wire _32045_;
  wire _32046_;
  wire _32047_;
  wire _32048_;
  wire _32049_;
  wire _32050_;
  wire _32051_;
  wire _32052_;
  wire _32053_;
  wire _32054_;
  wire _32055_;
  wire _32056_;
  wire _32057_;
  wire _32058_;
  wire _32059_;
  wire _32060_;
  wire _32061_;
  wire _32062_;
  wire _32063_;
  wire _32064_;
  wire _32065_;
  wire _32066_;
  wire _32067_;
  wire _32068_;
  wire _32069_;
  wire _32070_;
  wire _32071_;
  wire _32072_;
  wire _32073_;
  wire _32074_;
  wire _32075_;
  wire _32076_;
  wire _32077_;
  wire _32078_;
  wire _32079_;
  wire _32080_;
  wire _32081_;
  wire _32082_;
  wire _32083_;
  wire _32084_;
  wire _32085_;
  wire _32086_;
  wire _32087_;
  wire _32088_;
  wire _32089_;
  wire _32090_;
  wire _32091_;
  wire _32092_;
  wire _32093_;
  wire _32094_;
  wire _32095_;
  wire _32096_;
  wire _32097_;
  wire _32098_;
  wire _32099_;
  wire _32100_;
  wire _32101_;
  wire _32102_;
  wire _32103_;
  wire _32104_;
  wire _32105_;
  wire _32106_;
  wire _32107_;
  wire _32108_;
  wire _32109_;
  wire _32110_;
  wire _32111_;
  wire _32112_;
  wire _32113_;
  wire _32114_;
  wire _32115_;
  wire _32116_;
  wire _32117_;
  wire _32118_;
  wire _32119_;
  wire _32120_;
  wire _32121_;
  wire _32122_;
  wire _32123_;
  wire _32124_;
  wire _32125_;
  wire _32126_;
  wire _32127_;
  wire _32128_;
  wire _32129_;
  wire _32130_;
  wire _32131_;
  wire _32132_;
  wire _32133_;
  wire _32134_;
  wire _32135_;
  wire _32136_;
  wire _32137_;
  wire _32138_;
  wire _32139_;
  wire _32140_;
  wire _32141_;
  wire _32142_;
  wire _32143_;
  wire _32144_;
  wire _32145_;
  wire _32146_;
  wire _32147_;
  wire _32148_;
  wire _32149_;
  wire _32150_;
  wire _32151_;
  wire _32152_;
  wire _32153_;
  wire _32154_;
  wire _32155_;
  wire _32156_;
  wire _32157_;
  wire _32158_;
  wire _32159_;
  wire _32160_;
  wire _32161_;
  wire _32162_;
  wire _32163_;
  wire _32164_;
  wire _32165_;
  wire _32166_;
  wire _32167_;
  wire _32168_;
  wire _32169_;
  wire _32170_;
  wire _32171_;
  wire _32172_;
  wire _32173_;
  wire _32174_;
  wire _32175_;
  wire _32176_;
  wire _32177_;
  wire _32178_;
  wire _32179_;
  wire _32180_;
  wire _32181_;
  wire _32182_;
  wire _32183_;
  wire _32184_;
  wire _32185_;
  wire _32186_;
  wire _32187_;
  wire _32188_;
  wire _32189_;
  wire _32190_;
  wire _32191_;
  wire _32192_;
  wire _32193_;
  wire _32194_;
  wire _32195_;
  wire _32196_;
  wire _32197_;
  wire _32198_;
  wire _32199_;
  wire _32200_;
  wire _32201_;
  wire _32202_;
  wire _32203_;
  wire _32204_;
  wire _32205_;
  wire _32206_;
  wire _32207_;
  wire _32208_;
  wire _32209_;
  wire _32210_;
  wire _32211_;
  wire _32212_;
  wire _32213_;
  wire _32214_;
  wire _32215_;
  wire _32216_;
  wire _32217_;
  wire _32218_;
  wire _32219_;
  wire _32220_;
  wire _32221_;
  wire _32222_;
  wire _32223_;
  wire _32224_;
  wire _32225_;
  wire _32226_;
  wire _32227_;
  wire _32228_;
  wire _32229_;
  wire _32230_;
  wire _32231_;
  wire _32232_;
  wire _32233_;
  wire _32234_;
  wire _32235_;
  wire _32236_;
  wire _32237_;
  wire _32238_;
  wire _32239_;
  wire _32240_;
  wire _32241_;
  wire _32242_;
  wire _32243_;
  wire _32244_;
  wire _32245_;
  wire _32246_;
  wire _32247_;
  wire _32248_;
  wire _32249_;
  wire _32250_;
  wire _32251_;
  wire _32252_;
  wire _32253_;
  wire _32254_;
  wire _32255_;
  wire _32256_;
  wire _32257_;
  wire _32258_;
  wire _32259_;
  wire _32260_;
  wire _32261_;
  wire _32262_;
  wire _32263_;
  wire _32264_;
  wire _32265_;
  wire _32266_;
  wire _32267_;
  wire _32268_;
  wire _32269_;
  wire _32270_;
  wire _32271_;
  wire _32272_;
  wire _32273_;
  wire _32274_;
  wire _32275_;
  wire _32276_;
  wire _32277_;
  wire _32278_;
  wire _32279_;
  wire _32280_;
  wire _32281_;
  wire _32282_;
  wire _32283_;
  wire _32284_;
  wire _32285_;
  wire _32286_;
  wire _32287_;
  wire _32288_;
  wire _32289_;
  wire _32290_;
  wire _32291_;
  wire _32292_;
  wire _32293_;
  wire _32294_;
  wire _32295_;
  wire _32296_;
  wire _32297_;
  wire _32298_;
  wire _32299_;
  wire _32300_;
  wire _32301_;
  wire _32302_;
  wire _32303_;
  wire _32304_;
  wire _32305_;
  wire _32306_;
  wire _32307_;
  wire _32308_;
  wire _32309_;
  wire _32310_;
  wire _32311_;
  wire _32312_;
  wire _32313_;
  wire _32314_;
  wire _32315_;
  wire _32316_;
  wire _32317_;
  wire _32318_;
  wire _32319_;
  wire _32320_;
  wire _32321_;
  wire _32322_;
  wire _32323_;
  wire _32324_;
  wire _32325_;
  wire _32326_;
  wire _32327_;
  wire _32328_;
  wire _32329_;
  wire _32330_;
  wire _32331_;
  wire _32332_;
  wire _32333_;
  wire _32334_;
  wire _32335_;
  wire _32336_;
  wire _32337_;
  wire _32338_;
  wire _32339_;
  wire _32340_;
  wire _32341_;
  wire _32342_;
  wire _32343_;
  wire _32344_;
  wire _32345_;
  wire _32346_;
  wire _32347_;
  wire _32348_;
  wire _32349_;
  wire _32350_;
  wire _32351_;
  wire _32352_;
  wire _32353_;
  wire _32354_;
  wire _32355_;
  wire _32356_;
  wire _32357_;
  wire _32358_;
  wire _32359_;
  wire _32360_;
  wire _32361_;
  wire _32362_;
  wire _32363_;
  wire _32364_;
  wire _32365_;
  wire _32366_;
  wire _32367_;
  wire _32368_;
  wire _32369_;
  wire _32370_;
  wire _32371_;
  wire _32372_;
  wire _32373_;
  wire _32374_;
  wire _32375_;
  wire _32376_;
  wire _32377_;
  wire _32378_;
  wire _32379_;
  wire _32380_;
  wire _32381_;
  wire _32382_;
  wire _32383_;
  wire _32384_;
  wire _32385_;
  wire _32386_;
  wire _32387_;
  wire _32388_;
  wire _32389_;
  wire _32390_;
  wire _32391_;
  wire _32392_;
  wire _32393_;
  wire _32394_;
  wire _32395_;
  wire _32396_;
  wire _32397_;
  wire _32398_;
  wire _32399_;
  wire _32400_;
  wire _32401_;
  wire _32402_;
  wire _32403_;
  wire _32404_;
  wire _32405_;
  wire _32406_;
  wire _32407_;
  wire _32408_;
  wire _32409_;
  wire _32410_;
  wire _32411_;
  wire _32412_;
  wire _32413_;
  wire _32414_;
  wire _32415_;
  wire _32416_;
  wire _32417_;
  wire _32418_;
  wire _32419_;
  wire _32420_;
  wire _32421_;
  wire _32422_;
  wire _32423_;
  wire _32424_;
  wire _32425_;
  wire _32426_;
  wire _32427_;
  wire _32428_;
  wire _32429_;
  wire _32430_;
  wire _32431_;
  wire _32432_;
  wire _32433_;
  wire _32434_;
  wire _32435_;
  wire _32436_;
  wire _32437_;
  wire _32438_;
  wire _32439_;
  wire _32440_;
  wire _32441_;
  wire _32442_;
  wire _32443_;
  wire _32444_;
  wire _32445_;
  wire _32446_;
  wire _32447_;
  wire _32448_;
  wire _32449_;
  wire _32450_;
  wire _32451_;
  wire _32452_;
  wire _32453_;
  wire _32454_;
  wire _32455_;
  wire _32456_;
  wire _32457_;
  wire _32458_;
  wire _32459_;
  wire _32460_;
  wire _32461_;
  wire _32462_;
  wire _32463_;
  wire _32464_;
  wire _32465_;
  wire _32466_;
  wire _32467_;
  wire _32468_;
  wire _32469_;
  wire _32470_;
  wire _32471_;
  wire _32472_;
  wire _32473_;
  wire _32474_;
  wire _32475_;
  wire _32476_;
  wire _32477_;
  wire _32478_;
  wire _32479_;
  wire _32480_;
  wire _32481_;
  wire _32482_;
  wire _32483_;
  wire _32484_;
  wire _32485_;
  wire _32486_;
  wire _32487_;
  wire _32488_;
  wire _32489_;
  wire _32490_;
  wire _32491_;
  wire _32492_;
  wire _32493_;
  wire _32494_;
  wire _32495_;
  wire _32496_;
  wire _32497_;
  wire _32498_;
  wire _32499_;
  wire _32500_;
  wire _32501_;
  wire _32502_;
  wire _32503_;
  wire _32504_;
  wire _32505_;
  wire _32506_;
  wire _32507_;
  wire _32508_;
  wire _32509_;
  wire _32510_;
  wire _32511_;
  wire _32512_;
  wire _32513_;
  wire _32514_;
  wire _32515_;
  wire _32516_;
  wire _32517_;
  wire _32518_;
  wire _32519_;
  wire _32520_;
  wire _32521_;
  wire _32522_;
  wire _32523_;
  wire _32524_;
  wire _32525_;
  wire _32526_;
  wire _32527_;
  wire _32528_;
  wire _32529_;
  wire _32530_;
  wire _32531_;
  wire _32532_;
  wire _32533_;
  wire _32534_;
  wire _32535_;
  wire _32536_;
  wire _32537_;
  wire _32538_;
  wire _32539_;
  wire _32540_;
  wire _32541_;
  wire _32542_;
  wire _32543_;
  wire _32544_;
  wire _32545_;
  wire _32546_;
  wire _32547_;
  wire _32548_;
  wire _32549_;
  wire _32550_;
  wire _32551_;
  wire _32552_;
  wire _32553_;
  wire _32554_;
  wire _32555_;
  wire _32556_;
  wire _32557_;
  wire _32558_;
  wire _32559_;
  wire _32560_;
  wire _32561_;
  wire _32562_;
  wire _32563_;
  wire _32564_;
  wire _32565_;
  wire _32566_;
  wire _32567_;
  wire _32568_;
  wire _32569_;
  wire _32570_;
  wire _32571_;
  wire _32572_;
  wire _32573_;
  wire _32574_;
  wire _32575_;
  wire _32576_;
  wire _32577_;
  wire _32578_;
  wire _32579_;
  wire _32580_;
  wire _32581_;
  wire _32582_;
  wire _32583_;
  wire _32584_;
  wire _32585_;
  wire _32586_;
  wire _32587_;
  wire _32588_;
  wire _32589_;
  wire _32590_;
  wire _32591_;
  wire _32592_;
  wire _32593_;
  wire _32594_;
  wire _32595_;
  wire _32596_;
  wire _32597_;
  wire _32598_;
  wire _32599_;
  wire _32600_;
  wire _32601_;
  wire _32602_;
  wire _32603_;
  wire _32604_;
  wire _32605_;
  wire _32606_;
  wire _32607_;
  wire _32608_;
  wire _32609_;
  wire _32610_;
  wire _32611_;
  wire _32612_;
  wire _32613_;
  wire _32614_;
  wire _32615_;
  wire _32616_;
  wire _32617_;
  wire _32618_;
  wire _32619_;
  wire _32620_;
  wire _32621_;
  wire _32622_;
  wire _32623_;
  wire _32624_;
  wire _32625_;
  wire _32626_;
  wire _32627_;
  wire _32628_;
  wire _32629_;
  wire _32630_;
  wire _32631_;
  wire _32632_;
  wire _32633_;
  wire _32634_;
  wire _32635_;
  wire _32636_;
  wire _32637_;
  wire _32638_;
  wire _32639_;
  wire _32640_;
  wire _32641_;
  wire _32642_;
  wire _32643_;
  wire _32644_;
  wire _32645_;
  wire _32646_;
  wire _32647_;
  wire _32648_;
  wire _32649_;
  wire _32650_;
  wire _32651_;
  wire _32652_;
  wire _32653_;
  wire _32654_;
  wire _32655_;
  wire _32656_;
  wire _32657_;
  wire _32658_;
  wire _32659_;
  wire _32660_;
  wire _32661_;
  wire _32662_;
  wire _32663_;
  wire _32664_;
  wire _32665_;
  wire _32666_;
  wire _32667_;
  wire _32668_;
  wire _32669_;
  wire _32670_;
  wire _32671_;
  wire _32672_;
  wire _32673_;
  wire _32674_;
  wire _32675_;
  wire _32676_;
  wire _32677_;
  wire _32678_;
  wire _32679_;
  wire _32680_;
  wire _32681_;
  wire _32682_;
  wire _32683_;
  wire _32684_;
  wire _32685_;
  wire _32686_;
  wire _32687_;
  wire _32688_;
  wire _32689_;
  wire _32690_;
  wire _32691_;
  wire _32692_;
  wire _32693_;
  wire _32694_;
  wire _32695_;
  wire _32696_;
  wire _32697_;
  wire _32698_;
  wire _32699_;
  wire _32700_;
  wire _32701_;
  wire _32702_;
  wire _32703_;
  wire _32704_;
  wire _32705_;
  wire _32706_;
  wire _32707_;
  wire _32708_;
  wire _32709_;
  wire _32710_;
  wire _32711_;
  wire _32712_;
  wire _32713_;
  wire _32714_;
  wire _32715_;
  wire _32716_;
  wire _32717_;
  wire _32718_;
  wire _32719_;
  wire _32720_;
  wire _32721_;
  wire _32722_;
  wire _32723_;
  wire _32724_;
  wire _32725_;
  wire _32726_;
  wire _32727_;
  wire _32728_;
  wire _32729_;
  wire _32730_;
  wire _32731_;
  wire _32732_;
  wire _32733_;
  wire _32734_;
  wire _32735_;
  wire _32736_;
  wire _32737_;
  wire _32738_;
  wire _32739_;
  wire _32740_;
  wire _32741_;
  wire _32742_;
  wire _32743_;
  wire _32744_;
  wire _32745_;
  wire _32746_;
  wire _32747_;
  wire _32748_;
  wire _32749_;
  wire _32750_;
  wire _32751_;
  wire _32752_;
  wire _32753_;
  wire _32754_;
  wire _32755_;
  wire _32756_;
  wire _32757_;
  wire _32758_;
  wire _32759_;
  wire _32760_;
  wire _32761_;
  wire _32762_;
  wire _32763_;
  wire _32764_;
  wire _32765_;
  wire _32766_;
  wire _32767_;
  wire _32768_;
  wire _32769_;
  wire _32770_;
  wire _32771_;
  wire _32772_;
  wire _32773_;
  wire _32774_;
  wire _32775_;
  wire _32776_;
  wire _32777_;
  wire _32778_;
  wire _32779_;
  wire _32780_;
  wire _32781_;
  wire _32782_;
  wire _32783_;
  wire _32784_;
  wire _32785_;
  wire _32786_;
  wire _32787_;
  wire _32788_;
  wire _32789_;
  wire _32790_;
  wire _32791_;
  wire _32792_;
  wire _32793_;
  wire _32794_;
  wire _32795_;
  wire _32796_;
  wire _32797_;
  wire _32798_;
  wire _32799_;
  wire _32800_;
  wire _32801_;
  wire _32802_;
  wire _32803_;
  wire _32804_;
  wire _32805_;
  wire _32806_;
  wire _32807_;
  wire _32808_;
  wire _32809_;
  wire _32810_;
  wire _32811_;
  wire _32812_;
  wire _32813_;
  wire _32814_;
  wire _32815_;
  wire _32816_;
  wire _32817_;
  wire _32818_;
  wire _32819_;
  wire _32820_;
  wire _32821_;
  wire _32822_;
  wire _32823_;
  wire _32824_;
  wire _32825_;
  wire _32826_;
  wire _32827_;
  wire _32828_;
  wire _32829_;
  wire _32830_;
  wire _32831_;
  wire _32832_;
  wire _32833_;
  wire _32834_;
  wire _32835_;
  wire _32836_;
  wire _32837_;
  wire _32838_;
  wire _32839_;
  wire _32840_;
  wire _32841_;
  wire _32842_;
  wire _32843_;
  wire _32844_;
  wire _32845_;
  wire _32846_;
  wire _32847_;
  wire _32848_;
  wire _32849_;
  wire _32850_;
  wire _32851_;
  wire _32852_;
  wire _32853_;
  wire _32854_;
  wire _32855_;
  wire _32856_;
  wire _32857_;
  wire _32858_;
  wire _32859_;
  wire _32860_;
  wire _32861_;
  wire _32862_;
  wire _32863_;
  wire _32864_;
  wire _32865_;
  wire _32866_;
  wire _32867_;
  wire _32868_;
  wire _32869_;
  wire _32870_;
  wire _32871_;
  wire _32872_;
  wire _32873_;
  wire _32874_;
  wire _32875_;
  wire _32876_;
  wire _32877_;
  wire _32878_;
  wire _32879_;
  wire _32880_;
  wire _32881_;
  wire _32882_;
  wire _32883_;
  wire _32884_;
  wire _32885_;
  wire _32886_;
  wire _32887_;
  wire _32888_;
  wire _32889_;
  wire _32890_;
  wire _32891_;
  wire _32892_;
  wire _32893_;
  wire _32894_;
  wire _32895_;
  wire _32896_;
  wire _32897_;
  wire _32898_;
  wire _32899_;
  wire _32900_;
  wire _32901_;
  wire _32902_;
  wire _32903_;
  wire _32904_;
  wire _32905_;
  wire _32906_;
  wire _32907_;
  wire _32908_;
  wire _32909_;
  wire _32910_;
  wire _32911_;
  wire _32912_;
  wire _32913_;
  wire _32914_;
  wire _32915_;
  wire _32916_;
  wire _32917_;
  wire _32918_;
  wire _32919_;
  wire _32920_;
  wire _32921_;
  wire _32922_;
  wire _32923_;
  wire _32924_;
  wire _32925_;
  wire _32926_;
  wire _32927_;
  wire _32928_;
  wire _32929_;
  wire _32930_;
  wire _32931_;
  wire _32932_;
  wire _32933_;
  wire _32934_;
  wire _32935_;
  wire _32936_;
  wire _32937_;
  wire _32938_;
  wire _32939_;
  wire _32940_;
  wire _32941_;
  wire _32942_;
  wire _32943_;
  wire _32944_;
  wire _32945_;
  wire _32946_;
  wire _32947_;
  wire _32948_;
  wire _32949_;
  wire _32950_;
  wire _32951_;
  wire _32952_;
  wire _32953_;
  wire _32954_;
  wire _32955_;
  wire _32956_;
  wire _32957_;
  wire _32958_;
  wire _32959_;
  wire _32960_;
  wire _32961_;
  wire _32962_;
  wire _32963_;
  wire _32964_;
  wire _32965_;
  wire _32966_;
  wire _32967_;
  wire _32968_;
  wire _32969_;
  wire _32970_;
  wire _32971_;
  wire _32972_;
  wire _32973_;
  wire _32974_;
  wire _32975_;
  wire _32976_;
  wire _32977_;
  wire _32978_;
  wire _32979_;
  wire _32980_;
  wire _32981_;
  wire _32982_;
  wire _32983_;
  wire _32984_;
  wire _32985_;
  wire _32986_;
  wire _32987_;
  wire _32988_;
  wire _32989_;
  wire _32990_;
  wire _32991_;
  wire _32992_;
  wire _32993_;
  wire _32994_;
  wire _32995_;
  wire _32996_;
  wire _32997_;
  wire _32998_;
  wire _32999_;
  wire _33000_;
  wire _33001_;
  wire _33002_;
  wire _33003_;
  wire _33004_;
  wire _33005_;
  wire _33006_;
  wire _33007_;
  wire _33008_;
  wire _33009_;
  wire _33010_;
  wire _33011_;
  wire _33012_;
  wire _33013_;
  wire _33014_;
  wire _33015_;
  wire _33016_;
  wire _33017_;
  wire _33018_;
  wire _33019_;
  wire _33020_;
  wire _33021_;
  wire _33022_;
  wire _33023_;
  wire _33024_;
  wire _33025_;
  wire _33026_;
  wire _33027_;
  wire _33028_;
  wire _33029_;
  wire _33030_;
  wire _33031_;
  wire _33032_;
  wire _33033_;
  wire _33034_;
  wire _33035_;
  wire _33036_;
  wire _33037_;
  wire _33038_;
  wire _33039_;
  wire _33040_;
  wire _33041_;
  wire _33042_;
  wire _33043_;
  wire _33044_;
  wire _33045_;
  wire _33046_;
  wire _33047_;
  wire _33048_;
  wire _33049_;
  wire _33050_;
  wire _33051_;
  wire _33052_;
  wire _33053_;
  wire _33054_;
  wire _33055_;
  wire _33056_;
  wire _33057_;
  wire _33058_;
  wire _33059_;
  wire _33060_;
  wire _33061_;
  wire _33062_;
  wire _33063_;
  wire _33064_;
  wire _33065_;
  wire _33066_;
  wire _33067_;
  wire _33068_;
  wire _33069_;
  wire _33070_;
  wire _33071_;
  wire _33072_;
  wire _33073_;
  wire _33074_;
  wire _33075_;
  wire _33076_;
  wire _33077_;
  wire _33078_;
  wire _33079_;
  wire _33080_;
  wire _33081_;
  wire _33082_;
  wire _33083_;
  wire _33084_;
  wire _33085_;
  wire _33086_;
  wire _33087_;
  wire _33088_;
  wire _33089_;
  wire _33090_;
  wire _33091_;
  wire _33092_;
  wire _33093_;
  wire _33094_;
  wire _33095_;
  wire _33096_;
  wire _33097_;
  wire _33098_;
  wire _33099_;
  wire _33100_;
  wire _33101_;
  wire _33102_;
  wire _33103_;
  wire _33104_;
  wire _33105_;
  wire _33106_;
  wire _33107_;
  wire _33108_;
  wire _33109_;
  wire _33110_;
  wire _33111_;
  wire _33112_;
  wire _33113_;
  wire _33114_;
  wire _33115_;
  wire _33116_;
  wire _33117_;
  wire _33118_;
  wire _33119_;
  wire _33120_;
  wire _33121_;
  wire _33122_;
  wire _33123_;
  wire _33124_;
  wire _33125_;
  wire _33126_;
  wire _33127_;
  wire _33128_;
  wire _33129_;
  wire _33130_;
  wire _33131_;
  wire _33132_;
  wire _33133_;
  wire _33134_;
  wire _33135_;
  wire _33136_;
  wire _33137_;
  wire _33138_;
  wire _33139_;
  wire _33140_;
  wire _33141_;
  wire _33142_;
  wire _33143_;
  wire _33144_;
  wire _33145_;
  wire _33146_;
  wire _33147_;
  wire _33148_;
  wire _33149_;
  wire _33150_;
  wire _33151_;
  wire _33152_;
  wire _33153_;
  wire _33154_;
  wire _33155_;
  wire _33156_;
  wire _33157_;
  wire _33158_;
  wire _33159_;
  wire _33160_;
  wire _33161_;
  wire _33162_;
  wire _33163_;
  wire _33164_;
  wire _33165_;
  wire _33166_;
  wire _33167_;
  wire _33168_;
  wire _33169_;
  wire _33170_;
  wire _33171_;
  wire _33172_;
  wire _33173_;
  wire _33174_;
  wire _33175_;
  wire _33176_;
  wire _33177_;
  wire _33178_;
  wire _33179_;
  wire _33180_;
  wire _33181_;
  wire _33182_;
  wire _33183_;
  wire _33184_;
  wire _33185_;
  wire _33186_;
  wire _33187_;
  wire _33188_;
  wire _33189_;
  wire _33190_;
  wire _33191_;
  wire _33192_;
  wire _33193_;
  wire _33194_;
  wire _33195_;
  wire _33196_;
  wire _33197_;
  wire _33198_;
  wire _33199_;
  wire _33200_;
  wire _33201_;
  wire _33202_;
  wire _33203_;
  wire _33204_;
  wire _33205_;
  wire _33206_;
  wire _33207_;
  wire _33208_;
  wire _33209_;
  wire _33210_;
  wire _33211_;
  wire _33212_;
  wire _33213_;
  wire _33214_;
  wire _33215_;
  wire _33216_;
  wire _33217_;
  wire _33218_;
  wire _33219_;
  wire _33220_;
  wire _33221_;
  wire _33222_;
  wire _33223_;
  wire _33224_;
  wire _33225_;
  wire _33226_;
  wire _33227_;
  wire _33228_;
  wire _33229_;
  wire _33230_;
  wire _33231_;
  wire _33232_;
  wire _33233_;
  wire _33234_;
  wire _33235_;
  wire _33236_;
  wire _33237_;
  wire _33238_;
  wire _33239_;
  wire _33240_;
  wire _33241_;
  wire _33242_;
  wire _33243_;
  wire _33244_;
  wire _33245_;
  wire _33246_;
  wire _33247_;
  wire _33248_;
  wire _33249_;
  wire _33250_;
  wire _33251_;
  wire _33252_;
  wire _33253_;
  wire _33254_;
  wire _33255_;
  wire _33256_;
  wire _33257_;
  wire _33258_;
  wire _33259_;
  wire _33260_;
  wire _33261_;
  wire _33262_;
  wire _33263_;
  wire _33264_;
  wire _33265_;
  wire _33266_;
  wire _33267_;
  wire _33268_;
  wire _33269_;
  wire _33270_;
  wire _33271_;
  wire _33272_;
  wire _33273_;
  wire _33274_;
  wire _33275_;
  wire _33276_;
  wire _33277_;
  wire _33278_;
  wire _33279_;
  wire _33280_;
  wire _33281_;
  wire _33282_;
  wire _33283_;
  wire _33284_;
  wire _33285_;
  wire _33286_;
  wire _33287_;
  wire _33288_;
  wire _33289_;
  wire _33290_;
  wire _33291_;
  wire _33292_;
  wire _33293_;
  wire _33294_;
  wire _33295_;
  wire _33296_;
  wire _33297_;
  wire _33298_;
  wire _33299_;
  wire _33300_;
  wire _33301_;
  wire _33302_;
  wire _33303_;
  wire _33304_;
  wire _33305_;
  wire _33306_;
  wire _33307_;
  wire _33308_;
  wire _33309_;
  wire _33310_;
  wire _33311_;
  wire _33312_;
  wire _33313_;
  wire _33314_;
  wire _33315_;
  wire _33316_;
  wire _33317_;
  wire _33318_;
  wire _33319_;
  wire _33320_;
  wire _33321_;
  wire _33322_;
  wire _33323_;
  wire _33324_;
  wire _33325_;
  wire _33326_;
  wire _33327_;
  wire _33328_;
  wire _33329_;
  wire _33330_;
  wire _33331_;
  wire _33332_;
  wire _33333_;
  wire _33334_;
  wire _33335_;
  wire _33336_;
  wire _33337_;
  wire _33338_;
  wire _33339_;
  wire _33340_;
  wire _33341_;
  wire _33342_;
  wire _33343_;
  wire _33344_;
  wire _33345_;
  wire _33346_;
  wire _33347_;
  wire _33348_;
  wire _33349_;
  wire _33350_;
  wire _33351_;
  wire _33352_;
  wire _33353_;
  wire _33354_;
  wire _33355_;
  wire _33356_;
  wire _33357_;
  wire _33358_;
  wire _33359_;
  wire _33360_;
  wire _33361_;
  wire _33362_;
  wire _33363_;
  wire _33364_;
  wire _33365_;
  wire _33366_;
  wire _33367_;
  wire _33368_;
  wire _33369_;
  wire _33370_;
  wire _33371_;
  wire _33372_;
  wire _33373_;
  wire _33374_;
  wire _33375_;
  wire _33376_;
  wire _33377_;
  wire _33378_;
  wire _33379_;
  wire _33380_;
  wire _33381_;
  wire _33382_;
  wire _33383_;
  wire _33384_;
  wire _33385_;
  wire _33386_;
  wire _33387_;
  wire _33388_;
  wire _33389_;
  wire _33390_;
  wire _33391_;
  wire _33392_;
  wire _33393_;
  wire _33394_;
  wire _33395_;
  wire _33396_;
  wire _33397_;
  wire _33398_;
  wire _33399_;
  wire _33400_;
  wire _33401_;
  wire _33402_;
  wire _33403_;
  wire _33404_;
  wire _33405_;
  wire _33406_;
  wire _33407_;
  wire _33408_;
  wire _33409_;
  wire _33410_;
  wire _33411_;
  wire _33412_;
  wire _33413_;
  wire _33414_;
  wire _33415_;
  wire _33416_;
  wire _33417_;
  wire _33418_;
  wire _33419_;
  wire _33420_;
  wire _33421_;
  wire _33422_;
  wire _33423_;
  wire _33424_;
  wire _33425_;
  wire _33426_;
  wire _33427_;
  wire _33428_;
  wire _33429_;
  wire _33430_;
  wire _33431_;
  wire _33432_;
  wire _33433_;
  wire _33434_;
  wire _33435_;
  wire _33436_;
  wire _33437_;
  wire _33438_;
  wire _33439_;
  wire _33440_;
  wire _33441_;
  wire _33442_;
  wire _33443_;
  wire _33444_;
  wire _33445_;
  wire _33446_;
  wire _33447_;
  wire _33448_;
  wire _33449_;
  wire _33450_;
  wire _33451_;
  wire _33452_;
  wire _33453_;
  wire _33454_;
  wire _33455_;
  wire _33456_;
  wire _33457_;
  wire _33458_;
  wire _33459_;
  wire _33460_;
  wire _33461_;
  wire _33462_;
  wire _33463_;
  wire _33464_;
  wire _33465_;
  wire _33466_;
  wire _33467_;
  wire _33468_;
  wire _33469_;
  wire _33470_;
  wire _33471_;
  wire _33472_;
  wire _33473_;
  wire _33474_;
  wire _33475_;
  wire _33476_;
  wire _33477_;
  wire _33478_;
  wire _33479_;
  wire _33480_;
  wire _33481_;
  wire _33482_;
  wire _33483_;
  wire _33484_;
  wire _33485_;
  wire _33486_;
  wire _33487_;
  wire _33488_;
  wire _33489_;
  wire _33490_;
  wire _33491_;
  wire _33492_;
  wire _33493_;
  wire _33494_;
  wire _33495_;
  wire _33496_;
  wire _33497_;
  wire _33498_;
  wire _33499_;
  wire _33500_;
  wire _33501_;
  wire _33502_;
  wire _33503_;
  wire _33504_;
  wire _33505_;
  wire _33506_;
  wire _33507_;
  wire _33508_;
  wire _33509_;
  wire _33510_;
  wire _33511_;
  wire _33512_;
  wire _33513_;
  wire _33514_;
  wire _33515_;
  wire _33516_;
  wire _33517_;
  wire _33518_;
  wire _33519_;
  wire _33520_;
  wire _33521_;
  wire _33522_;
  wire _33523_;
  wire _33524_;
  wire _33525_;
  wire _33526_;
  wire _33527_;
  wire _33528_;
  wire _33529_;
  wire _33530_;
  wire _33531_;
  wire _33532_;
  wire _33533_;
  wire _33534_;
  wire _33535_;
  wire _33536_;
  wire _33537_;
  wire _33538_;
  wire _33539_;
  wire _33540_;
  wire _33541_;
  wire _33542_;
  wire _33543_;
  wire _33544_;
  wire _33545_;
  wire _33546_;
  wire _33547_;
  wire _33548_;
  wire _33549_;
  wire _33550_;
  wire _33551_;
  wire _33552_;
  wire _33553_;
  wire _33554_;
  wire _33555_;
  wire _33556_;
  wire _33557_;
  wire _33558_;
  wire _33559_;
  wire _33560_;
  wire _33561_;
  wire _33562_;
  wire _33563_;
  wire _33564_;
  wire _33565_;
  wire _33566_;
  wire _33567_;
  wire _33568_;
  wire _33569_;
  wire _33570_;
  wire _33571_;
  wire _33572_;
  wire _33573_;
  wire _33574_;
  wire _33575_;
  wire _33576_;
  wire _33577_;
  wire _33578_;
  wire _33579_;
  wire _33580_;
  wire _33581_;
  wire _33582_;
  wire _33583_;
  wire _33584_;
  wire _33585_;
  wire _33586_;
  wire _33587_;
  wire _33588_;
  wire _33589_;
  wire _33590_;
  wire _33591_;
  wire _33592_;
  wire _33593_;
  wire _33594_;
  wire _33595_;
  wire _33596_;
  wire _33597_;
  wire _33598_;
  wire _33599_;
  wire _33600_;
  wire _33601_;
  wire _33602_;
  wire _33603_;
  wire _33604_;
  wire _33605_;
  wire _33606_;
  wire _33607_;
  wire _33608_;
  wire _33609_;
  wire _33610_;
  wire _33611_;
  wire _33612_;
  wire _33613_;
  wire _33614_;
  wire _33615_;
  wire _33616_;
  wire _33617_;
  wire _33618_;
  wire _33619_;
  wire _33620_;
  wire _33621_;
  wire _33622_;
  wire _33623_;
  wire _33624_;
  wire _33625_;
  wire _33626_;
  wire _33627_;
  wire _33628_;
  wire _33629_;
  wire _33630_;
  wire _33631_;
  wire _33632_;
  wire _33633_;
  wire _33634_;
  wire _33635_;
  wire _33636_;
  wire _33637_;
  wire _33638_;
  wire _33639_;
  wire _33640_;
  wire _33641_;
  wire _33642_;
  wire _33643_;
  wire _33644_;
  wire _33645_;
  wire _33646_;
  wire _33647_;
  wire _33648_;
  wire _33649_;
  wire _33650_;
  wire _33651_;
  wire _33652_;
  wire _33653_;
  wire _33654_;
  wire _33655_;
  wire _33656_;
  wire _33657_;
  wire _33658_;
  wire _33659_;
  wire _33660_;
  wire _33661_;
  wire _33662_;
  wire _33663_;
  wire _33664_;
  wire _33665_;
  wire _33666_;
  wire _33667_;
  wire _33668_;
  wire _33669_;
  wire _33670_;
  wire _33671_;
  wire _33672_;
  wire _33673_;
  wire _33674_;
  wire _33675_;
  wire _33676_;
  wire _33677_;
  wire _33678_;
  wire _33679_;
  wire _33680_;
  wire _33681_;
  wire _33682_;
  wire _33683_;
  wire _33684_;
  wire _33685_;
  wire _33686_;
  wire _33687_;
  wire _33688_;
  wire _33689_;
  wire _33690_;
  wire _33691_;
  wire _33692_;
  wire _33693_;
  wire _33694_;
  wire _33695_;
  wire _33696_;
  wire _33697_;
  wire _33698_;
  wire _33699_;
  wire _33700_;
  wire _33701_;
  wire _33702_;
  wire _33703_;
  wire _33704_;
  wire _33705_;
  wire _33706_;
  wire _33707_;
  wire _33708_;
  wire _33709_;
  wire _33710_;
  wire _33711_;
  wire _33712_;
  wire _33713_;
  wire _33714_;
  wire _33715_;
  wire _33716_;
  wire _33717_;
  wire _33718_;
  wire _33719_;
  wire _33720_;
  wire _33721_;
  wire _33722_;
  wire _33723_;
  wire _33724_;
  wire _33725_;
  wire _33726_;
  wire _33727_;
  wire _33728_;
  wire _33729_;
  wire _33730_;
  wire _33731_;
  wire _33732_;
  wire _33733_;
  wire _33734_;
  wire _33735_;
  wire _33736_;
  wire _33737_;
  wire _33738_;
  wire _33739_;
  wire _33740_;
  wire _33741_;
  wire _33742_;
  wire _33743_;
  wire _33744_;
  wire _33745_;
  wire _33746_;
  wire _33747_;
  wire _33748_;
  wire _33749_;
  wire _33750_;
  wire _33751_;
  wire _33752_;
  wire _33753_;
  wire _33754_;
  wire _33755_;
  wire _33756_;
  wire _33757_;
  wire _33758_;
  wire _33759_;
  wire _33760_;
  wire _33761_;
  wire _33762_;
  wire _33763_;
  wire _33764_;
  wire _33765_;
  wire _33766_;
  wire _33767_;
  wire _33768_;
  wire _33769_;
  wire _33770_;
  wire _33771_;
  wire _33772_;
  wire _33773_;
  wire _33774_;
  wire _33775_;
  wire _33776_;
  wire _33777_;
  wire _33778_;
  wire _33779_;
  wire _33780_;
  wire _33781_;
  wire _33782_;
  wire _33783_;
  wire _33784_;
  wire _33785_;
  wire _33786_;
  wire _33787_;
  wire _33788_;
  wire _33789_;
  wire _33790_;
  wire _33791_;
  wire _33792_;
  wire _33793_;
  wire _33794_;
  wire _33795_;
  wire _33796_;
  wire _33797_;
  wire _33798_;
  wire _33799_;
  wire _33800_;
  wire _33801_;
  wire _33802_;
  wire _33803_;
  wire _33804_;
  wire _33805_;
  wire _33806_;
  wire _33807_;
  wire _33808_;
  wire _33809_;
  wire _33810_;
  wire _33811_;
  wire _33812_;
  wire _33813_;
  wire _33814_;
  wire _33815_;
  wire _33816_;
  wire _33817_;
  wire _33818_;
  wire _33819_;
  wire _33820_;
  wire _33821_;
  wire _33822_;
  wire _33823_;
  wire _33824_;
  wire _33825_;
  wire _33826_;
  wire _33827_;
  wire _33828_;
  wire _33829_;
  wire _33830_;
  wire _33831_;
  wire _33832_;
  wire _33833_;
  wire _33834_;
  wire _33835_;
  wire _33836_;
  wire _33837_;
  wire _33838_;
  wire _33839_;
  wire _33840_;
  wire _33841_;
  wire _33842_;
  wire _33843_;
  wire _33844_;
  wire _33845_;
  wire _33846_;
  wire _33847_;
  wire _33848_;
  wire _33849_;
  wire _33850_;
  wire _33851_;
  wire _33852_;
  wire _33853_;
  wire _33854_;
  wire _33855_;
  wire _33856_;
  wire _33857_;
  wire _33858_;
  wire _33859_;
  wire _33860_;
  wire _33861_;
  wire _33862_;
  wire _33863_;
  wire _33864_;
  wire _33865_;
  wire _33866_;
  wire _33867_;
  wire _33868_;
  wire _33869_;
  wire _33870_;
  wire _33871_;
  wire _33872_;
  wire _33873_;
  wire _33874_;
  wire _33875_;
  wire _33876_;
  wire _33877_;
  wire _33878_;
  wire _33879_;
  wire _33880_;
  wire _33881_;
  wire _33882_;
  wire _33883_;
  wire _33884_;
  wire _33885_;
  wire _33886_;
  wire _33887_;
  wire _33888_;
  wire _33889_;
  wire _33890_;
  wire _33891_;
  wire _33892_;
  wire _33893_;
  wire _33894_;
  wire _33895_;
  wire _33896_;
  wire _33897_;
  wire _33898_;
  wire _33899_;
  wire _33900_;
  wire _33901_;
  wire _33902_;
  wire _33903_;
  wire _33904_;
  wire _33905_;
  wire _33906_;
  wire _33907_;
  wire _33908_;
  wire _33909_;
  wire _33910_;
  wire _33911_;
  wire _33912_;
  wire _33913_;
  wire _33914_;
  wire _33915_;
  wire _33916_;
  wire _33917_;
  wire _33918_;
  wire _33919_;
  wire _33920_;
  wire _33921_;
  wire _33922_;
  wire _33923_;
  wire _33924_;
  wire _33925_;
  wire _33926_;
  wire _33927_;
  wire _33928_;
  wire _33929_;
  wire _33930_;
  wire _33931_;
  wire _33932_;
  wire _33933_;
  wire _33934_;
  wire _33935_;
  wire _33936_;
  wire _33937_;
  wire _33938_;
  wire _33939_;
  wire _33940_;
  wire _33941_;
  wire _33942_;
  wire _33943_;
  wire _33944_;
  wire _33945_;
  wire _33946_;
  wire _33947_;
  wire _33948_;
  wire _33949_;
  wire _33950_;
  wire _33951_;
  wire _33952_;
  wire _33953_;
  wire _33954_;
  wire _33955_;
  wire _33956_;
  wire _33957_;
  wire _33958_;
  wire _33959_;
  wire _33960_;
  wire _33961_;
  wire _33962_;
  wire _33963_;
  wire _33964_;
  wire _33965_;
  wire _33966_;
  wire _33967_;
  wire _33968_;
  wire _33969_;
  wire _33970_;
  wire _33971_;
  wire _33972_;
  wire _33973_;
  wire _33974_;
  wire _33975_;
  wire _33976_;
  wire _33977_;
  wire _33978_;
  wire _33979_;
  wire _33980_;
  wire _33981_;
  wire _33982_;
  wire _33983_;
  wire _33984_;
  wire _33985_;
  wire _33986_;
  wire _33987_;
  wire _33988_;
  wire _33989_;
  wire _33990_;
  wire _33991_;
  wire _33992_;
  wire _33993_;
  wire _33994_;
  wire _33995_;
  wire _33996_;
  wire _33997_;
  wire _33998_;
  wire _33999_;
  wire _34000_;
  wire _34001_;
  wire _34002_;
  wire _34003_;
  wire _34004_;
  wire _34005_;
  wire _34006_;
  wire _34007_;
  wire _34008_;
  wire _34009_;
  wire _34010_;
  wire _34011_;
  wire _34012_;
  wire _34013_;
  wire _34014_;
  wire _34015_;
  wire _34016_;
  wire _34017_;
  wire _34018_;
  wire _34019_;
  wire _34020_;
  wire _34021_;
  wire _34022_;
  wire _34023_;
  wire _34024_;
  wire _34025_;
  wire _34026_;
  wire _34027_;
  wire _34028_;
  wire _34029_;
  wire _34030_;
  wire _34031_;
  wire _34032_;
  wire _34033_;
  wire _34034_;
  wire _34035_;
  wire _34036_;
  wire _34037_;
  wire _34038_;
  wire _34039_;
  wire _34040_;
  wire _34041_;
  wire _34042_;
  wire _34043_;
  wire _34044_;
  wire _34045_;
  wire _34046_;
  wire _34047_;
  wire _34048_;
  wire _34049_;
  wire _34050_;
  wire _34051_;
  wire _34052_;
  wire _34053_;
  wire _34054_;
  wire _34055_;
  wire _34056_;
  wire _34057_;
  wire _34058_;
  wire _34059_;
  wire _34060_;
  wire _34061_;
  wire _34062_;
  wire _34063_;
  wire _34064_;
  wire _34065_;
  wire _34066_;
  wire _34067_;
  wire _34068_;
  wire _34069_;
  wire _34070_;
  wire _34071_;
  wire _34072_;
  wire _34073_;
  wire _34074_;
  wire _34075_;
  wire _34076_;
  wire _34077_;
  wire _34078_;
  wire _34079_;
  wire _34080_;
  wire _34081_;
  wire _34082_;
  wire _34083_;
  wire _34084_;
  wire _34085_;
  wire _34086_;
  wire _34087_;
  wire _34088_;
  wire _34089_;
  wire _34090_;
  wire _34091_;
  wire _34092_;
  wire _34093_;
  wire _34094_;
  wire _34095_;
  wire _34096_;
  wire _34097_;
  wire _34098_;
  wire _34099_;
  wire _34100_;
  wire _34101_;
  wire _34102_;
  wire _34103_;
  wire _34104_;
  wire _34105_;
  wire _34106_;
  wire _34107_;
  wire _34108_;
  wire _34109_;
  wire _34110_;
  wire _34111_;
  wire _34112_;
  wire _34113_;
  wire _34114_;
  wire _34115_;
  wire _34116_;
  wire _34117_;
  wire _34118_;
  wire _34119_;
  wire _34120_;
  wire _34121_;
  wire _34122_;
  wire _34123_;
  wire _34124_;
  wire _34125_;
  wire _34126_;
  wire _34127_;
  wire _34128_;
  wire _34129_;
  wire _34130_;
  wire _34131_;
  wire _34132_;
  wire _34133_;
  wire _34134_;
  wire _34135_;
  wire _34136_;
  wire _34137_;
  wire _34138_;
  wire _34139_;
  wire _34140_;
  wire _34141_;
  wire _34142_;
  wire _34143_;
  wire _34144_;
  wire _34145_;
  wire _34146_;
  wire _34147_;
  wire _34148_;
  wire _34149_;
  wire _34150_;
  wire _34151_;
  wire _34152_;
  wire _34153_;
  wire _34154_;
  wire _34155_;
  wire _34156_;
  wire _34157_;
  wire _34158_;
  wire _34159_;
  wire _34160_;
  wire _34161_;
  wire _34162_;
  wire _34163_;
  wire _34164_;
  wire _34165_;
  wire _34166_;
  wire _34167_;
  wire _34168_;
  wire _34169_;
  wire _34170_;
  wire _34171_;
  wire _34172_;
  wire _34173_;
  wire _34174_;
  wire _34175_;
  wire _34176_;
  wire _34177_;
  wire _34178_;
  wire _34179_;
  wire _34180_;
  wire _34181_;
  wire _34182_;
  wire _34183_;
  wire _34184_;
  wire _34185_;
  wire _34186_;
  wire _34187_;
  wire _34188_;
  wire _34189_;
  wire _34190_;
  wire _34191_;
  wire _34192_;
  wire _34193_;
  wire _34194_;
  wire _34195_;
  wire _34196_;
  wire _34197_;
  wire _34198_;
  wire _34199_;
  wire _34200_;
  wire _34201_;
  wire _34202_;
  wire _34203_;
  wire _34204_;
  wire _34205_;
  wire _34206_;
  wire _34207_;
  wire _34208_;
  wire _34209_;
  wire _34210_;
  wire _34211_;
  wire _34212_;
  wire _34213_;
  wire _34214_;
  wire _34215_;
  wire _34216_;
  wire _34217_;
  wire _34218_;
  wire _34219_;
  wire _34220_;
  wire _34221_;
  wire _34222_;
  wire _34223_;
  wire _34224_;
  wire _34225_;
  wire _34226_;
  wire _34227_;
  wire _34228_;
  wire _34229_;
  wire _34230_;
  wire _34231_;
  wire _34232_;
  wire _34233_;
  wire _34234_;
  wire _34235_;
  wire _34236_;
  wire _34237_;
  wire _34238_;
  wire _34239_;
  wire _34240_;
  wire _34241_;
  wire _34242_;
  wire _34243_;
  wire _34244_;
  wire _34245_;
  wire _34246_;
  wire _34247_;
  wire _34248_;
  wire _34249_;
  wire _34250_;
  wire _34251_;
  wire _34252_;
  wire _34253_;
  wire _34254_;
  wire _34255_;
  wire _34256_;
  wire _34257_;
  wire _34258_;
  wire _34259_;
  wire _34260_;
  wire _34261_;
  wire _34262_;
  wire _34263_;
  wire _34264_;
  wire _34265_;
  wire _34266_;
  wire _34267_;
  wire _34268_;
  wire _34269_;
  wire _34270_;
  wire _34271_;
  wire _34272_;
  wire _34273_;
  wire _34274_;
  wire _34275_;
  wire _34276_;
  wire _34277_;
  wire _34278_;
  wire _34279_;
  wire _34280_;
  wire _34281_;
  wire _34282_;
  wire _34283_;
  wire _34284_;
  wire _34285_;
  wire _34286_;
  wire _34287_;
  wire _34288_;
  wire _34289_;
  wire _34290_;
  wire _34291_;
  wire _34292_;
  wire _34293_;
  wire _34294_;
  wire _34295_;
  wire _34296_;
  wire _34297_;
  wire _34298_;
  wire _34299_;
  wire _34300_;
  wire _34301_;
  wire _34302_;
  wire _34303_;
  wire _34304_;
  wire _34305_;
  wire _34306_;
  wire _34307_;
  wire _34308_;
  wire _34309_;
  wire _34310_;
  wire _34311_;
  wire _34312_;
  wire _34313_;
  wire _34314_;
  wire _34315_;
  wire _34316_;
  wire _34317_;
  wire _34318_;
  wire _34319_;
  wire _34320_;
  wire _34321_;
  wire _34322_;
  wire _34323_;
  wire _34324_;
  wire _34325_;
  wire _34326_;
  wire _34327_;
  wire _34328_;
  wire _34329_;
  wire _34330_;
  wire _34331_;
  wire _34332_;
  wire _34333_;
  wire _34334_;
  wire _34335_;
  wire _34336_;
  wire _34337_;
  wire _34338_;
  wire _34339_;
  wire _34340_;
  wire _34341_;
  wire _34342_;
  wire _34343_;
  wire _34344_;
  wire _34345_;
  wire _34346_;
  wire _34347_;
  wire _34348_;
  wire _34349_;
  wire _34350_;
  wire _34351_;
  wire _34352_;
  wire _34353_;
  wire _34354_;
  wire _34355_;
  wire _34356_;
  wire _34357_;
  wire _34358_;
  wire _34359_;
  wire _34360_;
  wire _34361_;
  wire _34362_;
  wire _34363_;
  wire _34364_;
  wire _34365_;
  wire _34366_;
  wire _34367_;
  wire _34368_;
  wire _34369_;
  wire _34370_;
  wire _34371_;
  wire _34372_;
  wire _34373_;
  wire _34374_;
  wire _34375_;
  wire _34376_;
  wire _34377_;
  wire _34378_;
  wire _34379_;
  wire _34380_;
  wire _34381_;
  wire _34382_;
  wire _34383_;
  wire _34384_;
  wire _34385_;
  wire _34386_;
  wire _34387_;
  wire _34388_;
  wire _34389_;
  wire _34390_;
  wire _34391_;
  wire _34392_;
  wire _34393_;
  wire _34394_;
  wire _34395_;
  wire _34396_;
  wire _34397_;
  wire _34398_;
  wire _34399_;
  wire _34400_;
  wire _34401_;
  wire _34402_;
  wire _34403_;
  wire _34404_;
  wire _34405_;
  wire _34406_;
  wire _34407_;
  wire _34408_;
  wire _34409_;
  wire _34410_;
  wire _34411_;
  wire _34412_;
  wire _34413_;
  wire _34414_;
  wire _34415_;
  wire _34416_;
  wire _34417_;
  wire _34418_;
  wire _34419_;
  wire _34420_;
  wire _34421_;
  wire _34422_;
  wire _34423_;
  wire _34424_;
  wire _34425_;
  wire _34426_;
  wire _34427_;
  wire _34428_;
  wire _34429_;
  wire _34430_;
  wire _34431_;
  wire _34432_;
  wire _34433_;
  wire _34434_;
  wire _34435_;
  wire _34436_;
  wire _34437_;
  wire _34438_;
  wire _34439_;
  wire _34440_;
  wire _34441_;
  wire _34442_;
  wire _34443_;
  wire _34444_;
  wire _34445_;
  wire _34446_;
  wire _34447_;
  wire _34448_;
  wire _34449_;
  wire _34450_;
  wire _34451_;
  wire _34452_;
  wire _34453_;
  wire _34454_;
  wire _34455_;
  wire _34456_;
  wire _34457_;
  wire _34458_;
  wire _34459_;
  wire _34460_;
  wire _34461_;
  wire _34462_;
  wire _34463_;
  wire _34464_;
  wire _34465_;
  wire _34466_;
  wire _34467_;
  wire _34468_;
  wire _34469_;
  wire _34470_;
  wire _34471_;
  wire _34472_;
  wire _34473_;
  wire _34474_;
  wire _34475_;
  wire _34476_;
  wire _34477_;
  wire _34478_;
  wire _34479_;
  wire _34480_;
  wire _34481_;
  wire _34482_;
  wire _34483_;
  wire _34484_;
  wire _34485_;
  wire _34486_;
  wire _34487_;
  wire _34488_;
  wire _34489_;
  wire _34490_;
  wire _34491_;
  wire _34492_;
  wire _34493_;
  wire _34494_;
  wire _34495_;
  wire _34496_;
  wire _34497_;
  wire _34498_;
  wire _34499_;
  wire _34500_;
  wire _34501_;
  wire _34502_;
  wire _34503_;
  wire _34504_;
  wire _34505_;
  wire _34506_;
  wire _34507_;
  wire _34508_;
  wire _34509_;
  wire _34510_;
  wire _34511_;
  wire _34512_;
  wire _34513_;
  wire _34514_;
  wire _34515_;
  wire _34516_;
  wire _34517_;
  wire _34518_;
  wire _34519_;
  wire _34520_;
  wire _34521_;
  wire _34522_;
  wire _34523_;
  wire _34524_;
  wire _34525_;
  wire _34526_;
  wire _34527_;
  wire _34528_;
  wire _34529_;
  wire _34530_;
  wire _34531_;
  wire _34532_;
  wire _34533_;
  wire _34534_;
  wire _34535_;
  wire _34536_;
  wire _34537_;
  wire _34538_;
  wire _34539_;
  wire _34540_;
  wire _34541_;
  wire _34542_;
  wire _34543_;
  wire _34544_;
  wire _34545_;
  wire _34546_;
  wire _34547_;
  wire _34548_;
  wire _34549_;
  wire _34550_;
  wire _34551_;
  wire _34552_;
  wire _34553_;
  wire _34554_;
  wire _34555_;
  wire _34556_;
  wire _34557_;
  wire _34558_;
  wire _34559_;
  wire _34560_;
  wire _34561_;
  wire _34562_;
  wire _34563_;
  wire _34564_;
  wire _34565_;
  wire _34566_;
  wire _34567_;
  wire _34568_;
  wire _34569_;
  wire _34570_;
  wire _34571_;
  wire _34572_;
  wire _34573_;
  wire _34574_;
  wire _34575_;
  wire _34576_;
  wire _34577_;
  wire _34578_;
  wire _34579_;
  wire _34580_;
  wire _34581_;
  wire _34582_;
  wire _34583_;
  wire _34584_;
  wire _34585_;
  wire _34586_;
  wire _34587_;
  wire _34588_;
  wire _34589_;
  wire _34590_;
  wire _34591_;
  wire _34592_;
  wire _34593_;
  wire _34594_;
  wire _34595_;
  wire _34596_;
  wire _34597_;
  wire _34598_;
  wire _34599_;
  wire _34600_;
  wire _34601_;
  wire _34602_;
  wire _34603_;
  wire _34604_;
  wire _34605_;
  wire _34606_;
  wire _34607_;
  wire _34608_;
  wire _34609_;
  wire _34610_;
  wire _34611_;
  wire _34612_;
  wire _34613_;
  wire _34614_;
  wire _34615_;
  wire _34616_;
  wire _34617_;
  wire _34618_;
  wire _34619_;
  wire _34620_;
  wire _34621_;
  wire _34622_;
  wire _34623_;
  wire _34624_;
  wire _34625_;
  wire _34626_;
  wire _34627_;
  wire _34628_;
  wire _34629_;
  wire _34630_;
  wire _34631_;
  wire _34632_;
  wire _34633_;
  wire _34634_;
  wire _34635_;
  wire _34636_;
  wire _34637_;
  wire _34638_;
  wire _34639_;
  wire _34640_;
  wire _34641_;
  wire _34642_;
  wire _34643_;
  wire _34644_;
  wire _34645_;
  wire _34646_;
  wire _34647_;
  wire _34648_;
  wire _34649_;
  wire _34650_;
  wire _34651_;
  wire _34652_;
  wire _34653_;
  wire _34654_;
  wire _34655_;
  wire _34656_;
  wire _34657_;
  wire _34658_;
  wire _34659_;
  wire _34660_;
  wire _34661_;
  wire _34662_;
  wire _34663_;
  wire _34664_;
  wire _34665_;
  wire _34666_;
  wire _34667_;
  wire _34668_;
  wire _34669_;
  wire _34670_;
  wire _34671_;
  wire _34672_;
  wire _34673_;
  wire _34674_;
  wire _34675_;
  wire _34676_;
  wire _34677_;
  wire _34678_;
  wire _34679_;
  wire _34680_;
  wire _34681_;
  wire _34682_;
  wire _34683_;
  wire _34684_;
  wire _34685_;
  wire _34686_;
  wire _34687_;
  wire _34688_;
  wire _34689_;
  wire _34690_;
  wire _34691_;
  wire _34692_;
  wire _34693_;
  wire _34694_;
  wire _34695_;
  wire _34696_;
  wire _34697_;
  wire _34698_;
  wire _34699_;
  wire _34700_;
  wire _34701_;
  wire _34702_;
  wire _34703_;
  wire _34704_;
  wire _34705_;
  wire _34706_;
  wire _34707_;
  wire _34708_;
  wire _34709_;
  wire _34710_;
  wire _34711_;
  wire _34712_;
  wire _34713_;
  wire _34714_;
  wire _34715_;
  wire _34716_;
  wire _34717_;
  wire _34718_;
  wire _34719_;
  wire _34720_;
  wire _34721_;
  wire _34722_;
  wire _34723_;
  wire _34724_;
  wire _34725_;
  wire _34726_;
  wire _34727_;
  wire _34728_;
  wire _34729_;
  wire _34730_;
  wire _34731_;
  wire _34732_;
  wire _34733_;
  wire _34734_;
  wire _34735_;
  wire _34736_;
  wire _34737_;
  wire _34738_;
  wire _34739_;
  wire _34740_;
  wire _34741_;
  wire _34742_;
  wire _34743_;
  wire _34744_;
  wire _34745_;
  wire _34746_;
  wire _34747_;
  wire _34748_;
  wire _34749_;
  wire _34750_;
  wire _34751_;
  wire _34752_;
  wire _34753_;
  wire _34754_;
  wire _34755_;
  wire _34756_;
  wire _34757_;
  wire _34758_;
  wire _34759_;
  wire _34760_;
  wire _34761_;
  wire _34762_;
  wire _34763_;
  wire _34764_;
  wire _34765_;
  wire _34766_;
  wire _34767_;
  wire _34768_;
  wire _34769_;
  wire _34770_;
  wire _34771_;
  wire _34772_;
  wire _34773_;
  wire _34774_;
  wire _34775_;
  wire _34776_;
  wire _34777_;
  wire _34778_;
  wire _34779_;
  wire _34780_;
  wire _34781_;
  wire _34782_;
  wire _34783_;
  wire _34784_;
  wire _34785_;
  wire _34786_;
  wire _34787_;
  wire _34788_;
  wire _34789_;
  wire _34790_;
  wire _34791_;
  wire _34792_;
  wire _34793_;
  wire _34794_;
  wire _34795_;
  wire _34796_;
  wire _34797_;
  wire _34798_;
  wire _34799_;
  wire _34800_;
  wire _34801_;
  wire _34802_;
  wire _34803_;
  wire _34804_;
  wire _34805_;
  wire _34806_;
  wire _34807_;
  wire _34808_;
  wire _34809_;
  wire _34810_;
  wire _34811_;
  wire _34812_;
  wire _34813_;
  wire _34814_;
  wire _34815_;
  wire _34816_;
  wire _34817_;
  wire _34818_;
  wire _34819_;
  wire _34820_;
  wire _34821_;
  wire _34822_;
  wire _34823_;
  wire _34824_;
  wire _34825_;
  wire _34826_;
  wire _34827_;
  wire _34828_;
  wire _34829_;
  wire _34830_;
  wire _34831_;
  wire _34832_;
  wire _34833_;
  wire _34834_;
  wire _34835_;
  wire _34836_;
  wire _34837_;
  wire _34838_;
  wire _34839_;
  wire _34840_;
  wire _34841_;
  wire _34842_;
  wire _34843_;
  wire _34844_;
  wire _34845_;
  wire _34846_;
  wire _34847_;
  wire _34848_;
  wire _34849_;
  wire _34850_;
  wire _34851_;
  wire _34852_;
  wire _34853_;
  wire _34854_;
  wire _34855_;
  wire _34856_;
  wire _34857_;
  wire _34858_;
  wire _34859_;
  wire _34860_;
  wire _34861_;
  wire _34862_;
  wire _34863_;
  wire _34864_;
  wire _34865_;
  wire _34866_;
  wire _34867_;
  wire _34868_;
  wire _34869_;
  wire _34870_;
  wire _34871_;
  wire _34872_;
  wire _34873_;
  wire _34874_;
  wire _34875_;
  wire _34876_;
  wire _34877_;
  wire _34878_;
  wire _34879_;
  wire _34880_;
  wire _34881_;
  wire _34882_;
  wire _34883_;
  wire _34884_;
  wire _34885_;
  wire _34886_;
  wire _34887_;
  wire _34888_;
  wire _34889_;
  wire _34890_;
  wire _34891_;
  wire _34892_;
  wire _34893_;
  wire _34894_;
  wire _34895_;
  wire _34896_;
  wire _34897_;
  wire _34898_;
  wire _34899_;
  wire _34900_;
  wire _34901_;
  wire _34902_;
  wire _34903_;
  wire _34904_;
  wire _34905_;
  wire _34906_;
  wire _34907_;
  wire _34908_;
  wire _34909_;
  wire _34910_;
  wire _34911_;
  wire _34912_;
  wire _34913_;
  wire _34914_;
  wire _34915_;
  wire _34916_;
  wire _34917_;
  wire _34918_;
  wire _34919_;
  wire _34920_;
  wire _34921_;
  wire _34922_;
  wire _34923_;
  wire _34924_;
  wire _34925_;
  wire _34926_;
  wire _34927_;
  wire _34928_;
  wire _34929_;
  wire _34930_;
  wire _34931_;
  wire _34932_;
  wire _34933_;
  wire _34934_;
  wire _34935_;
  wire _34936_;
  wire _34937_;
  wire _34938_;
  wire _34939_;
  wire _34940_;
  wire _34941_;
  wire _34942_;
  wire _34943_;
  wire _34944_;
  wire _34945_;
  wire _34946_;
  wire _34947_;
  wire _34948_;
  wire _34949_;
  wire _34950_;
  wire _34951_;
  wire _34952_;
  wire _34953_;
  wire _34954_;
  wire _34955_;
  wire _34956_;
  wire _34957_;
  wire _34958_;
  wire _34959_;
  wire _34960_;
  wire _34961_;
  wire _34962_;
  wire _34963_;
  wire _34964_;
  wire _34965_;
  wire _34966_;
  wire _34967_;
  wire _34968_;
  wire _34969_;
  wire _34970_;
  wire _34971_;
  wire _34972_;
  wire _34973_;
  wire _34974_;
  wire _34975_;
  wire _34976_;
  wire _34977_;
  wire _34978_;
  wire _34979_;
  wire _34980_;
  wire _34981_;
  wire _34982_;
  wire _34983_;
  wire _34984_;
  wire _34985_;
  wire _34986_;
  wire _34987_;
  wire _34988_;
  wire _34989_;
  wire _34990_;
  wire _34991_;
  wire _34992_;
  wire _34993_;
  wire _34994_;
  wire _34995_;
  wire _34996_;
  wire _34997_;
  wire _34998_;
  wire _34999_;
  wire _35000_;
  wire _35001_;
  wire _35002_;
  wire _35003_;
  wire _35004_;
  wire _35005_;
  wire _35006_;
  wire _35007_;
  wire _35008_;
  wire _35009_;
  wire _35010_;
  wire _35011_;
  wire _35012_;
  wire _35013_;
  wire _35014_;
  wire _35015_;
  wire _35016_;
  wire _35017_;
  wire _35018_;
  wire _35019_;
  wire _35020_;
  wire _35021_;
  wire _35022_;
  wire _35023_;
  wire _35024_;
  wire _35025_;
  wire _35026_;
  wire _35027_;
  wire _35028_;
  wire _35029_;
  wire _35030_;
  wire _35031_;
  wire _35032_;
  wire _35033_;
  wire _35034_;
  wire _35035_;
  wire _35036_;
  wire _35037_;
  wire _35038_;
  wire _35039_;
  wire _35040_;
  wire _35041_;
  wire _35042_;
  wire _35043_;
  wire _35044_;
  wire _35045_;
  wire _35046_;
  wire _35047_;
  wire _35048_;
  wire _35049_;
  wire _35050_;
  wire _35051_;
  wire _35052_;
  wire _35053_;
  wire _35054_;
  wire _35055_;
  wire _35056_;
  wire _35057_;
  wire _35058_;
  wire _35059_;
  wire _35060_;
  wire _35061_;
  wire _35062_;
  wire _35063_;
  wire _35064_;
  wire _35065_;
  wire _35066_;
  wire _35067_;
  wire _35068_;
  wire _35069_;
  wire _35070_;
  wire _35071_;
  wire _35072_;
  wire _35073_;
  wire _35074_;
  wire _35075_;
  wire _35076_;
  wire _35077_;
  wire _35078_;
  wire _35079_;
  wire _35080_;
  wire _35081_;
  wire _35082_;
  wire _35083_;
  wire _35084_;
  wire _35085_;
  wire _35086_;
  wire _35087_;
  wire _35088_;
  wire _35089_;
  wire _35090_;
  wire _35091_;
  wire _35092_;
  wire _35093_;
  wire _35094_;
  wire _35095_;
  wire _35096_;
  wire _35097_;
  wire _35098_;
  wire _35099_;
  wire _35100_;
  wire _35101_;
  wire _35102_;
  wire _35103_;
  wire _35104_;
  wire _35105_;
  wire _35106_;
  wire _35107_;
  wire _35108_;
  wire _35109_;
  wire _35110_;
  wire _35111_;
  wire _35112_;
  wire _35113_;
  wire _35114_;
  wire _35115_;
  wire _35116_;
  wire _35117_;
  wire _35118_;
  wire _35119_;
  wire _35120_;
  wire _35121_;
  wire _35122_;
  wire _35123_;
  wire _35124_;
  wire _35125_;
  wire _35126_;
  wire _35127_;
  wire _35128_;
  wire _35129_;
  wire _35130_;
  wire _35131_;
  wire _35132_;
  wire _35133_;
  wire _35134_;
  wire _35135_;
  wire _35136_;
  wire _35137_;
  wire _35138_;
  wire _35139_;
  wire _35140_;
  wire _35141_;
  wire _35142_;
  wire _35143_;
  wire _35144_;
  wire _35145_;
  wire _35146_;
  wire _35147_;
  wire _35148_;
  wire _35149_;
  wire _35150_;
  wire _35151_;
  wire _35152_;
  wire _35153_;
  wire _35154_;
  wire _35155_;
  wire _35156_;
  wire _35157_;
  wire _35158_;
  wire _35159_;
  wire _35160_;
  wire _35161_;
  wire _35162_;
  wire _35163_;
  wire _35164_;
  wire _35165_;
  wire _35166_;
  wire _35167_;
  wire _35168_;
  wire _35169_;
  wire _35170_;
  wire _35171_;
  wire _35172_;
  wire _35173_;
  wire _35174_;
  wire _35175_;
  wire _35176_;
  wire _35177_;
  wire _35178_;
  wire _35179_;
  wire _35180_;
  wire _35181_;
  wire _35182_;
  wire _35183_;
  wire _35184_;
  wire _35185_;
  wire _35186_;
  wire _35187_;
  wire _35188_;
  wire _35189_;
  wire _35190_;
  wire _35191_;
  wire _35192_;
  wire _35193_;
  wire _35194_;
  wire _35195_;
  wire _35196_;
  wire _35197_;
  wire _35198_;
  wire _35199_;
  wire _35200_;
  wire _35201_;
  wire _35202_;
  wire _35203_;
  wire _35204_;
  wire _35205_;
  wire _35206_;
  wire _35207_;
  wire _35208_;
  wire _35209_;
  wire _35210_;
  wire _35211_;
  wire _35212_;
  wire _35213_;
  wire _35214_;
  wire _35215_;
  wire _35216_;
  wire _35217_;
  wire _35218_;
  wire _35219_;
  wire _35220_;
  wire _35221_;
  wire _35222_;
  wire _35223_;
  wire _35224_;
  wire _35225_;
  wire _35226_;
  wire _35227_;
  wire _35228_;
  wire _35229_;
  wire _35230_;
  wire _35231_;
  wire _35232_;
  wire _35233_;
  wire _35234_;
  wire _35235_;
  wire _35236_;
  wire _35237_;
  wire _35238_;
  wire _35239_;
  wire _35240_;
  wire _35241_;
  wire _35242_;
  wire _35243_;
  wire _35244_;
  wire _35245_;
  wire _35246_;
  wire _35247_;
  wire _35248_;
  wire _35249_;
  wire _35250_;
  wire _35251_;
  wire _35252_;
  wire _35253_;
  wire _35254_;
  wire _35255_;
  wire _35256_;
  wire _35257_;
  wire _35258_;
  wire _35259_;
  wire _35260_;
  wire _35261_;
  wire _35262_;
  wire _35263_;
  wire _35264_;
  wire _35265_;
  wire _35266_;
  wire _35267_;
  wire _35268_;
  wire _35269_;
  wire _35270_;
  wire _35271_;
  wire _35272_;
  wire _35273_;
  wire _35274_;
  wire _35275_;
  wire _35276_;
  wire _35277_;
  wire _35278_;
  wire _35279_;
  wire _35280_;
  wire _35281_;
  wire _35282_;
  wire _35283_;
  wire _35284_;
  wire _35285_;
  wire _35286_;
  wire _35287_;
  wire _35288_;
  wire _35289_;
  wire _35290_;
  wire _35291_;
  wire _35292_;
  wire _35293_;
  wire _35294_;
  wire _35295_;
  wire _35296_;
  wire _35297_;
  wire _35298_;
  wire _35299_;
  wire _35300_;
  wire _35301_;
  wire _35302_;
  wire _35303_;
  wire _35304_;
  wire _35305_;
  wire _35306_;
  wire _35307_;
  wire _35308_;
  wire _35309_;
  wire _35310_;
  wire _35311_;
  wire _35312_;
  wire _35313_;
  wire _35314_;
  wire _35315_;
  wire _35316_;
  wire _35317_;
  wire _35318_;
  wire _35319_;
  wire _35320_;
  wire _35321_;
  wire _35322_;
  wire _35323_;
  wire _35324_;
  wire _35325_;
  wire _35326_;
  wire _35327_;
  wire _35328_;
  wire _35329_;
  wire _35330_;
  wire _35331_;
  wire _35332_;
  wire _35333_;
  wire _35334_;
  wire _35335_;
  wire _35336_;
  wire _35337_;
  wire _35338_;
  wire _35339_;
  wire _35340_;
  wire _35341_;
  wire _35342_;
  wire _35343_;
  wire _35344_;
  wire _35345_;
  wire _35346_;
  wire _35347_;
  wire _35348_;
  wire _35349_;
  wire _35350_;
  wire _35351_;
  wire _35352_;
  wire _35353_;
  wire _35354_;
  wire _35355_;
  wire _35356_;
  wire _35357_;
  wire _35358_;
  wire _35359_;
  wire _35360_;
  wire _35361_;
  wire _35362_;
  wire _35363_;
  wire _35364_;
  wire _35365_;
  wire _35366_;
  wire _35367_;
  wire _35368_;
  wire _35369_;
  wire _35370_;
  wire _35371_;
  wire _35372_;
  wire _35373_;
  wire _35374_;
  wire _35375_;
  wire _35376_;
  wire _35377_;
  wire _35378_;
  wire _35379_;
  wire _35380_;
  wire _35381_;
  wire _35382_;
  wire _35383_;
  wire _35384_;
  wire _35385_;
  wire _35386_;
  wire _35387_;
  wire _35388_;
  wire _35389_;
  wire _35390_;
  wire _35391_;
  wire _35392_;
  wire _35393_;
  wire _35394_;
  wire _35395_;
  wire _35396_;
  wire _35397_;
  wire _35398_;
  wire _35399_;
  wire _35400_;
  wire _35401_;
  wire _35402_;
  wire _35403_;
  wire _35404_;
  wire _35405_;
  wire _35406_;
  wire _35407_;
  wire _35408_;
  wire _35409_;
  wire _35410_;
  wire _35411_;
  wire _35412_;
  wire _35413_;
  wire _35414_;
  wire _35415_;
  wire _35416_;
  wire _35417_;
  wire _35418_;
  wire _35419_;
  wire _35420_;
  wire _35421_;
  wire _35422_;
  wire _35423_;
  wire _35424_;
  wire _35425_;
  wire _35426_;
  wire _35427_;
  wire _35428_;
  wire _35429_;
  wire _35430_;
  wire _35431_;
  wire _35432_;
  wire _35433_;
  wire _35434_;
  wire _35435_;
  wire _35436_;
  wire _35437_;
  wire _35438_;
  wire _35439_;
  wire _35440_;
  wire _35441_;
  wire _35442_;
  wire _35443_;
  wire _35444_;
  wire _35445_;
  wire _35446_;
  wire _35447_;
  wire _35448_;
  wire _35449_;
  wire _35450_;
  wire _35451_;
  wire _35452_;
  wire _35453_;
  wire _35454_;
  wire _35455_;
  wire _35456_;
  wire _35457_;
  wire _35458_;
  wire _35459_;
  wire _35460_;
  wire _35461_;
  wire _35462_;
  wire _35463_;
  wire _35464_;
  wire _35465_;
  wire _35466_;
  wire _35467_;
  wire _35468_;
  wire _35469_;
  wire _35470_;
  wire _35471_;
  wire _35472_;
  wire _35473_;
  wire _35474_;
  wire _35475_;
  wire _35476_;
  wire _35477_;
  wire _35478_;
  wire _35479_;
  wire _35480_;
  wire _35481_;
  wire _35482_;
  wire _35483_;
  wire _35484_;
  wire _35485_;
  wire _35486_;
  wire _35487_;
  wire _35488_;
  wire _35489_;
  wire _35490_;
  wire _35491_;
  wire _35492_;
  wire _35493_;
  wire _35494_;
  wire _35495_;
  wire _35496_;
  wire _35497_;
  wire _35498_;
  wire _35499_;
  wire _35500_;
  wire _35501_;
  wire _35502_;
  wire _35503_;
  wire _35504_;
  wire _35505_;
  wire _35506_;
  wire _35507_;
  wire _35508_;
  wire _35509_;
  wire _35510_;
  wire _35511_;
  wire _35512_;
  wire _35513_;
  wire _35514_;
  wire _35515_;
  wire _35516_;
  wire _35517_;
  wire _35518_;
  wire _35519_;
  wire _35520_;
  wire _35521_;
  wire _35522_;
  wire _35523_;
  wire _35524_;
  wire _35525_;
  wire _35526_;
  wire _35527_;
  wire _35528_;
  wire _35529_;
  wire _35530_;
  wire _35531_;
  wire _35532_;
  wire _35533_;
  wire _35534_;
  wire _35535_;
  wire _35536_;
  wire _35537_;
  wire _35538_;
  wire _35539_;
  wire _35540_;
  wire _35541_;
  wire _35542_;
  wire _35543_;
  wire _35544_;
  wire _35545_;
  wire _35546_;
  wire _35547_;
  wire _35548_;
  wire _35549_;
  wire _35550_;
  wire _35551_;
  wire _35552_;
  wire _35553_;
  wire _35554_;
  wire _35555_;
  wire _35556_;
  wire _35557_;
  wire _35558_;
  wire _35559_;
  wire _35560_;
  wire _35561_;
  wire _35562_;
  wire _35563_;
  wire _35564_;
  wire _35565_;
  wire _35566_;
  wire _35567_;
  wire _35568_;
  wire _35569_;
  wire _35570_;
  wire _35571_;
  wire _35572_;
  wire _35573_;
  wire _35574_;
  wire _35575_;
  wire _35576_;
  wire _35577_;
  wire _35578_;
  wire _35579_;
  wire _35580_;
  wire _35581_;
  wire _35582_;
  wire _35583_;
  wire _35584_;
  wire _35585_;
  wire _35586_;
  wire _35587_;
  wire _35588_;
  wire _35589_;
  wire _35590_;
  wire _35591_;
  wire _35592_;
  wire _35593_;
  wire _35594_;
  wire _35595_;
  wire _35596_;
  wire _35597_;
  wire _35598_;
  wire _35599_;
  wire _35600_;
  wire _35601_;
  wire _35602_;
  wire _35603_;
  wire _35604_;
  wire _35605_;
  wire _35606_;
  wire _35607_;
  wire _35608_;
  wire _35609_;
  wire _35610_;
  wire _35611_;
  wire _35612_;
  wire _35613_;
  wire _35614_;
  wire _35615_;
  wire _35616_;
  wire _35617_;
  wire _35618_;
  wire _35619_;
  wire _35620_;
  wire _35621_;
  wire _35622_;
  wire _35623_;
  wire _35624_;
  wire _35625_;
  wire _35626_;
  wire _35627_;
  wire _35628_;
  wire _35629_;
  wire _35630_;
  wire _35631_;
  wire _35632_;
  wire _35633_;
  wire _35634_;
  wire _35635_;
  wire _35636_;
  wire _35637_;
  wire _35638_;
  wire _35639_;
  wire _35640_;
  wire _35641_;
  wire _35642_;
  wire _35643_;
  wire _35644_;
  wire _35645_;
  wire _35646_;
  wire _35647_;
  wire _35648_;
  wire _35649_;
  wire _35650_;
  wire _35651_;
  wire _35652_;
  wire _35653_;
  wire _35654_;
  wire _35655_;
  wire _35656_;
  wire _35657_;
  wire _35658_;
  wire _35659_;
  wire _35660_;
  wire _35661_;
  wire _35662_;
  wire _35663_;
  wire _35664_;
  wire _35665_;
  wire _35666_;
  wire _35667_;
  wire _35668_;
  wire _35669_;
  wire _35670_;
  wire _35671_;
  wire _35672_;
  wire _35673_;
  wire _35674_;
  wire _35675_;
  wire _35676_;
  wire _35677_;
  wire _35678_;
  wire _35679_;
  wire _35680_;
  wire _35681_;
  wire _35682_;
  wire _35683_;
  wire _35684_;
  wire _35685_;
  wire _35686_;
  wire _35687_;
  wire _35688_;
  wire _35689_;
  wire _35690_;
  wire _35691_;
  wire _35692_;
  wire _35693_;
  wire _35694_;
  wire _35695_;
  wire _35696_;
  wire _35697_;
  wire _35698_;
  wire _35699_;
  wire _35700_;
  wire _35701_;
  wire _35702_;
  wire _35703_;
  wire _35704_;
  wire _35705_;
  wire _35706_;
  wire _35707_;
  wire _35708_;
  wire _35709_;
  wire _35710_;
  wire _35711_;
  wire _35712_;
  wire _35713_;
  wire _35714_;
  wire _35715_;
  wire _35716_;
  wire _35717_;
  wire _35718_;
  wire _35719_;
  wire _35720_;
  wire _35721_;
  wire _35722_;
  wire _35723_;
  wire _35724_;
  wire _35725_;
  wire _35726_;
  wire _35727_;
  wire _35728_;
  wire _35729_;
  wire _35730_;
  wire _35731_;
  wire _35732_;
  wire _35733_;
  wire _35734_;
  wire _35735_;
  wire _35736_;
  wire _35737_;
  wire _35738_;
  wire _35739_;
  wire _35740_;
  wire _35741_;
  wire _35742_;
  wire _35743_;
  wire _35744_;
  wire _35745_;
  wire _35746_;
  wire _35747_;
  wire _35748_;
  wire _35749_;
  wire _35750_;
  wire _35751_;
  wire _35752_;
  wire _35753_;
  wire _35754_;
  wire _35755_;
  wire _35756_;
  wire _35757_;
  wire _35758_;
  wire _35759_;
  wire _35760_;
  wire _35761_;
  wire _35762_;
  wire _35763_;
  wire _35764_;
  wire _35765_;
  wire _35766_;
  wire _35767_;
  wire _35768_;
  wire _35769_;
  wire _35770_;
  wire _35771_;
  wire _35772_;
  wire _35773_;
  wire _35774_;
  wire _35775_;
  wire _35776_;
  wire _35777_;
  wire _35778_;
  wire _35779_;
  wire _35780_;
  wire _35781_;
  wire _35782_;
  wire _35783_;
  wire _35784_;
  wire _35785_;
  wire _35786_;
  wire _35787_;
  wire _35788_;
  wire _35789_;
  wire _35790_;
  wire _35791_;
  wire _35792_;
  wire _35793_;
  wire _35794_;
  wire _35795_;
  wire _35796_;
  wire _35797_;
  wire _35798_;
  wire _35799_;
  wire _35800_;
  wire _35801_;
  wire _35802_;
  wire _35803_;
  wire _35804_;
  wire _35805_;
  wire _35806_;
  wire _35807_;
  wire _35808_;
  wire _35809_;
  wire _35810_;
  wire _35811_;
  wire _35812_;
  wire _35813_;
  wire _35814_;
  wire _35815_;
  wire _35816_;
  wire _35817_;
  wire _35818_;
  wire _35819_;
  wire _35820_;
  wire _35821_;
  wire _35822_;
  wire _35823_;
  wire _35824_;
  wire _35825_;
  wire _35826_;
  wire _35827_;
  wire _35828_;
  wire _35829_;
  wire _35830_;
  wire _35831_;
  wire _35832_;
  wire _35833_;
  wire _35834_;
  wire _35835_;
  wire _35836_;
  wire _35837_;
  wire _35838_;
  wire _35839_;
  wire _35840_;
  wire _35841_;
  wire _35842_;
  wire _35843_;
  wire _35844_;
  wire _35845_;
  wire _35846_;
  wire _35847_;
  wire _35848_;
  wire _35849_;
  wire _35850_;
  wire _35851_;
  wire _35852_;
  wire _35853_;
  wire _35854_;
  wire _35855_;
  wire _35856_;
  wire _35857_;
  wire _35858_;
  wire _35859_;
  wire _35860_;
  wire _35861_;
  wire _35862_;
  wire _35863_;
  wire _35864_;
  wire _35865_;
  wire _35866_;
  wire _35867_;
  wire _35868_;
  wire _35869_;
  wire _35870_;
  wire _35871_;
  wire _35872_;
  wire _35873_;
  wire _35874_;
  wire _35875_;
  wire _35876_;
  wire _35877_;
  wire _35878_;
  wire _35879_;
  wire _35880_;
  wire _35881_;
  wire _35882_;
  wire _35883_;
  wire _35884_;
  wire _35885_;
  wire _35886_;
  wire _35887_;
  wire _35888_;
  wire _35889_;
  wire _35890_;
  wire _35891_;
  wire _35892_;
  wire _35893_;
  wire _35894_;
  wire _35895_;
  wire _35896_;
  wire _35897_;
  wire _35898_;
  wire _35899_;
  wire _35900_;
  wire _35901_;
  wire _35902_;
  wire _35903_;
  wire _35904_;
  wire _35905_;
  wire _35906_;
  wire _35907_;
  wire _35908_;
  wire _35909_;
  wire _35910_;
  wire _35911_;
  wire _35912_;
  wire _35913_;
  wire _35914_;
  wire _35915_;
  wire _35916_;
  wire _35917_;
  wire _35918_;
  wire _35919_;
  wire _35920_;
  wire _35921_;
  wire _35922_;
  wire _35923_;
  wire _35924_;
  wire _35925_;
  wire _35926_;
  wire _35927_;
  wire _35928_;
  wire _35929_;
  wire _35930_;
  wire _35931_;
  wire _35932_;
  wire _35933_;
  wire _35934_;
  wire _35935_;
  wire _35936_;
  wire _35937_;
  wire _35938_;
  wire _35939_;
  wire _35940_;
  wire _35941_;
  wire _35942_;
  wire _35943_;
  wire _35944_;
  wire _35945_;
  wire _35946_;
  wire _35947_;
  wire _35948_;
  wire _35949_;
  wire _35950_;
  wire _35951_;
  wire _35952_;
  wire _35953_;
  wire _35954_;
  wire _35955_;
  wire _35956_;
  wire _35957_;
  wire _35958_;
  wire _35959_;
  wire _35960_;
  wire _35961_;
  wire _35962_;
  wire _35963_;
  wire _35964_;
  wire _35965_;
  wire _35966_;
  wire _35967_;
  wire _35968_;
  wire _35969_;
  wire _35970_;
  wire _35971_;
  wire _35972_;
  wire _35973_;
  wire _35974_;
  wire _35975_;
  wire _35976_;
  wire _35977_;
  wire _35978_;
  wire _35979_;
  wire _35980_;
  wire _35981_;
  wire _35982_;
  wire _35983_;
  wire _35984_;
  wire _35985_;
  wire _35986_;
  wire _35987_;
  wire _35988_;
  wire _35989_;
  wire _35990_;
  wire _35991_;
  wire _35992_;
  wire _35993_;
  wire _35994_;
  wire _35995_;
  wire _35996_;
  wire _35997_;
  wire _35998_;
  wire _35999_;
  wire _36000_;
  wire _36001_;
  wire _36002_;
  wire _36003_;
  wire _36004_;
  wire _36005_;
  wire _36006_;
  wire _36007_;
  wire _36008_;
  wire _36009_;
  wire _36010_;
  wire _36011_;
  wire _36012_;
  wire _36013_;
  wire _36014_;
  wire _36015_;
  wire _36016_;
  wire _36017_;
  wire _36018_;
  wire _36019_;
  wire _36020_;
  wire _36021_;
  wire _36022_;
  wire _36023_;
  wire _36024_;
  wire _36025_;
  wire _36026_;
  wire _36027_;
  wire _36028_;
  wire _36029_;
  wire _36030_;
  wire _36031_;
  wire _36032_;
  wire _36033_;
  wire _36034_;
  wire _36035_;
  wire _36036_;
  wire _36037_;
  wire _36038_;
  wire _36039_;
  wire _36040_;
  wire _36041_;
  wire _36042_;
  wire _36043_;
  wire _36044_;
  wire _36045_;
  wire _36046_;
  wire _36047_;
  wire _36048_;
  wire _36049_;
  wire _36050_;
  wire _36051_;
  wire _36052_;
  wire _36053_;
  wire _36054_;
  wire _36055_;
  wire _36056_;
  wire _36057_;
  wire _36058_;
  wire _36059_;
  wire _36060_;
  wire _36061_;
  wire _36062_;
  wire _36063_;
  wire _36064_;
  wire _36065_;
  wire _36066_;
  wire _36067_;
  wire _36068_;
  wire _36069_;
  wire _36070_;
  wire _36071_;
  wire _36072_;
  wire _36073_;
  wire _36074_;
  wire _36075_;
  wire _36076_;
  wire _36077_;
  wire _36078_;
  wire _36079_;
  wire _36080_;
  wire _36081_;
  wire _36082_;
  wire _36083_;
  wire _36084_;
  wire _36085_;
  wire _36086_;
  wire _36087_;
  wire _36088_;
  wire _36089_;
  wire _36090_;
  wire _36091_;
  wire _36092_;
  wire _36093_;
  wire _36094_;
  wire _36095_;
  wire _36096_;
  wire _36097_;
  wire _36098_;
  wire _36099_;
  wire _36100_;
  wire _36101_;
  wire _36102_;
  wire _36103_;
  wire _36104_;
  wire _36105_;
  wire _36106_;
  wire _36107_;
  wire _36108_;
  wire _36109_;
  wire _36110_;
  wire _36111_;
  wire _36112_;
  wire _36113_;
  wire _36114_;
  wire _36115_;
  wire _36116_;
  wire _36117_;
  wire _36118_;
  wire _36119_;
  wire _36120_;
  wire _36121_;
  wire _36122_;
  wire _36123_;
  wire _36124_;
  wire _36125_;
  wire _36126_;
  wire _36127_;
  wire _36128_;
  wire _36129_;
  wire _36130_;
  wire _36131_;
  wire _36132_;
  wire _36133_;
  wire _36134_;
  wire _36135_;
  wire _36136_;
  wire _36137_;
  wire _36138_;
  wire _36139_;
  wire _36140_;
  wire _36141_;
  wire _36142_;
  wire _36143_;
  wire _36144_;
  wire _36145_;
  wire _36146_;
  wire _36147_;
  wire _36148_;
  wire _36149_;
  wire _36150_;
  wire _36151_;
  wire _36152_;
  wire _36153_;
  wire _36154_;
  wire _36155_;
  wire _36156_;
  wire _36157_;
  wire _36158_;
  wire _36159_;
  wire _36160_;
  wire _36161_;
  wire _36162_;
  wire _36163_;
  wire _36164_;
  wire _36165_;
  wire _36166_;
  wire _36167_;
  wire _36168_;
  wire _36169_;
  wire _36170_;
  wire _36171_;
  wire _36172_;
  wire _36173_;
  wire _36174_;
  wire _36175_;
  wire _36176_;
  wire _36177_;
  wire _36178_;
  wire _36179_;
  wire _36180_;
  wire _36181_;
  wire _36182_;
  wire _36183_;
  wire _36184_;
  wire _36185_;
  wire _36186_;
  wire _36187_;
  wire _36188_;
  wire _36189_;
  wire _36190_;
  wire _36191_;
  wire _36192_;
  wire _36193_;
  wire _36194_;
  wire _36195_;
  wire _36196_;
  wire _36197_;
  wire _36198_;
  wire _36199_;
  wire _36200_;
  wire _36201_;
  wire _36202_;
  wire _36203_;
  wire _36204_;
  wire _36205_;
  wire _36206_;
  wire _36207_;
  wire _36208_;
  wire _36209_;
  wire _36210_;
  wire _36211_;
  wire _36212_;
  wire _36213_;
  wire _36214_;
  wire _36215_;
  wire _36216_;
  wire _36217_;
  wire _36218_;
  wire _36219_;
  wire _36220_;
  wire _36221_;
  wire _36222_;
  wire _36223_;
  wire _36224_;
  wire _36225_;
  wire _36226_;
  wire _36227_;
  wire _36228_;
  wire _36229_;
  wire _36230_;
  wire _36231_;
  wire _36232_;
  wire _36233_;
  wire _36234_;
  wire _36235_;
  wire _36236_;
  wire _36237_;
  wire _36238_;
  wire _36239_;
  wire _36240_;
  wire _36241_;
  wire _36242_;
  wire _36243_;
  wire _36244_;
  wire _36245_;
  wire _36246_;
  wire _36247_;
  wire _36248_;
  wire _36249_;
  wire _36250_;
  wire _36251_;
  wire _36252_;
  wire _36253_;
  wire _36254_;
  wire _36255_;
  wire _36256_;
  wire _36257_;
  wire _36258_;
  wire _36259_;
  wire _36260_;
  wire _36261_;
  wire _36262_;
  wire _36263_;
  wire _36264_;
  wire _36265_;
  wire _36266_;
  wire _36267_;
  wire _36268_;
  wire _36269_;
  wire _36270_;
  wire _36271_;
  wire _36272_;
  wire _36273_;
  wire _36274_;
  wire _36275_;
  wire _36276_;
  wire _36277_;
  wire _36278_;
  wire _36279_;
  wire _36280_;
  wire _36281_;
  wire _36282_;
  wire _36283_;
  wire _36284_;
  wire _36285_;
  wire _36286_;
  wire _36287_;
  wire _36288_;
  wire _36289_;
  wire _36290_;
  wire _36291_;
  wire _36292_;
  wire _36293_;
  wire _36294_;
  wire _36295_;
  wire _36296_;
  wire _36297_;
  wire _36298_;
  wire _36299_;
  wire _36300_;
  wire _36301_;
  wire _36302_;
  wire _36303_;
  wire _36304_;
  wire _36305_;
  wire _36306_;
  wire _36307_;
  wire _36308_;
  wire _36309_;
  wire _36310_;
  wire _36311_;
  wire _36312_;
  wire _36313_;
  wire _36314_;
  wire _36315_;
  wire _36316_;
  wire _36317_;
  wire _36318_;
  wire _36319_;
  wire _36320_;
  wire _36321_;
  wire _36322_;
  wire _36323_;
  wire _36324_;
  wire _36325_;
  wire _36326_;
  wire _36327_;
  wire _36328_;
  wire _36329_;
  wire _36330_;
  wire _36331_;
  wire _36332_;
  wire _36333_;
  wire _36334_;
  wire _36335_;
  wire _36336_;
  wire _36337_;
  wire _36338_;
  wire _36339_;
  wire _36340_;
  wire _36341_;
  wire _36342_;
  wire _36343_;
  wire _36344_;
  wire _36345_;
  wire _36346_;
  wire _36347_;
  wire _36348_;
  wire _36349_;
  wire _36350_;
  wire _36351_;
  wire _36352_;
  wire _36353_;
  wire _36354_;
  wire _36355_;
  wire _36356_;
  wire _36357_;
  wire _36358_;
  wire _36359_;
  wire _36360_;
  wire _36361_;
  wire _36362_;
  wire _36363_;
  wire _36364_;
  wire _36365_;
  wire _36366_;
  wire _36367_;
  wire _36368_;
  wire _36369_;
  wire _36370_;
  wire _36371_;
  wire _36372_;
  wire _36373_;
  wire _36374_;
  wire _36375_;
  wire _36376_;
  wire _36377_;
  wire _36378_;
  wire _36379_;
  wire _36380_;
  wire _36381_;
  wire _36382_;
  wire _36383_;
  wire _36384_;
  wire _36385_;
  wire _36386_;
  wire _36387_;
  wire _36388_;
  wire _36389_;
  wire _36390_;
  wire _36391_;
  wire _36392_;
  wire _36393_;
  wire _36394_;
  wire _36395_;
  wire _36396_;
  wire _36397_;
  wire _36398_;
  wire _36399_;
  wire _36400_;
  wire _36401_;
  wire _36402_;
  wire _36403_;
  wire _36404_;
  wire _36405_;
  wire _36406_;
  wire _36407_;
  wire _36408_;
  wire _36409_;
  wire _36410_;
  wire _36411_;
  wire _36412_;
  wire _36413_;
  wire _36414_;
  wire _36415_;
  wire _36416_;
  wire _36417_;
  wire _36418_;
  wire _36419_;
  wire _36420_;
  wire _36421_;
  wire _36422_;
  wire _36423_;
  wire _36424_;
  wire _36425_;
  wire _36426_;
  wire _36427_;
  wire _36428_;
  wire _36429_;
  wire _36430_;
  wire _36431_;
  wire _36432_;
  wire _36433_;
  wire _36434_;
  wire _36435_;
  wire _36436_;
  wire _36437_;
  wire _36438_;
  wire _36439_;
  wire _36440_;
  wire _36441_;
  wire _36442_;
  wire _36443_;
  wire _36444_;
  wire _36445_;
  wire _36446_;
  wire _36447_;
  wire _36448_;
  wire _36449_;
  wire _36450_;
  wire _36451_;
  wire _36452_;
  wire _36453_;
  wire _36454_;
  wire _36455_;
  wire _36456_;
  wire _36457_;
  wire _36458_;
  wire _36459_;
  wire _36460_;
  wire _36461_;
  wire _36462_;
  wire _36463_;
  wire _36464_;
  wire _36465_;
  wire _36466_;
  wire _36467_;
  wire _36468_;
  wire _36469_;
  wire _36470_;
  wire _36471_;
  wire _36472_;
  wire _36473_;
  wire _36474_;
  wire _36475_;
  wire _36476_;
  wire _36477_;
  wire _36478_;
  wire _36479_;
  wire _36480_;
  wire _36481_;
  wire _36482_;
  wire _36483_;
  wire _36484_;
  wire _36485_;
  wire _36486_;
  wire _36487_;
  wire _36488_;
  wire _36489_;
  wire _36490_;
  wire _36491_;
  wire _36492_;
  wire _36493_;
  wire _36494_;
  wire _36495_;
  wire _36496_;
  wire _36497_;
  wire _36498_;
  wire _36499_;
  wire _36500_;
  wire _36501_;
  wire _36502_;
  wire _36503_;
  wire _36504_;
  wire _36505_;
  wire _36506_;
  wire _36507_;
  wire _36508_;
  wire _36509_;
  wire _36510_;
  wire _36511_;
  wire _36512_;
  wire _36513_;
  wire _36514_;
  wire _36515_;
  wire _36516_;
  wire _36517_;
  wire _36518_;
  wire _36519_;
  wire _36520_;
  wire _36521_;
  wire _36522_;
  wire _36523_;
  wire _36524_;
  wire _36525_;
  wire _36526_;
  wire _36527_;
  wire _36528_;
  wire _36529_;
  wire _36530_;
  wire _36531_;
  wire _36532_;
  wire _36533_;
  wire _36534_;
  wire _36535_;
  wire _36536_;
  wire _36537_;
  wire _36538_;
  wire _36539_;
  wire _36540_;
  wire _36541_;
  wire _36542_;
  wire _36543_;
  wire _36544_;
  wire _36545_;
  wire _36546_;
  wire _36547_;
  wire _36548_;
  wire _36549_;
  wire _36550_;
  wire _36551_;
  wire _36552_;
  wire _36553_;
  wire _36554_;
  wire _36555_;
  wire _36556_;
  wire _36557_;
  wire _36558_;
  wire _36559_;
  wire _36560_;
  wire _36561_;
  wire _36562_;
  wire _36563_;
  wire _36564_;
  wire _36565_;
  wire _36566_;
  wire _36567_;
  wire _36568_;
  wire _36569_;
  wire _36570_;
  wire _36571_;
  wire _36572_;
  wire _36573_;
  wire _36574_;
  wire _36575_;
  wire _36576_;
  wire _36577_;
  wire _36578_;
  wire _36579_;
  wire _36580_;
  wire _36581_;
  wire _36582_;
  wire _36583_;
  wire _36584_;
  wire _36585_;
  wire _36586_;
  wire _36587_;
  wire _36588_;
  wire _36589_;
  wire _36590_;
  wire _36591_;
  wire _36592_;
  wire _36593_;
  wire _36594_;
  wire _36595_;
  wire _36596_;
  wire _36597_;
  wire _36598_;
  wire _36599_;
  wire _36600_;
  wire _36601_;
  wire _36602_;
  wire _36603_;
  wire _36604_;
  wire _36605_;
  wire _36606_;
  wire _36607_;
  wire _36608_;
  wire _36609_;
  wire _36610_;
  wire _36611_;
  wire _36612_;
  wire _36613_;
  wire _36614_;
  wire _36615_;
  wire _36616_;
  wire _36617_;
  wire _36618_;
  wire _36619_;
  wire _36620_;
  wire _36621_;
  wire _36622_;
  wire _36623_;
  wire _36624_;
  wire _36625_;
  wire _36626_;
  wire _36627_;
  wire _36628_;
  wire _36629_;
  wire _36630_;
  wire _36631_;
  wire _36632_;
  wire _36633_;
  wire _36634_;
  wire _36635_;
  wire _36636_;
  wire _36637_;
  wire _36638_;
  wire _36639_;
  wire _36640_;
  wire _36641_;
  wire _36642_;
  wire _36643_;
  wire _36644_;
  wire _36645_;
  wire _36646_;
  wire _36647_;
  wire _36648_;
  wire _36649_;
  wire _36650_;
  wire _36651_;
  wire _36652_;
  wire _36653_;
  wire _36654_;
  wire _36655_;
  wire _36656_;
  wire _36657_;
  wire _36658_;
  wire _36659_;
  wire _36660_;
  wire _36661_;
  wire _36662_;
  wire _36663_;
  wire _36664_;
  wire _36665_;
  wire _36666_;
  wire _36667_;
  wire _36668_;
  wire _36669_;
  wire _36670_;
  wire _36671_;
  wire _36672_;
  wire _36673_;
  wire _36674_;
  wire _36675_;
  wire _36676_;
  wire _36677_;
  wire _36678_;
  wire _36679_;
  wire _36680_;
  wire _36681_;
  wire _36682_;
  wire _36683_;
  wire _36684_;
  wire _36685_;
  wire _36686_;
  wire _36687_;
  wire _36688_;
  wire _36689_;
  wire _36690_;
  wire _36691_;
  wire _36692_;
  wire _36693_;
  wire _36694_;
  wire _36695_;
  wire _36696_;
  wire _36697_;
  wire _36698_;
  wire _36699_;
  wire _36700_;
  wire _36701_;
  wire _36702_;
  wire _36703_;
  wire _36704_;
  wire _36705_;
  wire _36706_;
  wire _36707_;
  wire _36708_;
  wire _36709_;
  wire _36710_;
  wire _36711_;
  wire _36712_;
  wire _36713_;
  wire _36714_;
  wire _36715_;
  wire _36716_;
  wire _36717_;
  wire _36718_;
  wire _36719_;
  wire _36720_;
  wire _36721_;
  wire _36722_;
  wire _36723_;
  wire _36724_;
  wire _36725_;
  wire _36726_;
  wire _36727_;
  wire _36728_;
  wire _36729_;
  wire _36730_;
  wire _36731_;
  wire _36732_;
  wire _36733_;
  wire _36734_;
  wire _36735_;
  wire _36736_;
  wire _36737_;
  wire _36738_;
  wire _36739_;
  wire _36740_;
  wire _36741_;
  wire _36742_;
  wire _36743_;
  wire _36744_;
  wire _36745_;
  wire _36746_;
  wire _36747_;
  wire _36748_;
  wire _36749_;
  wire _36750_;
  wire _36751_;
  wire _36752_;
  wire _36753_;
  wire _36754_;
  wire _36755_;
  wire _36756_;
  wire _36757_;
  wire _36758_;
  wire _36759_;
  wire _36760_;
  wire _36761_;
  wire _36762_;
  wire _36763_;
  wire _36764_;
  wire _36765_;
  wire _36766_;
  wire _36767_;
  wire _36768_;
  wire _36769_;
  wire _36770_;
  wire _36771_;
  wire _36772_;
  wire _36773_;
  wire _36774_;
  wire _36775_;
  wire _36776_;
  wire _36777_;
  wire _36778_;
  wire _36779_;
  wire _36780_;
  wire _36781_;
  wire _36782_;
  wire _36783_;
  wire _36784_;
  wire _36785_;
  wire _36786_;
  wire _36787_;
  wire _36788_;
  wire _36789_;
  wire _36790_;
  wire _36791_;
  wire _36792_;
  wire _36793_;
  wire _36794_;
  wire _36795_;
  wire _36796_;
  wire _36797_;
  wire _36798_;
  wire _36799_;
  wire _36800_;
  wire _36801_;
  wire _36802_;
  wire _36803_;
  wire _36804_;
  wire _36805_;
  wire _36806_;
  wire _36807_;
  wire _36808_;
  wire _36809_;
  wire _36810_;
  wire _36811_;
  wire _36812_;
  wire _36813_;
  wire _36814_;
  wire _36815_;
  wire _36816_;
  wire _36817_;
  wire _36818_;
  wire _36819_;
  wire _36820_;
  wire _36821_;
  wire _36822_;
  wire _36823_;
  wire _36824_;
  wire _36825_;
  wire _36826_;
  wire _36827_;
  wire _36828_;
  wire _36829_;
  wire _36830_;
  wire _36831_;
  wire _36832_;
  wire _36833_;
  wire _36834_;
  wire _36835_;
  wire _36836_;
  wire _36837_;
  wire _36838_;
  wire _36839_;
  wire _36840_;
  wire _36841_;
  wire _36842_;
  wire _36843_;
  wire _36844_;
  wire _36845_;
  wire _36846_;
  wire _36847_;
  wire _36848_;
  wire _36849_;
  wire _36850_;
  wire _36851_;
  wire _36852_;
  wire _36853_;
  wire _36854_;
  wire _36855_;
  wire _36856_;
  wire _36857_;
  wire _36858_;
  wire _36859_;
  wire _36860_;
  wire _36861_;
  wire _36862_;
  wire _36863_;
  wire _36864_;
  wire _36865_;
  wire _36866_;
  wire _36867_;
  wire _36868_;
  wire _36869_;
  wire _36870_;
  wire _36871_;
  wire _36872_;
  wire _36873_;
  wire _36874_;
  wire _36875_;
  wire _36876_;
  wire _36877_;
  wire _36878_;
  wire _36879_;
  wire _36880_;
  wire _36881_;
  wire _36882_;
  wire _36883_;
  wire _36884_;
  wire _36885_;
  wire _36886_;
  wire _36887_;
  wire _36888_;
  wire _36889_;
  wire _36890_;
  wire _36891_;
  wire _36892_;
  wire _36893_;
  wire _36894_;
  wire _36895_;
  wire _36896_;
  wire _36897_;
  wire _36898_;
  wire _36899_;
  wire _36900_;
  wire _36901_;
  wire _36902_;
  wire _36903_;
  wire _36904_;
  wire _36905_;
  wire _36906_;
  wire _36907_;
  wire _36908_;
  wire _36909_;
  wire _36910_;
  wire _36911_;
  wire _36912_;
  wire _36913_;
  wire _36914_;
  wire _36915_;
  wire _36916_;
  wire _36917_;
  wire _36918_;
  wire _36919_;
  wire _36920_;
  wire _36921_;
  wire _36922_;
  wire _36923_;
  wire _36924_;
  wire _36925_;
  wire _36926_;
  wire _36927_;
  wire _36928_;
  wire _36929_;
  wire _36930_;
  wire _36931_;
  wire _36932_;
  wire _36933_;
  wire _36934_;
  wire _36935_;
  wire _36936_;
  wire _36937_;
  wire _36938_;
  wire _36939_;
  wire _36940_;
  wire _36941_;
  wire _36942_;
  wire _36943_;
  wire _36944_;
  wire _36945_;
  wire _36946_;
  wire _36947_;
  wire _36948_;
  wire _36949_;
  wire _36950_;
  wire _36951_;
  wire _36952_;
  wire _36953_;
  wire _36954_;
  wire _36955_;
  wire _36956_;
  wire _36957_;
  wire _36958_;
  wire _36959_;
  wire _36960_;
  wire _36961_;
  wire _36962_;
  wire _36963_;
  wire _36964_;
  wire _36965_;
  wire _36966_;
  wire _36967_;
  wire _36968_;
  wire _36969_;
  wire _36970_;
  wire _36971_;
  wire _36972_;
  wire _36973_;
  wire _36974_;
  wire _36975_;
  wire _36976_;
  wire _36977_;
  wire _36978_;
  wire _36979_;
  wire _36980_;
  wire _36981_;
  wire _36982_;
  wire _36983_;
  wire _36984_;
  wire _36985_;
  wire _36986_;
  wire _36987_;
  wire _36988_;
  wire _36989_;
  wire _36990_;
  wire _36991_;
  wire _36992_;
  wire _36993_;
  wire _36994_;
  wire _36995_;
  wire _36996_;
  wire _36997_;
  wire _36998_;
  wire _36999_;
  wire _37000_;
  wire _37001_;
  wire _37002_;
  wire _37003_;
  wire _37004_;
  wire _37005_;
  wire _37006_;
  wire _37007_;
  wire _37008_;
  wire _37009_;
  wire _37010_;
  wire _37011_;
  wire _37012_;
  wire _37013_;
  wire _37014_;
  wire _37015_;
  wire _37016_;
  wire _37017_;
  wire _37018_;
  wire _37019_;
  wire _37020_;
  wire _37021_;
  wire _37022_;
  wire _37023_;
  wire _37024_;
  wire _37025_;
  wire _37026_;
  wire _37027_;
  wire _37028_;
  wire _37029_;
  wire _37030_;
  wire _37031_;
  wire _37032_;
  wire _37033_;
  wire _37034_;
  wire _37035_;
  wire _37036_;
  wire _37037_;
  wire _37038_;
  wire _37039_;
  wire _37040_;
  wire _37041_;
  wire _37042_;
  wire _37043_;
  wire _37044_;
  wire _37045_;
  wire _37046_;
  wire _37047_;
  wire _37048_;
  wire _37049_;
  wire _37050_;
  wire _37051_;
  wire _37052_;
  wire _37053_;
  wire _37054_;
  wire _37055_;
  wire _37056_;
  wire _37057_;
  wire _37058_;
  wire _37059_;
  wire _37060_;
  wire _37061_;
  wire _37062_;
  wire _37063_;
  wire _37064_;
  wire _37065_;
  wire _37066_;
  wire _37067_;
  wire _37068_;
  wire _37069_;
  wire _37070_;
  wire _37071_;
  wire _37072_;
  wire _37073_;
  wire _37074_;
  wire _37075_;
  wire _37076_;
  wire _37077_;
  wire _37078_;
  wire _37079_;
  wire _37080_;
  wire _37081_;
  wire _37082_;
  wire _37083_;
  wire _37084_;
  wire _37085_;
  wire _37086_;
  wire _37087_;
  wire _37088_;
  wire _37089_;
  wire _37090_;
  wire _37091_;
  wire _37092_;
  wire _37093_;
  wire _37094_;
  wire _37095_;
  wire _37096_;
  wire _37097_;
  wire _37098_;
  wire _37099_;
  wire _37100_;
  wire _37101_;
  wire _37102_;
  wire _37103_;
  wire _37104_;
  wire _37105_;
  wire _37106_;
  wire _37107_;
  wire _37108_;
  wire _37109_;
  wire _37110_;
  wire _37111_;
  wire _37112_;
  wire _37113_;
  wire _37114_;
  wire _37115_;
  wire _37116_;
  wire _37117_;
  wire _37118_;
  wire _37119_;
  wire _37120_;
  wire _37121_;
  wire _37122_;
  wire _37123_;
  wire _37124_;
  wire _37125_;
  wire _37126_;
  wire _37127_;
  wire _37128_;
  wire _37129_;
  wire _37130_;
  wire _37131_;
  wire _37132_;
  wire _37133_;
  wire _37134_;
  wire _37135_;
  wire _37136_;
  wire _37137_;
  wire _37138_;
  wire _37139_;
  wire _37140_;
  wire _37141_;
  wire _37142_;
  wire _37143_;
  wire _37144_;
  wire _37145_;
  wire _37146_;
  wire _37147_;
  wire _37148_;
  wire _37149_;
  wire _37150_;
  wire _37151_;
  wire _37152_;
  wire _37153_;
  wire _37154_;
  wire _37155_;
  wire _37156_;
  wire _37157_;
  wire _37158_;
  wire _37159_;
  wire _37160_;
  wire _37161_;
  wire _37162_;
  wire _37163_;
  wire _37164_;
  wire _37165_;
  wire _37166_;
  wire _37167_;
  wire _37168_;
  wire _37169_;
  wire _37170_;
  wire _37171_;
  wire _37172_;
  wire _37173_;
  wire _37174_;
  wire _37175_;
  wire _37176_;
  wire _37177_;
  wire _37178_;
  wire _37179_;
  wire _37180_;
  wire _37181_;
  wire _37182_;
  wire _37183_;
  wire _37184_;
  wire _37185_;
  wire _37186_;
  wire _37187_;
  wire _37188_;
  wire _37189_;
  wire _37190_;
  wire _37191_;
  wire _37192_;
  wire _37193_;
  wire _37194_;
  wire _37195_;
  wire _37196_;
  wire _37197_;
  wire _37198_;
  wire _37199_;
  wire _37200_;
  wire _37201_;
  wire _37202_;
  wire _37203_;
  wire _37204_;
  wire _37205_;
  wire _37206_;
  wire _37207_;
  wire _37208_;
  wire _37209_;
  wire _37210_;
  wire _37211_;
  wire _37212_;
  wire _37213_;
  wire _37214_;
  wire _37215_;
  wire _37216_;
  wire _37217_;
  wire _37218_;
  wire _37219_;
  wire _37220_;
  wire _37221_;
  wire _37222_;
  wire _37223_;
  wire _37224_;
  wire _37225_;
  wire _37226_;
  wire _37227_;
  wire _37228_;
  wire _37229_;
  wire _37230_;
  wire _37231_;
  wire _37232_;
  wire _37233_;
  wire _37234_;
  wire _37235_;
  wire _37236_;
  wire _37237_;
  wire _37238_;
  wire _37239_;
  wire _37240_;
  wire _37241_;
  wire _37242_;
  wire _37243_;
  wire _37244_;
  wire _37245_;
  wire _37246_;
  wire _37247_;
  wire _37248_;
  wire _37249_;
  wire _37250_;
  wire _37251_;
  wire _37252_;
  wire _37253_;
  wire _37254_;
  wire _37255_;
  wire _37256_;
  wire _37257_;
  wire _37258_;
  wire _37259_;
  wire _37260_;
  wire _37261_;
  wire _37262_;
  wire _37263_;
  wire _37264_;
  wire _37265_;
  wire _37266_;
  wire _37267_;
  wire _37268_;
  wire _37269_;
  wire _37270_;
  wire _37271_;
  wire _37272_;
  wire _37273_;
  wire _37274_;
  wire _37275_;
  wire _37276_;
  wire _37277_;
  wire _37278_;
  wire _37279_;
  wire _37280_;
  wire _37281_;
  wire _37282_;
  wire _37283_;
  wire _37284_;
  wire _37285_;
  wire _37286_;
  wire _37287_;
  wire _37288_;
  wire _37289_;
  wire _37290_;
  wire _37291_;
  wire _37292_;
  wire _37293_;
  wire _37294_;
  wire _37295_;
  wire _37296_;
  wire _37297_;
  wire _37298_;
  wire _37299_;
  wire _37300_;
  wire _37301_;
  wire _37302_;
  wire _37303_;
  wire _37304_;
  wire _37305_;
  wire _37306_;
  wire _37307_;
  wire _37308_;
  wire _37309_;
  wire _37310_;
  wire _37311_;
  wire _37312_;
  wire _37313_;
  wire _37314_;
  wire _37315_;
  wire _37316_;
  wire _37317_;
  wire _37318_;
  wire _37319_;
  wire _37320_;
  wire _37321_;
  wire _37322_;
  wire _37323_;
  wire _37324_;
  wire _37325_;
  wire _37326_;
  wire _37327_;
  wire _37328_;
  wire _37329_;
  wire _37330_;
  wire _37331_;
  wire _37332_;
  wire _37333_;
  wire _37334_;
  wire _37335_;
  wire _37336_;
  wire _37337_;
  wire _37338_;
  wire _37339_;
  wire _37340_;
  wire _37341_;
  wire _37342_;
  wire _37343_;
  wire _37344_;
  wire _37345_;
  wire _37346_;
  wire _37347_;
  wire _37348_;
  wire _37349_;
  wire _37350_;
  wire _37351_;
  wire _37352_;
  wire _37353_;
  wire _37354_;
  wire _37355_;
  wire _37356_;
  wire _37357_;
  wire _37358_;
  wire _37359_;
  wire _37360_;
  wire _37361_;
  wire _37362_;
  wire _37363_;
  wire _37364_;
  wire _37365_;
  wire _37366_;
  wire _37367_;
  wire _37368_;
  wire _37369_;
  wire _37370_;
  wire _37371_;
  wire _37372_;
  wire _37373_;
  wire _37374_;
  wire _37375_;
  wire _37376_;
  wire _37377_;
  wire _37378_;
  wire _37379_;
  wire _37380_;
  wire _37381_;
  wire _37382_;
  wire _37383_;
  wire _37384_;
  wire _37385_;
  wire _37386_;
  wire _37387_;
  wire _37388_;
  wire _37389_;
  wire _37390_;
  wire _37391_;
  wire _37392_;
  wire _37393_;
  wire _37394_;
  wire _37395_;
  wire _37396_;
  wire _37397_;
  wire _37398_;
  wire _37399_;
  wire _37400_;
  wire _37401_;
  wire _37402_;
  wire _37403_;
  wire _37404_;
  wire _37405_;
  wire _37406_;
  wire _37407_;
  wire _37408_;
  wire _37409_;
  wire _37410_;
  wire _37411_;
  wire _37412_;
  wire _37413_;
  wire _37414_;
  wire _37415_;
  wire _37416_;
  wire _37417_;
  wire _37418_;
  wire _37419_;
  wire _37420_;
  wire _37421_;
  wire _37422_;
  wire _37423_;
  wire _37424_;
  wire _37425_;
  wire _37426_;
  wire _37427_;
  wire _37428_;
  wire _37429_;
  wire _37430_;
  wire _37431_;
  wire _37432_;
  wire _37433_;
  wire _37434_;
  wire _37435_;
  wire _37436_;
  wire _37437_;
  wire _37438_;
  wire _37439_;
  wire _37440_;
  wire _37441_;
  wire _37442_;
  wire _37443_;
  wire _37444_;
  wire _37445_;
  wire _37446_;
  wire _37447_;
  wire _37448_;
  wire _37449_;
  wire _37450_;
  wire _37451_;
  wire _37452_;
  wire _37453_;
  wire _37454_;
  wire _37455_;
  wire _37456_;
  wire _37457_;
  wire _37458_;
  wire _37459_;
  wire _37460_;
  wire _37461_;
  wire _37462_;
  wire _37463_;
  wire _37464_;
  wire _37465_;
  wire _37466_;
  wire _37467_;
  wire _37468_;
  wire _37469_;
  wire _37470_;
  wire _37471_;
  wire _37472_;
  wire _37473_;
  wire _37474_;
  wire _37475_;
  wire _37476_;
  wire _37477_;
  wire _37478_;
  wire _37479_;
  wire _37480_;
  wire _37481_;
  wire _37482_;
  wire _37483_;
  wire _37484_;
  wire _37485_;
  wire _37486_;
  wire _37487_;
  wire _37488_;
  wire _37489_;
  wire _37490_;
  wire _37491_;
  wire _37492_;
  wire _37493_;
  wire _37494_;
  wire _37495_;
  wire _37496_;
  wire _37497_;
  wire _37498_;
  wire _37499_;
  wire _37500_;
  wire _37501_;
  wire _37502_;
  wire _37503_;
  wire _37504_;
  wire _37505_;
  wire _37506_;
  wire _37507_;
  wire _37508_;
  wire _37509_;
  wire _37510_;
  wire _37511_;
  wire _37512_;
  wire _37513_;
  wire _37514_;
  wire _37515_;
  wire _37516_;
  wire _37517_;
  wire _37518_;
  wire _37519_;
  wire _37520_;
  wire _37521_;
  wire _37522_;
  wire _37523_;
  wire _37524_;
  wire _37525_;
  wire _37526_;
  wire _37527_;
  wire _37528_;
  wire _37529_;
  wire _37530_;
  wire _37531_;
  wire _37532_;
  wire _37533_;
  wire _37534_;
  wire _37535_;
  wire _37536_;
  wire _37537_;
  wire _37538_;
  wire _37539_;
  wire _37540_;
  wire _37541_;
  wire _37542_;
  wire _37543_;
  wire _37544_;
  wire _37545_;
  wire _37546_;
  wire _37547_;
  wire _37548_;
  wire _37549_;
  wire _37550_;
  wire _37551_;
  wire _37552_;
  wire _37553_;
  wire _37554_;
  wire _37555_;
  wire _37556_;
  wire _37557_;
  wire _37558_;
  wire _37559_;
  wire _37560_;
  wire _37561_;
  wire _37562_;
  wire _37563_;
  wire _37564_;
  wire _37565_;
  wire _37566_;
  wire _37567_;
  wire _37568_;
  wire _37569_;
  wire _37570_;
  wire _37571_;
  wire _37572_;
  wire _37573_;
  wire _37574_;
  wire _37575_;
  wire _37576_;
  wire _37577_;
  wire _37578_;
  wire _37579_;
  wire _37580_;
  wire _37581_;
  wire _37582_;
  wire _37583_;
  wire _37584_;
  wire _37585_;
  wire _37586_;
  wire _37587_;
  wire _37588_;
  wire _37589_;
  wire _37590_;
  wire _37591_;
  wire _37592_;
  wire _37593_;
  wire _37594_;
  wire _37595_;
  wire _37596_;
  wire _37597_;
  wire _37598_;
  wire _37599_;
  wire _37600_;
  wire _37601_;
  wire _37602_;
  wire _37603_;
  wire _37604_;
  wire _37605_;
  wire _37606_;
  wire _37607_;
  wire _37608_;
  wire _37609_;
  wire _37610_;
  wire _37611_;
  wire _37612_;
  wire _37613_;
  wire _37614_;
  wire _37615_;
  wire _37616_;
  wire _37617_;
  wire _37618_;
  wire _37619_;
  wire _37620_;
  wire _37621_;
  wire _37622_;
  wire _37623_;
  wire _37624_;
  wire _37625_;
  wire _37626_;
  wire _37627_;
  wire _37628_;
  wire _37629_;
  wire _37630_;
  wire _37631_;
  wire _37632_;
  wire _37633_;
  wire _37634_;
  wire _37635_;
  wire _37636_;
  wire _37637_;
  wire _37638_;
  wire _37639_;
  wire _37640_;
  wire _37641_;
  wire _37642_;
  wire _37643_;
  wire _37644_;
  wire _37645_;
  wire _37646_;
  wire _37647_;
  wire _37648_;
  wire _37649_;
  wire _37650_;
  wire _37651_;
  wire _37652_;
  wire _37653_;
  wire _37654_;
  wire _37655_;
  wire _37656_;
  wire _37657_;
  wire _37658_;
  wire _37659_;
  wire _37660_;
  wire _37661_;
  wire _37662_;
  wire _37663_;
  wire _37664_;
  wire _37665_;
  wire _37666_;
  wire _37667_;
  wire _37668_;
  wire _37669_;
  wire _37670_;
  wire _37671_;
  wire _37672_;
  wire _37673_;
  wire _37674_;
  wire _37675_;
  wire _37676_;
  wire _37677_;
  wire _37678_;
  wire _37679_;
  wire _37680_;
  wire _37681_;
  wire _37682_;
  wire _37683_;
  wire _37684_;
  wire _37685_;
  wire _37686_;
  wire _37687_;
  wire _37688_;
  wire _37689_;
  wire _37690_;
  wire _37691_;
  wire _37692_;
  wire _37693_;
  wire _37694_;
  wire _37695_;
  wire _37696_;
  wire _37697_;
  wire _37698_;
  wire _37699_;
  wire _37700_;
  wire _37701_;
  wire _37702_;
  wire _37703_;
  wire _37704_;
  wire _37705_;
  wire _37706_;
  wire _37707_;
  wire _37708_;
  wire _37709_;
  wire _37710_;
  wire _37711_;
  wire _37712_;
  wire _37713_;
  wire _37714_;
  wire _37715_;
  wire _37716_;
  wire _37717_;
  wire _37718_;
  wire _37719_;
  wire _37720_;
  wire _37721_;
  wire _37722_;
  wire _37723_;
  wire _37724_;
  wire _37725_;
  wire _37726_;
  wire _37727_;
  wire _37728_;
  wire _37729_;
  wire _37730_;
  wire _37731_;
  wire _37732_;
  wire _37733_;
  wire _37734_;
  wire _37735_;
  wire _37736_;
  wire _37737_;
  wire _37738_;
  wire _37739_;
  wire _37740_;
  wire _37741_;
  wire _37742_;
  wire _37743_;
  wire _37744_;
  wire _37745_;
  wire _37746_;
  wire _37747_;
  wire _37748_;
  wire _37749_;
  wire _37750_;
  wire _37751_;
  wire _37752_;
  wire _37753_;
  wire _37754_;
  wire _37755_;
  wire _37756_;
  wire _37757_;
  wire _37758_;
  wire _37759_;
  wire _37760_;
  wire _37761_;
  wire _37762_;
  wire _37763_;
  wire _37764_;
  wire _37765_;
  wire _37766_;
  wire _37767_;
  wire _37768_;
  wire _37769_;
  wire _37770_;
  wire _37771_;
  wire _37772_;
  wire _37773_;
  wire _37774_;
  wire _37775_;
  wire _37776_;
  wire _37777_;
  wire _37778_;
  wire _37779_;
  wire _37780_;
  wire _37781_;
  wire _37782_;
  wire _37783_;
  wire _37784_;
  wire _37785_;
  wire _37786_;
  wire _37787_;
  wire _37788_;
  wire _37789_;
  wire _37790_;
  wire _37791_;
  wire _37792_;
  wire _37793_;
  wire _37794_;
  wire _37795_;
  wire _37796_;
  wire _37797_;
  wire _37798_;
  wire _37799_;
  wire _37800_;
  wire _37801_;
  wire _37802_;
  wire _37803_;
  wire _37804_;
  wire _37805_;
  wire _37806_;
  wire _37807_;
  wire _37808_;
  wire _37809_;
  wire _37810_;
  wire _37811_;
  wire _37812_;
  wire _37813_;
  wire _37814_;
  wire _37815_;
  wire _37816_;
  wire _37817_;
  wire _37818_;
  wire _37819_;
  wire _37820_;
  wire _37821_;
  wire _37822_;
  wire _37823_;
  wire _37824_;
  wire _37825_;
  wire _37826_;
  wire _37827_;
  wire _37828_;
  wire _37829_;
  wire _37830_;
  wire _37831_;
  wire _37832_;
  wire _37833_;
  wire _37834_;
  wire _37835_;
  wire _37836_;
  wire _37837_;
  wire _37838_;
  wire _37839_;
  wire _37840_;
  wire _37841_;
  wire _37842_;
  wire _37843_;
  wire _37844_;
  wire _37845_;
  wire _37846_;
  wire _37847_;
  wire _37848_;
  wire _37849_;
  wire _37850_;
  wire _37851_;
  wire _37852_;
  wire _37853_;
  wire _37854_;
  wire _37855_;
  wire _37856_;
  wire _37857_;
  wire _37858_;
  wire _37859_;
  wire _37860_;
  wire _37861_;
  wire _37862_;
  wire _37863_;
  wire _37864_;
  wire _37865_;
  wire _37866_;
  wire _37867_;
  wire _37868_;
  wire _37869_;
  wire _37870_;
  wire _37871_;
  wire _37872_;
  wire _37873_;
  wire _37874_;
  wire _37875_;
  wire _37876_;
  wire _37877_;
  wire _37878_;
  wire _37879_;
  wire _37880_;
  wire _37881_;
  wire _37882_;
  wire _37883_;
  wire _37884_;
  wire _37885_;
  wire _37886_;
  wire _37887_;
  wire _37888_;
  wire _37889_;
  wire _37890_;
  wire _37891_;
  wire _37892_;
  wire _37893_;
  wire _37894_;
  wire _37895_;
  wire _37896_;
  wire _37897_;
  wire _37898_;
  wire _37899_;
  wire _37900_;
  wire _37901_;
  wire _37902_;
  wire _37903_;
  wire _37904_;
  wire _37905_;
  wire _37906_;
  wire _37907_;
  wire _37908_;
  wire _37909_;
  wire _37910_;
  wire _37911_;
  wire _37912_;
  wire _37913_;
  wire _37914_;
  wire _37915_;
  wire _37916_;
  wire _37917_;
  wire _37918_;
  wire _37919_;
  wire _37920_;
  wire _37921_;
  wire _37922_;
  wire _37923_;
  wire _37924_;
  wire _37925_;
  wire _37926_;
  wire _37927_;
  wire _37928_;
  wire _37929_;
  wire _37930_;
  wire _37931_;
  wire _37932_;
  wire _37933_;
  wire _37934_;
  wire _37935_;
  wire _37936_;
  wire _37937_;
  wire _37938_;
  wire _37939_;
  wire _37940_;
  wire _37941_;
  wire _37942_;
  wire _37943_;
  wire _37944_;
  wire _37945_;
  wire _37946_;
  wire _37947_;
  wire _37948_;
  wire _37949_;
  wire _37950_;
  wire _37951_;
  wire _37952_;
  wire _37953_;
  wire _37954_;
  wire _37955_;
  wire _37956_;
  wire _37957_;
  wire _37958_;
  wire _37959_;
  wire _37960_;
  wire _37961_;
  wire _37962_;
  wire _37963_;
  wire _37964_;
  wire _37965_;
  wire _37966_;
  wire _37967_;
  wire _37968_;
  wire _37969_;
  wire _37970_;
  wire _37971_;
  wire _37972_;
  wire _37973_;
  wire _37974_;
  wire _37975_;
  wire _37976_;
  wire _37977_;
  wire _37978_;
  wire _37979_;
  wire _37980_;
  wire _37981_;
  wire _37982_;
  wire _37983_;
  wire _37984_;
  wire _37985_;
  wire _37986_;
  wire _37987_;
  wire _37988_;
  wire _37989_;
  wire _37990_;
  wire _37991_;
  wire _37992_;
  wire _37993_;
  wire _37994_;
  wire _37995_;
  wire _37996_;
  wire _37997_;
  wire _37998_;
  wire _37999_;
  wire _38000_;
  wire _38001_;
  wire _38002_;
  wire _38003_;
  wire _38004_;
  wire _38005_;
  wire _38006_;
  wire _38007_;
  wire _38008_;
  wire _38009_;
  wire _38010_;
  wire _38011_;
  wire _38012_;
  wire _38013_;
  wire _38014_;
  wire _38015_;
  wire _38016_;
  wire _38017_;
  wire _38018_;
  wire _38019_;
  wire _38020_;
  wire _38021_;
  wire _38022_;
  wire _38023_;
  wire _38024_;
  wire _38025_;
  wire _38026_;
  wire _38027_;
  wire _38028_;
  wire _38029_;
  wire _38030_;
  wire _38031_;
  wire _38032_;
  wire _38033_;
  wire _38034_;
  wire _38035_;
  wire _38036_;
  wire _38037_;
  wire _38038_;
  wire _38039_;
  wire _38040_;
  wire _38041_;
  wire _38042_;
  wire _38043_;
  wire _38044_;
  wire _38045_;
  wire _38046_;
  wire _38047_;
  wire _38048_;
  wire _38049_;
  wire _38050_;
  wire _38051_;
  wire _38052_;
  wire _38053_;
  wire _38054_;
  wire _38055_;
  wire _38056_;
  wire _38057_;
  wire _38058_;
  wire _38059_;
  wire _38060_;
  wire _38061_;
  wire _38062_;
  wire _38063_;
  wire _38064_;
  wire _38065_;
  wire _38066_;
  wire _38067_;
  wire _38068_;
  wire _38069_;
  wire _38070_;
  wire _38071_;
  wire _38072_;
  wire _38073_;
  wire _38074_;
  wire _38075_;
  wire _38076_;
  wire _38077_;
  wire _38078_;
  wire _38079_;
  wire _38080_;
  wire _38081_;
  wire _38082_;
  wire _38083_;
  wire _38084_;
  wire _38085_;
  wire _38086_;
  wire _38087_;
  wire _38088_;
  wire _38089_;
  wire _38090_;
  wire _38091_;
  wire _38092_;
  wire _38093_;
  wire _38094_;
  wire _38095_;
  wire _38096_;
  wire _38097_;
  wire _38098_;
  wire _38099_;
  wire _38100_;
  wire _38101_;
  wire _38102_;
  wire _38103_;
  wire _38104_;
  wire _38105_;
  wire _38106_;
  wire _38107_;
  wire _38108_;
  wire _38109_;
  wire _38110_;
  wire _38111_;
  wire _38112_;
  wire _38113_;
  wire _38114_;
  wire _38115_;
  wire _38116_;
  wire _38117_;
  wire _38118_;
  wire _38119_;
  wire _38120_;
  wire _38121_;
  wire _38122_;
  wire _38123_;
  wire _38124_;
  wire _38125_;
  wire _38126_;
  wire _38127_;
  wire _38128_;
  wire _38129_;
  wire _38130_;
  wire _38131_;
  wire _38132_;
  wire _38133_;
  wire _38134_;
  wire _38135_;
  wire _38136_;
  wire _38137_;
  wire _38138_;
  wire _38139_;
  wire _38140_;
  wire _38141_;
  wire _38142_;
  wire _38143_;
  wire _38144_;
  wire _38145_;
  wire _38146_;
  wire _38147_;
  wire _38148_;
  wire _38149_;
  wire _38150_;
  wire _38151_;
  wire _38152_;
  wire _38153_;
  wire _38154_;
  wire _38155_;
  wire _38156_;
  wire _38157_;
  wire _38158_;
  wire _38159_;
  wire _38160_;
  wire _38161_;
  wire _38162_;
  wire _38163_;
  wire _38164_;
  wire _38165_;
  wire _38166_;
  wire _38167_;
  wire _38168_;
  wire _38169_;
  wire _38170_;
  wire _38171_;
  wire _38172_;
  wire _38173_;
  wire _38174_;
  wire _38175_;
  wire _38176_;
  wire _38177_;
  wire _38178_;
  wire _38179_;
  wire _38180_;
  wire _38181_;
  wire _38182_;
  wire _38183_;
  wire _38184_;
  wire _38185_;
  wire _38186_;
  wire _38187_;
  wire _38188_;
  wire _38189_;
  wire _38190_;
  wire _38191_;
  wire _38192_;
  wire _38193_;
  wire _38194_;
  wire _38195_;
  wire _38196_;
  wire _38197_;
  wire _38198_;
  wire _38199_;
  wire _38200_;
  wire _38201_;
  wire _38202_;
  wire _38203_;
  wire _38204_;
  wire _38205_;
  wire _38206_;
  wire _38207_;
  wire _38208_;
  wire _38209_;
  wire _38210_;
  wire _38211_;
  wire _38212_;
  wire _38213_;
  wire _38214_;
  wire _38215_;
  wire _38216_;
  wire _38217_;
  wire _38218_;
  wire _38219_;
  wire _38220_;
  wire _38221_;
  wire _38222_;
  wire _38223_;
  wire _38224_;
  wire _38225_;
  wire _38226_;
  wire _38227_;
  wire _38228_;
  wire _38229_;
  wire _38230_;
  wire _38231_;
  wire _38232_;
  wire _38233_;
  wire _38234_;
  wire _38235_;
  wire _38236_;
  wire _38237_;
  wire _38238_;
  wire _38239_;
  wire _38240_;
  wire _38241_;
  wire _38242_;
  wire _38243_;
  wire _38244_;
  wire _38245_;
  wire _38246_;
  wire _38247_;
  wire _38248_;
  wire _38249_;
  wire _38250_;
  wire _38251_;
  wire _38252_;
  wire _38253_;
  wire _38254_;
  wire _38255_;
  wire _38256_;
  wire _38257_;
  wire _38258_;
  wire _38259_;
  wire _38260_;
  wire _38261_;
  wire _38262_;
  wire _38263_;
  wire _38264_;
  wire _38265_;
  wire _38266_;
  wire _38267_;
  wire _38268_;
  wire _38269_;
  wire _38270_;
  wire _38271_;
  wire _38272_;
  wire _38273_;
  wire _38274_;
  wire _38275_;
  wire _38276_;
  wire _38277_;
  wire _38278_;
  wire _38279_;
  wire _38280_;
  wire _38281_;
  wire _38282_;
  wire _38283_;
  wire _38284_;
  wire _38285_;
  wire _38286_;
  wire _38287_;
  wire _38288_;
  wire _38289_;
  wire _38290_;
  wire _38291_;
  wire _38292_;
  wire _38293_;
  wire _38294_;
  wire _38295_;
  wire _38296_;
  wire _38297_;
  wire _38298_;
  wire _38299_;
  wire _38300_;
  wire _38301_;
  wire _38302_;
  wire _38303_;
  wire _38304_;
  wire _38305_;
  wire _38306_;
  wire _38307_;
  wire _38308_;
  wire _38309_;
  wire _38310_;
  wire _38311_;
  wire _38312_;
  wire _38313_;
  wire _38314_;
  wire _38315_;
  wire _38316_;
  wire _38317_;
  wire _38318_;
  wire _38319_;
  wire _38320_;
  wire _38321_;
  wire _38322_;
  wire _38323_;
  wire _38324_;
  wire _38325_;
  wire _38326_;
  wire _38327_;
  wire _38328_;
  wire _38329_;
  wire _38330_;
  wire _38331_;
  wire _38332_;
  wire _38333_;
  wire _38334_;
  wire _38335_;
  wire _38336_;
  wire _38337_;
  wire _38338_;
  wire _38339_;
  wire _38340_;
  wire _38341_;
  wire _38342_;
  wire _38343_;
  wire _38344_;
  wire _38345_;
  wire _38346_;
  wire _38347_;
  wire _38348_;
  wire _38349_;
  wire _38350_;
  wire _38351_;
  wire _38352_;
  wire _38353_;
  wire _38354_;
  wire _38355_;
  wire _38356_;
  wire _38357_;
  wire _38358_;
  wire _38359_;
  wire _38360_;
  wire _38361_;
  wire _38362_;
  wire _38363_;
  wire _38364_;
  wire _38365_;
  wire _38366_;
  wire _38367_;
  wire _38368_;
  wire _38369_;
  wire _38370_;
  wire _38371_;
  wire _38372_;
  wire _38373_;
  wire _38374_;
  wire _38375_;
  wire _38376_;
  wire _38377_;
  wire _38378_;
  wire _38379_;
  wire _38380_;
  wire _38381_;
  wire _38382_;
  wire _38383_;
  wire _38384_;
  wire _38385_;
  wire _38386_;
  wire _38387_;
  wire _38388_;
  wire _38389_;
  wire _38390_;
  wire _38391_;
  wire _38392_;
  wire _38393_;
  wire _38394_;
  wire _38395_;
  wire _38396_;
  wire _38397_;
  wire _38398_;
  wire _38399_;
  wire _38400_;
  wire _38401_;
  wire _38402_;
  wire _38403_;
  wire _38404_;
  wire _38405_;
  wire _38406_;
  wire _38407_;
  wire _38408_;
  wire _38409_;
  wire _38410_;
  wire _38411_;
  wire _38412_;
  wire _38413_;
  wire _38414_;
  wire _38415_;
  wire _38416_;
  wire _38417_;
  wire _38418_;
  wire _38419_;
  wire _38420_;
  wire _38421_;
  wire _38422_;
  wire _38423_;
  wire _38424_;
  wire _38425_;
  wire _38426_;
  wire _38427_;
  wire _38428_;
  wire _38429_;
  wire _38430_;
  wire _38431_;
  wire _38432_;
  wire _38433_;
  wire _38434_;
  wire _38435_;
  wire _38436_;
  wire _38437_;
  wire _38438_;
  wire _38439_;
  wire _38440_;
  wire _38441_;
  wire _38442_;
  wire _38443_;
  wire _38444_;
  wire _38445_;
  wire _38446_;
  wire _38447_;
  wire _38448_;
  wire _38449_;
  wire _38450_;
  wire _38451_;
  wire _38452_;
  wire _38453_;
  wire _38454_;
  wire _38455_;
  wire _38456_;
  wire _38457_;
  wire _38458_;
  wire _38459_;
  wire _38460_;
  wire _38461_;
  wire _38462_;
  wire _38463_;
  wire _38464_;
  wire _38465_;
  wire _38466_;
  wire _38467_;
  wire _38468_;
  wire _38469_;
  wire _38470_;
  wire _38471_;
  wire _38472_;
  wire _38473_;
  wire _38474_;
  wire _38475_;
  wire _38476_;
  wire _38477_;
  wire _38478_;
  wire _38479_;
  wire _38480_;
  wire _38481_;
  wire _38482_;
  wire _38483_;
  wire _38484_;
  wire _38485_;
  wire _38486_;
  wire _38487_;
  wire _38488_;
  wire _38489_;
  wire _38490_;
  wire _38491_;
  wire _38492_;
  wire _38493_;
  wire _38494_;
  wire _38495_;
  wire _38496_;
  wire _38497_;
  wire _38498_;
  wire _38499_;
  wire _38500_;
  wire _38501_;
  wire _38502_;
  wire _38503_;
  wire _38504_;
  wire _38505_;
  wire _38506_;
  wire _38507_;
  wire _38508_;
  wire _38509_;
  wire _38510_;
  wire _38511_;
  wire _38512_;
  wire _38513_;
  wire _38514_;
  wire _38515_;
  wire _38516_;
  wire _38517_;
  wire _38518_;
  wire _38519_;
  wire _38520_;
  wire _38521_;
  wire _38522_;
  wire _38523_;
  wire _38524_;
  wire _38525_;
  wire _38526_;
  wire _38527_;
  wire _38528_;
  wire _38529_;
  wire _38530_;
  wire _38531_;
  wire _38532_;
  wire _38533_;
  wire _38534_;
  wire _38535_;
  wire _38536_;
  wire _38537_;
  wire _38538_;
  wire _38539_;
  wire _38540_;
  wire _38541_;
  wire _38542_;
  wire _38543_;
  wire _38544_;
  wire _38545_;
  wire _38546_;
  wire _38547_;
  wire _38548_;
  wire _38549_;
  wire _38550_;
  wire _38551_;
  wire _38552_;
  wire _38553_;
  wire _38554_;
  wire _38555_;
  wire _38556_;
  wire _38557_;
  wire _38558_;
  wire _38559_;
  wire _38560_;
  wire _38561_;
  wire _38562_;
  wire _38563_;
  wire _38564_;
  wire _38565_;
  wire _38566_;
  wire _38567_;
  wire _38568_;
  wire _38569_;
  wire _38570_;
  wire _38571_;
  wire _38572_;
  wire _38573_;
  wire _38574_;
  wire _38575_;
  wire _38576_;
  wire _38577_;
  wire _38578_;
  wire _38579_;
  wire _38580_;
  wire _38581_;
  wire _38582_;
  wire _38583_;
  wire _38584_;
  wire _38585_;
  wire _38586_;
  wire _38587_;
  wire _38588_;
  wire _38589_;
  wire _38590_;
  wire _38591_;
  wire _38592_;
  wire _38593_;
  wire _38594_;
  wire _38595_;
  wire _38596_;
  wire _38597_;
  wire _38598_;
  wire _38599_;
  wire _38600_;
  wire _38601_;
  wire _38602_;
  wire _38603_;
  wire _38604_;
  wire _38605_;
  wire _38606_;
  wire _38607_;
  wire _38608_;
  wire _38609_;
  wire _38610_;
  wire _38611_;
  wire _38612_;
  wire _38613_;
  wire _38614_;
  wire _38615_;
  wire _38616_;
  wire _38617_;
  wire _38618_;
  wire _38619_;
  wire _38620_;
  wire _38621_;
  wire _38622_;
  wire _38623_;
  wire _38624_;
  wire _38625_;
  wire _38626_;
  wire _38627_;
  wire _38628_;
  wire _38629_;
  wire _38630_;
  wire _38631_;
  wire _38632_;
  wire _38633_;
  wire _38634_;
  wire _38635_;
  wire _38636_;
  wire _38637_;
  wire _38638_;
  wire _38639_;
  wire _38640_;
  wire _38641_;
  wire _38642_;
  wire _38643_;
  wire _38644_;
  wire _38645_;
  wire _38646_;
  wire _38647_;
  wire _38648_;
  wire _38649_;
  wire _38650_;
  wire _38651_;
  wire _38652_;
  wire _38653_;
  wire _38654_;
  wire _38655_;
  wire _38656_;
  wire _38657_;
  wire _38658_;
  wire _38659_;
  wire _38660_;
  wire _38661_;
  wire _38662_;
  wire _38663_;
  wire _38664_;
  wire _38665_;
  wire _38666_;
  wire _38667_;
  wire _38668_;
  wire _38669_;
  wire _38670_;
  wire _38671_;
  wire _38672_;
  wire _38673_;
  wire _38674_;
  wire _38675_;
  wire _38676_;
  wire _38677_;
  wire _38678_;
  wire _38679_;
  wire _38680_;
  wire _38681_;
  wire _38682_;
  wire _38683_;
  wire _38684_;
  wire _38685_;
  wire _38686_;
  wire _38687_;
  wire _38688_;
  wire _38689_;
  wire _38690_;
  wire _38691_;
  wire _38692_;
  wire _38693_;
  wire _38694_;
  wire _38695_;
  wire _38696_;
  wire _38697_;
  wire _38698_;
  wire _38699_;
  wire _38700_;
  wire _38701_;
  wire _38702_;
  wire _38703_;
  wire _38704_;
  wire _38705_;
  wire _38706_;
  wire _38707_;
  wire _38708_;
  wire _38709_;
  wire _38710_;
  wire _38711_;
  wire _38712_;
  wire _38713_;
  wire _38714_;
  wire _38715_;
  wire _38716_;
  wire _38717_;
  wire _38718_;
  wire _38719_;
  wire _38720_;
  wire _38721_;
  wire _38722_;
  wire _38723_;
  wire _38724_;
  wire _38725_;
  wire _38726_;
  wire _38727_;
  wire _38728_;
  wire _38729_;
  wire _38730_;
  wire _38731_;
  wire _38732_;
  wire _38733_;
  wire _38734_;
  wire _38735_;
  wire _38736_;
  wire _38737_;
  wire _38738_;
  wire _38739_;
  wire _38740_;
  wire _38741_;
  wire _38742_;
  wire _38743_;
  wire _38744_;
  wire _38745_;
  wire _38746_;
  wire _38747_;
  wire _38748_;
  wire _38749_;
  wire _38750_;
  wire _38751_;
  wire _38752_;
  wire _38753_;
  wire _38754_;
  wire _38755_;
  wire _38756_;
  wire _38757_;
  wire _38758_;
  wire _38759_;
  wire _38760_;
  wire _38761_;
  wire _38762_;
  wire _38763_;
  wire _38764_;
  wire _38765_;
  wire _38766_;
  wire _38767_;
  wire _38768_;
  wire _38769_;
  wire _38770_;
  wire _38771_;
  wire _38772_;
  wire _38773_;
  wire _38774_;
  wire _38775_;
  wire _38776_;
  wire _38777_;
  wire _38778_;
  wire _38779_;
  wire _38780_;
  wire _38781_;
  wire _38782_;
  wire _38783_;
  wire _38784_;
  wire _38785_;
  wire _38786_;
  wire _38787_;
  wire _38788_;
  wire _38789_;
  wire _38790_;
  wire _38791_;
  wire _38792_;
  wire _38793_;
  wire _38794_;
  wire _38795_;
  wire _38796_;
  wire _38797_;
  wire _38798_;
  wire _38799_;
  wire _38800_;
  wire _38801_;
  wire _38802_;
  wire _38803_;
  wire _38804_;
  wire _38805_;
  wire _38806_;
  wire _38807_;
  wire _38808_;
  wire _38809_;
  wire _38810_;
  wire _38811_;
  wire _38812_;
  wire _38813_;
  wire _38814_;
  wire _38815_;
  wire _38816_;
  wire _38817_;
  wire _38818_;
  wire _38819_;
  wire _38820_;
  wire _38821_;
  wire _38822_;
  wire _38823_;
  wire _38824_;
  wire _38825_;
  wire _38826_;
  wire _38827_;
  wire _38828_;
  wire _38829_;
  wire _38830_;
  wire _38831_;
  wire _38832_;
  wire _38833_;
  wire _38834_;
  wire _38835_;
  wire _38836_;
  wire _38837_;
  wire _38838_;
  wire _38839_;
  wire _38840_;
  wire _38841_;
  wire _38842_;
  wire _38843_;
  wire _38844_;
  wire _38845_;
  wire _38846_;
  wire _38847_;
  wire _38848_;
  wire _38849_;
  wire _38850_;
  wire _38851_;
  wire _38852_;
  wire _38853_;
  wire _38854_;
  wire _38855_;
  wire _38856_;
  wire _38857_;
  wire _38858_;
  wire _38859_;
  wire _38860_;
  wire _38861_;
  wire _38862_;
  wire _38863_;
  wire _38864_;
  wire _38865_;
  wire _38866_;
  wire _38867_;
  wire _38868_;
  wire _38869_;
  wire _38870_;
  wire _38871_;
  wire _38872_;
  wire _38873_;
  wire _38874_;
  wire _38875_;
  wire _38876_;
  wire _38877_;
  wire _38878_;
  wire _38879_;
  wire _38880_;
  wire _38881_;
  wire _38882_;
  wire _38883_;
  wire _38884_;
  wire _38885_;
  wire _38886_;
  wire _38887_;
  wire _38888_;
  wire _38889_;
  wire _38890_;
  wire _38891_;
  wire _38892_;
  wire _38893_;
  wire _38894_;
  wire _38895_;
  wire _38896_;
  wire _38897_;
  wire _38898_;
  wire _38899_;
  wire _38900_;
  wire _38901_;
  wire _38902_;
  wire _38903_;
  wire _38904_;
  wire _38905_;
  wire _38906_;
  wire _38907_;
  wire _38908_;
  wire _38909_;
  wire _38910_;
  wire _38911_;
  wire _38912_;
  wire _38913_;
  wire _38914_;
  wire _38915_;
  wire _38916_;
  wire _38917_;
  wire _38918_;
  wire _38919_;
  wire _38920_;
  wire _38921_;
  wire _38922_;
  wire _38923_;
  wire _38924_;
  wire _38925_;
  wire _38926_;
  wire _38927_;
  wire _38928_;
  wire _38929_;
  wire _38930_;
  wire _38931_;
  wire _38932_;
  wire _38933_;
  wire _38934_;
  wire _38935_;
  wire _38936_;
  wire _38937_;
  wire _38938_;
  wire _38939_;
  wire _38940_;
  wire _38941_;
  wire _38942_;
  wire _38943_;
  wire _38944_;
  wire _38945_;
  wire _38946_;
  wire _38947_;
  wire _38948_;
  wire _38949_;
  wire _38950_;
  wire _38951_;
  wire _38952_;
  wire _38953_;
  wire _38954_;
  wire _38955_;
  wire _38956_;
  wire _38957_;
  wire _38958_;
  wire _38959_;
  wire _38960_;
  wire _38961_;
  wire _38962_;
  wire _38963_;
  wire _38964_;
  wire _38965_;
  wire _38966_;
  wire _38967_;
  wire _38968_;
  wire _38969_;
  wire _38970_;
  wire _38971_;
  wire _38972_;
  wire _38973_;
  wire _38974_;
  wire _38975_;
  wire _38976_;
  wire _38977_;
  wire _38978_;
  wire _38979_;
  wire _38980_;
  wire _38981_;
  wire _38982_;
  wire _38983_;
  wire _38984_;
  wire _38985_;
  wire _38986_;
  wire _38987_;
  wire _38988_;
  wire _38989_;
  wire _38990_;
  wire _38991_;
  wire _38992_;
  wire _38993_;
  wire _38994_;
  wire _38995_;
  wire _38996_;
  wire _38997_;
  wire _38998_;
  wire _38999_;
  wire _39000_;
  wire _39001_;
  wire _39002_;
  wire _39003_;
  wire _39004_;
  wire _39005_;
  wire _39006_;
  wire _39007_;
  wire _39008_;
  wire _39009_;
  wire _39010_;
  wire _39011_;
  wire _39012_;
  wire _39013_;
  wire _39014_;
  wire _39015_;
  wire _39016_;
  wire _39017_;
  wire _39018_;
  wire _39019_;
  wire _39020_;
  wire _39021_;
  wire _39022_;
  wire _39023_;
  wire _39024_;
  wire _39025_;
  wire _39026_;
  wire _39027_;
  wire _39028_;
  wire _39029_;
  wire _39030_;
  wire _39031_;
  wire _39032_;
  wire _39033_;
  wire _39034_;
  wire _39035_;
  wire _39036_;
  wire _39037_;
  wire _39038_;
  wire _39039_;
  wire _39040_;
  wire _39041_;
  wire _39042_;
  wire _39043_;
  wire _39044_;
  wire _39045_;
  wire _39046_;
  wire _39047_;
  wire _39048_;
  wire _39049_;
  wire _39050_;
  wire _39051_;
  wire _39052_;
  wire _39053_;
  wire _39054_;
  wire _39055_;
  wire _39056_;
  wire _39057_;
  wire _39058_;
  wire _39059_;
  wire _39060_;
  wire _39061_;
  wire _39062_;
  wire _39063_;
  wire _39064_;
  wire _39065_;
  wire _39066_;
  wire _39067_;
  wire _39068_;
  wire _39069_;
  wire _39070_;
  wire _39071_;
  wire _39072_;
  wire _39073_;
  wire _39074_;
  wire _39075_;
  wire _39076_;
  wire _39077_;
  wire _39078_;
  wire _39079_;
  wire _39080_;
  wire _39081_;
  wire _39082_;
  wire _39083_;
  wire _39084_;
  wire _39085_;
  wire _39086_;
  wire _39087_;
  wire _39088_;
  wire _39089_;
  wire _39090_;
  wire _39091_;
  wire _39092_;
  wire _39093_;
  wire _39094_;
  wire _39095_;
  wire _39096_;
  wire _39097_;
  wire _39098_;
  wire _39099_;
  wire _39100_;
  wire _39101_;
  wire _39102_;
  wire _39103_;
  wire _39104_;
  wire _39105_;
  wire _39106_;
  wire _39107_;
  wire _39108_;
  wire _39109_;
  wire _39110_;
  wire _39111_;
  wire _39112_;
  wire _39113_;
  wire _39114_;
  wire _39115_;
  wire _39116_;
  wire _39117_;
  wire _39118_;
  wire _39119_;
  wire _39120_;
  wire _39121_;
  wire _39122_;
  wire _39123_;
  wire _39124_;
  wire _39125_;
  wire _39126_;
  wire _39127_;
  wire _39128_;
  wire _39129_;
  wire _39130_;
  wire _39131_;
  wire _39132_;
  wire _39133_;
  wire _39134_;
  wire _39135_;
  wire _39136_;
  wire _39137_;
  wire _39138_;
  wire _39139_;
  wire _39140_;
  wire _39141_;
  wire _39142_;
  wire _39143_;
  wire _39144_;
  wire _39145_;
  wire _39146_;
  wire _39147_;
  wire _39148_;
  wire _39149_;
  wire _39150_;
  wire _39151_;
  wire _39152_;
  wire _39153_;
  wire _39154_;
  wire _39155_;
  wire _39156_;
  wire _39157_;
  wire _39158_;
  wire _39159_;
  wire _39160_;
  wire _39161_;
  wire _39162_;
  wire _39163_;
  wire _39164_;
  wire _39165_;
  wire _39166_;
  wire _39167_;
  wire _39168_;
  wire _39169_;
  wire _39170_;
  wire _39171_;
  wire _39172_;
  wire _39173_;
  wire _39174_;
  wire _39175_;
  wire _39176_;
  wire _39177_;
  wire _39178_;
  wire _39179_;
  wire _39180_;
  wire _39181_;
  wire _39182_;
  wire _39183_;
  wire _39184_;
  wire _39185_;
  wire _39186_;
  wire _39187_;
  wire _39188_;
  wire _39189_;
  wire _39190_;
  wire _39191_;
  wire _39192_;
  wire _39193_;
  wire _39194_;
  wire _39195_;
  wire _39196_;
  wire _39197_;
  wire _39198_;
  wire _39199_;
  wire _39200_;
  wire _39201_;
  wire _39202_;
  wire _39203_;
  wire _39204_;
  wire _39205_;
  wire _39206_;
  wire _39207_;
  wire _39208_;
  wire _39209_;
  wire _39210_;
  wire _39211_;
  wire _39212_;
  wire _39213_;
  wire _39214_;
  wire _39215_;
  wire _39216_;
  wire _39217_;
  wire _39218_;
  wire _39219_;
  wire _39220_;
  wire _39221_;
  wire _39222_;
  wire _39223_;
  wire _39224_;
  wire _39225_;
  wire _39226_;
  wire _39227_;
  wire _39228_;
  wire _39229_;
  wire _39230_;
  wire _39231_;
  wire _39232_;
  wire _39233_;
  wire _39234_;
  wire _39235_;
  wire _39236_;
  wire _39237_;
  wire _39238_;
  wire _39239_;
  wire _39240_;
  wire _39241_;
  wire _39242_;
  wire _39243_;
  wire _39244_;
  wire _39245_;
  wire _39246_;
  wire _39247_;
  wire _39248_;
  wire _39249_;
  wire _39250_;
  wire _39251_;
  wire _39252_;
  wire _39253_;
  wire _39254_;
  wire _39255_;
  wire _39256_;
  wire _39257_;
  wire _39258_;
  wire _39259_;
  wire _39260_;
  wire _39261_;
  wire _39262_;
  wire _39263_;
  wire _39264_;
  wire _39265_;
  wire _39266_;
  wire _39267_;
  wire _39268_;
  wire _39269_;
  wire _39270_;
  wire _39271_;
  wire _39272_;
  wire _39273_;
  wire _39274_;
  wire _39275_;
  wire _39276_;
  wire _39277_;
  wire _39278_;
  wire _39279_;
  wire _39280_;
  wire _39281_;
  wire _39282_;
  wire _39283_;
  wire _39284_;
  wire _39285_;
  wire _39286_;
  wire _39287_;
  wire _39288_;
  wire _39289_;
  wire _39290_;
  wire _39291_;
  wire _39292_;
  wire _39293_;
  wire _39294_;
  wire _39295_;
  wire _39296_;
  wire _39297_;
  wire _39298_;
  wire _39299_;
  wire _39300_;
  wire _39301_;
  wire _39302_;
  wire _39303_;
  wire _39304_;
  wire _39305_;
  wire _39306_;
  wire _39307_;
  wire _39308_;
  wire _39309_;
  wire _39310_;
  wire _39311_;
  wire _39312_;
  wire _39313_;
  wire _39314_;
  wire _39315_;
  wire _39316_;
  wire _39317_;
  wire _39318_;
  wire _39319_;
  wire _39320_;
  wire _39321_;
  wire _39322_;
  wire _39323_;
  wire _39324_;
  wire _39325_;
  wire _39326_;
  wire _39327_;
  wire _39328_;
  wire _39329_;
  wire _39330_;
  wire _39331_;
  wire _39332_;
  wire _39333_;
  wire _39334_;
  wire _39335_;
  wire _39336_;
  wire _39337_;
  wire _39338_;
  wire _39339_;
  wire _39340_;
  wire _39341_;
  wire _39342_;
  wire _39343_;
  wire _39344_;
  wire _39345_;
  wire _39346_;
  wire _39347_;
  wire _39348_;
  wire _39349_;
  wire _39350_;
  wire _39351_;
  wire _39352_;
  wire _39353_;
  wire _39354_;
  wire _39355_;
  wire _39356_;
  wire _39357_;
  wire _39358_;
  wire _39359_;
  wire _39360_;
  wire _39361_;
  wire _39362_;
  wire _39363_;
  wire _39364_;
  wire _39365_;
  wire _39366_;
  wire _39367_;
  wire _39368_;
  wire _39369_;
  wire _39370_;
  wire _39371_;
  wire _39372_;
  wire _39373_;
  wire _39374_;
  wire _39375_;
  wire _39376_;
  wire _39377_;
  wire _39378_;
  wire _39379_;
  wire _39380_;
  wire _39381_;
  wire _39382_;
  wire _39383_;
  wire _39384_;
  wire _39385_;
  wire _39386_;
  wire _39387_;
  wire _39388_;
  wire _39389_;
  wire _39390_;
  wire _39391_;
  wire _39392_;
  wire _39393_;
  wire _39394_;
  wire _39395_;
  wire _39396_;
  wire _39397_;
  wire _39398_;
  wire _39399_;
  wire _39400_;
  wire _39401_;
  wire _39402_;
  wire _39403_;
  wire _39404_;
  wire _39405_;
  wire _39406_;
  wire _39407_;
  wire _39408_;
  wire _39409_;
  wire _39410_;
  wire _39411_;
  wire _39412_;
  wire _39413_;
  wire _39414_;
  wire _39415_;
  wire _39416_;
  wire _39417_;
  wire _39418_;
  wire _39419_;
  wire _39420_;
  wire _39421_;
  wire _39422_;
  wire _39423_;
  wire _39424_;
  wire _39425_;
  wire _39426_;
  wire _39427_;
  wire _39428_;
  wire _39429_;
  wire _39430_;
  wire _39431_;
  wire _39432_;
  wire _39433_;
  wire _39434_;
  wire _39435_;
  wire _39436_;
  wire _39437_;
  wire _39438_;
  wire _39439_;
  wire _39440_;
  wire _39441_;
  wire _39442_;
  wire _39443_;
  wire _39444_;
  wire _39445_;
  wire _39446_;
  wire _39447_;
  wire _39448_;
  wire _39449_;
  wire _39450_;
  wire _39451_;
  wire _39452_;
  wire _39453_;
  wire _39454_;
  wire _39455_;
  wire _39456_;
  wire _39457_;
  wire _39458_;
  wire _39459_;
  wire _39460_;
  wire _39461_;
  wire _39462_;
  wire _39463_;
  wire _39464_;
  wire _39465_;
  wire _39466_;
  wire _39467_;
  wire _39468_;
  wire _39469_;
  wire _39470_;
  wire _39471_;
  wire _39472_;
  wire _39473_;
  wire _39474_;
  wire _39475_;
  wire _39476_;
  wire _39477_;
  wire _39478_;
  wire _39479_;
  wire _39480_;
  wire _39481_;
  wire _39482_;
  wire _39483_;
  wire _39484_;
  wire _39485_;
  wire _39486_;
  wire _39487_;
  wire _39488_;
  wire _39489_;
  wire _39490_;
  wire _39491_;
  wire _39492_;
  wire _39493_;
  wire _39494_;
  wire _39495_;
  wire _39496_;
  wire _39497_;
  wire _39498_;
  wire _39499_;
  wire _39500_;
  wire _39501_;
  wire _39502_;
  wire _39503_;
  wire _39504_;
  wire _39505_;
  wire _39506_;
  wire _39507_;
  wire _39508_;
  wire _39509_;
  wire _39510_;
  wire _39511_;
  wire _39512_;
  wire _39513_;
  wire _39514_;
  wire _39515_;
  wire _39516_;
  wire _39517_;
  wire _39518_;
  wire _39519_;
  wire _39520_;
  wire _39521_;
  wire _39522_;
  wire _39523_;
  wire _39524_;
  wire _39525_;
  wire _39526_;
  wire _39527_;
  wire _39528_;
  wire _39529_;
  wire _39530_;
  wire _39531_;
  wire _39532_;
  wire _39533_;
  wire _39534_;
  wire _39535_;
  wire _39536_;
  wire _39537_;
  wire _39538_;
  wire _39539_;
  wire _39540_;
  wire _39541_;
  wire _39542_;
  wire _39543_;
  wire _39544_;
  wire _39545_;
  wire _39546_;
  wire _39547_;
  wire _39548_;
  wire _39549_;
  wire _39550_;
  wire _39551_;
  wire _39552_;
  wire _39553_;
  wire _39554_;
  wire _39555_;
  wire _39556_;
  wire _39557_;
  wire _39558_;
  wire _39559_;
  wire _39560_;
  wire _39561_;
  wire _39562_;
  wire _39563_;
  wire _39564_;
  wire _39565_;
  wire _39566_;
  wire _39567_;
  wire _39568_;
  wire _39569_;
  wire _39570_;
  wire _39571_;
  wire _39572_;
  wire _39573_;
  wire _39574_;
  wire _39575_;
  wire _39576_;
  wire _39577_;
  wire _39578_;
  wire _39579_;
  wire _39580_;
  wire _39581_;
  wire _39582_;
  wire _39583_;
  wire _39584_;
  wire _39585_;
  wire _39586_;
  wire _39587_;
  wire _39588_;
  wire _39589_;
  wire _39590_;
  wire _39591_;
  wire _39592_;
  wire _39593_;
  wire _39594_;
  wire _39595_;
  wire _39596_;
  wire _39597_;
  wire _39598_;
  wire _39599_;
  wire _39600_;
  wire _39601_;
  wire _39602_;
  wire _39603_;
  wire _39604_;
  wire _39605_;
  wire _39606_;
  wire _39607_;
  wire _39608_;
  wire _39609_;
  wire _39610_;
  wire _39611_;
  wire _39612_;
  wire _39613_;
  wire _39614_;
  wire _39615_;
  wire _39616_;
  wire _39617_;
  wire _39618_;
  wire _39619_;
  wire _39620_;
  wire _39621_;
  wire _39622_;
  wire _39623_;
  wire _39624_;
  wire _39625_;
  wire _39626_;
  wire _39627_;
  wire _39628_;
  wire _39629_;
  wire _39630_;
  wire _39631_;
  wire _39632_;
  wire _39633_;
  wire _39634_;
  wire _39635_;
  wire _39636_;
  wire _39637_;
  wire _39638_;
  wire _39639_;
  wire _39640_;
  wire _39641_;
  wire _39642_;
  wire _39643_;
  wire _39644_;
  wire _39645_;
  wire _39646_;
  wire _39647_;
  wire _39648_;
  wire _39649_;
  wire _39650_;
  wire _39651_;
  wire _39652_;
  wire _39653_;
  wire _39654_;
  wire _39655_;
  wire _39656_;
  wire _39657_;
  wire _39658_;
  wire _39659_;
  wire _39660_;
  wire _39661_;
  wire _39662_;
  wire _39663_;
  wire _39664_;
  wire _39665_;
  wire _39666_;
  wire _39667_;
  wire _39668_;
  wire _39669_;
  wire _39670_;
  wire _39671_;
  wire _39672_;
  wire _39673_;
  wire _39674_;
  wire _39675_;
  wire _39676_;
  wire _39677_;
  wire _39678_;
  wire _39679_;
  wire _39680_;
  wire _39681_;
  wire _39682_;
  wire _39683_;
  wire _39684_;
  wire _39685_;
  wire _39686_;
  wire _39687_;
  wire _39688_;
  wire _39689_;
  wire _39690_;
  wire _39691_;
  wire _39692_;
  wire _39693_;
  wire _39694_;
  wire _39695_;
  wire _39696_;
  wire _39697_;
  wire _39698_;
  wire _39699_;
  wire _39700_;
  wire _39701_;
  wire _39702_;
  wire _39703_;
  wire _39704_;
  wire _39705_;
  wire _39706_;
  wire _39707_;
  wire _39708_;
  wire _39709_;
  wire _39710_;
  wire _39711_;
  wire _39712_;
  wire _39713_;
  wire _39714_;
  wire _39715_;
  wire _39716_;
  wire _39717_;
  wire _39718_;
  wire _39719_;
  wire _39720_;
  wire _39721_;
  wire _39722_;
  wire _39723_;
  wire _39724_;
  wire _39725_;
  wire _39726_;
  wire _39727_;
  wire _39728_;
  wire _39729_;
  wire _39730_;
  wire _39731_;
  wire _39732_;
  wire _39733_;
  wire _39734_;
  wire _39735_;
  wire _39736_;
  wire _39737_;
  wire _39738_;
  wire _39739_;
  wire _39740_;
  wire _39741_;
  wire _39742_;
  wire _39743_;
  wire _39744_;
  wire _39745_;
  wire _39746_;
  wire _39747_;
  wire _39748_;
  wire _39749_;
  wire _39750_;
  wire _39751_;
  wire _39752_;
  wire _39753_;
  wire _39754_;
  wire _39755_;
  wire _39756_;
  wire _39757_;
  wire _39758_;
  wire _39759_;
  wire _39760_;
  wire _39761_;
  wire _39762_;
  wire _39763_;
  wire _39764_;
  wire _39765_;
  wire _39766_;
  wire _39767_;
  wire _39768_;
  wire _39769_;
  wire _39770_;
  wire _39771_;
  wire _39772_;
  wire _39773_;
  wire _39774_;
  wire _39775_;
  wire _39776_;
  wire _39777_;
  wire _39778_;
  wire _39779_;
  wire _39780_;
  wire _39781_;
  wire _39782_;
  wire _39783_;
  wire _39784_;
  wire _39785_;
  wire _39786_;
  wire _39787_;
  wire _39788_;
  wire _39789_;
  wire _39790_;
  wire _39791_;
  wire _39792_;
  wire _39793_;
  wire _39794_;
  wire _39795_;
  wire _39796_;
  wire _39797_;
  wire _39798_;
  wire _39799_;
  wire _39800_;
  wire _39801_;
  wire _39802_;
  wire _39803_;
  wire _39804_;
  wire _39805_;
  wire _39806_;
  wire _39807_;
  wire _39808_;
  wire _39809_;
  wire _39810_;
  wire _39811_;
  wire _39812_;
  wire _39813_;
  wire _39814_;
  wire _39815_;
  wire _39816_;
  wire _39817_;
  wire _39818_;
  wire _39819_;
  wire _39820_;
  wire _39821_;
  wire _39822_;
  wire _39823_;
  wire _39824_;
  wire _39825_;
  wire _39826_;
  wire _39827_;
  wire _39828_;
  wire _39829_;
  wire _39830_;
  wire _39831_;
  wire _39832_;
  wire _39833_;
  wire _39834_;
  wire _39835_;
  wire _39836_;
  wire _39837_;
  wire _39838_;
  wire _39839_;
  wire _39840_;
  wire _39841_;
  wire _39842_;
  wire _39843_;
  wire _39844_;
  wire _39845_;
  wire _39846_;
  wire _39847_;
  wire _39848_;
  wire _39849_;
  wire _39850_;
  wire _39851_;
  wire _39852_;
  wire _39853_;
  wire _39854_;
  wire _39855_;
  wire _39856_;
  wire _39857_;
  wire _39858_;
  wire _39859_;
  wire _39860_;
  wire _39861_;
  wire _39862_;
  wire _39863_;
  wire _39864_;
  wire _39865_;
  wire _39866_;
  wire _39867_;
  wire _39868_;
  wire _39869_;
  wire _39870_;
  wire _39871_;
  wire _39872_;
  wire _39873_;
  wire _39874_;
  wire _39875_;
  wire _39876_;
  wire _39877_;
  wire _39878_;
  wire _39879_;
  wire _39880_;
  wire _39881_;
  wire _39882_;
  wire _39883_;
  wire _39884_;
  wire _39885_;
  wire _39886_;
  wire _39887_;
  wire _39888_;
  wire _39889_;
  wire _39890_;
  wire _39891_;
  wire _39892_;
  wire _39893_;
  wire _39894_;
  wire _39895_;
  wire _39896_;
  wire _39897_;
  wire _39898_;
  wire _39899_;
  wire _39900_;
  wire _39901_;
  wire _39902_;
  wire _39903_;
  wire _39904_;
  wire _39905_;
  wire _39906_;
  wire _39907_;
  wire _39908_;
  wire _39909_;
  wire _39910_;
  wire _39911_;
  wire _39912_;
  wire _39913_;
  wire _39914_;
  wire _39915_;
  wire _39916_;
  wire _39917_;
  wire _39918_;
  wire _39919_;
  wire _39920_;
  wire _39921_;
  wire _39922_;
  wire _39923_;
  wire _39924_;
  wire _39925_;
  wire _39926_;
  wire _39927_;
  wire _39928_;
  wire _39929_;
  wire _39930_;
  wire _39931_;
  wire _39932_;
  wire _39933_;
  wire _39934_;
  wire _39935_;
  wire _39936_;
  wire _39937_;
  wire _39938_;
  wire _39939_;
  wire _39940_;
  wire _39941_;
  wire _39942_;
  wire _39943_;
  wire _39944_;
  wire _39945_;
  wire _39946_;
  wire _39947_;
  wire _39948_;
  wire _39949_;
  wire _39950_;
  wire _39951_;
  wire _39952_;
  wire _39953_;
  wire _39954_;
  wire _39955_;
  wire _39956_;
  wire _39957_;
  wire _39958_;
  wire _39959_;
  wire _39960_;
  wire _39961_;
  wire _39962_;
  wire _39963_;
  wire _39964_;
  wire _39965_;
  wire _39966_;
  wire _39967_;
  wire _39968_;
  wire _39969_;
  wire _39970_;
  wire _39971_;
  wire _39972_;
  wire _39973_;
  wire _39974_;
  wire _39975_;
  wire _39976_;
  wire _39977_;
  wire _39978_;
  wire _39979_;
  wire _39980_;
  wire _39981_;
  wire _39982_;
  wire _39983_;
  wire _39984_;
  wire _39985_;
  wire _39986_;
  wire _39987_;
  wire _39988_;
  wire _39989_;
  wire _39990_;
  wire _39991_;
  wire _39992_;
  wire _39993_;
  wire _39994_;
  wire _39995_;
  wire _39996_;
  wire _39997_;
  wire _39998_;
  wire _39999_;
  wire _40000_;
  wire _40001_;
  wire _40002_;
  wire _40003_;
  wire _40004_;
  wire _40005_;
  wire _40006_;
  wire _40007_;
  wire _40008_;
  wire _40009_;
  wire _40010_;
  wire _40011_;
  wire _40012_;
  wire _40013_;
  wire _40014_;
  wire _40015_;
  wire _40016_;
  wire _40017_;
  wire _40018_;
  wire _40019_;
  wire _40020_;
  wire _40021_;
  wire _40022_;
  wire _40023_;
  wire _40024_;
  wire _40025_;
  wire _40026_;
  wire _40027_;
  wire _40028_;
  wire _40029_;
  wire _40030_;
  wire _40031_;
  wire _40032_;
  wire _40033_;
  wire _40034_;
  wire _40035_;
  wire _40036_;
  wire _40037_;
  wire _40038_;
  wire _40039_;
  wire _40040_;
  wire _40041_;
  wire _40042_;
  wire _40043_;
  wire _40044_;
  wire _40045_;
  wire _40046_;
  wire _40047_;
  wire _40048_;
  wire _40049_;
  wire _40050_;
  wire _40051_;
  wire _40052_;
  wire _40053_;
  wire _40054_;
  wire _40055_;
  wire _40056_;
  wire _40057_;
  wire _40058_;
  wire _40059_;
  wire _40060_;
  wire _40061_;
  wire _40062_;
  wire _40063_;
  wire _40064_;
  wire _40065_;
  wire _40066_;
  wire _40067_;
  wire _40068_;
  wire _40069_;
  wire _40070_;
  wire _40071_;
  wire _40072_;
  wire _40073_;
  wire _40074_;
  wire _40075_;
  wire _40076_;
  wire _40077_;
  wire _40078_;
  wire _40079_;
  wire _40080_;
  wire _40081_;
  wire _40082_;
  wire _40083_;
  wire _40084_;
  wire _40085_;
  wire _40086_;
  wire _40087_;
  wire _40088_;
  wire _40089_;
  wire _40090_;
  wire _40091_;
  wire _40092_;
  wire _40093_;
  wire _40094_;
  wire _40095_;
  wire _40096_;
  wire _40097_;
  wire _40098_;
  wire _40099_;
  wire _40100_;
  wire _40101_;
  wire _40102_;
  wire _40103_;
  wire _40104_;
  wire _40105_;
  wire _40106_;
  wire _40107_;
  wire _40108_;
  wire _40109_;
  wire _40110_;
  wire _40111_;
  wire _40112_;
  wire _40113_;
  wire _40114_;
  wire _40115_;
  wire _40116_;
  wire _40117_;
  wire _40118_;
  wire _40119_;
  wire _40120_;
  wire _40121_;
  wire _40122_;
  wire _40123_;
  wire _40124_;
  wire _40125_;
  wire _40126_;
  wire _40127_;
  wire _40128_;
  wire _40129_;
  wire _40130_;
  wire _40131_;
  wire _40132_;
  wire _40133_;
  wire _40134_;
  wire _40135_;
  wire _40136_;
  wire _40137_;
  wire _40138_;
  wire _40139_;
  wire _40140_;
  wire _40141_;
  wire _40142_;
  wire _40143_;
  wire _40144_;
  wire _40145_;
  wire _40146_;
  wire _40147_;
  wire _40148_;
  wire _40149_;
  wire _40150_;
  wire _40151_;
  wire _40152_;
  wire _40153_;
  wire _40154_;
  wire _40155_;
  wire _40156_;
  wire _40157_;
  wire _40158_;
  wire _40159_;
  wire _40160_;
  wire _40161_;
  wire _40162_;
  wire _40163_;
  wire _40164_;
  wire _40165_;
  wire _40166_;
  wire _40167_;
  wire _40168_;
  wire _40169_;
  wire _40170_;
  wire _40171_;
  wire _40172_;
  wire _40173_;
  wire _40174_;
  wire _40175_;
  wire _40176_;
  wire _40177_;
  wire _40178_;
  wire _40179_;
  wire _40180_;
  wire _40181_;
  wire _40182_;
  wire _40183_;
  wire _40184_;
  wire _40185_;
  wire _40186_;
  wire _40187_;
  wire _40188_;
  wire _40189_;
  wire _40190_;
  wire _40191_;
  wire _40192_;
  wire _40193_;
  wire _40194_;
  wire _40195_;
  wire _40196_;
  wire _40197_;
  wire _40198_;
  wire _40199_;
  wire _40200_;
  wire _40201_;
  wire _40202_;
  wire _40203_;
  wire _40204_;
  wire _40205_;
  wire _40206_;
  wire _40207_;
  wire _40208_;
  wire _40209_;
  wire _40210_;
  wire _40211_;
  wire _40212_;
  wire _40213_;
  wire _40214_;
  wire _40215_;
  wire _40216_;
  wire _40217_;
  wire _40218_;
  wire _40219_;
  wire _40220_;
  wire _40221_;
  wire _40222_;
  wire _40223_;
  wire _40224_;
  wire _40225_;
  wire _40226_;
  wire _40227_;
  wire _40228_;
  wire _40229_;
  wire _40230_;
  wire _40231_;
  wire _40232_;
  wire _40233_;
  wire _40234_;
  wire _40235_;
  wire _40236_;
  wire _40237_;
  wire _40238_;
  wire _40239_;
  wire _40240_;
  wire _40241_;
  wire _40242_;
  wire _40243_;
  wire _40244_;
  wire _40245_;
  wire _40246_;
  wire _40247_;
  wire _40248_;
  wire _40249_;
  wire _40250_;
  wire _40251_;
  wire _40252_;
  wire _40253_;
  wire _40254_;
  wire _40255_;
  wire _40256_;
  wire _40257_;
  wire _40258_;
  wire _40259_;
  wire _40260_;
  wire _40261_;
  wire _40262_;
  wire _40263_;
  wire _40264_;
  wire _40265_;
  wire _40266_;
  wire _40267_;
  wire _40268_;
  wire _40269_;
  wire _40270_;
  wire _40271_;
  wire _40272_;
  wire _40273_;
  wire _40274_;
  wire _40275_;
  wire _40276_;
  wire _40277_;
  wire _40278_;
  wire _40279_;
  wire _40280_;
  wire _40281_;
  wire _40282_;
  wire _40283_;
  wire _40284_;
  wire _40285_;
  wire _40286_;
  wire _40287_;
  wire _40288_;
  wire _40289_;
  wire _40290_;
  wire _40291_;
  wire _40292_;
  wire _40293_;
  wire _40294_;
  wire _40295_;
  wire _40296_;
  wire _40297_;
  wire _40298_;
  wire _40299_;
  wire _40300_;
  wire _40301_;
  wire _40302_;
  wire _40303_;
  wire _40304_;
  wire _40305_;
  wire _40306_;
  wire _40307_;
  wire _40308_;
  wire _40309_;
  wire _40310_;
  wire _40311_;
  wire _40312_;
  wire _40313_;
  wire _40314_;
  wire _40315_;
  wire _40316_;
  wire _40317_;
  wire _40318_;
  wire _40319_;
  wire _40320_;
  wire _40321_;
  wire _40322_;
  wire _40323_;
  wire _40324_;
  wire _40325_;
  wire _40326_;
  wire _40327_;
  wire _40328_;
  wire _40329_;
  wire _40330_;
  wire _40331_;
  wire _40332_;
  wire _40333_;
  wire _40334_;
  wire _40335_;
  wire _40336_;
  wire _40337_;
  wire _40338_;
  wire _40339_;
  wire _40340_;
  wire _40341_;
  wire _40342_;
  wire _40343_;
  wire _40344_;
  wire _40345_;
  wire _40346_;
  wire _40347_;
  wire _40348_;
  wire _40349_;
  wire _40350_;
  wire _40351_;
  wire _40352_;
  wire _40353_;
  wire _40354_;
  wire _40355_;
  wire _40356_;
  wire _40357_;
  wire _40358_;
  wire _40359_;
  wire _40360_;
  wire _40361_;
  wire _40362_;
  wire _40363_;
  wire _40364_;
  wire _40365_;
  wire _40366_;
  wire _40367_;
  wire _40368_;
  wire _40369_;
  wire _40370_;
  wire _40371_;
  wire _40372_;
  wire _40373_;
  wire _40374_;
  wire _40375_;
  wire _40376_;
  wire _40377_;
  wire _40378_;
  wire _40379_;
  wire _40380_;
  wire _40381_;
  wire _40382_;
  wire _40383_;
  wire _40384_;
  wire _40385_;
  wire _40386_;
  wire _40387_;
  wire _40388_;
  wire _40389_;
  wire _40390_;
  wire _40391_;
  wire _40392_;
  wire _40393_;
  wire _40394_;
  wire _40395_;
  wire _40396_;
  wire _40397_;
  wire _40398_;
  wire _40399_;
  wire _40400_;
  wire _40401_;
  wire _40402_;
  wire _40403_;
  wire _40404_;
  wire _40405_;
  wire _40406_;
  wire _40407_;
  wire _40408_;
  wire _40409_;
  wire _40410_;
  wire _40411_;
  wire _40412_;
  wire _40413_;
  wire _40414_;
  wire _40415_;
  wire _40416_;
  wire _40417_;
  wire _40418_;
  wire _40419_;
  wire _40420_;
  wire _40421_;
  wire _40422_;
  wire _40423_;
  wire _40424_;
  wire _40425_;
  wire _40426_;
  wire _40427_;
  wire _40428_;
  wire _40429_;
  wire _40430_;
  wire _40431_;
  wire _40432_;
  wire _40433_;
  wire _40434_;
  wire _40435_;
  wire _40436_;
  wire _40437_;
  wire _40438_;
  wire _40439_;
  wire _40440_;
  wire _40441_;
  wire _40442_;
  wire _40443_;
  wire _40444_;
  wire _40445_;
  wire _40446_;
  wire _40447_;
  wire _40448_;
  wire _40449_;
  wire _40450_;
  wire _40451_;
  wire _40452_;
  wire _40453_;
  wire _40454_;
  wire _40455_;
  wire _40456_;
  wire _40457_;
  wire _40458_;
  wire _40459_;
  wire _40460_;
  wire _40461_;
  wire _40462_;
  wire _40463_;
  wire _40464_;
  wire _40465_;
  wire _40466_;
  wire _40467_;
  wire _40468_;
  wire _40469_;
  wire _40470_;
  wire _40471_;
  wire _40472_;
  wire _40473_;
  wire _40474_;
  wire _40475_;
  wire _40476_;
  wire _40477_;
  wire _40478_;
  wire _40479_;
  wire _40480_;
  wire _40481_;
  wire _40482_;
  wire _40483_;
  wire _40484_;
  wire _40485_;
  wire _40486_;
  wire _40487_;
  wire _40488_;
  wire _40489_;
  wire _40490_;
  wire _40491_;
  wire _40492_;
  wire _40493_;
  wire _40494_;
  wire _40495_;
  wire _40496_;
  wire _40497_;
  wire _40498_;
  wire _40499_;
  wire _40500_;
  wire _40501_;
  wire _40502_;
  wire _40503_;
  wire _40504_;
  wire _40505_;
  wire _40506_;
  wire _40507_;
  wire _40508_;
  wire _40509_;
  wire _40510_;
  wire _40511_;
  wire _40512_;
  wire _40513_;
  wire _40514_;
  wire _40515_;
  wire _40516_;
  wire _40517_;
  wire _40518_;
  wire _40519_;
  wire _40520_;
  wire _40521_;
  wire _40522_;
  wire _40523_;
  wire _40524_;
  wire _40525_;
  wire _40526_;
  wire _40527_;
  wire _40528_;
  wire _40529_;
  wire _40530_;
  wire _40531_;
  wire _40532_;
  wire _40533_;
  wire _40534_;
  wire _40535_;
  wire _40536_;
  wire _40537_;
  wire _40538_;
  wire _40539_;
  wire _40540_;
  wire _40541_;
  wire _40542_;
  wire _40543_;
  wire _40544_;
  wire _40545_;
  wire _40546_;
  wire _40547_;
  wire _40548_;
  wire _40549_;
  wire _40550_;
  wire _40551_;
  wire _40552_;
  wire _40553_;
  wire _40554_;
  wire _40555_;
  wire _40556_;
  wire _40557_;
  wire _40558_;
  wire _40559_;
  wire _40560_;
  wire _40561_;
  wire _40562_;
  wire _40563_;
  wire _40564_;
  wire _40565_;
  wire _40566_;
  wire _40567_;
  wire _40568_;
  wire _40569_;
  wire _40570_;
  wire _40571_;
  wire _40572_;
  wire _40573_;
  wire _40574_;
  wire _40575_;
  wire _40576_;
  wire _40577_;
  wire _40578_;
  wire _40579_;
  wire _40580_;
  wire _40581_;
  wire _40582_;
  wire _40583_;
  wire _40584_;
  wire _40585_;
  wire _40586_;
  wire _40587_;
  wire _40588_;
  wire _40589_;
  wire _40590_;
  wire _40591_;
  wire _40592_;
  wire _40593_;
  wire _40594_;
  wire _40595_;
  wire _40596_;
  wire _40597_;
  wire _40598_;
  wire _40599_;
  wire _40600_;
  wire _40601_;
  wire _40602_;
  wire _40603_;
  wire _40604_;
  wire _40605_;
  wire _40606_;
  wire _40607_;
  wire _40608_;
  wire _40609_;
  wire _40610_;
  wire _40611_;
  wire _40612_;
  wire _40613_;
  wire _40614_;
  wire _40615_;
  wire _40616_;
  wire _40617_;
  wire _40618_;
  wire _40619_;
  wire _40620_;
  wire _40621_;
  wire _40622_;
  wire _40623_;
  wire _40624_;
  wire _40625_;
  wire _40626_;
  wire _40627_;
  wire _40628_;
  wire _40629_;
  wire _40630_;
  wire _40631_;
  wire _40632_;
  wire _40633_;
  wire _40634_;
  wire _40635_;
  wire _40636_;
  wire _40637_;
  wire _40638_;
  wire _40639_;
  wire _40640_;
  wire _40641_;
  wire _40642_;
  wire _40643_;
  wire _40644_;
  wire _40645_;
  wire _40646_;
  wire _40647_;
  wire _40648_;
  wire _40649_;
  wire _40650_;
  wire _40651_;
  wire _40652_;
  wire _40653_;
  wire _40654_;
  wire _40655_;
  wire _40656_;
  wire _40657_;
  wire _40658_;
  wire _40659_;
  wire _40660_;
  wire _40661_;
  wire _40662_;
  wire _40663_;
  wire _40664_;
  wire _40665_;
  wire _40666_;
  wire _40667_;
  wire _40668_;
  wire _40669_;
  wire _40670_;
  wire _40671_;
  wire _40672_;
  wire _40673_;
  wire _40674_;
  wire _40675_;
  wire _40676_;
  wire _40677_;
  wire _40678_;
  wire _40679_;
  wire _40680_;
  wire _40681_;
  wire _40682_;
  wire _40683_;
  wire _40684_;
  wire _40685_;
  wire _40686_;
  wire _40687_;
  wire _40688_;
  wire _40689_;
  wire _40690_;
  wire _40691_;
  wire _40692_;
  wire _40693_;
  wire _40694_;
  wire _40695_;
  wire _40696_;
  wire _40697_;
  wire _40698_;
  wire _40699_;
  wire _40700_;
  wire _40701_;
  wire _40702_;
  wire _40703_;
  wire _40704_;
  wire _40705_;
  wire _40706_;
  wire _40707_;
  wire _40708_;
  wire _40709_;
  wire _40710_;
  wire _40711_;
  wire _40712_;
  wire _40713_;
  wire _40714_;
  wire _40715_;
  wire _40716_;
  wire _40717_;
  wire _40718_;
  wire _40719_;
  wire _40720_;
  wire _40721_;
  wire _40722_;
  wire _40723_;
  wire _40724_;
  wire _40725_;
  wire _40726_;
  wire _40727_;
  wire _40728_;
  wire _40729_;
  wire _40730_;
  wire _40731_;
  wire _40732_;
  wire _40733_;
  wire _40734_;
  wire _40735_;
  wire _40736_;
  wire _40737_;
  wire _40738_;
  wire _40739_;
  wire _40740_;
  wire _40741_;
  wire _40742_;
  wire _40743_;
  wire _40744_;
  wire _40745_;
  wire _40746_;
  wire _40747_;
  wire _40748_;
  wire _40749_;
  wire _40750_;
  wire _40751_;
  wire _40752_;
  wire _40753_;
  wire _40754_;
  wire _40755_;
  wire _40756_;
  wire _40757_;
  wire _40758_;
  wire _40759_;
  wire _40760_;
  wire _40761_;
  wire _40762_;
  wire _40763_;
  wire _40764_;
  wire _40765_;
  wire _40766_;
  wire _40767_;
  wire _40768_;
  wire _40769_;
  wire _40770_;
  wire _40771_;
  wire _40772_;
  wire _40773_;
  wire _40774_;
  wire _40775_;
  wire _40776_;
  wire _40777_;
  wire _40778_;
  wire _40779_;
  wire _40780_;
  wire _40781_;
  wire _40782_;
  wire _40783_;
  wire _40784_;
  wire _40785_;
  wire _40786_;
  wire _40787_;
  wire _40788_;
  wire _40789_;
  wire _40790_;
  wire _40791_;
  wire _40792_;
  wire _40793_;
  wire _40794_;
  wire _40795_;
  wire _40796_;
  wire _40797_;
  wire _40798_;
  wire _40799_;
  wire _40800_;
  wire _40801_;
  wire _40802_;
  wire _40803_;
  wire _40804_;
  wire _40805_;
  wire _40806_;
  wire _40807_;
  wire _40808_;
  wire _40809_;
  wire _40810_;
  wire _40811_;
  wire _40812_;
  wire _40813_;
  wire _40814_;
  wire _40815_;
  wire _40816_;
  wire _40817_;
  wire _40818_;
  wire _40819_;
  wire _40820_;
  wire _40821_;
  wire _40822_;
  wire _40823_;
  wire _40824_;
  wire _40825_;
  wire _40826_;
  wire _40827_;
  wire _40828_;
  wire _40829_;
  wire _40830_;
  wire _40831_;
  wire _40832_;
  wire _40833_;
  wire _40834_;
  wire _40835_;
  wire _40836_;
  wire _40837_;
  wire _40838_;
  wire _40839_;
  wire _40840_;
  wire _40841_;
  wire _40842_;
  wire _40843_;
  wire _40844_;
  wire _40845_;
  wire _40846_;
  wire _40847_;
  wire _40848_;
  wire _40849_;
  wire _40850_;
  wire _40851_;
  wire _40852_;
  wire _40853_;
  wire _40854_;
  wire _40855_;
  wire _40856_;
  wire _40857_;
  wire _40858_;
  wire _40859_;
  wire _40860_;
  wire _40861_;
  wire _40862_;
  wire _40863_;
  wire _40864_;
  wire _40865_;
  wire _40866_;
  wire _40867_;
  wire _40868_;
  wire _40869_;
  wire _40870_;
  wire _40871_;
  wire _40872_;
  wire _40873_;
  wire _40874_;
  wire _40875_;
  wire _40876_;
  wire _40877_;
  wire _40878_;
  wire _40879_;
  wire _40880_;
  wire _40881_;
  wire _40882_;
  wire _40883_;
  wire _40884_;
  wire _40885_;
  wire _40886_;
  wire _40887_;
  wire _40888_;
  wire _40889_;
  wire _40890_;
  wire _40891_;
  wire _40892_;
  wire _40893_;
  wire _40894_;
  wire _40895_;
  wire _40896_;
  wire _40897_;
  wire _40898_;
  wire _40899_;
  wire _40900_;
  wire _40901_;
  wire _40902_;
  wire _40903_;
  wire _40904_;
  wire _40905_;
  wire _40906_;
  wire _40907_;
  wire _40908_;
  wire _40909_;
  wire _40910_;
  wire _40911_;
  wire _40912_;
  wire _40913_;
  wire _40914_;
  wire _40915_;
  wire _40916_;
  wire _40917_;
  wire _40918_;
  wire _40919_;
  wire _40920_;
  wire _40921_;
  wire _40922_;
  wire _40923_;
  wire _40924_;
  wire _40925_;
  wire _40926_;
  wire _40927_;
  wire _40928_;
  wire _40929_;
  wire _40930_;
  wire _40931_;
  wire _40932_;
  wire _40933_;
  wire _40934_;
  wire _40935_;
  wire _40936_;
  wire _40937_;
  wire _40938_;
  wire _40939_;
  wire _40940_;
  wire _40941_;
  wire _40942_;
  wire _40943_;
  wire _40944_;
  wire _40945_;
  wire _40946_;
  wire _40947_;
  wire _40948_;
  wire _40949_;
  wire _40950_;
  wire _40951_;
  wire _40952_;
  wire _40953_;
  wire _40954_;
  wire _40955_;
  wire _40956_;
  wire _40957_;
  wire _40958_;
  wire _40959_;
  wire _40960_;
  wire _40961_;
  wire _40962_;
  wire _40963_;
  wire _40964_;
  wire _40965_;
  wire _40966_;
  wire _40967_;
  wire _40968_;
  wire _40969_;
  wire _40970_;
  wire _40971_;
  wire _40972_;
  wire _40973_;
  wire _40974_;
  wire _40975_;
  wire _40976_;
  wire _40977_;
  wire _40978_;
  wire _40979_;
  wire _40980_;
  wire _40981_;
  wire _40982_;
  wire _40983_;
  wire _40984_;
  wire _40985_;
  wire _40986_;
  wire _40987_;
  wire _40988_;
  wire _40989_;
  wire _40990_;
  wire _40991_;
  wire _40992_;
  wire _40993_;
  wire _40994_;
  wire _40995_;
  wire _40996_;
  wire _40997_;
  wire _40998_;
  wire _40999_;
  wire _41000_;
  wire _41001_;
  wire _41002_;
  wire _41003_;
  wire _41004_;
  wire _41005_;
  wire _41006_;
  wire _41007_;
  wire _41008_;
  wire _41009_;
  wire _41010_;
  wire _41011_;
  wire _41012_;
  wire _41013_;
  wire _41014_;
  wire _41015_;
  wire _41016_;
  wire _41017_;
  wire _41018_;
  wire _41019_;
  wire _41020_;
  wire _41021_;
  wire _41022_;
  wire _41023_;
  wire _41024_;
  wire _41025_;
  wire _41026_;
  wire _41027_;
  wire _41028_;
  wire _41029_;
  wire _41030_;
  wire _41031_;
  wire _41032_;
  wire _41033_;
  wire _41034_;
  wire _41035_;
  wire _41036_;
  wire _41037_;
  wire _41038_;
  wire _41039_;
  wire _41040_;
  wire _41041_;
  wire _41042_;
  wire _41043_;
  wire _41044_;
  wire _41045_;
  wire _41046_;
  wire _41047_;
  wire _41048_;
  wire _41049_;
  wire _41050_;
  wire _41051_;
  wire _41052_;
  wire _41053_;
  wire _41054_;
  wire _41055_;
  wire _41056_;
  wire _41057_;
  wire _41058_;
  wire _41059_;
  wire _41060_;
  wire _41061_;
  wire _41062_;
  wire _41063_;
  wire _41064_;
  wire _41065_;
  wire _41066_;
  wire _41067_;
  wire _41068_;
  wire _41069_;
  wire _41070_;
  wire _41071_;
  wire _41072_;
  wire _41073_;
  wire _41074_;
  wire _41075_;
  wire _41076_;
  wire _41077_;
  wire _41078_;
  wire _41079_;
  wire _41080_;
  wire _41081_;
  wire _41082_;
  wire _41083_;
  wire _41084_;
  wire _41085_;
  wire _41086_;
  wire _41087_;
  wire _41088_;
  wire _41089_;
  wire _41090_;
  wire _41091_;
  wire _41092_;
  wire _41093_;
  wire _41094_;
  wire _41095_;
  wire _41096_;
  wire _41097_;
  wire _41098_;
  wire _41099_;
  wire _41100_;
  wire _41101_;
  wire _41102_;
  wire _41103_;
  wire _41104_;
  wire _41105_;
  wire _41106_;
  wire _41107_;
  wire _41108_;
  wire _41109_;
  wire _41110_;
  wire _41111_;
  wire _41112_;
  wire _41113_;
  wire _41114_;
  wire _41115_;
  wire _41116_;
  wire _41117_;
  wire _41118_;
  wire _41119_;
  wire _41120_;
  wire _41121_;
  wire _41122_;
  wire _41123_;
  wire _41124_;
  wire _41125_;
  wire _41126_;
  wire _41127_;
  wire _41128_;
  wire _41129_;
  wire _41130_;
  wire _41131_;
  wire _41132_;
  wire _41133_;
  wire _41134_;
  wire _41135_;
  wire _41136_;
  wire _41137_;
  wire _41138_;
  wire _41139_;
  wire _41140_;
  wire _41141_;
  wire _41142_;
  wire _41143_;
  wire _41144_;
  wire _41145_;
  wire _41146_;
  wire _41147_;
  wire _41148_;
  wire _41149_;
  wire _41150_;
  wire _41151_;
  wire _41152_;
  wire _41153_;
  wire _41154_;
  wire _41155_;
  wire _41156_;
  wire _41157_;
  wire _41158_;
  wire _41159_;
  wire _41160_;
  wire _41161_;
  wire _41162_;
  wire _41163_;
  wire _41164_;
  wire _41165_;
  wire _41166_;
  wire _41167_;
  wire _41168_;
  wire _41169_;
  wire _41170_;
  wire _41171_;
  wire _41172_;
  wire _41173_;
  wire _41174_;
  wire _41175_;
  wire _41176_;
  wire _41177_;
  wire _41178_;
  wire _41179_;
  wire _41180_;
  wire _41181_;
  wire _41182_;
  wire _41183_;
  wire _41184_;
  wire _41185_;
  wire _41186_;
  wire _41187_;
  wire _41188_;
  wire _41189_;
  wire _41190_;
  wire _41191_;
  wire _41192_;
  wire _41193_;
  wire _41194_;
  wire _41195_;
  wire _41196_;
  wire _41197_;
  wire _41198_;
  wire _41199_;
  wire _41200_;
  wire _41201_;
  wire _41202_;
  wire _41203_;
  wire _41204_;
  wire _41205_;
  wire _41206_;
  wire _41207_;
  wire _41208_;
  wire _41209_;
  wire _41210_;
  wire _41211_;
  wire _41212_;
  wire _41213_;
  wire _41214_;
  wire _41215_;
  wire _41216_;
  wire _41217_;
  wire _41218_;
  wire _41219_;
  wire _41220_;
  wire _41221_;
  wire _41222_;
  wire _41223_;
  wire _41224_;
  wire _41225_;
  wire _41226_;
  wire _41227_;
  wire _41228_;
  wire _41229_;
  wire _41230_;
  wire _41231_;
  wire _41232_;
  wire _41233_;
  wire _41234_;
  wire _41235_;
  wire _41236_;
  wire _41237_;
  wire _41238_;
  wire _41239_;
  wire _41240_;
  wire _41241_;
  wire _41242_;
  wire _41243_;
  wire _41244_;
  wire _41245_;
  wire _41246_;
  wire _41247_;
  wire _41248_;
  wire _41249_;
  wire _41250_;
  wire _41251_;
  wire _41252_;
  wire _41253_;
  wire _41254_;
  input [34:0] ABINPUT;
  wire [7:0] ACC_gm;
  wire [7:0] B_gm;
  wire [7:0] DPH_gm;
  wire [7:0] DPL_gm;
  wire [7:0] IE_gm;
  wire [7:0] IP_gm;
  wire [7:0] P0_gm;
  wire [7:0] P1_gm;
  wire [7:0] P2_gm;
  wire [7:0] P3_gm;
  wire [7:0] PCON_gm;
  wire [7:0] PSW_gm;
  wire [7:0] SBUF_gm;
  wire [7:0] SCON_gm;
  wire [7:0] SP_gm;
  wire [7:0] TCON_gm;
  wire [7:0] TH0_gm;
  wire [7:0] TH1_gm;
  wire [7:0] TL0_gm;
  wire [7:0] TL1_gm;
  wire [7:0] TMOD_gm;
  wire [7:0] acc_impl;
  wire [7:0] b_reg_impl;
  input clk;
  wire [31:0] cxrom_data_out;
  wire [15:0] dptr_impl;
  wire \oc8051_gm_cxrom_1.cell0.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell0.data ;
  wire \oc8051_gm_cxrom_1.cell0.rst ;
  wire \oc8051_gm_cxrom_1.cell0.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell0.word ;
  wire \oc8051_gm_cxrom_1.cell1.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell1.data ;
  wire \oc8051_gm_cxrom_1.cell1.rst ;
  wire \oc8051_gm_cxrom_1.cell1.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell1.word ;
  wire \oc8051_gm_cxrom_1.cell10.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell10.data ;
  wire \oc8051_gm_cxrom_1.cell10.rst ;
  wire \oc8051_gm_cxrom_1.cell10.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell10.word ;
  wire \oc8051_gm_cxrom_1.cell11.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell11.data ;
  wire \oc8051_gm_cxrom_1.cell11.rst ;
  wire \oc8051_gm_cxrom_1.cell11.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell11.word ;
  wire \oc8051_gm_cxrom_1.cell12.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell12.data ;
  wire \oc8051_gm_cxrom_1.cell12.rst ;
  wire \oc8051_gm_cxrom_1.cell12.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell12.word ;
  wire \oc8051_gm_cxrom_1.cell13.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell13.data ;
  wire \oc8051_gm_cxrom_1.cell13.rst ;
  wire \oc8051_gm_cxrom_1.cell13.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell13.word ;
  wire \oc8051_gm_cxrom_1.cell14.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell14.data ;
  wire \oc8051_gm_cxrom_1.cell14.rst ;
  wire \oc8051_gm_cxrom_1.cell14.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell14.word ;
  wire \oc8051_gm_cxrom_1.cell15.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell15.data ;
  wire \oc8051_gm_cxrom_1.cell15.rst ;
  wire \oc8051_gm_cxrom_1.cell15.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell15.word ;
  wire \oc8051_gm_cxrom_1.cell2.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell2.data ;
  wire \oc8051_gm_cxrom_1.cell2.rst ;
  wire \oc8051_gm_cxrom_1.cell2.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell2.word ;
  wire \oc8051_gm_cxrom_1.cell3.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell3.data ;
  wire \oc8051_gm_cxrom_1.cell3.rst ;
  wire \oc8051_gm_cxrom_1.cell3.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell3.word ;
  wire \oc8051_gm_cxrom_1.cell4.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell4.data ;
  wire \oc8051_gm_cxrom_1.cell4.rst ;
  wire \oc8051_gm_cxrom_1.cell4.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell4.word ;
  wire \oc8051_gm_cxrom_1.cell5.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell5.data ;
  wire \oc8051_gm_cxrom_1.cell5.rst ;
  wire \oc8051_gm_cxrom_1.cell5.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell5.word ;
  wire \oc8051_gm_cxrom_1.cell6.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell6.data ;
  wire \oc8051_gm_cxrom_1.cell6.rst ;
  wire \oc8051_gm_cxrom_1.cell6.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell6.word ;
  wire \oc8051_gm_cxrom_1.cell7.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell7.data ;
  wire \oc8051_gm_cxrom_1.cell7.rst ;
  wire \oc8051_gm_cxrom_1.cell7.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell7.word ;
  wire \oc8051_gm_cxrom_1.cell8.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell8.data ;
  wire \oc8051_gm_cxrom_1.cell8.rst ;
  wire \oc8051_gm_cxrom_1.cell8.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell8.word ;
  wire \oc8051_gm_cxrom_1.cell9.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell9.data ;
  wire \oc8051_gm_cxrom_1.cell9.rst ;
  wire \oc8051_gm_cxrom_1.cell9.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell9.word ;
  wire \oc8051_gm_cxrom_1.clk ;
  wire [31:0] \oc8051_gm_cxrom_1.cxrom_data_out ;
  wire [15:0] \oc8051_gm_cxrom_1.rd_addr_0 ;
  wire \oc8051_gm_cxrom_1.rst ;
  wire [127:0] \oc8051_gm_cxrom_1.word_in ;
  wire [7:0] \oc8051_golden_model_1.ACC ;
  wire [7:0] \oc8051_golden_model_1.ACC_03 ;
  wire [7:0] \oc8051_golden_model_1.ACC_13 ;
  wire [7:0] \oc8051_golden_model_1.ACC_23 ;
  wire [7:0] \oc8051_golden_model_1.ACC_33 ;
  wire [7:0] \oc8051_golden_model_1.ACC_c4 ;
  wire [7:0] \oc8051_golden_model_1.ACC_d6 ;
  wire [7:0] \oc8051_golden_model_1.ACC_d7 ;
  wire [7:0] \oc8051_golden_model_1.ACC_e6 ;
  wire [7:0] \oc8051_golden_model_1.ACC_e7 ;
  wire [7:0] \oc8051_golden_model_1.B ;
  wire [7:0] \oc8051_golden_model_1.DPH ;
  wire [7:0] \oc8051_golden_model_1.DPL ;
  wire [7:0] \oc8051_golden_model_1.IE ;
  wire [7:0] \oc8051_golden_model_1.IP ;
  wire [7:0] \oc8051_golden_model_1.IRAM[0] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[10] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[11] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[12] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[13] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[14] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[15] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[1] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[2] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[3] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[4] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[5] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[6] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[7] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[8] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[9] ;
  wire [7:0] \oc8051_golden_model_1.P0 ;
  wire [7:0] \oc8051_golden_model_1.P0INREG ;
  wire [7:0] \oc8051_golden_model_1.P1 ;
  wire [7:0] \oc8051_golden_model_1.P1INREG ;
  wire [7:0] \oc8051_golden_model_1.P2 ;
  wire [7:0] \oc8051_golden_model_1.P2INREG ;
  wire [7:0] \oc8051_golden_model_1.P3 ;
  wire [7:0] \oc8051_golden_model_1.P3INREG ;
  wire [15:0] \oc8051_golden_model_1.PC ;
  wire [7:0] \oc8051_golden_model_1.PCON ;
  wire [15:0] \oc8051_golden_model_1.PC_22 ;
  wire [15:0] \oc8051_golden_model_1.PC_32 ;
  wire [7:0] \oc8051_golden_model_1.PSW ;
  wire [7:0] \oc8051_golden_model_1.PSW_00 ;
  wire [7:0] \oc8051_golden_model_1.PSW_01 ;
  wire [7:0] \oc8051_golden_model_1.PSW_02 ;
  wire [7:0] \oc8051_golden_model_1.PSW_03 ;
  wire [7:0] \oc8051_golden_model_1.PSW_04 ;
  wire [7:0] \oc8051_golden_model_1.PSW_06 ;
  wire [7:0] \oc8051_golden_model_1.PSW_07 ;
  wire [7:0] \oc8051_golden_model_1.PSW_08 ;
  wire [7:0] \oc8051_golden_model_1.PSW_09 ;
  wire [7:0] \oc8051_golden_model_1.PSW_0a ;
  wire [7:0] \oc8051_golden_model_1.PSW_0b ;
  wire [7:0] \oc8051_golden_model_1.PSW_0c ;
  wire [7:0] \oc8051_golden_model_1.PSW_0d ;
  wire [7:0] \oc8051_golden_model_1.PSW_0e ;
  wire [7:0] \oc8051_golden_model_1.PSW_0f ;
  wire [7:0] \oc8051_golden_model_1.PSW_11 ;
  wire [7:0] \oc8051_golden_model_1.PSW_12 ;
  wire [7:0] \oc8051_golden_model_1.PSW_13 ;
  wire [7:0] \oc8051_golden_model_1.PSW_14 ;
  wire [7:0] \oc8051_golden_model_1.PSW_16 ;
  wire [7:0] \oc8051_golden_model_1.PSW_17 ;
  wire [7:0] \oc8051_golden_model_1.PSW_18 ;
  wire [7:0] \oc8051_golden_model_1.PSW_19 ;
  wire [7:0] \oc8051_golden_model_1.PSW_1a ;
  wire [7:0] \oc8051_golden_model_1.PSW_1b ;
  wire [7:0] \oc8051_golden_model_1.PSW_1c ;
  wire [7:0] \oc8051_golden_model_1.PSW_1d ;
  wire [7:0] \oc8051_golden_model_1.PSW_1e ;
  wire [7:0] \oc8051_golden_model_1.PSW_1f ;
  wire [7:0] \oc8051_golden_model_1.PSW_20 ;
  wire [7:0] \oc8051_golden_model_1.PSW_21 ;
  wire [7:0] \oc8051_golden_model_1.PSW_22 ;
  wire [7:0] \oc8051_golden_model_1.PSW_23 ;
  wire [7:0] \oc8051_golden_model_1.PSW_24 ;
  wire [7:0] \oc8051_golden_model_1.PSW_25 ;
  wire [7:0] \oc8051_golden_model_1.PSW_26 ;
  wire [7:0] \oc8051_golden_model_1.PSW_27 ;
  wire [7:0] \oc8051_golden_model_1.PSW_28 ;
  wire [7:0] \oc8051_golden_model_1.PSW_29 ;
  wire [7:0] \oc8051_golden_model_1.PSW_2a ;
  wire [7:0] \oc8051_golden_model_1.PSW_2b ;
  wire [7:0] \oc8051_golden_model_1.PSW_2c ;
  wire [7:0] \oc8051_golden_model_1.PSW_2d ;
  wire [7:0] \oc8051_golden_model_1.PSW_2e ;
  wire [7:0] \oc8051_golden_model_1.PSW_2f ;
  wire [7:0] \oc8051_golden_model_1.PSW_30 ;
  wire [7:0] \oc8051_golden_model_1.PSW_31 ;
  wire [7:0] \oc8051_golden_model_1.PSW_32 ;
  wire [7:0] \oc8051_golden_model_1.PSW_33 ;
  wire [7:0] \oc8051_golden_model_1.PSW_34 ;
  wire [7:0] \oc8051_golden_model_1.PSW_35 ;
  wire [7:0] \oc8051_golden_model_1.PSW_36 ;
  wire [7:0] \oc8051_golden_model_1.PSW_37 ;
  wire [7:0] \oc8051_golden_model_1.PSW_38 ;
  wire [7:0] \oc8051_golden_model_1.PSW_39 ;
  wire [7:0] \oc8051_golden_model_1.PSW_3a ;
  wire [7:0] \oc8051_golden_model_1.PSW_3b ;
  wire [7:0] \oc8051_golden_model_1.PSW_3c ;
  wire [7:0] \oc8051_golden_model_1.PSW_3d ;
  wire [7:0] \oc8051_golden_model_1.PSW_3e ;
  wire [7:0] \oc8051_golden_model_1.PSW_3f ;
  wire [7:0] \oc8051_golden_model_1.PSW_40 ;
  wire [7:0] \oc8051_golden_model_1.PSW_41 ;
  wire [7:0] \oc8051_golden_model_1.PSW_42 ;
  wire [7:0] \oc8051_golden_model_1.PSW_44 ;
  wire [7:0] \oc8051_golden_model_1.PSW_45 ;
  wire [7:0] \oc8051_golden_model_1.PSW_46 ;
  wire [7:0] \oc8051_golden_model_1.PSW_47 ;
  wire [7:0] \oc8051_golden_model_1.PSW_48 ;
  wire [7:0] \oc8051_golden_model_1.PSW_49 ;
  wire [7:0] \oc8051_golden_model_1.PSW_4a ;
  wire [7:0] \oc8051_golden_model_1.PSW_4b ;
  wire [7:0] \oc8051_golden_model_1.PSW_4c ;
  wire [7:0] \oc8051_golden_model_1.PSW_4d ;
  wire [7:0] \oc8051_golden_model_1.PSW_4e ;
  wire [7:0] \oc8051_golden_model_1.PSW_4f ;
  wire [7:0] \oc8051_golden_model_1.PSW_50 ;
  wire [7:0] \oc8051_golden_model_1.PSW_51 ;
  wire [7:0] \oc8051_golden_model_1.PSW_52 ;
  wire [7:0] \oc8051_golden_model_1.PSW_54 ;
  wire [7:0] \oc8051_golden_model_1.PSW_55 ;
  wire [7:0] \oc8051_golden_model_1.PSW_56 ;
  wire [7:0] \oc8051_golden_model_1.PSW_57 ;
  wire [7:0] \oc8051_golden_model_1.PSW_58 ;
  wire [7:0] \oc8051_golden_model_1.PSW_59 ;
  wire [7:0] \oc8051_golden_model_1.PSW_5a ;
  wire [7:0] \oc8051_golden_model_1.PSW_5b ;
  wire [7:0] \oc8051_golden_model_1.PSW_5c ;
  wire [7:0] \oc8051_golden_model_1.PSW_5d ;
  wire [7:0] \oc8051_golden_model_1.PSW_5e ;
  wire [7:0] \oc8051_golden_model_1.PSW_5f ;
  wire [7:0] \oc8051_golden_model_1.PSW_60 ;
  wire [7:0] \oc8051_golden_model_1.PSW_61 ;
  wire [7:0] \oc8051_golden_model_1.PSW_64 ;
  wire [7:0] \oc8051_golden_model_1.PSW_65 ;
  wire [7:0] \oc8051_golden_model_1.PSW_66 ;
  wire [7:0] \oc8051_golden_model_1.PSW_67 ;
  wire [7:0] \oc8051_golden_model_1.PSW_68 ;
  wire [7:0] \oc8051_golden_model_1.PSW_69 ;
  wire [7:0] \oc8051_golden_model_1.PSW_6a ;
  wire [7:0] \oc8051_golden_model_1.PSW_6b ;
  wire [7:0] \oc8051_golden_model_1.PSW_6c ;
  wire [7:0] \oc8051_golden_model_1.PSW_6d ;
  wire [7:0] \oc8051_golden_model_1.PSW_6e ;
  wire [7:0] \oc8051_golden_model_1.PSW_6f ;
  wire [7:0] \oc8051_golden_model_1.PSW_70 ;
  wire [7:0] \oc8051_golden_model_1.PSW_71 ;
  wire [7:0] \oc8051_golden_model_1.PSW_72 ;
  wire [7:0] \oc8051_golden_model_1.PSW_73 ;
  wire [7:0] \oc8051_golden_model_1.PSW_74 ;
  wire [7:0] \oc8051_golden_model_1.PSW_76 ;
  wire [7:0] \oc8051_golden_model_1.PSW_77 ;
  wire [7:0] \oc8051_golden_model_1.PSW_78 ;
  wire [7:0] \oc8051_golden_model_1.PSW_79 ;
  wire [7:0] \oc8051_golden_model_1.PSW_7a ;
  wire [7:0] \oc8051_golden_model_1.PSW_7b ;
  wire [7:0] \oc8051_golden_model_1.PSW_7c ;
  wire [7:0] \oc8051_golden_model_1.PSW_7d ;
  wire [7:0] \oc8051_golden_model_1.PSW_7e ;
  wire [7:0] \oc8051_golden_model_1.PSW_7f ;
  wire [7:0] \oc8051_golden_model_1.PSW_80 ;
  wire [7:0] \oc8051_golden_model_1.PSW_81 ;
  wire [7:0] \oc8051_golden_model_1.PSW_82 ;
  wire [7:0] \oc8051_golden_model_1.PSW_83 ;
  wire [7:0] \oc8051_golden_model_1.PSW_84 ;
  wire [7:0] \oc8051_golden_model_1.PSW_90 ;
  wire [7:0] \oc8051_golden_model_1.PSW_91 ;
  wire [7:0] \oc8051_golden_model_1.PSW_93 ;
  wire [7:0] \oc8051_golden_model_1.PSW_94 ;
  wire [7:0] \oc8051_golden_model_1.PSW_95 ;
  wire [7:0] \oc8051_golden_model_1.PSW_96 ;
  wire [7:0] \oc8051_golden_model_1.PSW_97 ;
  wire [7:0] \oc8051_golden_model_1.PSW_98 ;
  wire [7:0] \oc8051_golden_model_1.PSW_99 ;
  wire [7:0] \oc8051_golden_model_1.PSW_9a ;
  wire [7:0] \oc8051_golden_model_1.PSW_9b ;
  wire [7:0] \oc8051_golden_model_1.PSW_9c ;
  wire [7:0] \oc8051_golden_model_1.PSW_9d ;
  wire [7:0] \oc8051_golden_model_1.PSW_9e ;
  wire [7:0] \oc8051_golden_model_1.PSW_9f ;
  wire [7:0] \oc8051_golden_model_1.PSW_a0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a2 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_aa ;
  wire [7:0] \oc8051_golden_model_1.PSW_ab ;
  wire [7:0] \oc8051_golden_model_1.PSW_ac ;
  wire [7:0] \oc8051_golden_model_1.PSW_ad ;
  wire [7:0] \oc8051_golden_model_1.PSW_ae ;
  wire [7:0] \oc8051_golden_model_1.PSW_af ;
  wire [7:0] \oc8051_golden_model_1.PSW_b0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_ba ;
  wire [7:0] \oc8051_golden_model_1.PSW_bb ;
  wire [7:0] \oc8051_golden_model_1.PSW_bc ;
  wire [7:0] \oc8051_golden_model_1.PSW_bd ;
  wire [7:0] \oc8051_golden_model_1.PSW_be ;
  wire [7:0] \oc8051_golden_model_1.PSW_bf ;
  wire [7:0] \oc8051_golden_model_1.PSW_c0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_ca ;
  wire [7:0] \oc8051_golden_model_1.PSW_cb ;
  wire [7:0] \oc8051_golden_model_1.PSW_cc ;
  wire [7:0] \oc8051_golden_model_1.PSW_cd ;
  wire [7:0] \oc8051_golden_model_1.PSW_ce ;
  wire [7:0] \oc8051_golden_model_1.PSW_cf ;
  wire [7:0] \oc8051_golden_model_1.PSW_d1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_da ;
  wire [7:0] \oc8051_golden_model_1.PSW_db ;
  wire [7:0] \oc8051_golden_model_1.PSW_dc ;
  wire [7:0] \oc8051_golden_model_1.PSW_dd ;
  wire [7:0] \oc8051_golden_model_1.PSW_de ;
  wire [7:0] \oc8051_golden_model_1.PSW_df ;
  wire [7:0] \oc8051_golden_model_1.PSW_e1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_ea ;
  wire [7:0] \oc8051_golden_model_1.PSW_eb ;
  wire [7:0] \oc8051_golden_model_1.PSW_ec ;
  wire [7:0] \oc8051_golden_model_1.PSW_ed ;
  wire [7:0] \oc8051_golden_model_1.PSW_ee ;
  wire [7:0] \oc8051_golden_model_1.PSW_ef ;
  wire [7:0] \oc8051_golden_model_1.PSW_f1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_fa ;
  wire [7:0] \oc8051_golden_model_1.PSW_fb ;
  wire [7:0] \oc8051_golden_model_1.PSW_fc ;
  wire [7:0] \oc8051_golden_model_1.PSW_fd ;
  wire [7:0] \oc8051_golden_model_1.PSW_fe ;
  wire [7:0] \oc8051_golden_model_1.PSW_ff ;
  wire [7:0] \oc8051_golden_model_1.RD_IRAM_0 ;
  wire [7:0] \oc8051_golden_model_1.RD_IRAM_1 ;
  wire [15:0] \oc8051_golden_model_1.RD_ROM_0_ADDR ;
  wire [7:0] \oc8051_golden_model_1.SBUF ;
  wire [7:0] \oc8051_golden_model_1.SCON ;
  wire [7:0] \oc8051_golden_model_1.SP ;
  wire [7:0] \oc8051_golden_model_1.TCON ;
  wire [7:0] \oc8051_golden_model_1.TH0 ;
  wire [7:0] \oc8051_golden_model_1.TH1 ;
  wire [7:0] \oc8051_golden_model_1.TL0 ;
  wire [7:0] \oc8051_golden_model_1.TL1 ;
  wire [7:0] \oc8051_golden_model_1.TMOD ;
  wire \oc8051_golden_model_1.clk ;
  wire [1:0] \oc8051_golden_model_1.n0006 ;
  wire [7:0] \oc8051_golden_model_1.n0007 ;
  wire [7:0] \oc8051_golden_model_1.n0011 ;
  wire [7:0] \oc8051_golden_model_1.n0019 ;
  wire [7:0] \oc8051_golden_model_1.n0023 ;
  wire [7:0] \oc8051_golden_model_1.n0027 ;
  wire [7:0] \oc8051_golden_model_1.n0031 ;
  wire [7:0] \oc8051_golden_model_1.n0035 ;
  wire [7:0] \oc8051_golden_model_1.n0039 ;
  wire [7:0] \oc8051_golden_model_1.n0573 ;
  wire [7:0] \oc8051_golden_model_1.n0606 ;
  wire [15:0] \oc8051_golden_model_1.n0713 ;
  wire [15:0] \oc8051_golden_model_1.n0745 ;
  wire [15:0] \oc8051_golden_model_1.n1004 ;
  wire [6:0] \oc8051_golden_model_1.n1008 ;
  wire \oc8051_golden_model_1.n1009 ;
  wire \oc8051_golden_model_1.n1010 ;
  wire \oc8051_golden_model_1.n1011 ;
  wire \oc8051_golden_model_1.n1012 ;
  wire \oc8051_golden_model_1.n1013 ;
  wire \oc8051_golden_model_1.n1014 ;
  wire \oc8051_golden_model_1.n1015 ;
  wire \oc8051_golden_model_1.n1016 ;
  wire \oc8051_golden_model_1.n1023 ;
  wire [7:0] \oc8051_golden_model_1.n1024 ;
  wire [7:0] \oc8051_golden_model_1.n1031 ;
  wire \oc8051_golden_model_1.n1032 ;
  wire \oc8051_golden_model_1.n1033 ;
  wire \oc8051_golden_model_1.n1034 ;
  wire \oc8051_golden_model_1.n1035 ;
  wire \oc8051_golden_model_1.n1036 ;
  wire \oc8051_golden_model_1.n1037 ;
  wire \oc8051_golden_model_1.n1038 ;
  wire \oc8051_golden_model_1.n1039 ;
  wire \oc8051_golden_model_1.n1046 ;
  wire [7:0] \oc8051_golden_model_1.n1047 ;
  wire \oc8051_golden_model_1.n1063 ;
  wire [7:0] \oc8051_golden_model_1.n1064 ;
  wire [3:0] \oc8051_golden_model_1.n1157 ;
  wire [3:0] \oc8051_golden_model_1.n1159 ;
  wire [3:0] \oc8051_golden_model_1.n1161 ;
  wire [3:0] \oc8051_golden_model_1.n1162 ;
  wire [3:0] \oc8051_golden_model_1.n1163 ;
  wire [3:0] \oc8051_golden_model_1.n1164 ;
  wire [3:0] \oc8051_golden_model_1.n1165 ;
  wire [3:0] \oc8051_golden_model_1.n1166 ;
  wire [3:0] \oc8051_golden_model_1.n1167 ;
  wire \oc8051_golden_model_1.n1214 ;
  wire \oc8051_golden_model_1.n1259 ;
  wire [8:0] \oc8051_golden_model_1.n1260 ;
  wire [8:0] \oc8051_golden_model_1.n1261 ;
  wire [7:0] \oc8051_golden_model_1.n1262 ;
  wire \oc8051_golden_model_1.n1263 ;
  wire [2:0] \oc8051_golden_model_1.n1264 ;
  wire \oc8051_golden_model_1.n1265 ;
  wire [1:0] \oc8051_golden_model_1.n1266 ;
  wire [7:0] \oc8051_golden_model_1.n1267 ;
  wire [6:0] \oc8051_golden_model_1.n1268 ;
  wire \oc8051_golden_model_1.n1269 ;
  wire \oc8051_golden_model_1.n1270 ;
  wire \oc8051_golden_model_1.n1271 ;
  wire \oc8051_golden_model_1.n1272 ;
  wire \oc8051_golden_model_1.n1273 ;
  wire \oc8051_golden_model_1.n1274 ;
  wire \oc8051_golden_model_1.n1275 ;
  wire \oc8051_golden_model_1.n1276 ;
  wire \oc8051_golden_model_1.n1283 ;
  wire [7:0] \oc8051_golden_model_1.n1284 ;
  wire \oc8051_golden_model_1.n1300 ;
  wire [7:0] \oc8051_golden_model_1.n1301 ;
  wire [15:0] \oc8051_golden_model_1.n1343 ;
  wire [7:0] \oc8051_golden_model_1.n1345 ;
  wire \oc8051_golden_model_1.n1346 ;
  wire \oc8051_golden_model_1.n1347 ;
  wire \oc8051_golden_model_1.n1348 ;
  wire \oc8051_golden_model_1.n1349 ;
  wire \oc8051_golden_model_1.n1350 ;
  wire \oc8051_golden_model_1.n1351 ;
  wire \oc8051_golden_model_1.n1352 ;
  wire \oc8051_golden_model_1.n1353 ;
  wire \oc8051_golden_model_1.n1360 ;
  wire [7:0] \oc8051_golden_model_1.n1361 ;
  wire [8:0] \oc8051_golden_model_1.n1363 ;
  wire [8:0] \oc8051_golden_model_1.n1367 ;
  wire \oc8051_golden_model_1.n1368 ;
  wire [3:0] \oc8051_golden_model_1.n1369 ;
  wire [4:0] \oc8051_golden_model_1.n1370 ;
  wire [4:0] \oc8051_golden_model_1.n1374 ;
  wire \oc8051_golden_model_1.n1375 ;
  wire [8:0] \oc8051_golden_model_1.n1376 ;
  wire \oc8051_golden_model_1.n1384 ;
  wire [7:0] \oc8051_golden_model_1.n1385 ;
  wire [6:0] \oc8051_golden_model_1.n1386 ;
  wire \oc8051_golden_model_1.n1401 ;
  wire [7:0] \oc8051_golden_model_1.n1402 ;
  wire [8:0] \oc8051_golden_model_1.n1424 ;
  wire \oc8051_golden_model_1.n1425 ;
  wire [4:0] \oc8051_golden_model_1.n1430 ;
  wire \oc8051_golden_model_1.n1431 ;
  wire \oc8051_golden_model_1.n1439 ;
  wire [7:0] \oc8051_golden_model_1.n1440 ;
  wire [6:0] \oc8051_golden_model_1.n1441 ;
  wire \oc8051_golden_model_1.n1456 ;
  wire [7:0] \oc8051_golden_model_1.n1457 ;
  wire [8:0] \oc8051_golden_model_1.n1459 ;
  wire [8:0] \oc8051_golden_model_1.n1461 ;
  wire \oc8051_golden_model_1.n1462 ;
  wire [3:0] \oc8051_golden_model_1.n1463 ;
  wire [4:0] \oc8051_golden_model_1.n1464 ;
  wire [4:0] \oc8051_golden_model_1.n1466 ;
  wire \oc8051_golden_model_1.n1467 ;
  wire [8:0] \oc8051_golden_model_1.n1468 ;
  wire \oc8051_golden_model_1.n1475 ;
  wire [7:0] \oc8051_golden_model_1.n1476 ;
  wire [6:0] \oc8051_golden_model_1.n1477 ;
  wire \oc8051_golden_model_1.n1492 ;
  wire [7:0] \oc8051_golden_model_1.n1493 ;
  wire [8:0] \oc8051_golden_model_1.n1496 ;
  wire \oc8051_golden_model_1.n1497 ;
  wire \oc8051_golden_model_1.n1504 ;
  wire [7:0] \oc8051_golden_model_1.n1505 ;
  wire [6:0] \oc8051_golden_model_1.n1506 ;
  wire [7:0] \oc8051_golden_model_1.n1507 ;
  wire [8:0] \oc8051_golden_model_1.n1509 ;
  wire [8:0] \oc8051_golden_model_1.n1511 ;
  wire \oc8051_golden_model_1.n1512 ;
  wire [4:0] \oc8051_golden_model_1.n1513 ;
  wire [4:0] \oc8051_golden_model_1.n1515 ;
  wire \oc8051_golden_model_1.n1516 ;
  wire [8:0] \oc8051_golden_model_1.n1517 ;
  wire \oc8051_golden_model_1.n1524 ;
  wire [7:0] \oc8051_golden_model_1.n1525 ;
  wire [6:0] \oc8051_golden_model_1.n1526 ;
  wire \oc8051_golden_model_1.n1541 ;
  wire [7:0] \oc8051_golden_model_1.n1542 ;
  wire [4:0] \oc8051_golden_model_1.n1544 ;
  wire \oc8051_golden_model_1.n1545 ;
  wire [7:0] \oc8051_golden_model_1.n1546 ;
  wire [6:0] \oc8051_golden_model_1.n1547 ;
  wire [7:0] \oc8051_golden_model_1.n1548 ;
  wire [8:0] \oc8051_golden_model_1.n1550 ;
  wire \oc8051_golden_model_1.n1551 ;
  wire \oc8051_golden_model_1.n1558 ;
  wire [7:0] \oc8051_golden_model_1.n1559 ;
  wire [6:0] \oc8051_golden_model_1.n1560 ;
  wire [7:0] \oc8051_golden_model_1.n1561 ;
  wire [7:0] \oc8051_golden_model_1.n1562 ;
  wire [6:0] \oc8051_golden_model_1.n1563 ;
  wire [7:0] \oc8051_golden_model_1.n1564 ;
  wire [8:0] \oc8051_golden_model_1.n1567 ;
  wire [8:0] \oc8051_golden_model_1.n1568 ;
  wire [7:0] \oc8051_golden_model_1.n1569 ;
  wire [7:0] \oc8051_golden_model_1.n1570 ;
  wire [6:0] \oc8051_golden_model_1.n1571 ;
  wire \oc8051_golden_model_1.n1572 ;
  wire \oc8051_golden_model_1.n1573 ;
  wire \oc8051_golden_model_1.n1574 ;
  wire \oc8051_golden_model_1.n1575 ;
  wire \oc8051_golden_model_1.n1576 ;
  wire \oc8051_golden_model_1.n1577 ;
  wire \oc8051_golden_model_1.n1578 ;
  wire \oc8051_golden_model_1.n1579 ;
  wire \oc8051_golden_model_1.n1586 ;
  wire [7:0] \oc8051_golden_model_1.n1587 ;
  wire [7:0] \oc8051_golden_model_1.n1588 ;
  wire [8:0] \oc8051_golden_model_1.n1591 ;
  wire [8:0] \oc8051_golden_model_1.n1593 ;
  wire \oc8051_golden_model_1.n1594 ;
  wire [4:0] \oc8051_golden_model_1.n1595 ;
  wire [4:0] \oc8051_golden_model_1.n1597 ;
  wire \oc8051_golden_model_1.n1598 ;
  wire \oc8051_golden_model_1.n1605 ;
  wire [7:0] \oc8051_golden_model_1.n1606 ;
  wire [6:0] \oc8051_golden_model_1.n1607 ;
  wire \oc8051_golden_model_1.n1622 ;
  wire [7:0] \oc8051_golden_model_1.n1623 ;
  wire [8:0] \oc8051_golden_model_1.n1627 ;
  wire \oc8051_golden_model_1.n1628 ;
  wire [4:0] \oc8051_golden_model_1.n1630 ;
  wire \oc8051_golden_model_1.n1631 ;
  wire \oc8051_golden_model_1.n1638 ;
  wire [7:0] \oc8051_golden_model_1.n1639 ;
  wire [6:0] \oc8051_golden_model_1.n1640 ;
  wire \oc8051_golden_model_1.n1655 ;
  wire [7:0] \oc8051_golden_model_1.n1656 ;
  wire [8:0] \oc8051_golden_model_1.n1660 ;
  wire \oc8051_golden_model_1.n1661 ;
  wire [4:0] \oc8051_golden_model_1.n1663 ;
  wire \oc8051_golden_model_1.n1664 ;
  wire \oc8051_golden_model_1.n1671 ;
  wire [7:0] \oc8051_golden_model_1.n1672 ;
  wire [6:0] \oc8051_golden_model_1.n1673 ;
  wire \oc8051_golden_model_1.n1688 ;
  wire [7:0] \oc8051_golden_model_1.n1689 ;
  wire [8:0] \oc8051_golden_model_1.n1693 ;
  wire \oc8051_golden_model_1.n1694 ;
  wire [4:0] \oc8051_golden_model_1.n1696 ;
  wire \oc8051_golden_model_1.n1697 ;
  wire \oc8051_golden_model_1.n1704 ;
  wire [7:0] \oc8051_golden_model_1.n1705 ;
  wire [6:0] \oc8051_golden_model_1.n1706 ;
  wire \oc8051_golden_model_1.n1721 ;
  wire [7:0] \oc8051_golden_model_1.n1722 ;
  wire [7:0] \oc8051_golden_model_1.n1747 ;
  wire [6:0] \oc8051_golden_model_1.n1748 ;
  wire [7:0] \oc8051_golden_model_1.n1749 ;
  wire \oc8051_golden_model_1.n1804 ;
  wire [7:0] \oc8051_golden_model_1.n1805 ;
  wire \oc8051_golden_model_1.n1821 ;
  wire [7:0] \oc8051_golden_model_1.n1822 ;
  wire \oc8051_golden_model_1.n1838 ;
  wire [7:0] \oc8051_golden_model_1.n1839 ;
  wire \oc8051_golden_model_1.n1855 ;
  wire [7:0] \oc8051_golden_model_1.n1856 ;
  wire [7:0] \oc8051_golden_model_1.n1879 ;
  wire [6:0] \oc8051_golden_model_1.n1880 ;
  wire [7:0] \oc8051_golden_model_1.n1881 ;
  wire \oc8051_golden_model_1.n1936 ;
  wire [7:0] \oc8051_golden_model_1.n1937 ;
  wire \oc8051_golden_model_1.n1953 ;
  wire [7:0] \oc8051_golden_model_1.n1954 ;
  wire \oc8051_golden_model_1.n1970 ;
  wire [7:0] \oc8051_golden_model_1.n1971 ;
  wire \oc8051_golden_model_1.n1987 ;
  wire [7:0] \oc8051_golden_model_1.n1988 ;
  wire \oc8051_golden_model_1.n2085 ;
  wire [7:0] \oc8051_golden_model_1.n2086 ;
  wire \oc8051_golden_model_1.n2102 ;
  wire [7:0] \oc8051_golden_model_1.n2103 ;
  wire \oc8051_golden_model_1.n2119 ;
  wire [7:0] \oc8051_golden_model_1.n2120 ;
  wire \oc8051_golden_model_1.n2136 ;
  wire [7:0] \oc8051_golden_model_1.n2137 ;
  wire \oc8051_golden_model_1.n2141 ;
  wire [6:0] \oc8051_golden_model_1.n2142 ;
  wire [7:0] \oc8051_golden_model_1.n2143 ;
  wire [6:0] \oc8051_golden_model_1.n2144 ;
  wire [7:0] \oc8051_golden_model_1.n2145 ;
  wire \oc8051_golden_model_1.n2160 ;
  wire [7:0] \oc8051_golden_model_1.n2161 ;
  wire \oc8051_golden_model_1.n2200 ;
  wire [7:0] \oc8051_golden_model_1.n2201 ;
  wire [6:0] \oc8051_golden_model_1.n2202 ;
  wire [7:0] \oc8051_golden_model_1.n2203 ;
  wire [3:0] \oc8051_golden_model_1.n2210 ;
  wire \oc8051_golden_model_1.n2211 ;
  wire [7:0] \oc8051_golden_model_1.n2212 ;
  wire [6:0] \oc8051_golden_model_1.n2213 ;
  wire \oc8051_golden_model_1.n2228 ;
  wire [7:0] \oc8051_golden_model_1.n2229 ;
  wire [7:0] \oc8051_golden_model_1.n2441 ;
  wire \oc8051_golden_model_1.n2444 ;
  wire \oc8051_golden_model_1.n2446 ;
  wire \oc8051_golden_model_1.n2452 ;
  wire [7:0] \oc8051_golden_model_1.n2453 ;
  wire [6:0] \oc8051_golden_model_1.n2454 ;
  wire \oc8051_golden_model_1.n2469 ;
  wire [7:0] \oc8051_golden_model_1.n2470 ;
  wire \oc8051_golden_model_1.n2474 ;
  wire \oc8051_golden_model_1.n2476 ;
  wire \oc8051_golden_model_1.n2482 ;
  wire [7:0] \oc8051_golden_model_1.n2483 ;
  wire [6:0] \oc8051_golden_model_1.n2484 ;
  wire \oc8051_golden_model_1.n2499 ;
  wire [7:0] \oc8051_golden_model_1.n2500 ;
  wire \oc8051_golden_model_1.n2504 ;
  wire \oc8051_golden_model_1.n2506 ;
  wire \oc8051_golden_model_1.n2512 ;
  wire [7:0] \oc8051_golden_model_1.n2513 ;
  wire [6:0] \oc8051_golden_model_1.n2514 ;
  wire \oc8051_golden_model_1.n2529 ;
  wire [7:0] \oc8051_golden_model_1.n2530 ;
  wire \oc8051_golden_model_1.n2534 ;
  wire \oc8051_golden_model_1.n2536 ;
  wire \oc8051_golden_model_1.n2542 ;
  wire [7:0] \oc8051_golden_model_1.n2543 ;
  wire [6:0] \oc8051_golden_model_1.n2544 ;
  wire \oc8051_golden_model_1.n2559 ;
  wire [7:0] \oc8051_golden_model_1.n2560 ;
  wire \oc8051_golden_model_1.n2562 ;
  wire [7:0] \oc8051_golden_model_1.n2563 ;
  wire [6:0] \oc8051_golden_model_1.n2564 ;
  wire [7:0] \oc8051_golden_model_1.n2565 ;
  wire [7:0] \oc8051_golden_model_1.n2566 ;
  wire [6:0] \oc8051_golden_model_1.n2567 ;
  wire [7:0] \oc8051_golden_model_1.n2568 ;
  wire [15:0] \oc8051_golden_model_1.n2572 ;
  wire \oc8051_golden_model_1.n2578 ;
  wire [7:0] \oc8051_golden_model_1.n2579 ;
  wire [6:0] \oc8051_golden_model_1.n2580 ;
  wire \oc8051_golden_model_1.n2595 ;
  wire [7:0] \oc8051_golden_model_1.n2596 ;
  wire \oc8051_golden_model_1.n2599 ;
  wire [7:0] \oc8051_golden_model_1.n2600 ;
  wire [6:0] \oc8051_golden_model_1.n2601 ;
  wire [7:0] \oc8051_golden_model_1.n2602 ;
  wire \oc8051_golden_model_1.n2634 ;
  wire [7:0] \oc8051_golden_model_1.n2635 ;
  wire [6:0] \oc8051_golden_model_1.n2636 ;
  wire [7:0] \oc8051_golden_model_1.n2637 ;
  wire \oc8051_golden_model_1.n2642 ;
  wire [7:0] \oc8051_golden_model_1.n2643 ;
  wire [6:0] \oc8051_golden_model_1.n2644 ;
  wire [7:0] \oc8051_golden_model_1.n2645 ;
  wire \oc8051_golden_model_1.n2650 ;
  wire [7:0] \oc8051_golden_model_1.n2651 ;
  wire [6:0] \oc8051_golden_model_1.n2652 ;
  wire [7:0] \oc8051_golden_model_1.n2653 ;
  wire \oc8051_golden_model_1.n2658 ;
  wire [7:0] \oc8051_golden_model_1.n2659 ;
  wire [6:0] \oc8051_golden_model_1.n2660 ;
  wire [7:0] \oc8051_golden_model_1.n2661 ;
  wire \oc8051_golden_model_1.n2666 ;
  wire [7:0] \oc8051_golden_model_1.n2667 ;
  wire [6:0] \oc8051_golden_model_1.n2668 ;
  wire [7:0] \oc8051_golden_model_1.n2669 ;
  wire [7:0] \oc8051_golden_model_1.n2694 ;
  wire [6:0] \oc8051_golden_model_1.n2695 ;
  wire [7:0] \oc8051_golden_model_1.n2696 ;
  wire [3:0] \oc8051_golden_model_1.n2697 ;
  wire [7:0] \oc8051_golden_model_1.n2698 ;
  wire \oc8051_golden_model_1.n2699 ;
  wire \oc8051_golden_model_1.n2700 ;
  wire \oc8051_golden_model_1.n2701 ;
  wire \oc8051_golden_model_1.n2702 ;
  wire \oc8051_golden_model_1.n2703 ;
  wire \oc8051_golden_model_1.n2704 ;
  wire \oc8051_golden_model_1.n2705 ;
  wire \oc8051_golden_model_1.n2706 ;
  wire \oc8051_golden_model_1.n2713 ;
  wire [7:0] \oc8051_golden_model_1.n2714 ;
  wire [7:0] \oc8051_golden_model_1.n2734 ;
  wire [6:0] \oc8051_golden_model_1.n2735 ;
  wire \oc8051_golden_model_1.n2750 ;
  wire [7:0] \oc8051_golden_model_1.n2751 ;
  wire \oc8051_golden_model_1.n2752 ;
  wire \oc8051_golden_model_1.n2753 ;
  wire \oc8051_golden_model_1.n2754 ;
  wire \oc8051_golden_model_1.n2755 ;
  wire \oc8051_golden_model_1.n2756 ;
  wire \oc8051_golden_model_1.n2757 ;
  wire \oc8051_golden_model_1.n2758 ;
  wire \oc8051_golden_model_1.n2759 ;
  wire \oc8051_golden_model_1.n2766 ;
  wire [7:0] \oc8051_golden_model_1.n2767 ;
  wire \oc8051_golden_model_1.n2768 ;
  wire \oc8051_golden_model_1.n2769 ;
  wire \oc8051_golden_model_1.n2770 ;
  wire \oc8051_golden_model_1.n2771 ;
  wire \oc8051_golden_model_1.n2772 ;
  wire \oc8051_golden_model_1.n2773 ;
  wire \oc8051_golden_model_1.n2774 ;
  wire \oc8051_golden_model_1.n2775 ;
  wire \oc8051_golden_model_1.n2782 ;
  wire [7:0] \oc8051_golden_model_1.n2783 ;
  wire [7:0] \oc8051_golden_model_1.n2815 ;
  wire [6:0] \oc8051_golden_model_1.n2816 ;
  wire [7:0] \oc8051_golden_model_1.n2817 ;
  wire \oc8051_golden_model_1.n2836 ;
  wire [7:0] \oc8051_golden_model_1.n2837 ;
  wire [6:0] \oc8051_golden_model_1.n2838 ;
  wire \oc8051_golden_model_1.n2853 ;
  wire [7:0] \oc8051_golden_model_1.n2854 ;
  wire [7:0] \oc8051_golden_model_1.n2858 ;
  wire [3:0] \oc8051_golden_model_1.n2859 ;
  wire [7:0] \oc8051_golden_model_1.n2860 ;
  wire \oc8051_golden_model_1.n2861 ;
  wire \oc8051_golden_model_1.n2862 ;
  wire \oc8051_golden_model_1.n2863 ;
  wire \oc8051_golden_model_1.n2864 ;
  wire \oc8051_golden_model_1.n2865 ;
  wire \oc8051_golden_model_1.n2866 ;
  wire \oc8051_golden_model_1.n2867 ;
  wire \oc8051_golden_model_1.n2868 ;
  wire \oc8051_golden_model_1.n2875 ;
  wire [7:0] \oc8051_golden_model_1.n2876 ;
  wire \oc8051_golden_model_1.n2894 ;
  wire [7:0] \oc8051_golden_model_1.n2895 ;
  wire [7:0] \oc8051_golden_model_1.n2896 ;
  wire \oc8051_golden_model_1.n2912 ;
  wire [7:0] \oc8051_golden_model_1.n2913 ;
  wire [7:0] \oc8051_golden_model_1.n2914 ;
  wire \oc8051_golden_model_1.rst ;
  wire [34:0] \oc8051_top_1.ABINPUT ;
  wire [7:0] \oc8051_top_1.acc ;
  wire [7:0] \oc8051_top_1.b_reg ;
  wire [31:0] \oc8051_top_1.cxrom_data_out ;
  wire \oc8051_top_1.cy ;
  wire [1:0] \oc8051_top_1.cy_sel ;
  wire [7:0] \oc8051_top_1.des1 ;
  wire [7:0] \oc8051_top_1.des2 ;
  wire \oc8051_top_1.desAc ;
  wire \oc8051_top_1.desCy ;
  wire \oc8051_top_1.desOv ;
  wire [7:0] \oc8051_top_1.des_acc ;
  wire [15:0] \oc8051_top_1.dptr ;
  wire [7:0] \oc8051_top_1.dptr_hi ;
  wire [7:0] \oc8051_top_1.dptr_lo ;
  wire \oc8051_top_1.ea_int ;
  wire [31:0] \oc8051_top_1.idat_onchip ;
  wire [7:0] \oc8051_top_1.ie ;
  wire \oc8051_top_1.int_ack ;
  wire [7:0] \oc8051_top_1.int_src ;
  wire \oc8051_top_1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.acc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.clk ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.dptr ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op1_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op2_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op3_r ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.pc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_alu_src_sel1.sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_alu_src_sel1.sel2 ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.sel3 ;
  wire [7:0] \oc8051_top_1.oc8051_comp1.acc ;
  wire \oc8051_top_1.oc8051_comp1.cy ;
  wire [7:0] \oc8051_top_1.oc8051_comp1.des ;
  wire \oc8051_top_1.oc8051_cy_select1.cy_in ;
  wire [1:0] \oc8051_top_1.oc8051_cy_select1.cy_sel ;
  wire [3:0] \oc8051_top_1.oc8051_decoder1.alu_op ;
  wire \oc8051_top_1.oc8051_decoder1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.cy_sel ;
  wire \oc8051_top_1.oc8051_decoder1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_decoder1.op ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.psw_set ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_wr_sel ;
  wire \oc8051_top_1.oc8051_decoder1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.src_sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.src_sel2 ;
  wire \oc8051_top_1.oc8051_decoder1.src_sel3 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.state ;
  wire \oc8051_top_1.oc8051_decoder1.wait_data ;
  wire \oc8051_top_1.oc8051_decoder1.wr ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.wr_sfr ;
  wire \oc8051_top_1.oc8051_indi_addr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.data_in ;
  wire \oc8051_top_1.oc8051_indi_addr1.rst ;
  wire \oc8051_top_1.oc8051_indi_addr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.acc ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.alu ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.cdata ;
  wire \oc8051_top_1.oc8051_memory_interface1.cdone ;
  wire \oc8051_top_1.oc8051_memory_interface1.clk ;
  wire \oc8051_top_1.oc8051_memory_interface1.dack_ir ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dadr_o ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dadr_ot ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_ir ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_o ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.des1 ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.des2 ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.des_acc ;
  wire \oc8051_top_1.oc8051_memory_interface1.dmem_wait ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dptr ;
  wire \oc8051_top_1.oc8051_memory_interface1.dstb_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.dwe_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.ea_int ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.iadr_t ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_cur ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_old ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_onchip ;
  wire \oc8051_top_1.oc8051_memory_interface1.imem_wait ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm2_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_t ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_v ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_vec_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.istb_t ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op2_buff ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op3_buff ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.op_pos ;
  wire \oc8051_top_1.oc8051_memory_interface1.out_of_rst ;
  wire [3:0] \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_buf ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log_prev ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_addr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_ind ;
  wire \oc8051_top_1.oc8051_memory_interface1.reti ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ri_r ;
  wire [4:0] \oc8051_top_1.oc8051_memory_interface1.rn_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.sfr ;
  wire \oc8051_top_1.oc8051_memory_interface1.sfr_bit ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.wr_dat ;
  wire \oc8051_top_1.oc8051_ram_top1.bit_addr_r ;
  wire \oc8051_top_1.oc8051_ram_top1.bit_data_in ;
  wire [2:0] \oc8051_top_1.oc8051_ram_top1.bit_select ;
  wire \oc8051_top_1.oc8051_ram_top1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.rd_data_m ;
  wire \oc8051_top_1.oc8051_ram_top1.rd_en_r ;
  wire \oc8051_top_1.oc8051_ram_top1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.wr_data ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.wr_data_r ;
  wire \oc8051_top_1.oc8051_rom1.clk ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.cxrom_data_out ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.data_o ;
  wire \oc8051_top_1.oc8051_rom1.ea_int ;
  wire \oc8051_top_1.oc8051_rom1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.b_reg ;
  wire \oc8051_top_1.oc8051_sfr1.bit_in ;
  wire \oc8051_top_1.oc8051_sfr1.bit_out ;
  wire \oc8051_top_1.oc8051_sfr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.cy ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat2 ;
  wire \oc8051_top_1.oc8051_sfr1.desAc ;
  wire \oc8051_top_1.oc8051_sfr1.desOv ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.des_acc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_lo ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.int_ack ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ip ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.bit_in ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.p ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.bit_in ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ack ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.bit_in ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.data_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie1_buff ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.bit_in ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.data_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.ac_in ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.cy_in ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.ov_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.set ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.data_in ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.p ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw_next ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.psw_set ;
  wire \oc8051_top_1.oc8051_sfr1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.srcAc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.wait_data ;
  wire \oc8051_top_1.oc8051_sfr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.p0_o ;
  wire [7:0] \oc8051_top_1.p1_o ;
  wire [7:0] \oc8051_top_1.p2_o ;
  wire [7:0] \oc8051_top_1.p3_o ;
  wire [15:0] \oc8051_top_1.pc ;
  wire [15:0] \oc8051_top_1.pc_log ;
  wire [15:0] \oc8051_top_1.pc_log_prev ;
  wire [7:0] \oc8051_top_1.psw ;
  wire [1:0] \oc8051_top_1.psw_set ;
  wire \oc8051_top_1.rd_ind ;
  wire \oc8051_top_1.reti ;
  wire \oc8051_top_1.sfr_bit ;
  wire [7:0] \oc8051_top_1.sfr_out ;
  wire \oc8051_top_1.srcAc ;
  wire [2:0] \oc8051_top_1.src_sel1 ;
  wire [1:0] \oc8051_top_1.src_sel2 ;
  wire \oc8051_top_1.src_sel3 ;
  wire [7:0] \oc8051_top_1.sub_result ;
  wire \oc8051_top_1.wait_data ;
  wire \oc8051_top_1.wb_clk_i ;
  wire \oc8051_top_1.wb_rst_i ;
  wire [15:0] \oc8051_top_1.wbd_adr_o ;
  wire \oc8051_top_1.wbd_cyc_o ;
  wire [7:0] \oc8051_top_1.wbd_dat_o ;
  wire \oc8051_top_1.wbd_stb_o ;
  wire \oc8051_top_1.wbd_we_o ;
  wire [7:0] \oc8051_top_1.wr_dat ;
  input [7:0] p0_in;
  wire [7:0] p0_out;
  wire [7:0] p0in_reg;
  input [7:0] p1_in;
  wire [7:0] p1_out;
  wire [7:0] p1in_reg;
  input [7:0] p2_in;
  wire [7:0] p2_out;
  wire [7:0] p2in_reg;
  input [7:0] p3_in;
  wire [7:0] p3_out;
  wire [7:0] p3in_reg;
  wire [15:0] pc_impl;
  output property_invalid_rom_pc;
  wire [7:0] psw_impl;
  wire [15:0] rd_rom_0_addr;
  input rst;
  wire [15:0] wbd_adr_o;
  wire wbd_cyc_o;
  wire [7:0] wbd_dat_o;
  wire wbd_stb_o;
  wire wbd_we_o;
  input [127:0] word_in;
  not (_37580_, rst);
  not (_15554_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  not (_15565_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_15576_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _15565_);
  and (_15596_, _15576_, _15554_);
  and (_15597_, \oc8051_top_1.oc8051_decoder1.wr , _15565_);
  not (_15608_, _15597_);
  nor (_15619_, _15608_, _15596_);
  and (_15630_, _15619_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_15641_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and (_15652_, _15641_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  and (_15663_, _15652_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  and (_15674_, _15663_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  and (_15684_, _15674_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  not (_15695_, _15684_);
  and (_15706_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _15565_);
  and (_15717_, _15706_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  and (_15728_, _15717_, _15554_);
  not (_15739_, _15728_);
  nor (_15750_, _15674_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor (_15761_, _15750_, _15739_);
  and (_15772_, _15761_, _15695_);
  not (_15782_, _15772_);
  not (_15793_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  and (_15804_, _15706_, _15793_);
  and (_15815_, _15804_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_15826_, _15815_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [5]);
  and (_15837_, _15804_, _15554_);
  and (_15848_, _15837_, \oc8051_top_1.oc8051_memory_interface1.imm_r [5]);
  nor (_15859_, _15848_, _15826_);
  and (_15869_, _15717_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  nor (_15880_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_15891_, _15880_, _15576_);
  and (_15902_, _15891_, \oc8051_top_1.oc8051_memory_interface1.ri_r [5]);
  nor (_15913_, _15902_, _15869_);
  and (_15924_, _15913_, _15859_);
  and (_15935_, _15924_, _15782_);
  and (_15946_, _15684_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  not (_15957_, _15946_);
  nor (_15967_, _15684_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor (_15978_, _15967_, _15739_);
  and (_15989_, _15978_, _15957_);
  not (_16000_, _15989_);
  and (_16011_, _15837_, \oc8051_top_1.oc8051_memory_interface1.imm_r [6]);
  nor (_16022_, _16011_, _15869_);
  and (_16043_, _15891_, \oc8051_top_1.oc8051_memory_interface1.ri_r [6]);
  and (_16044_, _15815_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [6]);
  nor (_16055_, _16044_, _16043_);
  and (_16065_, _16055_, _16022_);
  and (_16076_, _16065_, _16000_);
  nor (_16087_, _16076_, _15935_);
  not (_16098_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  nor (_16109_, _15946_, _16098_);
  and (_16120_, _15946_, _16098_);
  nor (_16131_, _16120_, _16109_);
  nor (_16142_, _16131_, _15739_);
  not (_16152_, _16142_);
  and (_16163_, _15891_, \oc8051_top_1.oc8051_memory_interface1.ri_r [7]);
  not (_16174_, _16163_);
  not (_16185_, _15869_);
  and (_16196_, _15837_, \oc8051_top_1.oc8051_memory_interface1.imm_r [7]);
  and (_16207_, _15815_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [7]);
  nor (_16218_, _16207_, _16196_);
  and (_16229_, _16218_, _16185_);
  and (_16239_, _16229_, _16174_);
  and (_16250_, _16239_, _16152_);
  not (_16261_, _16250_);
  not (_16272_, _15663_);
  nor (_16283_, _15652_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor (_16294_, _16283_, _15739_);
  and (_16305_, _16294_, _16272_);
  not (_16316_, _16305_);
  and (_16327_, _15815_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [3]);
  nor (_16337_, _15880_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_16348_, _16337_, _15576_);
  and (_16359_, _16348_, \oc8051_top_1.oc8051_memory_interface1.rn_r [3]);
  nor (_16370_, _16359_, _16327_);
  and (_16381_, _15837_, \oc8051_top_1.oc8051_memory_interface1.imm_r [3]);
  and (_16392_, _15891_, \oc8051_top_1.oc8051_memory_interface1.ri_r [3]);
  nor (_16403_, _16392_, _16381_);
  and (_16414_, _16403_, _16370_);
  and (_16425_, _16414_, _16316_);
  not (_16435_, _16425_);
  and (_16446_, _15815_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [4]);
  not (_16457_, _16446_);
  and (_16468_, _15891_, \oc8051_top_1.oc8051_memory_interface1.ri_r [4]);
  nor (_16479_, _16468_, _15869_);
  and (_16490_, _16479_, _16457_);
  nor (_16501_, _15663_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  not (_16512_, _16501_);
  nor (_16522_, _15739_, _15674_);
  and (_16533_, _16522_, _16512_);
  and (_16544_, _16348_, \oc8051_top_1.oc8051_memory_interface1.rn_r [4]);
  and (_16555_, _15837_, \oc8051_top_1.oc8051_memory_interface1.imm_r [4]);
  nor (_16566_, _16555_, _16544_);
  not (_16577_, _16566_);
  nor (_16588_, _16577_, _16533_);
  and (_16599_, _16588_, _16490_);
  nor (_16610_, _16599_, _16435_);
  and (_16620_, _16610_, _16261_);
  and (_16631_, _16620_, _16087_);
  nor (_16642_, _15641_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_16653_, _16642_, _15652_);
  and (_16674_, _16653_, _15728_);
  and (_16675_, _15891_, \oc8051_top_1.oc8051_memory_interface1.ri_r [2]);
  nor (_16686_, _16675_, _16674_);
  and (_16697_, _15815_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [2]);
  and (_16707_, _15837_, \oc8051_top_1.oc8051_memory_interface1.imm_r [2]);
  and (_16718_, _16348_, \oc8051_top_1.oc8051_memory_interface1.rn_r [2]);
  or (_16729_, _16718_, _16707_);
  nor (_16740_, _16729_, _16697_);
  and (_16751_, _16740_, _16686_);
  not (_16762_, _16751_);
  and (_16773_, _15837_, \oc8051_top_1.oc8051_memory_interface1.imm_r [0]);
  and (_16784_, _15891_, \oc8051_top_1.oc8051_memory_interface1.ri_r [0]);
  nor (_16795_, _16784_, _16773_);
  and (_16805_, _15815_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [0]);
  not (_16816_, _16805_);
  not (_16827_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and (_16838_, _15728_, _16827_);
  and (_16849_, _16348_, \oc8051_top_1.oc8051_memory_interface1.rn_r [0]);
  nor (_16860_, _16849_, _16838_);
  and (_16871_, _16860_, _16816_);
  and (_16882_, _16871_, _16795_);
  and (_16893_, _15815_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [1]);
  nor (_16904_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  nor (_16914_, _16904_, _15641_);
  and (_16925_, _16914_, _15728_);
  nor (_16936_, _16925_, _16893_);
  and (_16947_, _15891_, \oc8051_top_1.oc8051_memory_interface1.ri_r [1]);
  and (_16958_, _16348_, \oc8051_top_1.oc8051_memory_interface1.rn_r [1]);
  and (_16969_, _15837_, \oc8051_top_1.oc8051_memory_interface1.imm_r [1]);
  or (_16980_, _16969_, _16958_);
  nor (_16991_, _16980_, _16947_);
  and (_17002_, _16991_, _16936_);
  nor (_17013_, _17002_, _16882_);
  and (_17023_, _17013_, _16762_);
  and (_17034_, _17023_, _16631_);
  or (_17055_, _17034_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  not (_17056_, ABINPUT[0]);
  nand (_17067_, _17034_, _17056_);
  and (_17078_, _17067_, _17055_);
  and (_17089_, _17078_, _15630_);
  not (_17100_, _15619_);
  and (_17111_, _17100_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  not (_17122_, ABINPUT[26]);
  and (_17132_, _17002_, _16882_);
  and (_17143_, _17132_, _16751_);
  and (_17154_, _17143_, _16631_);
  nand (_17165_, _17154_, _17122_);
  not (_17176_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_17187_, _15619_, _17176_);
  or (_17198_, _17154_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_17209_, _17198_, _17187_);
  and (_17220_, _17209_, _17165_);
  or (_17231_, _17220_, _17111_);
  or (_17241_, _17231_, _17089_);
  and (_05323_, _17241_, _37580_);
  not (_17262_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nor (_17273_, _17154_, _17262_);
  and (_17284_, _17143_, ABINPUT[0]);
  and (_17295_, _17284_, _16631_);
  or (_17306_, _17295_, _17273_);
  and (_17317_, _17306_, _15630_);
  nor (_17328_, _15619_, _17262_);
  and (_17339_, _17154_, ABINPUT[19]);
  or (_17350_, _17339_, _17273_);
  and (_17360_, _17350_, _17187_);
  or (_17371_, _17360_, _17328_);
  or (_17382_, _17371_, _17317_);
  and (_29076_, _17382_, _37580_);
  not (_17403_, _16882_);
  and (_17414_, _17002_, _17403_);
  and (_17425_, _17414_, _16751_);
  nand (_17436_, _17425_, _16631_);
  and (_17447_, _17436_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_17467_, _17425_, ABINPUT[0]);
  and (_17468_, _17467_, _16631_);
  or (_17479_, _17468_, _17447_);
  and (_17490_, _17479_, _15630_);
  and (_17501_, _17100_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  not (_17512_, ABINPUT[20]);
  nand (_17523_, _17154_, _17512_);
  or (_17534_, _17154_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_17545_, _17534_, _17187_);
  and (_17556_, _17545_, _17523_);
  or (_17567_, _17556_, _17501_);
  or (_17577_, _17567_, _17490_);
  and (_29184_, _17577_, _37580_);
  not (_17598_, _17002_);
  and (_17609_, _17598_, _16882_);
  and (_17620_, _17609_, _16751_);
  nand (_17631_, _17620_, _16631_);
  and (_17642_, _17631_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_17653_, _17620_, ABINPUT[0]);
  and (_17664_, _17653_, _16631_);
  or (_17675_, _17664_, _17642_);
  and (_17685_, _17675_, _15630_);
  and (_17696_, _17100_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  not (_17707_, ABINPUT[21]);
  nand (_17718_, _17154_, _17707_);
  or (_17729_, _17154_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_17740_, _17729_, _17187_);
  and (_17751_, _17740_, _17718_);
  or (_17762_, _17751_, _17696_);
  or (_17773_, _17762_, _17685_);
  and (_29294_, _17773_, _37580_);
  and (_17793_, _17013_, _16751_);
  nand (_17804_, _17793_, _16631_);
  and (_17815_, _17804_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_17826_, _17793_, ABINPUT[0]);
  and (_17837_, _17826_, _16631_);
  or (_17848_, _17837_, _17815_);
  and (_17859_, _17848_, _15630_);
  and (_17870_, _17100_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  not (_17891_, ABINPUT[22]);
  nand (_17892_, _17154_, _17891_);
  or (_17902_, _17154_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_17913_, _17902_, _17187_);
  and (_17924_, _17913_, _17892_);
  or (_17935_, _17924_, _17870_);
  or (_17946_, _17935_, _17859_);
  and (_29403_, _17946_, _37580_);
  and (_17967_, _17132_, _16762_);
  nand (_17978_, _17967_, _16631_);
  and (_17989_, _17978_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_18000_, _17967_, ABINPUT[0]);
  and (_18010_, _18000_, _16631_);
  or (_18021_, _18010_, _17989_);
  and (_18032_, _18021_, _15630_);
  and (_18043_, _17100_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  not (_18054_, ABINPUT[23]);
  nand (_18065_, _17154_, _18054_);
  or (_18076_, _17154_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_18087_, _18076_, _17187_);
  and (_18098_, _18087_, _18065_);
  or (_18109_, _18098_, _18043_);
  or (_18119_, _18109_, _18032_);
  and (_29511_, _18119_, _37580_);
  and (_18140_, _17414_, _16762_);
  nand (_18151_, _18140_, _16631_);
  and (_18162_, _18151_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_18173_, _18140_, ABINPUT[0]);
  and (_18184_, _18173_, _16631_);
  or (_18195_, _18184_, _18162_);
  and (_18206_, _18195_, _15630_);
  and (_18217_, _17100_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  not (_18228_, ABINPUT[24]);
  nand (_18238_, _17154_, _18228_);
  or (_18249_, _17154_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_18260_, _18249_, _17187_);
  and (_18271_, _18260_, _18238_);
  or (_18282_, _18271_, _18217_);
  or (_18293_, _18282_, _18206_);
  and (_29620_, _18293_, _37580_);
  and (_18314_, _17609_, _16762_);
  nand (_18325_, _18314_, _16631_);
  and (_18345_, _18325_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_18346_, _18314_, ABINPUT[0]);
  and (_18357_, _18346_, _16631_);
  or (_18368_, _18357_, _18345_);
  and (_18379_, _18368_, _15630_);
  and (_18390_, _17100_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  not (_18401_, ABINPUT[25]);
  nand (_18412_, _17154_, _18401_);
  or (_18423_, _17154_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_18434_, _18423_, _17187_);
  and (_18445_, _18434_, _18412_);
  or (_18456_, _18445_, _18390_);
  or (_18466_, _18456_, _18379_);
  and (_29730_, _18466_, _37580_);
  and (_18487_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_18498_, \oc8051_top_1.oc8051_decoder1.state [0], \oc8051_top_1.oc8051_decoder1.state [1]);
  nor (_18509_, _18498_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_18520_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  nor (_18531_, \oc8051_top_1.oc8051_memory_interface1.imem_wait , \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and (_18542_, _18531_, _18520_);
  and (_18553_, _18498_, _15565_);
  and (_18564_, _18553_, _18542_);
  and (_18575_, _18542_, \oc8051_top_1.oc8051_decoder1.op [2]);
  nor (_18585_, _18575_, _18564_);
  and (_18596_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_18607_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], \oc8051_top_1.oc8051_memory_interface1.cdone );
  not (_18618_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_18629_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_18640_, _18629_, _18618_);
  and (_18651_, _18640_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  not (_18662_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_18673_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], _18662_);
  and (_18684_, _18673_, _18618_);
  and (_18695_, _18684_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_18706_, _18695_, _18651_);
  nor (_18716_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_18727_, _18716_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_18738_, _18727_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  not (_18749_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_18760_, _18749_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_18771_, _18760_, _18618_);
  and (_18782_, _18771_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  nor (_18793_, _18782_, _18738_);
  and (_18804_, _18793_, _18706_);
  nor (_18825_, _18716_, _18618_);
  and (_18826_, _18825_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_18836_, _18716_, _18618_);
  and (_18847_, _18836_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  nor (_18858_, _18847_, _18826_);
  and (_18869_, _18858_, _18804_);
  and (_18880_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  or (_18891_, _18880_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor (_18902_, _18891_, _18869_);
  nor (_18913_, _18902_, _18607_);
  nor (_18924_, _18913_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_18935_, _18924_, _18596_);
  and (_18946_, _18935_, _18564_);
  nor (_18957_, _18946_, _18585_);
  and (_18967_, _18542_, \oc8051_top_1.oc8051_decoder1.op [3]);
  nor (_18978_, _18967_, _18564_);
  and (_18989_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_19000_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], \oc8051_top_1.oc8051_memory_interface1.cdone );
  not (_19011_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_19022_, _18727_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_19033_, _18771_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor (_19044_, _19033_, _19022_);
  and (_19055_, _18640_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  and (_19066_, _18684_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_19077_, _19066_, _19055_);
  and (_19088_, _18825_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_19098_, _18836_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  nor (_19109_, _19098_, _19088_);
  and (_19120_, _19109_, _19077_);
  and (_19131_, _19120_, _19044_);
  nor (_19142_, _19131_, _18880_);
  and (_19153_, _19142_, _19011_);
  nor (_19164_, _19153_, _19000_);
  nor (_19175_, _19164_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_19186_, _19175_, _18989_);
  and (_19197_, _19186_, _18564_);
  nor (_19208_, _19197_, _18978_);
  nor (_19218_, _19208_, _18957_);
  and (_19229_, _18542_, \oc8051_top_1.oc8051_decoder1.op [1]);
  nor (_19240_, _19229_, _18564_);
  and (_19251_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  not (_19262_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_19273_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], \oc8051_top_1.oc8051_memory_interface1.cdone );
  not (_19284_, _18880_);
  and (_19295_, _18836_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  and (_19306_, _18727_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nor (_19327_, _19306_, _19295_);
  and (_19328_, _18640_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  and (_19350_, _18684_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_19351_, _19350_, _19328_);
  and (_19373_, _18825_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_19374_, _18771_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor (_19396_, _19374_, _19373_);
  and (_19397_, _19396_, _19351_);
  and (_19408_, _19397_, _19327_);
  and (_19419_, _19408_, _19284_);
  nor (_19430_, _19419_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  or (_19440_, _19430_, _19273_);
  and (_19451_, _19440_, _19262_);
  nor (_19462_, _19451_, _19251_);
  and (_19473_, _19462_, _18564_);
  nor (_19484_, _19473_, _19240_);
  and (_19495_, _18542_, \oc8051_top_1.oc8051_decoder1.op [0]);
  nor (_19506_, _19495_, _18564_);
  and (_19517_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_19528_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_19539_, _18640_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  and (_19549_, _18684_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_19560_, _19549_, _19539_);
  and (_19571_, _18727_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_19582_, _18771_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor (_19593_, _19582_, _19571_);
  and (_19604_, _19593_, _19560_);
  and (_19615_, _18825_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_19626_, _18836_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  nor (_19637_, _19626_, _19615_);
  and (_19648_, _19637_, _19604_);
  nor (_19659_, _19648_, _18880_);
  and (_19669_, _19659_, _19011_);
  or (_19680_, _19669_, _19528_);
  and (_19691_, _19680_, _19262_);
  nor (_19702_, _19691_, _19517_);
  and (_19713_, _19702_, _18564_);
  nor (_19724_, _19713_, _19506_);
  nor (_19735_, _19724_, _19484_);
  and (_19746_, _19735_, _19218_);
  and (_19757_, _18542_, \oc8051_top_1.oc8051_decoder1.op [4]);
  nor (_19768_, _19757_, _18564_);
  and (_19778_, _18727_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_19789_, _18771_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  nor (_19800_, _19789_, _19778_);
  and (_19811_, _18640_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  and (_19822_, _18684_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_19833_, _19822_, _19811_);
  and (_19844_, _18825_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_19855_, _18836_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  nor (_19866_, _19855_, _19844_);
  and (_19877_, _19866_, _19833_);
  and (_19887_, _19877_, _19800_);
  not (_19898_, _19887_);
  nor (_19909_, _19898_, _18891_);
  nor (_19920_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], _19011_);
  nor (_19931_, _19920_, _19909_);
  nor (_19942_, _19931_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_19953_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _19262_);
  nor (_19964_, _19953_, _19942_);
  not (_19975_, _19964_);
  and (_19986_, _19975_, _18564_);
  nor (_19996_, _19986_, _19768_);
  and (_20007_, _18542_, \oc8051_top_1.oc8051_decoder1.op [7]);
  nor (_20018_, _20007_, _18564_);
  and (_20029_, \oc8051_top_1.oc8051_memory_interface1.dack_ir , \oc8051_top_1.oc8051_memory_interface1.ddat_ir [7]);
  and (_20040_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  and (_20051_, _18836_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  and (_20062_, _18727_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor (_20073_, _20062_, _20051_);
  and (_20084_, _18640_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  and (_20095_, _18684_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_20105_, _20095_, _20084_);
  and (_20116_, _18825_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_20127_, _18771_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  nor (_20138_, _20127_, _20116_);
  and (_20149_, _20138_, _20105_);
  and (_20160_, _20149_, _20073_);
  nor (_20171_, _20160_, _18880_);
  and (_20182_, _20171_, _19011_);
  or (_20193_, _20182_, _20040_);
  and (_20204_, _20193_, _19262_);
  nor (_20214_, _20204_, _20029_);
  and (_20225_, _20214_, _18564_);
  nor (_20236_, _20225_, _20018_);
  and (_20247_, _18542_, \oc8051_top_1.oc8051_decoder1.op [6]);
  nor (_20258_, _20247_, _18564_);
  and (_20269_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_20280_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_20291_, _18836_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  and (_20302_, _18727_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor (_20313_, _20302_, _20291_);
  and (_20323_, _18640_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  and (_20334_, _18684_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_20345_, _20334_, _20323_);
  and (_20356_, _18825_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_20367_, _18771_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor (_20378_, _20367_, _20356_);
  and (_20389_, _20378_, _20345_);
  and (_20400_, _20389_, _20313_);
  nor (_20411_, _20400_, _18880_);
  and (_20422_, _20411_, _19011_);
  or (_20432_, _20422_, _20280_);
  and (_20443_, _20432_, _19262_);
  nor (_20454_, _20443_, _20269_);
  and (_20465_, _20454_, _18564_);
  nor (_20476_, _20465_, _20258_);
  and (_20487_, _18542_, \oc8051_top_1.oc8051_decoder1.op [5]);
  nor (_20498_, _20487_, _18564_);
  and (_20509_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_20520_, \oc8051_top_1.oc8051_memory_interface1.cdata [5], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_20531_, _18640_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  and (_20542_, _18684_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_20552_, _20542_, _20531_);
  and (_20563_, _18727_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_20574_, _18771_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor (_20585_, _20574_, _20563_);
  and (_20596_, _20585_, _20552_);
  and (_20607_, _18825_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_20618_, _18836_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  nor (_20629_, _20618_, _20607_);
  and (_20640_, _20629_, _20596_);
  nor (_20651_, _20640_, _18880_);
  and (_20661_, _20651_, _19011_);
  or (_20672_, _20661_, _20520_);
  and (_20683_, _20672_, _19262_);
  nor (_20694_, _20683_, _20509_);
  and (_20705_, _20694_, _18564_);
  nor (_20716_, _20705_, _20498_);
  not (_20727_, _20716_);
  and (_20738_, _20727_, _20476_);
  and (_20749_, _20738_, _20236_);
  and (_20760_, _20749_, _19996_);
  and (_20770_, _20760_, _19746_);
  not (_20781_, _19724_);
  and (_20792_, _19218_, _19484_);
  and (_20803_, _20792_, _20781_);
  nor (_20814_, _20476_, _20236_);
  and (_20825_, _20814_, _20716_);
  and (_20836_, _20825_, _20803_);
  nor (_20847_, _20836_, _20770_);
  not (_20858_, _19996_);
  not (_20869_, _19208_);
  and (_20879_, _19484_, _18957_);
  and (_20890_, _20879_, _20869_);
  and (_20901_, _20890_, _20858_);
  not (_20912_, _20236_);
  and (_20923_, _20476_, _20912_);
  and (_20934_, _20923_, _20727_);
  and (_20945_, _20934_, _20901_);
  and (_20956_, _20716_, _20476_);
  and (_20967_, _20956_, _20236_);
  and (_20978_, _20967_, _20901_);
  or (_20988_, _20978_, _20945_);
  not (_20999_, _20988_);
  and (_21010_, _20999_, _20847_);
  and (_21021_, _19996_, _20869_);
  and (_21032_, _21021_, _20879_);
  and (_21043_, _21032_, _20934_);
  and (_21054_, _20890_, _20825_);
  or (_21065_, _21054_, _21043_);
  not (_21076_, _21065_);
  and (_21087_, _20956_, _20912_);
  and (_21097_, _21087_, _20858_);
  and (_21108_, _21097_, _20890_);
  nor (_21119_, _20476_, _20912_);
  and (_21130_, _21119_, _20727_);
  and (_21141_, _21130_, _20858_);
  and (_21152_, _21141_, _20890_);
  nor (_21163_, _21152_, _21108_);
  and (_21174_, _21163_, _21076_);
  and (_21185_, _21174_, _21010_);
  and (_21196_, _20792_, _19724_);
  nor (_21206_, _20727_, _19996_);
  and (_21217_, _21119_, _21206_);
  and (_21228_, _21217_, _21196_);
  and (_21239_, _21130_, _19996_);
  and (_21250_, _21087_, _19996_);
  or (_21261_, _21250_, _21239_);
  and (_21272_, _21261_, _21196_);
  nor (_21283_, _21272_, _21228_);
  and (_21294_, _21119_, _20716_);
  and (_21305_, _21294_, _19996_);
  and (_21316_, _21305_, _20890_);
  and (_21326_, _20890_, _20749_);
  and (_21337_, _20814_, _20727_);
  and (_21348_, _21337_, _20890_);
  or (_21359_, _21348_, _21326_);
  and (_21370_, _21239_, _20890_);
  or (_21381_, _21370_, _21359_);
  nor (_21392_, _21381_, _21316_);
  and (_21403_, _21392_, _21283_);
  and (_21414_, _21403_, _21185_);
  nor (_21425_, _21414_, _18509_);
  and (_21435_, \oc8051_top_1.oc8051_decoder1.state [1], _15565_);
  and (_21446_, _20836_, _21435_);
  and (_21457_, _21446_, \oc8051_top_1.oc8051_decoder1.state [0]);
  not (_21468_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and (_21479_, _21435_, _21468_);
  and (_21490_, _21479_, _21087_);
  and (_21501_, _21490_, _19746_);
  or (_21512_, _21501_, _21457_);
  nor (_21523_, _21512_, _21425_);
  nor (_21534_, _21523_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_21544_, _21534_, _18487_);
  and (_21555_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_21566_, _21305_, _19746_);
  not (_21577_, _21566_);
  and (_21588_, _21305_, _20803_);
  and (_21599_, _20749_, _20858_);
  and (_21610_, _21599_, _20803_);
  nor (_21621_, _21610_, _21588_);
  and (_21632_, _21621_, _21577_);
  and (_21643_, _21217_, _19746_);
  and (_21654_, _20869_, _18957_);
  not (_21665_, _19484_);
  and (_21676_, _19724_, _21665_);
  and (_21687_, _21676_, _21654_);
  and (_21698_, _20934_, _20858_);
  and (_21709_, _21698_, _21687_);
  nor (_21720_, _21709_, _21643_);
  and (_21731_, _21337_, _19996_);
  or (_21742_, _21731_, _20760_);
  and (_21753_, _21742_, _21687_);
  and (_21764_, _21250_, _20803_);
  and (_21775_, _21698_, _20792_);
  or (_21786_, _21775_, _21764_);
  nor (_21797_, _21786_, _21753_);
  and (_21808_, _21797_, _21720_);
  and (_21819_, _21808_, _21632_);
  and (_21830_, _21687_, _21097_);
  and (_21841_, _21654_, _21665_);
  and (_21852_, _21841_, _21599_);
  and (_21863_, _21852_, _19724_);
  nor (_21874_, _21863_, _21830_);
  and (_21885_, _20825_, _19746_);
  and (_21896_, _21885_, _20858_);
  and (_21907_, _20825_, _19996_);
  or (_21918_, _21731_, _21907_);
  and (_21929_, _21918_, _19746_);
  nor (_21940_, _21929_, _21896_);
  and (_21951_, _21294_, _20901_);
  not (_21962_, _21951_);
  and (_21973_, _21337_, _20858_);
  and (_21984_, _21973_, _21687_);
  and (_21995_, _21217_, _19208_);
  nor (_22006_, _21995_, _21984_);
  and (_22017_, _22006_, _21962_);
  and (_22028_, _22017_, _21940_);
  and (_22039_, _22028_, _21874_);
  and (_22050_, _20803_, _20760_);
  and (_22061_, _21217_, _20803_);
  nor (_22072_, _22061_, _22050_);
  and (_22083_, _21239_, _20803_);
  and (_22094_, _21687_, _21141_);
  or (_22105_, _22094_, _22083_);
  or (_22116_, _21305_, _21239_);
  and (_22127_, _22116_, _21687_);
  nor (_22138_, _22127_, _22105_);
  and (_22149_, _22138_, _22072_);
  and (_22160_, _20934_, _19996_);
  nor (_22171_, _22160_, _20825_);
  not (_22182_, _21687_);
  nor (_22193_, _22182_, _22171_);
  and (_22204_, _21141_, _20803_);
  and (_22215_, _22160_, _20792_);
  nor (_22226_, _22215_, _22204_);
  not (_22237_, _22226_);
  nor (_22248_, _22237_, _22193_);
  and (_22259_, _20749_, _19746_);
  and (_22270_, _21097_, _20792_);
  nor (_22281_, _22270_, _22259_);
  and (_22292_, _20967_, _20858_);
  and (_22303_, _22292_, _21687_);
  nor (_22314_, _22303_, _20836_);
  and (_22325_, _22314_, _22281_);
  and (_22336_, _22325_, _22248_);
  and (_22347_, _22336_, _22149_);
  and (_22358_, _22347_, _22039_);
  and (_22369_, _22358_, _21819_);
  nor (_22380_, _22369_, _18509_);
  and (_22391_, _21731_, _19746_);
  or (_22402_, _22391_, _21896_);
  and (_22413_, _22402_, _21479_);
  and (_22424_, _20923_, _19746_);
  and (_22435_, _22424_, _21479_);
  or (_22446_, _22435_, _21457_);
  or (_22457_, _22446_, _22413_);
  nor (_22468_, _22457_, _22380_);
  nor (_22479_, _22468_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_22490_, _22479_, _21555_);
  nor (_22501_, _22490_, _21544_);
  and (_22512_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_22523_, _21654_, _19735_);
  and (_22534_, _22523_, _21141_);
  and (_22545_, _22523_, _21217_);
  nor (_22556_, _22545_, _22534_);
  and (_22567_, _22556_, _21283_);
  nor (_22578_, _22567_, _18509_);
  nor (_22589_, _22578_, _22435_);
  not (_22600_, _18509_);
  nor (_22611_, _22556_, _22600_);
  not (_22622_, _22611_);
  and (_22633_, _22622_, _22589_);
  nor (_22644_, _22633_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_22655_, _22644_, _22512_);
  and (_22666_, _22655_, _37580_);
  and (_35258_, _22666_, _22501_);
  not (_22687_, _17187_);
  not (_22698_, _16076_);
  nor (_22709_, _16250_, _22698_);
  and (_22720_, _16599_, _15935_);
  and (_22731_, _22720_, _22709_);
  and (_22742_, _22731_, _16425_);
  nand (_22753_, _22742_, _17425_);
  nor (_22764_, _22753_, _22687_);
  and (_22775_, _22764_, ABINPUT[10]);
  nor (_22786_, _22764_, _16098_);
  nor (_22797_, _22786_, _22775_);
  not (_22808_, _22797_);
  not (_22819_, _22764_);
  and (_22830_, _22819_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  and (_22841_, _22764_, ABINPUT[9]);
  nor (_22852_, _22841_, _22830_);
  and (_22863_, _22819_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  and (_22874_, _22764_, ABINPUT[8]);
  nor (_22885_, _22874_, _22863_);
  and (_22896_, _22819_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  and (_22907_, _22764_, ABINPUT[7]);
  nor (_22918_, _22907_, _22896_);
  and (_22929_, _22819_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  and (_22940_, _22764_, ABINPUT[6]);
  nor (_22951_, _22940_, _22929_);
  and (_22962_, _22819_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  and (_22973_, _22764_, ABINPUT[5]);
  nor (_22984_, _22973_, _22962_);
  and (_22994_, _22819_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  and (_23005_, _22764_, ABINPUT[4]);
  nor (_23016_, _23005_, _22994_);
  nor (_23027_, _22764_, _16827_);
  and (_23038_, _22764_, ABINPUT[3]);
  nor (_23049_, _23038_, _23027_);
  and (_23060_, _23049_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and (_23071_, _23060_, _23016_);
  and (_23082_, _23071_, _22984_);
  and (_23093_, _23082_, _22951_);
  and (_23103_, _23093_, _22918_);
  and (_23114_, _23103_, _22885_);
  and (_23125_, _23114_, _22852_);
  and (_23136_, _23125_, _22808_);
  nor (_23147_, _23125_, _22808_);
  nor (_23158_, _23147_, _23136_);
  and (_23169_, _23158_, _15739_);
  nor (_23180_, _23169_, _16142_);
  nor (_23191_, _23180_, _22764_);
  nor (_23202_, _23191_, _22775_);
  nor (_35441_, _23202_, rst);
  not (_23223_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and (_23234_, _23049_, _23223_);
  nor (_23245_, _23049_, _23223_);
  nor (_23256_, _23245_, _23234_);
  and (_23267_, _23256_, _15739_);
  nor (_23278_, _23267_, _16838_);
  nor (_23289_, _23278_, _22764_);
  nor (_23300_, _23289_, _23038_);
  nand (_36625_, _23300_, _37580_);
  nor (_23321_, _23060_, _23016_);
  nor (_23332_, _23321_, _23071_);
  nor (_23342_, _23332_, _15728_);
  nor (_23353_, _23342_, _16925_);
  nor (_23364_, _23353_, _22764_);
  nor (_23375_, _23364_, _23005_);
  nand (_36633_, _23375_, _37580_);
  nor (_23396_, _23071_, _22984_);
  nor (_23407_, _23396_, _23082_);
  nor (_23418_, _23407_, _15728_);
  nor (_23429_, _23418_, _16674_);
  nor (_23440_, _23429_, _22764_);
  nor (_23450_, _23440_, _22973_);
  nand (_36641_, _23450_, _37580_);
  nor (_23471_, _23082_, _22951_);
  nor (_23482_, _23471_, _23093_);
  nor (_23493_, _23482_, _15728_);
  nor (_23504_, _23493_, _16305_);
  nor (_23515_, _23504_, _22764_);
  nor (_23526_, _23515_, _22940_);
  nor (_36649_, _23526_, rst);
  nor (_23547_, _23093_, _22918_);
  nor (_23557_, _23547_, _23103_);
  nor (_23568_, _23557_, _15728_);
  nor (_23579_, _23568_, _16533_);
  nor (_23590_, _23579_, _22764_);
  nor (_23601_, _23590_, _22907_);
  nor (_36657_, _23601_, rst);
  nor (_23622_, _23103_, _22885_);
  nor (_23633_, _23622_, _23114_);
  nor (_23644_, _23633_, _15728_);
  nor (_23655_, _23644_, _15772_);
  nor (_23665_, _23655_, _22764_);
  nor (_23676_, _23665_, _22874_);
  nor (_36665_, _23676_, rst);
  nor (_23697_, _23114_, _22852_);
  nor (_23708_, _23697_, _23125_);
  nor (_23719_, _23708_, _15728_);
  nor (_23730_, _23719_, _15989_);
  nor (_23741_, _23730_, _22764_);
  nor (_23752_, _23741_, _22841_);
  nor (_36672_, _23752_, rst);
  and (_23773_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], _15565_);
  and (_23784_, _23773_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_23795_, _17793_, _16425_);
  nand (_23806_, _23795_, _22731_);
  nor (_23817_, _23806_, _22687_);
  or (_23827_, _23817_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  nand (_23838_, _23817_, _17122_);
  and (_23849_, _23838_, _23827_);
  or (_23860_, _23849_, _23784_);
  not (_23871_, ABINPUT[18]);
  nand (_23882_, _23784_, _23871_);
  and (_23893_, _23882_, _37580_);
  and (_38754_, _23893_, _23860_);
  and (_23913_, _22742_, _17620_);
  and (_23924_, _23913_, _17187_);
  nor (_23935_, _23924_, _23784_);
  and (_23946_, _23935_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  nor (_23957_, _23935_, _17122_);
  or (_23968_, _23957_, _23946_);
  and (_38774_, _23968_, _37580_);
  or (_23989_, _23817_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  not (_23999_, ABINPUT[19]);
  nand (_24010_, _23817_, _23999_);
  and (_24021_, _24010_, _23989_);
  or (_24032_, _24021_, _23784_);
  not (_24043_, ABINPUT[11]);
  nand (_24054_, _23784_, _24043_);
  and (_24065_, _24054_, _37580_);
  and (_39759_, _24065_, _24032_);
  or (_24085_, _23817_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  nand (_24096_, _23817_, _17512_);
  and (_24107_, _24096_, _24085_);
  or (_24118_, _24107_, _23784_);
  not (_24129_, ABINPUT[12]);
  nand (_24140_, _23784_, _24129_);
  and (_24151_, _24140_, _37580_);
  and (_39767_, _24151_, _24118_);
  or (_24171_, _23817_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  nand (_24182_, _23817_, _17707_);
  and (_24193_, _24182_, _24171_);
  or (_24204_, _24193_, _23784_);
  not (_24215_, ABINPUT[13]);
  nand (_24226_, _23784_, _24215_);
  and (_24237_, _24226_, _37580_);
  and (_39776_, _24237_, _24204_);
  or (_24257_, _23817_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  nand (_24268_, _23817_, _17891_);
  and (_24279_, _24268_, _24257_);
  or (_24290_, _24279_, _23784_);
  not (_24301_, ABINPUT[14]);
  nand (_24312_, _23784_, _24301_);
  and (_24323_, _24312_, _37580_);
  and (_39785_, _24323_, _24290_);
  or (_24343_, _23817_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  nand (_24354_, _23817_, _18054_);
  and (_24365_, _24354_, _24343_);
  or (_24376_, _24365_, _23784_);
  not (_24387_, ABINPUT[15]);
  nand (_24398_, _23784_, _24387_);
  and (_24409_, _24398_, _37580_);
  and (_39793_, _24409_, _24376_);
  or (_24429_, _23817_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  nand (_24440_, _23817_, _18228_);
  and (_24451_, _24440_, _24429_);
  or (_24462_, _24451_, _23784_);
  not (_24473_, ABINPUT[16]);
  nand (_24484_, _23784_, _24473_);
  and (_24494_, _24484_, _37580_);
  and (_39802_, _24494_, _24462_);
  or (_24515_, _23817_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  nand (_24526_, _23817_, _18401_);
  and (_24537_, _24526_, _24515_);
  or (_24548_, _24537_, _23784_);
  not (_24559_, ABINPUT[17]);
  nand (_24570_, _23784_, _24559_);
  and (_24580_, _24570_, _37580_);
  and (_39810_, _24580_, _24548_);
  and (_24601_, _23935_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  nor (_24612_, _23935_, _23999_);
  or (_24623_, _24612_, _24601_);
  and (_39819_, _24623_, _37580_);
  and (_24644_, _23935_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  nor (_24654_, _23935_, _17512_);
  or (_24665_, _24654_, _24644_);
  and (_39827_, _24665_, _37580_);
  and (_24686_, _23935_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  nor (_24697_, _23935_, _17707_);
  or (_24708_, _24697_, _24686_);
  and (_39836_, _24708_, _37580_);
  and (_24729_, _23935_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  nor (_24739_, _23935_, _17891_);
  or (_24750_, _24739_, _24729_);
  and (_39844_, _24750_, _37580_);
  and (_24771_, _23935_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  nor (_24782_, _23935_, _18054_);
  or (_24793_, _24782_, _24771_);
  and (_39853_, _24793_, _37580_);
  and (_24814_, _23935_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  nor (_24824_, _23935_, _18228_);
  or (_24835_, _24824_, _24814_);
  and (_39861_, _24835_, _37580_);
  and (_24856_, _23935_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  nor (_24867_, _23935_, _18401_);
  or (_24878_, _24867_, _24856_);
  and (_39870_, _24878_, _37580_);
  and (_24899_, _16610_, _15935_);
  and (_24909_, _24899_, _22698_);
  not (_24920_, _15630_);
  nor (_24931_, _24920_, _16250_);
  and (_24942_, _24931_, _24909_);
  and (_24953_, _17023_, ABINPUT[0]);
  not (_24964_, _17023_);
  and (_24975_, _24964_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_24986_, _24975_, _24953_);
  nand (_24996_, _24986_, _24942_);
  nor (_25007_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  nor (_25018_, _25007_, _17056_);
  and (_25029_, _25007_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or (_25040_, _25029_, _25018_);
  or (_25051_, _25040_, _24942_);
  and (_25062_, _25051_, _24996_);
  and (_25073_, _17187_, _17143_);
  and (_25084_, _25073_, _16261_);
  and (_25094_, _25084_, _24909_);
  not (_25105_, _25094_);
  and (_25116_, _25105_, _25062_);
  and (_25127_, _25094_, ABINPUT[10]);
  or (_25138_, _25127_, _25116_);
  and (_01571_, _25138_, _37580_);
  and (_25159_, _24942_, _17425_);
  nand (_25170_, _25159_, _17056_);
  or (_25181_, _25159_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_25192_, _25181_, _25170_);
  or (_25203_, _25192_, _25094_);
  not (_25213_, ABINPUT[4]);
  nor (_25224_, _16250_, _16076_);
  and (_25235_, _25073_, _24899_);
  and (_25246_, _25235_, _25224_);
  nand (_25257_, _25246_, _25213_);
  and (_25268_, _25257_, _25203_);
  and (_06388_, _25268_, _37580_);
  not (_25289_, _17620_);
  and (_25300_, _25289_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  nor (_25311_, _25300_, _17653_);
  nand (_25321_, _25311_, _24942_);
  and (_25332_, ABINPUT[2], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  not (_25343_, \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  and (_25354_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], _25343_);
  or (_25365_, _25354_, _25332_);
  or (_25376_, _25365_, _24942_);
  and (_25387_, _25376_, _25321_);
  and (_25398_, _25387_, _25105_);
  and (_25409_, _25094_, ABINPUT[5]);
  or (_25420_, _25409_, _25398_);
  and (_06399_, _25420_, _37580_);
  not (_25440_, _25246_);
  nand (_25451_, _24942_, _17793_);
  and (_25462_, _25451_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_25473_, _24942_, _17826_);
  or (_25484_, _25473_, _25462_);
  and (_25495_, _25484_, _25440_);
  and (_25506_, _17143_, _16425_);
  not (_25517_, _25506_);
  not (_25528_, _15935_);
  nor (_25538_, _16599_, _25528_);
  nand (_25549_, _25538_, _25224_);
  nor (_25560_, _25549_, _25517_);
  and (_25571_, _25560_, _17187_);
  and (_25582_, _25571_, ABINPUT[6]);
  or (_25593_, _25582_, _25495_);
  and (_06409_, _25593_, _37580_);
  nand (_25614_, _24942_, _17967_);
  and (_25625_, _25614_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_25636_, _24942_, _18000_);
  or (_25646_, _25636_, _25625_);
  and (_25657_, _25646_, _25440_);
  and (_25668_, _25571_, ABINPUT[7]);
  or (_25679_, _25668_, _25657_);
  and (_06420_, _25679_, _37580_);
  nand (_25700_, _24942_, _18140_);
  and (_25711_, _25700_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_25722_, _24942_, _18173_);
  or (_25733_, _25722_, _25094_);
  or (_25744_, _25733_, _25711_);
  not (_25755_, ABINPUT[8]);
  nand (_25765_, _25094_, _25755_);
  and (_25776_, _25765_, _25744_);
  and (_06431_, _25776_, _37580_);
  not (_25797_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_25808_, _18314_, _25797_);
  nor (_25819_, _25808_, _18346_);
  nand (_25830_, _25819_, _24942_);
  and (_25840_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  and (_25851_, _25840_, ABINPUT[1]);
  nor (_25862_, _25840_, _25797_);
  or (_25873_, _25862_, _25851_);
  or (_25884_, _25873_, _24942_);
  and (_25895_, _25884_, _25830_);
  and (_25906_, _25895_, _25105_);
  and (_25917_, _25094_, ABINPUT[9]);
  or (_25928_, _25917_, _25906_);
  and (_06442_, _25928_, _37580_);
  not (_25948_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_25959_, _23773_, _25948_);
  and (_25970_, _25959_, ABINPUT[18]);
  not (_25981_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_25992_, _16599_, _16425_);
  and (_26003_, _25992_, _16087_);
  and (_26014_, _26003_, _24931_);
  and (_26025_, _26014_, _17023_);
  nor (_26036_, _26025_, _25981_);
  not (_26047_, _26036_);
  nor (_26058_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_26068_, _26058_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_26079_, _25992_, _25528_);
  and (_26090_, _26079_, _25073_);
  and (_26101_, _26090_, _25224_);
  nor (_26112_, _26101_, _26068_);
  and (_26123_, _26014_, _24953_);
  not (_26134_, _26123_);
  and (_26145_, _26134_, _26112_);
  and (_26156_, _26145_, _26047_);
  not (_26167_, _25959_);
  and (_26178_, _26112_, _26167_);
  nor (_26188_, _25959_, _17122_);
  nor (_26199_, _26188_, _26178_);
  nor (_26210_, _26199_, _26156_);
  nor (_26221_, _26210_, _25970_);
  nor (_07163_, _26221_, rst);
  not (_26242_, _26178_);
  not (_26253_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and (_26264_, _26014_, _17143_);
  nor (_26275_, _26264_, _26253_);
  and (_26286_, _26014_, _17284_);
  nor (_26297_, _26286_, _26275_);
  nor (_26307_, _26297_, _26242_);
  not (_26318_, _26307_);
  and (_26329_, _25959_, ABINPUT[11]);
  or (_26340_, _25959_, _23999_);
  nor (_26351_, _26340_, _26112_);
  nor (_26362_, _26351_, _26329_);
  and (_26373_, _26362_, _26318_);
  nor (_08869_, _26373_, rst);
  not (_26394_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_26405_, _26014_, _17425_);
  nor (_26416_, _26405_, _26394_);
  and (_26427_, _26014_, _17467_);
  nor (_26437_, _26427_, _26416_);
  nor (_26448_, _26437_, _26242_);
  not (_26459_, _26448_);
  and (_26470_, _25959_, ABINPUT[12]);
  or (_26481_, _25959_, _17512_);
  nor (_26492_, _26481_, _26112_);
  nor (_26503_, _26492_, _26470_);
  and (_26514_, _26503_, _26459_);
  nor (_08880_, _26514_, rst);
  and (_26535_, _25959_, ABINPUT[13]);
  not (_26546_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_26556_, _26014_, _17620_);
  nor (_26567_, _26556_, _26546_);
  not (_26578_, _26567_);
  and (_26589_, _26014_, _17653_);
  not (_26600_, _26589_);
  and (_26611_, _26600_, _26112_);
  and (_26622_, _26611_, _26578_);
  nor (_26633_, _25959_, _17707_);
  nor (_26644_, _26633_, _26178_);
  nor (_26655_, _26644_, _26622_);
  nor (_26665_, _26655_, _26535_);
  nor (_08891_, _26665_, rst);
  and (_26686_, _25959_, ABINPUT[14]);
  not (_26697_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_26708_, _26014_, _17793_);
  nor (_26719_, _26708_, _26697_);
  not (_26730_, _26719_);
  and (_26741_, _26014_, _17826_);
  not (_26752_, _26741_);
  and (_26763_, _26752_, _26112_);
  and (_26773_, _26763_, _26730_);
  nor (_26784_, _25959_, _17891_);
  nor (_26795_, _26784_, _26178_);
  nor (_26806_, _26795_, _26773_);
  nor (_26817_, _26806_, _26686_);
  nor (_08902_, _26817_, rst);
  and (_26838_, _25959_, ABINPUT[15]);
  not (_26849_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_26860_, _26014_, _17967_);
  nor (_26871_, _26860_, _26849_);
  not (_26881_, _26871_);
  and (_26892_, _26014_, _18000_);
  not (_26903_, _26892_);
  and (_26914_, _26903_, _26112_);
  and (_26925_, _26914_, _26881_);
  nor (_26936_, _25959_, _18054_);
  nor (_26947_, _26936_, _26178_);
  nor (_26958_, _26947_, _26925_);
  nor (_26969_, _26958_, _26838_);
  nor (_08913_, _26969_, rst);
  and (_26990_, _25959_, ABINPUT[16]);
  not (_27000_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_27011_, _26014_, _18140_);
  nor (_27022_, _27011_, _27000_);
  not (_27033_, _27022_);
  and (_27044_, _26014_, _18173_);
  not (_27055_, _27044_);
  and (_27066_, _27055_, _26112_);
  and (_27077_, _27066_, _27033_);
  nor (_27088_, _25959_, _18228_);
  nor (_27099_, _27088_, _26178_);
  nor (_27109_, _27099_, _27077_);
  nor (_27120_, _27109_, _26990_);
  nor (_08924_, _27120_, rst);
  and (_27141_, _25959_, ABINPUT[17]);
  not (_27152_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_27163_, _26014_, _18314_);
  nor (_27174_, _27163_, _27152_);
  and (_27185_, _26014_, _18346_);
  nor (_27196_, _27185_, _27174_);
  and (_27207_, _27196_, _26112_);
  nor (_27217_, _26112_, ABINPUT[25]);
  or (_27228_, _27217_, _27207_);
  nor (_27239_, _27228_, _25959_);
  nor (_27250_, _27239_, _27141_);
  nor (_08935_, _27250_, rst);
  and (_27271_, _22742_, _17023_);
  or (_27282_, _27271_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  nand (_27293_, _27271_, _17056_);
  and (_27304_, _27293_, _15630_);
  and (_27315_, _27304_, _27282_);
  not (_27325_, ABINPUT[10]);
  and (_27336_, _22731_, _25506_);
  nand (_27347_, _27336_, _27325_);
  or (_27358_, _27336_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_27369_, _27358_, _17187_);
  and (_27380_, _27369_, _27347_);
  and (_27391_, _17100_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  or (_27401_, _27391_, rst);
  or (_27412_, _27401_, _27380_);
  or (_19317_, _27412_, _27315_);
  and (_27433_, _24899_, _22709_);
  nand (_27444_, _27433_, _17023_);
  and (_27455_, _27444_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_27466_, _27433_, _24953_);
  or (_27477_, _27466_, _27455_);
  and (_27487_, _27477_, _15630_);
  and (_27498_, _27433_, _17143_);
  and (_27509_, _27498_, ABINPUT[10]);
  not (_27520_, _27498_);
  and (_27531_, _27520_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  or (_27542_, _27531_, _27509_);
  and (_27553_, _27542_, _17187_);
  and (_27564_, _17100_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  or (_27574_, _27564_, rst);
  or (_27585_, _27574_, _27553_);
  or (_19339_, _27585_, _27487_);
  and (_27606_, _16599_, _25528_);
  and (_27617_, _27606_, _22709_);
  and (_27628_, _27617_, _25506_);
  and (_27639_, _27628_, ABINPUT[10]);
  not (_27650_, _27628_);
  and (_27660_, _27650_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or (_27671_, _27660_, _27639_);
  and (_27682_, _27671_, _17187_);
  and (_27693_, _27617_, _16425_);
  and (_27704_, _24964_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or (_27715_, _27704_, _24953_);
  and (_27726_, _27715_, _27693_);
  not (_27737_, _27693_);
  and (_27747_, _27737_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or (_27758_, _27747_, _27726_);
  and (_27769_, _27758_, _15630_);
  and (_27780_, _17100_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or (_27791_, _27780_, rst);
  or (_27802_, _27791_, _27769_);
  or (_19362_, _27802_, _27682_);
  nor (_27823_, _16599_, _15935_);
  and (_27833_, _22709_, _27823_);
  and (_27844_, _27833_, _25506_);
  and (_27855_, _27844_, ABINPUT[10]);
  not (_27866_, _27844_);
  and (_27877_, _27866_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or (_27888_, _27877_, _27855_);
  and (_27899_, _27888_, _17187_);
  and (_27909_, _24964_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or (_27920_, _27909_, _24953_);
  and (_27931_, _16076_, _25528_);
  and (_27942_, _27931_, _16620_);
  and (_27953_, _27942_, _27920_);
  not (_27964_, _27942_);
  and (_27975_, _27964_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or (_27986_, _27975_, _27953_);
  and (_27996_, _27986_, _15630_);
  and (_28007_, _17100_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or (_28018_, _28007_, rst);
  or (_28029_, _28018_, _27996_);
  or (_19385_, _28029_, _27899_);
  not (_28050_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  nor (_28061_, _27336_, _28050_);
  and (_28072_, _22742_, _17284_);
  or (_28082_, _28072_, _28061_);
  and (_28093_, _28082_, _15630_);
  and (_28104_, _27336_, ABINPUT[3]);
  or (_28115_, _28104_, _28061_);
  and (_28126_, _28115_, _17187_);
  nor (_28137_, _15619_, _28050_);
  or (_28148_, _28137_, rst);
  or (_28158_, _28148_, _28126_);
  or (_36859_, _28158_, _28093_);
  and (_28179_, _22742_, _17467_);
  and (_28190_, _22753_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  or (_28201_, _28190_, _28179_);
  and (_28212_, _28201_, _15630_);
  nand (_28223_, _27336_, _25213_);
  or (_28234_, _27336_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_28244_, _28234_, _17187_);
  and (_28255_, _28244_, _28223_);
  and (_28266_, _17100_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  or (_28277_, _28266_, _28255_);
  or (_28288_, _28277_, _28212_);
  or (_36861_, _28288_, rst);
  not (_28309_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  nor (_28320_, _23913_, _28309_);
  and (_28330_, _22742_, _17653_);
  or (_28341_, _28330_, _28320_);
  and (_28352_, _28341_, _15630_);
  or (_28363_, _27336_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_28374_, _28363_, _17187_);
  not (_28385_, ABINPUT[5]);
  nand (_28396_, _27336_, _28385_);
  and (_28407_, _28396_, _28374_);
  nor (_28417_, _15619_, _28309_);
  or (_28428_, _28417_, rst);
  or (_28439_, _28428_, _28407_);
  or (_36863_, _28439_, _28352_);
  not (_28460_, ABINPUT[6]);
  nand (_28471_, _27336_, _28460_);
  or (_28482_, _27336_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_28493_, _28482_, _17187_);
  and (_28503_, _28493_, _28471_);
  and (_28514_, _23806_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_28525_, _22742_, _17826_);
  or (_28536_, _28525_, _28514_);
  and (_28547_, _28536_, _15630_);
  and (_28558_, _17100_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or (_28569_, _28558_, rst);
  or (_28579_, _28569_, _28547_);
  or (_36865_, _28579_, _28503_);
  nand (_28600_, _22742_, _17967_);
  and (_28611_, _28600_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_28622_, _22742_, _18000_);
  or (_28633_, _28622_, _28611_);
  and (_28644_, _28633_, _15630_);
  not (_28655_, ABINPUT[7]);
  nand (_28665_, _27336_, _28655_);
  or (_28676_, _27336_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_28687_, _28676_, _17187_);
  and (_28698_, _28687_, _28665_);
  and (_28709_, _17100_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or (_28720_, _28709_, rst);
  or (_28731_, _28720_, _28698_);
  or (_36867_, _28731_, _28644_);
  nand (_28751_, _22742_, _18140_);
  and (_28762_, _28751_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_28773_, _22742_, _18173_);
  or (_28784_, _28773_, _28762_);
  and (_28795_, _28784_, _15630_);
  nand (_28806_, _27336_, _25755_);
  or (_28817_, _27336_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_28828_, _28817_, _17187_);
  and (_28838_, _28828_, _28806_);
  and (_28849_, _17100_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  or (_28860_, _28849_, rst);
  or (_28871_, _28860_, _28838_);
  or (_36869_, _28871_, _28795_);
  nand (_28892_, _22742_, _18314_);
  and (_28903_, _28892_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_28913_, _22742_, _18346_);
  or (_28924_, _28913_, _28903_);
  and (_28935_, _28924_, _15630_);
  not (_28946_, ABINPUT[9]);
  nand (_28957_, _27336_, _28946_);
  or (_28968_, _27336_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_28979_, _28968_, _17187_);
  and (_28990_, _28979_, _28957_);
  and (_29000_, _17100_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  or (_29011_, _29000_, rst);
  or (_29022_, _29011_, _28990_);
  or (_36871_, _29022_, _28935_);
  not (_29043_, ABINPUT[3]);
  nand (_29054_, _27498_, _29043_);
  or (_29065_, _27498_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and (_29077_, _29065_, _17187_);
  and (_29087_, _29077_, _29054_);
  nand (_29098_, _27498_, _17056_);
  and (_29109_, _29098_, _15630_);
  and (_29120_, _29109_, _29065_);
  and (_29131_, _17100_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  or (_29142_, _29131_, rst);
  or (_29153_, _29142_, _29120_);
  or (_36873_, _29153_, _29087_);
  nand (_29173_, _27433_, _17425_);
  and (_29185_, _29173_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_29196_, _27433_, _17467_);
  or (_29207_, _29196_, _29185_);
  and (_29218_, _29207_, _15630_);
  and (_29229_, _27498_, ABINPUT[4]);
  and (_29240_, _27520_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  or (_29250_, _29240_, _29229_);
  and (_29261_, _29250_, _17187_);
  and (_29272_, _17100_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  or (_29283_, _29272_, rst);
  or (_29295_, _29283_, _29261_);
  or (_36875_, _29295_, _29218_);
  and (_29316_, _27433_, _17620_);
  nor (_29327_, _29316_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_29337_, _29316_, _17056_);
  or (_29348_, _29337_, _24920_);
  nor (_29359_, _29348_, _29327_);
  or (_29370_, _27498_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  nand (_29381_, _27498_, _28385_);
  and (_29392_, _29381_, _17187_);
  and (_29404_, _29392_, _29370_);
  and (_29415_, _17100_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  or (_29425_, _29415_, rst);
  or (_29436_, _29425_, _29404_);
  or (_36877_, _29436_, _29359_);
  nand (_29457_, _27433_, _17793_);
  and (_29468_, _29457_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_29479_, _27433_, _17826_);
  or (_29490_, _29479_, _29468_);
  and (_29501_, _29490_, _15630_);
  and (_29512_, _27498_, ABINPUT[6]);
  and (_29523_, _27520_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or (_29534_, _29523_, _29512_);
  and (_29545_, _29534_, _17187_);
  and (_29556_, _17100_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or (_29567_, _29556_, rst);
  or (_29578_, _29567_, _29545_);
  or (_36879_, _29578_, _29501_);
  and (_29598_, _27433_, _17967_);
  nor (_29609_, _29598_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_29621_, _29598_, _17056_);
  or (_29632_, _29621_, _24920_);
  nor (_29643_, _29632_, _29609_);
  and (_29654_, _27520_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_29665_, _27498_, ABINPUT[7]);
  or (_29675_, _29665_, _29654_);
  and (_29686_, _29675_, _17187_);
  and (_29697_, _17100_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  or (_29708_, _29697_, rst);
  or (_29719_, _29708_, _29686_);
  or (_36881_, _29719_, _29643_);
  and (_29741_, _27433_, _18140_);
  nor (_29751_, _29741_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_29762_, _29741_, _17056_);
  or (_29773_, _29762_, _24920_);
  nor (_29784_, _29773_, _29751_);
  and (_29795_, _27520_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_29806_, _27498_, ABINPUT[8]);
  or (_29817_, _29806_, _29795_);
  and (_29828_, _29817_, _17187_);
  and (_29838_, _17100_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  or (_29849_, _29838_, rst);
  or (_29860_, _29849_, _29828_);
  or (_36883_, _29860_, _29784_);
  nand (_29881_, _27433_, _18314_);
  and (_29892_, _29881_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_29903_, _27433_, _18346_);
  or (_29914_, _29903_, _29892_);
  and (_29924_, _29914_, _15630_);
  and (_29935_, _27520_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_29946_, _27498_, ABINPUT[9]);
  or (_29957_, _29946_, _29935_);
  and (_29968_, _29957_, _17187_);
  and (_29979_, _17100_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  or (_29990_, _29979_, rst);
  or (_30001_, _29990_, _29968_);
  or (_36885_, _30001_, _29924_);
  and (_30021_, _27628_, ABINPUT[3]);
  and (_30032_, _27650_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  or (_30043_, _30032_, _30021_);
  and (_30054_, _30043_, _17187_);
  and (_30065_, _27737_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  not (_30076_, _17143_);
  and (_30087_, _30076_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  or (_30097_, _30087_, _17284_);
  and (_30108_, _30097_, _27693_);
  or (_30119_, _30108_, _30065_);
  and (_30130_, _30119_, _15630_);
  and (_30141_, _17100_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  or (_30152_, _30141_, rst);
  or (_30163_, _30152_, _30130_);
  or (_36887_, _30163_, _30054_);
  and (_30183_, _27628_, ABINPUT[4]);
  and (_30194_, _27650_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or (_30205_, _30194_, _30183_);
  and (_30216_, _30205_, _17187_);
  not (_30227_, _17425_);
  and (_30238_, _30227_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or (_30249_, _30238_, _17467_);
  and (_30259_, _30249_, _27693_);
  and (_30270_, _27737_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or (_30281_, _30270_, _30259_);
  and (_30292_, _30281_, _15630_);
  and (_30303_, _17100_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or (_30314_, _30303_, rst);
  or (_30325_, _30314_, _30292_);
  or (_36888_, _30325_, _30216_);
  and (_30346_, _27628_, ABINPUT[5]);
  and (_30357_, _27650_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or (_30368_, _30357_, _30346_);
  and (_30379_, _30368_, _17187_);
  and (_30390_, _25289_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or (_30401_, _30390_, _17653_);
  and (_30412_, _30401_, _27693_);
  and (_30423_, _27737_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or (_30434_, _30423_, _30412_);
  and (_30445_, _30434_, _15630_);
  and (_30456_, _17100_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or (_30467_, _30456_, rst);
  or (_30478_, _30467_, _30445_);
  or (_36890_, _30478_, _30379_);
  and (_30498_, _27628_, ABINPUT[6]);
  and (_30509_, _27650_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_30520_, _30509_, _30498_);
  and (_30531_, _30520_, _17187_);
  not (_30542_, _17793_);
  and (_30553_, _30542_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_30564_, _30553_, _17826_);
  and (_30575_, _30564_, _27693_);
  and (_30586_, _27737_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_30597_, _30586_, _30575_);
  and (_30608_, _30597_, _15630_);
  and (_30619_, _17100_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_30630_, _30619_, rst);
  or (_30641_, _30630_, _30608_);
  or (_36892_, _30641_, _30531_);
  and (_30662_, _27628_, ABINPUT[7]);
  and (_30673_, _27650_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or (_30684_, _30673_, _30662_);
  and (_30695_, _30684_, _17187_);
  not (_30706_, _17967_);
  and (_30717_, _30706_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or (_30728_, _30717_, _18000_);
  and (_30739_, _30728_, _27693_);
  and (_30750_, _27737_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or (_30761_, _30750_, _30739_);
  and (_30772_, _30761_, _15630_);
  and (_30783_, _17100_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or (_30794_, _30783_, rst);
  or (_30805_, _30794_, _30772_);
  or (_36894_, _30805_, _30695_);
  and (_30826_, _27628_, ABINPUT[8]);
  and (_30837_, _27650_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or (_30848_, _30837_, _30826_);
  and (_30859_, _30848_, _17187_);
  not (_30870_, _18140_);
  and (_30881_, _30870_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or (_30891_, _30881_, _18173_);
  and (_30902_, _30891_, _27693_);
  and (_30913_, _27737_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or (_30924_, _30913_, _30902_);
  and (_30935_, _30924_, _15630_);
  and (_30946_, _17100_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or (_30957_, _30946_, rst);
  or (_30968_, _30957_, _30935_);
  or (_36896_, _30968_, _30859_);
  and (_30989_, _27628_, ABINPUT[9]);
  and (_31000_, _27650_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or (_31011_, _31000_, _30989_);
  and (_31022_, _31011_, _17187_);
  not (_31033_, _18314_);
  and (_31044_, _31033_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or (_31055_, _31044_, _18346_);
  and (_31066_, _31055_, _27693_);
  and (_31077_, _27737_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or (_31088_, _31077_, _31066_);
  and (_31099_, _31088_, _15630_);
  and (_31110_, _17100_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or (_31121_, _31110_, rst);
  or (_31132_, _31121_, _31099_);
  or (_36898_, _31132_, _31022_);
  and (_31153_, _27844_, ABINPUT[3]);
  and (_31164_, _27866_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  or (_31175_, _31164_, _31153_);
  and (_31186_, _31175_, _17187_);
  and (_31197_, _30076_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  or (_31208_, _31197_, _17284_);
  and (_31219_, _31208_, _27942_);
  and (_31230_, _27964_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  or (_31241_, _31230_, _31219_);
  and (_31252_, _31241_, _15630_);
  and (_31263_, _17100_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  or (_31273_, _31263_, rst);
  or (_31284_, _31273_, _31252_);
  or (_36900_, _31284_, _31186_);
  and (_31305_, _27844_, ABINPUT[4]);
  and (_31316_, _27866_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or (_31327_, _31316_, _31305_);
  and (_31338_, _31327_, _17187_);
  and (_31349_, _30227_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or (_31360_, _31349_, _17467_);
  and (_31371_, _31360_, _27942_);
  and (_31382_, _27964_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or (_31393_, _31382_, _31371_);
  and (_31404_, _31393_, _15630_);
  and (_31415_, _17100_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or (_31426_, _31415_, rst);
  or (_31437_, _31426_, _31404_);
  or (_36902_, _31437_, _31338_);
  and (_31458_, _27844_, ABINPUT[5]);
  and (_31469_, _27866_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or (_31480_, _31469_, _31458_);
  and (_31491_, _31480_, _17187_);
  and (_31502_, _25289_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or (_31513_, _31502_, _17653_);
  and (_31524_, _31513_, _27942_);
  and (_31535_, _27964_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or (_31546_, _31535_, _31524_);
  and (_31557_, _31546_, _15630_);
  and (_31568_, _17100_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or (_31579_, _31568_, rst);
  or (_31590_, _31579_, _31557_);
  or (_36904_, _31590_, _31491_);
  and (_31611_, _27844_, ABINPUT[6]);
  and (_31621_, _27866_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_31632_, _31621_, _31611_);
  and (_31643_, _31632_, _17187_);
  and (_31654_, _30542_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_31665_, _31654_, _17826_);
  and (_31676_, _31665_, _27942_);
  and (_31687_, _27964_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_31698_, _31687_, _31676_);
  and (_31709_, _31698_, _15630_);
  and (_31720_, _17100_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_31731_, _31720_, rst);
  or (_31742_, _31731_, _31709_);
  or (_36906_, _31742_, _31643_);
  and (_31763_, _27844_, ABINPUT[7]);
  and (_31774_, _27866_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or (_31785_, _31774_, _31763_);
  and (_31796_, _31785_, _17187_);
  and (_31807_, _30706_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or (_31818_, _31807_, _18000_);
  and (_31829_, _31818_, _27942_);
  and (_31840_, _27964_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or (_31851_, _31840_, _31829_);
  and (_31862_, _31851_, _15630_);
  and (_31873_, _17100_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or (_31884_, _31873_, rst);
  or (_31895_, _31884_, _31862_);
  or (_36908_, _31895_, _31796_);
  and (_31916_, _27844_, ABINPUT[8]);
  and (_31927_, _27866_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or (_31938_, _31927_, _31916_);
  and (_31949_, _31938_, _17187_);
  and (_31960_, _30870_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or (_31971_, _31960_, _18173_);
  and (_31981_, _31971_, _27942_);
  and (_31992_, _27964_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or (_32003_, _31992_, _31981_);
  and (_32014_, _32003_, _15630_);
  and (_32025_, _17100_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or (_32036_, _32025_, rst);
  or (_32047_, _32036_, _32014_);
  or (_36910_, _32047_, _31949_);
  and (_32068_, _27844_, ABINPUT[9]);
  and (_32079_, _27866_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or (_32090_, _32079_, _32068_);
  and (_32101_, _32090_, _17187_);
  and (_32112_, _31033_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or (_32123_, _32112_, _18346_);
  and (_32134_, _32123_, _27942_);
  and (_32145_, _27964_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or (_32156_, _32145_, _32134_);
  and (_32167_, _32156_, _15630_);
  and (_32178_, _17100_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or (_32189_, _32178_, rst);
  or (_32200_, _32189_, _32167_);
  or (_36912_, _32200_, _32101_);
  and (_32221_, _25073_, _16435_);
  and (_32232_, _32221_, _27617_);
  nor (_32243_, _24920_, _16425_);
  and (_32254_, _32243_, _27617_);
  and (_32265_, _32254_, _17023_);
  nand (_32276_, _32265_, _17056_);
  or (_32287_, _32265_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_32298_, _32287_, _32276_);
  or (_32309_, _32298_, _32232_);
  nand (_32320_, _32232_, _27325_);
  and (_32330_, _32320_, _37580_);
  and (_37492_, _32330_, _32309_);
  and (_32351_, _32221_, _27833_);
  not (_32362_, _16599_);
  and (_32373_, _32243_, _32362_);
  and (_32384_, _32373_, _16261_);
  and (_32395_, _32384_, _27931_);
  and (_32406_, _32395_, _17023_);
  nand (_32417_, _32406_, _17056_);
  or (_32428_, _32406_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and (_32439_, _32428_, _32417_);
  or (_32450_, _32439_, _32351_);
  nand (_32461_, _32351_, _27325_);
  and (_32472_, _32461_, _37580_);
  and (_37528_, _32472_, _32450_);
  and (_32513_, \oc8051_top_1.oc8051_memory_interface1.reti , \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  and (_32524_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _37580_);
  and (_37547_, _32524_, _32513_);
  not (_32545_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_32556_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and (_32567_, _32556_, _32545_);
  not (_32578_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_32589_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_32600_, _32589_, _32578_);
  nor (_32611_, _32600_, _32567_);
  not (_32622_, _32611_);
  not (_32633_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_32644_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and (_32655_, _32644_, _32633_);
  not (_32666_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and (_32677_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and (_32687_, _32677_, _32666_);
  or (_32698_, _32687_, _32655_);
  or (_32709_, _32698_, _32622_);
  and (_32720_, _32709_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  not (_32731_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  and (_32742_, _32556_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_32753_, _32589_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  nor (_32764_, _32753_, _32742_);
  not (_32775_, _32764_);
  and (_32786_, _32644_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_32797_, _32677_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_32808_, _32797_, _32786_);
  nor (_32819_, _32808_, _32775_);
  nand (_32830_, _32819_, _32731_);
  or (_32841_, _32830_, _32720_);
  not (_32852_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_32863_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _32852_);
  nand (_32874_, _32863_, _32513_);
  and (_32885_, _32874_, _37580_);
  and (_37549_, _32885_, _32841_);
  and (_32906_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_32917_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _32852_);
  nor (_32928_, _32917_, _32906_);
  and (_32939_, _32928_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  nor (_32950_, _32939_, _32731_);
  nor (_32961_, _32950_, _32819_);
  not (_32972_, _32797_);
  and (_32983_, _32972_, _32764_);
  and (_32994_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], _32852_);
  or (_33005_, _32994_, _32983_);
  and (_33016_, _32786_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_33027_, _32775_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  or (_33038_, _33027_, _33016_);
  and (_33048_, _33038_, _33005_);
  and (_33059_, _33048_, _32961_);
  or (_33070_, _33059_, _32513_);
  and (_33081_, _32655_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_33092_, _33081_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  and (_33103_, _32687_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_33114_, _33103_, _32622_);
  and (_33125_, _33114_, _33092_);
  and (_33136_, _32994_, _32622_);
  or (_33147_, _33136_, _33125_);
  and (_33158_, _32720_, _32731_);
  and (_33169_, _33158_, _32819_);
  and (_33180_, _33169_, _33147_);
  nor (_33191_, _33158_, _32961_);
  and (_33202_, _33191_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  or (_33213_, _33202_, _33180_);
  or (_33224_, _33213_, _33070_);
  not (_33235_, _32513_);
  or (_33246_, _33235_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  and (_33257_, _33246_, _37580_);
  and (_37551_, _33257_, _33224_);
  and (_33278_, _32243_, _22731_);
  and (_33289_, _33278_, _17793_);
  nand (_33300_, _33289_, _17056_);
  and (_33311_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and (_33322_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _32852_);
  and (_33333_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_33344_, _33333_, _33322_);
  nor (_33355_, _33344_, _32731_);
  nand (_33365_, _33355_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  and (_33376_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _32852_);
  and (_33387_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_33398_, _33387_, _33376_);
  nor (_33409_, _33398_, _32731_);
  and (_33420_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_33431_, _33420_, _32994_);
  nand (_33442_, _33431_, _33409_);
  or (_33453_, _33442_, _33365_);
  and (_33464_, _33453_, _33311_);
  or (_33475_, _33464_, _33289_);
  and (_33486_, _33475_, _33300_);
  and (_33497_, _32221_, _22731_);
  or (_33508_, _33497_, _33486_);
  nand (_33519_, _33497_, _28460_);
  and (_33530_, _33519_, _37580_);
  and (_37571_, _33530_, _33508_);
  not (_33551_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  or (_33562_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff , _33551_);
  nor (_33573_, _33431_, _32731_);
  or (_33584_, _33573_, _33409_);
  or (_33595_, _33584_, _33365_);
  and (_33606_, _33595_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or (_33617_, _33606_, _33562_);
  nand (_33628_, _33278_, _17425_);
  and (_33639_, _33628_, _33617_);
  nor (_33650_, _33628_, _17056_);
  or (_33661_, _33650_, _33497_);
  or (_33672_, _33661_, _33639_);
  nand (_33683_, _33497_, _25213_);
  and (_33693_, _33683_, _37580_);
  and (_37573_, _33693_, _33672_);
  not (_33714_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  or (_33725_, _33355_, _33714_);
  or (_33736_, _33725_, _33442_);
  and (_33747_, _33736_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  nand (_33758_, _33278_, _18140_);
  and (_33769_, _33758_, _33747_);
  and (_33780_, _33278_, _18173_);
  or (_33791_, _33780_, _33497_);
  or (_33802_, _33791_, _33769_);
  nand (_33813_, _33497_, _25755_);
  and (_33824_, _33813_, _37580_);
  and (_37575_, _33824_, _33802_);
  nand (_33845_, _33573_, _33398_);
  or (_33856_, _33845_, _33725_);
  and (_33867_, _33856_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  nand (_33878_, _33278_, _17023_);
  and (_33889_, _33878_, _33867_);
  and (_33900_, _33278_, _24953_);
  or (_33911_, _33900_, _33497_);
  or (_33922_, _33911_, _33889_);
  nand (_33933_, _33497_, _27325_);
  and (_33944_, _33933_, _37580_);
  and (_37576_, _33944_, _33922_);
  nand (_33965_, _33278_, _18314_);
  and (_33976_, _33965_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and (_33987_, _33278_, _18346_);
  or (_33997_, _33987_, _33497_);
  or (_34008_, _33997_, _33976_);
  nand (_34019_, _33497_, _28946_);
  and (_34030_, _34019_, _37580_);
  and (_37578_, _34030_, _34008_);
  and (_34051_, _33191_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  and (_34062_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _32852_);
  nor (_34073_, _34062_, _32863_);
  not (_34084_, _34073_);
  and (_34095_, _34084_, _32961_);
  or (_34106_, _34095_, _32513_);
  or (_34117_, _34106_, _34051_);
  or (_34128_, _34073_, _33235_);
  and (_34139_, _34128_, _37580_);
  and (_37582_, _34139_, _34117_);
  and (_34160_, _33191_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  or (_34171_, _33420_, _32983_);
  and (_34182_, _32786_, _32852_);
  or (_34193_, _32775_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  or (_34204_, _34193_, _34182_);
  and (_34215_, _34204_, _34171_);
  and (_34226_, _34215_, _32961_);
  or (_34237_, _34226_, _34160_);
  and (_34248_, _32655_, _32852_);
  or (_34259_, _34248_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  and (_34270_, _32687_, _32852_);
  nor (_34281_, _34270_, _32622_);
  and (_34292_, _34281_, _34259_);
  and (_34302_, _33420_, _32622_);
  or (_34313_, _34302_, _34292_);
  and (_34324_, _34313_, _33169_);
  or (_34335_, _34324_, _32513_);
  or (_34346_, _34335_, _34237_);
  or (_34357_, _33235_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  and (_34368_, _34357_, _37580_);
  and (_37584_, _34368_, _34346_);
  nor (_34389_, _32513_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_34400_, _34389_, _32961_);
  nand (_34411_, _33158_, _32852_);
  and (_34422_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [1], _37580_);
  nand (_34433_, _34422_, _34411_);
  nor (_37586_, _34433_, _34400_);
  nor (_34454_, _32513_, _32852_);
  and (_34465_, _34454_, _32961_);
  nand (_34476_, _33158_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_34487_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [1], _37580_);
  nand (_34498_, _34487_, _34476_);
  nor (_37588_, _34498_, _34465_);
  nor (_34529_, _33191_, _32513_);
  and (_34540_, _32513_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  or (_34551_, _34540_, _34529_);
  and (_38571_, _34551_, _37580_);
  and (_34572_, _32513_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  or (_34583_, _34572_, _34529_);
  and (_38573_, _34583_, _37580_);
  and (_34603_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _37580_);
  and (_38575_, _34603_, _32513_);
  not (_34624_, _32600_);
  nor (_34635_, _32655_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nor (_34646_, _34635_, _32687_);
  or (_34657_, _34646_, _32567_);
  and (_34668_, _34657_, _34624_);
  and (_34679_, _34668_, _33169_);
  not (_34690_, _32753_);
  or (_34701_, _32786_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_34712_, _34701_, _32972_);
  or (_34723_, _34712_, _32742_);
  and (_34734_, _34723_, _34690_);
  and (_34745_, _34734_, _32961_);
  or (_34756_, _34745_, _32513_);
  or (_34767_, _34756_, _34679_);
  or (_34778_, _33235_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_34789_, _34778_, _37580_);
  and (_38577_, _34789_, _34767_);
  or (_34810_, _32698_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and (_34821_, _34810_, _32611_);
  and (_34832_, _34821_, _33169_);
  or (_34843_, _32808_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and (_34854_, _34843_, _32764_);
  and (_34865_, _34854_, _32961_);
  or (_34876_, _34865_, _32513_);
  or (_34887_, _34876_, _34832_);
  or (_34898_, _33235_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and (_34908_, _34898_, _37580_);
  and (_38579_, _34908_, _34887_);
  and (_34929_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], _37580_);
  and (_38581_, _34929_, _32513_);
  and (_34950_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _37580_);
  and (_38583_, _34950_, _32513_);
  nand (_34971_, _34389_, _33191_);
  nor (_34982_, _32961_, _32513_);
  or (_34993_, _34982_, _32852_);
  and (_35004_, _34993_, _37580_);
  and (_38585_, _35004_, _34971_);
  not (_35025_, _34529_);
  and (_35036_, _35025_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  not (_35047_, _34182_);
  and (_35058_, _35047_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  and (_35069_, _32797_, _32852_);
  or (_35080_, _35069_, _32742_);
  or (_35091_, _35080_, _35058_);
  not (_35102_, _32742_);
  or (_35113_, _33333_, _35102_);
  and (_35124_, _35113_, _35091_);
  or (_35135_, _35124_, _32753_);
  or (_35146_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _32852_);
  or (_35157_, _35146_, _34690_);
  and (_35168_, _35157_, _32961_);
  and (_35179_, _35168_, _35135_);
  not (_35190_, _34248_);
  and (_35201_, _35190_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  or (_35212_, _34270_, _32567_);
  or (_35219_, _35212_, _35201_);
  not (_35227_, _32567_);
  or (_35235_, _33333_, _35227_);
  and (_35242_, _35235_, _34624_);
  and (_35250_, _35242_, _35219_);
  and (_35259_, _35146_, _32600_);
  or (_35266_, _35259_, _35250_);
  and (_35274_, _35266_, _33169_);
  or (_35278_, _35274_, _35179_);
  and (_35279_, _35278_, _33235_);
  or (_35280_, _35279_, _35036_);
  and (_38587_, _35280_, _37580_);
  and (_35298_, _35047_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  or (_35309_, _35298_, _35080_);
  or (_35320_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _32852_);
  or (_35331_, _35320_, _35102_);
  and (_35342_, _35331_, _35309_);
  or (_35353_, _35342_, _32753_);
  or (_35364_, _33387_, _34690_);
  and (_35375_, _35364_, _32961_);
  and (_35386_, _35375_, _35353_);
  and (_35397_, _33191_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  or (_35408_, _35397_, _35386_);
  and (_35419_, _35408_, _33235_);
  and (_35430_, _32513_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_35442_, _35190_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  or (_35453_, _35442_, _35212_);
  or (_35464_, _35320_, _35227_);
  and (_35475_, _35464_, _34624_);
  and (_35486_, _35475_, _35453_);
  and (_35497_, _33387_, _32600_);
  or (_35508_, _35497_, _35486_);
  and (_35519_, _35508_, _33169_);
  or (_35530_, _35519_, _35430_);
  or (_35541_, _35530_, _35419_);
  and (_38589_, _35541_, _37580_);
  and (_35562_, _35025_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  not (_35573_, _33016_);
  and (_35584_, _35573_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  and (_35595_, _32797_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_35606_, _35595_, _32742_);
  or (_35617_, _35606_, _35584_);
  or (_35628_, _33322_, _35102_);
  and (_35639_, _35628_, _35617_);
  or (_35650_, _35639_, _32753_);
  or (_35651_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_35652_, _35651_, _34690_);
  and (_35653_, _35652_, _32961_);
  and (_35654_, _35653_, _35650_);
  not (_35655_, _33081_);
  and (_35656_, _35655_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  or (_35657_, _33103_, _32567_);
  or (_35658_, _35657_, _35656_);
  or (_35659_, _33322_, _35227_);
  and (_35660_, _35659_, _34624_);
  and (_35661_, _35660_, _35658_);
  and (_35662_, _35651_, _32600_);
  or (_35663_, _35662_, _35661_);
  and (_35664_, _35663_, _33169_);
  or (_35665_, _35664_, _35654_);
  and (_35666_, _35665_, _33235_);
  or (_35667_, _35666_, _35562_);
  and (_38591_, _35667_, _37580_);
  and (_35668_, _35573_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  or (_35669_, _35668_, _35606_);
  or (_35670_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_35671_, _35670_, _35102_);
  and (_35672_, _35671_, _35669_);
  or (_35673_, _35672_, _32753_);
  or (_35674_, _33376_, _34690_);
  and (_35675_, _35674_, _32961_);
  and (_35676_, _35675_, _35673_);
  and (_35677_, _33191_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  or (_35678_, _35677_, _35676_);
  and (_35679_, _35678_, _33235_);
  and (_35680_, _32513_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_35681_, _35655_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  or (_35682_, _35681_, _35657_);
  or (_35683_, _35670_, _35227_);
  and (_35684_, _35683_, _34624_);
  and (_35685_, _35684_, _35682_);
  and (_35686_, _33376_, _32600_);
  or (_35687_, _35686_, _35685_);
  and (_35688_, _35687_, _33169_);
  or (_35689_, _35688_, _35680_);
  or (_35690_, _35689_, _35679_);
  and (_38593_, _35690_, _37580_);
  and (_35691_, _34411_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0]);
  or (_35692_, _35691_, _34400_);
  and (_38595_, _35692_, _37580_);
  and (_35693_, _34476_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0]);
  or (_35694_, _35693_, _34465_);
  and (_38597_, _35694_, _37580_);
  and (_35695_, _33278_, _17143_);
  nand (_35696_, _35695_, _17056_);
  or (_35697_, _35695_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and (_35698_, _35697_, _35696_);
  or (_35699_, _35698_, _33497_);
  nand (_35700_, _33497_, _29043_);
  and (_35701_, _35700_, _37580_);
  and (_38599_, _35701_, _35699_);
  nand (_35702_, _33278_, _17620_);
  and (_35703_, _35702_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and (_35704_, _33278_, _17653_);
  or (_35705_, _35704_, _33497_);
  or (_35706_, _35705_, _35703_);
  nand (_35707_, _33497_, _28385_);
  and (_35708_, _35707_, _37580_);
  and (_38601_, _35708_, _35706_);
  nand (_35709_, _33278_, _17967_);
  and (_35710_, _35709_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and (_35711_, _33278_, _18000_);
  or (_35712_, _35711_, _33497_);
  or (_35713_, _35712_, _35710_);
  nand (_35714_, _33497_, _28655_);
  and (_35715_, _35714_, _37580_);
  and (_38603_, _35715_, _35713_);
  nand (_35716_, _32254_, _17143_);
  and (_35717_, _35716_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_35718_, _32254_, _17284_);
  or (_35719_, _35718_, _32232_);
  or (_35720_, _35719_, _35717_);
  nand (_35721_, _32232_, _29043_);
  and (_35722_, _35721_, _37580_);
  and (_38605_, _35722_, _35720_);
  nand (_35723_, _32254_, _17425_);
  and (_35724_, _35723_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_35725_, _32254_, _17467_);
  or (_35726_, _35725_, _32232_);
  or (_35727_, _35726_, _35724_);
  nand (_35728_, _32232_, _25213_);
  and (_35729_, _35728_, _37580_);
  and (_38607_, _35729_, _35727_);
  nand (_35730_, _32254_, _17620_);
  and (_35731_, _35730_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and (_35732_, _32254_, _17653_);
  or (_35733_, _35732_, _32232_);
  or (_35734_, _35733_, _35731_);
  nand (_35735_, _32232_, _28385_);
  and (_35736_, _35735_, _37580_);
  and (_38609_, _35736_, _35734_);
  nand (_35737_, _32254_, _17793_);
  and (_35738_, _35737_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_35739_, _32254_, _17826_);
  or (_35740_, _35739_, _32232_);
  or (_35741_, _35740_, _35738_);
  nand (_35742_, _32232_, _28460_);
  and (_35743_, _35742_, _37580_);
  and (_38611_, _35743_, _35741_);
  and (_35744_, _32254_, _17967_);
  or (_35745_, _35744_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  nand (_35746_, _35744_, _17056_);
  and (_35747_, _35746_, _35745_);
  or (_35748_, _35747_, _32232_);
  nand (_35749_, _32232_, _28655_);
  and (_35750_, _35749_, _37580_);
  and (_38613_, _35750_, _35748_);
  nand (_35751_, _32254_, _18140_);
  and (_35752_, _35751_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and (_35753_, _32254_, _18173_);
  or (_35754_, _35753_, _32232_);
  or (_35755_, _35754_, _35752_);
  nand (_35756_, _32232_, _25755_);
  and (_35757_, _35756_, _37580_);
  and (_38615_, _35757_, _35755_);
  nand (_35758_, _32254_, _18314_);
  and (_35759_, _35758_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_35760_, _32254_, _18346_);
  or (_35761_, _35760_, _32232_);
  or (_35762_, _35761_, _35759_);
  nand (_35763_, _32232_, _28946_);
  and (_35764_, _35763_, _37580_);
  and (_38617_, _35764_, _35762_);
  nand (_35765_, _32395_, _17143_);
  and (_35766_, _35765_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_35767_, _32395_, _17284_);
  or (_35768_, _35767_, _32351_);
  or (_35769_, _35768_, _35766_);
  nand (_35770_, _32351_, _29043_);
  and (_35771_, _35770_, _37580_);
  and (_38619_, _35771_, _35769_);
  nand (_35772_, _32395_, _17425_);
  and (_35773_, _35772_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_35774_, _32395_, _17467_);
  or (_35775_, _35774_, _32351_);
  or (_35776_, _35775_, _35773_);
  nand (_35777_, _32351_, _25213_);
  and (_35778_, _35777_, _37580_);
  and (_38621_, _35778_, _35776_);
  and (_35779_, _32395_, _17620_);
  or (_35780_, _35779_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  nand (_35791_, _35779_, _17056_);
  and (_35793_, _35791_, _35780_);
  or (_35794_, _35793_, _32351_);
  nand (_35795_, _32351_, _28385_);
  and (_35796_, _35795_, _37580_);
  and (_38623_, _35796_, _35794_);
  nand (_35797_, _32395_, _17793_);
  and (_35798_, _35797_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_35799_, _32395_, _17826_);
  or (_35800_, _35799_, _32351_);
  or (_35801_, _35800_, _35798_);
  nand (_35802_, _32351_, _28460_);
  and (_35803_, _35802_, _37580_);
  and (_38625_, _35803_, _35801_);
  and (_35804_, _32395_, _17967_);
  or (_35805_, _35804_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  nand (_35806_, _35804_, _17056_);
  and (_35807_, _35806_, _35805_);
  or (_35808_, _35807_, _32351_);
  nand (_35809_, _32351_, _28655_);
  and (_35810_, _35809_, _37580_);
  and (_38626_, _35810_, _35808_);
  nand (_35811_, _32395_, _18140_);
  and (_35812_, _35811_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_35813_, _32395_, _18173_);
  or (_35814_, _35813_, _32351_);
  or (_35815_, _35814_, _35812_);
  nand (_35816_, _32351_, _25755_);
  and (_35817_, _35816_, _37580_);
  and (_38628_, _35817_, _35815_);
  nand (_35818_, _32395_, _18314_);
  and (_35819_, _35818_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and (_35820_, _32395_, _18346_);
  or (_35821_, _35820_, _32351_);
  or (_35822_, _35821_, _35819_);
  nand (_35823_, _32351_, _28946_);
  and (_35824_, _35823_, _37580_);
  and (_38630_, _35824_, _35822_);
  and (_35825_, _22655_, _22501_);
  not (_35826_, _23202_);
  and (_35827_, _35826_, _35825_);
  not (_35828_, _35827_);
  and (_35829_, _22655_, _21544_);
  not (_35830_, _35829_);
  nor (_35831_, _35830_, _22490_);
  not (_35832_, _18553_);
  and (_35833_, _35832_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [7]);
  and (_35834_, _18640_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_35835_, _18684_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor (_35836_, _35835_, _35834_);
  and (_35837_, _18727_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_35838_, _18771_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_35839_, _35838_, _35837_);
  and (_35840_, _35839_, _35836_);
  and (_35841_, _18825_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_35842_, _18836_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  nor (_35843_, _35842_, _35841_);
  and (_35844_, _35843_, _35840_);
  and (_35845_, _19284_, _18553_);
  not (_35846_, _35845_);
  nor (_35847_, _35846_, _35844_);
  nor (_35848_, _35847_, _35833_);
  not (_35849_, _35848_);
  and (_35850_, _35849_, _35831_);
  not (_35851_, _35850_);
  not (_35852_, _22655_);
  not (_35853_, _21544_);
  and (_35854_, _22490_, _35853_);
  and (_35855_, _25440_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  nor (_35856_, _35855_, _25582_);
  nor (_35857_, _35856_, _16435_);
  and (_35858_, _35856_, _16435_);
  nor (_35859_, _35858_, _35857_);
  and (_35860_, _19724_, _16882_);
  not (_35861_, _35860_);
  nor (_35862_, _16762_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and (_35863_, _35862_, _17002_);
  nor (_35864_, _19724_, _16882_);
  and (_35865_, _15597_, _16229_);
  not (_35866_, _35865_);
  nor (_35867_, _35866_, _35864_);
  and (_35868_, _35867_, _35863_);
  and (_35869_, _35868_, _35861_);
  and (_35870_, _35869_, _35859_);
  and (_35871_, _35856_, _19724_);
  and (_35872_, _35871_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  nor (_35873_, _35856_, _19724_);
  and (_35874_, _35873_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  nor (_35875_, _35874_, _35872_);
  nor (_35876_, _35856_, _20781_);
  and (_35877_, _35876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  and (_35878_, _35856_, _20781_);
  and (_35879_, _35878_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  nor (_35880_, _35879_, _35877_);
  and (_35881_, _35880_, _35875_);
  nor (_35882_, _35881_, _35870_);
  and (_35883_, _35870_, ABINPUT[10]);
  nor (_35884_, _35883_, _35882_);
  not (_35885_, _35884_);
  and (_35886_, _35885_, _35854_);
  nor (_35887_, _35886_, _35852_);
  and (_35888_, _35887_, _35851_);
  and (_35889_, _35888_, _35828_);
  and (_35890_, _20825_, _20858_);
  and (_35891_, _35890_, _19746_);
  nor (_35892_, _35891_, _22083_);
  and (_35893_, _35892_, _22072_);
  and (_35894_, _21907_, _19746_);
  nor (_35895_, _22391_, _35894_);
  and (_35896_, _35895_, _21621_);
  nor (_35897_, _21764_, _21643_);
  nor (_35898_, _22204_, _21566_);
  and (_35899_, _35898_, _35897_);
  and (_35900_, _35899_, _35896_);
  and (_35901_, _35900_, _35893_);
  nor (_35902_, _35901_, _18509_);
  not (_35903_, _21479_);
  nor (_35904_, _35895_, _35903_);
  nor (_35905_, _35904_, _35902_);
  not (_35906_, _35905_);
  and (_35907_, _35906_, _35889_);
  not (_35908_, _23676_);
  and (_35909_, _35908_, _35825_);
  and (_35910_, _35832_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [5]);
  and (_35911_, _18836_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  and (_35912_, _18727_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  nor (_35913_, _35912_, _35911_);
  and (_35914_, _18640_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_35915_, _18684_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_35916_, _35915_, _35914_);
  and (_35917_, _18825_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_35918_, _18771_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_35919_, _35918_, _35917_);
  and (_35920_, _35919_, _35916_);
  and (_35921_, _35920_, _35913_);
  nor (_35922_, _35921_, _35846_);
  nor (_35923_, _35922_, _35910_);
  not (_35924_, _35923_);
  and (_35925_, _35924_, _35831_);
  nor (_35926_, _35925_, _35909_);
  and (_35927_, _35852_, _21544_);
  and (_35928_, _35927_, _22490_);
  and (_35929_, _35852_, _22501_);
  or (_35930_, _35929_, _35928_);
  and (_35931_, _35854_, _22655_);
  and (_35932_, _35871_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  and (_35933_, _35873_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  nor (_35934_, _35933_, _35932_);
  and (_35935_, _35876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  and (_35936_, _35878_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nor (_35937_, _35936_, _35935_);
  and (_35938_, _35937_, _35934_);
  nor (_35939_, _35938_, _35870_);
  and (_35940_, _35870_, ABINPUT[8]);
  nor (_35941_, _35940_, _35939_);
  not (_35942_, _35941_);
  and (_35943_, _35942_, _35931_);
  nor (_35944_, _35943_, _35930_);
  and (_35945_, _35944_, _35926_);
  not (_35946_, _35945_);
  and (_35947_, _35946_, _35907_);
  and (_35948_, _35871_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  and (_35949_, _35873_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  nor (_35950_, _35949_, _35948_);
  and (_35951_, _35876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  and (_35952_, _35878_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  nor (_35953_, _35952_, _35951_);
  and (_35954_, _35953_, _35950_);
  nor (_35955_, _35954_, _35870_);
  and (_35956_, _35870_, ABINPUT[5]);
  nor (_35957_, _35956_, _35955_);
  not (_35958_, _35957_);
  and (_35959_, _35958_, _35931_);
  not (_35960_, _35959_);
  and (_35961_, _35829_, _22490_);
  and (_35962_, _35961_, _18957_);
  not (_35963_, _23450_);
  and (_35964_, _35963_, _35825_);
  and (_35965_, _35832_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [2]);
  and (_35966_, _18640_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_35967_, _18684_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_35968_, _35967_, _35966_);
  and (_35969_, _18727_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_35970_, _18771_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_35971_, _35970_, _35969_);
  and (_35972_, _35971_, _35968_);
  and (_35973_, _18825_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_35974_, _18836_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  nor (_35975_, _35974_, _35973_);
  and (_35976_, _35975_, _35972_);
  nor (_35977_, _35976_, _35846_);
  nor (_35978_, _35977_, _35965_);
  not (_35979_, _35978_);
  and (_35980_, _35979_, _35831_);
  or (_35981_, _35980_, _35964_);
  nor (_35982_, _35981_, _35962_);
  and (_35983_, _35982_, _35960_);
  nor (_35984_, _35983_, _35906_);
  nor (_35985_, _35984_, _35947_);
  and (_35986_, _16250_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_35987_, _35986_, _25528_);
  nor (_35988_, _16751_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_35989_, _35988_, _35987_);
  not (_35990_, _35989_);
  and (_35991_, _35990_, _35985_);
  not (_35992_, _23526_);
  and (_35993_, _35992_, _35825_);
  not (_35994_, _35993_);
  not (_35995_, _35856_);
  and (_35996_, _35961_, _35995_);
  and (_35997_, _35871_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  and (_35998_, _35873_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  nor (_35999_, _35998_, _35997_);
  and (_36000_, _35876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  and (_36001_, _35878_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  nor (_36002_, _36001_, _36000_);
  and (_36003_, _36002_, _35999_);
  nor (_36004_, _36003_, _35870_);
  and (_36005_, _35870_, ABINPUT[6]);
  nor (_36006_, _36005_, _36004_);
  not (_36007_, _36006_);
  and (_36008_, _36007_, _35931_);
  and (_36009_, _35832_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [3]);
  and (_36010_, _18640_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_36011_, _18684_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_36012_, _36011_, _36010_);
  and (_36013_, _18727_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_36014_, _18771_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_36015_, _36014_, _36013_);
  and (_36016_, _36015_, _36012_);
  and (_36017_, _18825_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_36018_, _18836_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor (_36019_, _36018_, _36017_);
  and (_36020_, _36019_, _36016_);
  nor (_36021_, _36020_, _35846_);
  nor (_36022_, _36021_, _36009_);
  not (_36023_, _36022_);
  and (_36024_, _36023_, _35831_);
  or (_36025_, _36024_, _36008_);
  nor (_36026_, _36025_, _35996_);
  and (_36027_, _36026_, _35994_);
  not (_36028_, _36027_);
  and (_36029_, _36028_, _35907_);
  not (_36030_, _23300_);
  and (_36031_, _36030_, _35825_);
  not (_36032_, _36031_);
  and (_36033_, _35961_, _19724_);
  and (_36034_, _35873_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  and (_36035_, _35871_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  nor (_36036_, _36035_, _36034_);
  and (_36037_, _35876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  and (_36038_, _35878_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  nor (_36039_, _36038_, _36037_);
  and (_36040_, _36039_, _36036_);
  nor (_36041_, _36040_, _35870_);
  and (_36042_, _35870_, ABINPUT[3]);
  nor (_36043_, _36042_, _36041_);
  not (_36044_, _36043_);
  and (_36045_, _36044_, _35931_);
  and (_36046_, _35832_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [0]);
  and (_36047_, _18640_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_36048_, _18684_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_36049_, _36048_, _36047_);
  and (_36050_, _18727_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_36051_, _18771_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_36052_, _36051_, _36050_);
  and (_36053_, _36052_, _36049_);
  and (_36054_, _18825_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_36055_, _18836_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor (_36056_, _36055_, _36054_);
  and (_36057_, _36056_, _36053_);
  nor (_36058_, _36057_, _35846_);
  nor (_36059_, _36058_, _36046_);
  not (_36060_, _36059_);
  and (_36061_, _36060_, _35831_);
  or (_36062_, _36061_, _36045_);
  nor (_36063_, _36062_, _36033_);
  and (_36064_, _36063_, _36032_);
  nor (_36065_, _36064_, _35906_);
  nor (_36066_, _36065_, _36029_);
  and (_36067_, _35986_, _16435_);
  nor (_36068_, _16882_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_36069_, _36068_, _36067_);
  not (_36070_, _36069_);
  nor (_36071_, _36070_, _36066_);
  nor (_36072_, _36071_, _35991_);
  nor (_36073_, _35990_, _35985_);
  not (_36074_, _36073_);
  not (_36075_, _23752_);
  and (_36076_, _36075_, _35825_);
  and (_36077_, _35832_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [6]);
  and (_36078_, _18727_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_36079_, _18771_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_36080_, _36079_, _36078_);
  and (_36081_, _18640_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_36082_, _18684_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor (_36083_, _36082_, _36081_);
  and (_36084_, _18825_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_36085_, _18836_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor (_36086_, _36085_, _36084_);
  and (_36087_, _36086_, _36083_);
  and (_36088_, _36087_, _36080_);
  nor (_36089_, _36088_, _35846_);
  nor (_36090_, _36089_, _36077_);
  not (_36091_, _36090_);
  and (_36092_, _36091_, _35831_);
  nor (_36093_, _36092_, _36076_);
  nor (_36094_, _35854_, _22655_);
  and (_36095_, _35871_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  and (_36096_, _35873_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  nor (_36097_, _36096_, _36095_);
  and (_36098_, _35876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  and (_36099_, _35878_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  nor (_36100_, _36099_, _36098_);
  and (_36101_, _36100_, _36097_);
  nor (_36102_, _36101_, _35870_);
  and (_36103_, _35870_, ABINPUT[9]);
  nor (_36104_, _36103_, _36102_);
  not (_36105_, _36104_);
  and (_36106_, _36105_, _35931_);
  nor (_36107_, _36106_, _36094_);
  and (_36108_, _36107_, _36093_);
  and (_36109_, _36108_, _35907_);
  nor (_36110_, _36028_, _35907_);
  nor (_36111_, _36110_, _36109_);
  nor (_36112_, _35986_, _16435_);
  and (_36113_, _35986_, _16076_);
  nor (_36114_, _36113_, _36112_);
  not (_36115_, _36114_);
  and (_36116_, _36115_, _36111_);
  nor (_36117_, _36115_, _36111_);
  nor (_36118_, _36117_, _36116_);
  and (_36119_, _36118_, _36074_);
  and (_36120_, _35873_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  and (_36121_, _35878_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  nor (_36122_, _36121_, _36120_);
  and (_36123_, _35876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  and (_36124_, _35871_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  nor (_36125_, _36124_, _36123_);
  and (_36126_, _36125_, _36122_);
  nor (_36127_, _36126_, _35870_);
  and (_36128_, _35870_, ABINPUT[7]);
  nor (_36129_, _36128_, _36127_);
  not (_36130_, _36129_);
  and (_36131_, _36130_, _35931_);
  not (_36132_, _36131_);
  not (_36133_, _23601_);
  and (_36134_, _36133_, _35825_);
  nor (_36135_, _36134_, _35927_);
  and (_36136_, _25440_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  nor (_36137_, _36136_, _25668_);
  not (_36138_, _36137_);
  and (_36139_, _36138_, _35961_);
  and (_36140_, _35832_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [4]);
  and (_36141_, _18727_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_36142_, _18771_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_36143_, _36142_, _36141_);
  and (_36144_, _18640_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_36145_, _18684_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_36146_, _36145_, _36144_);
  and (_36147_, _18825_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_36148_, _18836_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  nor (_36149_, _36148_, _36147_);
  and (_36150_, _36149_, _36146_);
  and (_36151_, _36150_, _36143_);
  nor (_36152_, _36151_, _35846_);
  nor (_36153_, _36152_, _36140_);
  not (_36154_, _36153_);
  and (_36155_, _36154_, _35831_);
  nor (_36156_, _36155_, _36139_);
  and (_36157_, _36156_, _36135_);
  and (_36158_, _36157_, _36132_);
  not (_36159_, _36158_);
  and (_36160_, _36159_, _35907_);
  and (_36161_, _35961_, _19484_);
  not (_36162_, _36161_);
  and (_36163_, _35854_, _35852_);
  and (_36164_, _35832_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [1]);
  and (_36165_, _18640_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_36166_, _18684_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_36167_, _36166_, _36165_);
  and (_36168_, _18727_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_36169_, _18771_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_36170_, _36169_, _36168_);
  and (_36171_, _36170_, _36167_);
  and (_36172_, _18825_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_36173_, _18836_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor (_36174_, _36173_, _36172_);
  and (_36175_, _36174_, _36171_);
  nor (_36176_, _36175_, _35846_);
  nor (_36177_, _36176_, _36164_);
  not (_36178_, _36177_);
  and (_36179_, _36178_, _35831_);
  nor (_36180_, _36179_, _36163_);
  and (_36181_, _36180_, _36162_);
  not (_36182_, _23375_);
  and (_36183_, _36182_, _35825_);
  and (_36184_, _35871_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  and (_36185_, _35873_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  nor (_36186_, _36185_, _36184_);
  and (_36187_, _35876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  and (_36188_, _35878_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  nor (_36189_, _36188_, _36187_);
  and (_36190_, _36189_, _36186_);
  nor (_36191_, _36190_, _35870_);
  and (_36192_, _35870_, ABINPUT[4]);
  nor (_36193_, _36192_, _36191_);
  not (_36194_, _36193_);
  and (_36195_, _36194_, _35931_);
  nor (_36196_, _36195_, _36183_);
  and (_36197_, _36196_, _36181_);
  nor (_36198_, _36197_, _35906_);
  nor (_36199_, _36198_, _36160_);
  and (_36200_, _35986_, _32362_);
  nor (_36201_, _17002_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_36202_, _36201_, _36200_);
  nand (_36203_, _36202_, _36199_);
  or (_36204_, _36202_, _36199_);
  and (_36205_, _36204_, _36203_);
  not (_36206_, _36205_);
  and (_36207_, _36070_, _36066_);
  nor (_36208_, _36207_, _35866_);
  and (_36209_, _36208_, _36206_);
  and (_36210_, _36209_, _36119_);
  and (_36211_, _36210_, _36072_);
  not (_36212_, _35985_);
  and (_36213_, _36066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  not (_36214_, _36066_);
  and (_36215_, _36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  or (_36216_, _36215_, _36213_);
  and (_36217_, _36216_, _36199_);
  not (_36218_, _36199_);
  and (_36219_, _36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  and (_36220_, _36066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  or (_36221_, _36220_, _36219_);
  and (_36222_, _36221_, _36218_);
  or (_36223_, _36222_, _36217_);
  or (_36224_, _36223_, _36212_);
  not (_36225_, _36111_);
  and (_36226_, _36066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  and (_36227_, _36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  or (_36228_, _36227_, _36226_);
  and (_36229_, _36228_, _36199_);
  and (_36230_, _36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  and (_36231_, _36066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  or (_36232_, _36231_, _36230_);
  and (_36233_, _36232_, _36218_);
  or (_36234_, _36233_, _36229_);
  or (_36235_, _36234_, _35985_);
  and (_36236_, _36235_, _36225_);
  and (_36237_, _36236_, _36224_);
  or (_36238_, _36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  or (_36239_, _36066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  and (_36240_, _36239_, _36238_);
  and (_36241_, _36240_, _36199_);
  or (_36242_, _36066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  or (_36243_, _36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  and (_36244_, _36243_, _36242_);
  and (_36245_, _36244_, _36218_);
  or (_36246_, _36245_, _36241_);
  or (_36247_, _36246_, _36212_);
  or (_36248_, _36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  or (_36249_, _36066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  and (_36250_, _36249_, _36248_);
  and (_36251_, _36250_, _36199_);
  or (_36252_, _36066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  or (_36253_, _36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  and (_36254_, _36253_, _36252_);
  and (_36255_, _36254_, _36218_);
  or (_36256_, _36255_, _36251_);
  or (_36257_, _36256_, _35985_);
  and (_36258_, _36257_, _36111_);
  and (_36259_, _36258_, _36247_);
  or (_36260_, _36259_, _36237_);
  or (_36261_, _36260_, _36211_);
  not (_36262_, _36211_);
  or (_36263_, _36262_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  and (_36264_, _36263_, _37580_);
  and (_38712_, _36264_, _36261_);
  nor (_36265_, _36069_, _35866_);
  nor (_36266_, _36202_, _35866_);
  and (_36267_, _36266_, _36265_);
  and (_36268_, _36114_, _35865_);
  nor (_36269_, _35989_, _35866_);
  and (_36270_, _36269_, _36268_);
  and (_36271_, _36270_, _36267_);
  or (_36272_, _36271_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  not (_36273_, _36271_);
  and (_36274_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_36275_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_36276_, _36275_, _36274_);
  and (_36277_, _36276_, ABINPUT[0]);
  not (_36278_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_36279_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  not (_36280_, \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  nor (_36281_, _36280_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [7]);
  nor (_36282_, _36281_, _36279_);
  and (_36283_, _36274_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  not (_36284_, _36283_);
  and (_36285_, _36284_, _36282_);
  or (_36286_, _36285_, _36278_);
  or (_36287_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , ABINPUT[10]);
  and (_36288_, _36287_, _36286_);
  or (_36289_, _36288_, _36277_);
  and (_36290_, _36289_, _35865_);
  or (_36291_, _36290_, _36273_);
  and (_38724_, _36291_, _36272_);
  nor (_36292_, _36269_, _36268_);
  nor (_36293_, _36266_, _36265_);
  and (_36294_, _36293_, _35865_);
  and (_36295_, _36294_, _36292_);
  not (_36296_, _36295_);
  and (_36297_, _36296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  not (_36298_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_36299_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , _36298_);
  nor (_36300_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_36301_, _36300_, _36299_);
  and (_36302_, _36301_, ABINPUT[0]);
  and (_36303_, _36278_, ABINPUT[3]);
  or (_36304_, _36303_, _36302_);
  and (_36305_, _36300_, _36298_);
  nor (_36306_, _36305_, _36278_);
  nor (_36307_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  nor (_36308_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _36280_);
  nor (_36309_, _36308_, _36307_);
  and (_36310_, _36309_, _36306_);
  or (_36311_, _36310_, _36304_);
  and (_36312_, _36311_, _35865_);
  and (_36313_, _36312_, _36295_);
  or (_39004_, _36313_, _36297_);
  and (_36314_, _36296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  nor (_36315_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  nor (_36316_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _36280_);
  nor (_36317_, _36316_, _36315_);
  not (_36318_, \oc8051_top_1.oc8051_ram_top1.bit_select [0]);
  nor (_36319_, _36318_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_36320_, _36319_, _36298_);
  nor (_36321_, _36320_, _36278_);
  and (_36322_, _36321_, _36317_);
  and (_36323_, _36319_, _36299_);
  and (_36324_, _36323_, ABINPUT[0]);
  and (_36325_, _36278_, ABINPUT[4]);
  or (_36326_, _36325_, _36324_);
  or (_36327_, _36326_, _36322_);
  and (_36328_, _36327_, _35865_);
  and (_36329_, _36328_, _36295_);
  or (_39008_, _36329_, _36314_);
  and (_36330_, _36296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  nor (_36331_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  nor (_36332_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _36280_);
  nor (_36333_, _36332_, _36331_);
  and (_36334_, _36318_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_36335_, _36334_, _36298_);
  nor (_36336_, _36335_, _36278_);
  and (_36337_, _36336_, _36333_);
  and (_36338_, _36299_, _36334_);
  and (_36339_, _36338_, ABINPUT[0]);
  and (_36340_, _36278_, ABINPUT[5]);
  or (_36341_, _36340_, _36339_);
  or (_36342_, _36341_, _36337_);
  and (_36343_, _36342_, _35865_);
  and (_36344_, _36343_, _36295_);
  or (_39013_, _36344_, _36330_);
  and (_36345_, _36296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  and (_36346_, _36299_, _36274_);
  and (_36347_, _36346_, ABINPUT[0]);
  nor (_36348_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  nor (_36349_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _36280_);
  nor (_36350_, _36349_, _36348_);
  and (_36351_, _36274_, _36298_);
  not (_36352_, _36351_);
  and (_36353_, _36352_, _36350_);
  or (_36354_, _36353_, _36278_);
  or (_36355_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , ABINPUT[6]);
  and (_36356_, _36355_, _36354_);
  or (_36357_, _36356_, _36347_);
  and (_36358_, _36357_, _35865_);
  and (_36359_, _36358_, _36295_);
  or (_39019_, _36359_, _36345_);
  and (_36360_, _36296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  nor (_36361_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  nor (_36362_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _36280_);
  nor (_36363_, _36362_, _36361_);
  and (_36364_, _36300_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  nor (_36365_, _36364_, _36278_);
  and (_36366_, _36365_, _36363_);
  and (_36367_, _36300_, _36275_);
  and (_36368_, _36367_, ABINPUT[0]);
  and (_36369_, _36278_, ABINPUT[7]);
  or (_36370_, _36369_, _36368_);
  or (_36371_, _36370_, _36366_);
  and (_36372_, _36371_, _35865_);
  and (_36373_, _36372_, _36295_);
  or (_39025_, _36373_, _36360_);
  and (_36374_, _36296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nor (_36375_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  nor (_36376_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _36280_);
  nor (_36377_, _36376_, _36375_);
  and (_36378_, _36319_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  nor (_36379_, _36378_, _36278_);
  and (_36380_, _36379_, _36377_);
  and (_36381_, _36319_, _36275_);
  and (_36382_, _36381_, ABINPUT[0]);
  and (_36383_, _36278_, ABINPUT[8]);
  or (_36384_, _36383_, _36382_);
  or (_36385_, _36384_, _36380_);
  and (_36386_, _36385_, _35865_);
  and (_36387_, _36386_, _36295_);
  or (_39031_, _36387_, _36374_);
  and (_36388_, _36296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  nor (_36389_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  nor (_36390_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _36280_);
  nor (_36391_, _36390_, _36389_);
  and (_36392_, _36334_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  nor (_36393_, _36392_, _36278_);
  and (_36394_, _36393_, _36391_);
  and (_36395_, _36334_, _36275_);
  and (_36396_, _36395_, ABINPUT[0]);
  and (_36397_, _36278_, ABINPUT[9]);
  or (_36398_, _36397_, _36396_);
  or (_36399_, _36398_, _36394_);
  and (_36400_, _36399_, _35865_);
  and (_36401_, _36400_, _36295_);
  or (_39037_, _36401_, _36388_);
  and (_36402_, _36296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  and (_36403_, _36295_, _36290_);
  or (_39040_, _36403_, _36402_);
  and (_36404_, _36265_, _36202_);
  and (_36405_, _36404_, _36292_);
  or (_36406_, _36405_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  not (_36407_, _36405_);
  or (_36408_, _36407_, _36312_);
  and (_39048_, _36408_, _36406_);
  or (_36409_, _36405_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  or (_36410_, _36407_, _36328_);
  and (_39052_, _36410_, _36409_);
  or (_36411_, _36405_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  or (_36412_, _36407_, _36343_);
  and (_39056_, _36412_, _36411_);
  or (_36413_, _36405_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  or (_36414_, _36407_, _36358_);
  and (_39060_, _36414_, _36413_);
  or (_36415_, _36405_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  or (_36416_, _36407_, _36372_);
  and (_39064_, _36416_, _36415_);
  or (_36417_, _36405_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  or (_36418_, _36407_, _36386_);
  and (_39068_, _36418_, _36417_);
  or (_36419_, _36405_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  or (_36420_, _36407_, _36400_);
  and (_39072_, _36420_, _36419_);
  or (_36421_, _36405_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  or (_36422_, _36407_, _36290_);
  and (_39075_, _36422_, _36421_);
  and (_36423_, _36266_, _36069_);
  and (_36424_, _36423_, _36292_);
  or (_36425_, _36424_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  not (_36426_, _36424_);
  or (_36427_, _36426_, _36312_);
  and (_39083_, _36427_, _36425_);
  or (_36428_, _36424_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  or (_36429_, _36426_, _36328_);
  and (_39087_, _36429_, _36428_);
  or (_36430_, _36424_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  or (_36431_, _36426_, _36343_);
  and (_39091_, _36431_, _36430_);
  or (_36432_, _36424_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or (_36433_, _36426_, _36358_);
  and (_39095_, _36433_, _36432_);
  or (_36434_, _36424_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  or (_36435_, _36426_, _36372_);
  and (_39099_, _36435_, _36434_);
  or (_36436_, _36424_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  or (_36437_, _36426_, _36386_);
  and (_39103_, _36437_, _36436_);
  or (_36438_, _36424_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  or (_36439_, _36426_, _36400_);
  and (_39107_, _36439_, _36438_);
  or (_36440_, _36424_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  or (_36441_, _36426_, _36290_);
  and (_39110_, _36441_, _36440_);
  and (_36442_, _36292_, _36267_);
  or (_36443_, _36442_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  not (_36444_, _36442_);
  or (_36445_, _36444_, _36312_);
  and (_39116_, _36445_, _36443_);
  or (_36446_, _36442_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  or (_36447_, _36444_, _36328_);
  and (_39120_, _36447_, _36446_);
  or (_36448_, _36442_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  or (_36449_, _36444_, _36343_);
  and (_39124_, _36449_, _36448_);
  or (_36450_, _36442_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  or (_36451_, _36444_, _36358_);
  and (_39128_, _36451_, _36450_);
  or (_36452_, _36442_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  or (_36453_, _36444_, _36372_);
  and (_39132_, _36453_, _36452_);
  or (_36454_, _36442_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  or (_36455_, _36444_, _36386_);
  and (_39136_, _36455_, _36454_);
  or (_36456_, _36442_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  or (_36457_, _36444_, _36400_);
  and (_39140_, _36457_, _36456_);
  or (_36458_, _36442_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  or (_36459_, _36444_, _36290_);
  and (_39143_, _36459_, _36458_);
  and (_36460_, _36269_, _36115_);
  and (_36461_, _36460_, _36293_);
  or (_36462_, _36461_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  not (_36463_, _36461_);
  or (_36464_, _36463_, _36312_);
  and (_39151_, _36464_, _36462_);
  or (_36465_, _36461_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  or (_36466_, _36463_, _36328_);
  and (_39155_, _36466_, _36465_);
  or (_36467_, _36461_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  or (_36468_, _36463_, _36343_);
  and (_39159_, _36468_, _36467_);
  or (_36469_, _36461_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  or (_36470_, _36463_, _36358_);
  and (_39163_, _36470_, _36469_);
  or (_36471_, _36461_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  or (_36472_, _36463_, _36372_);
  and (_39167_, _36472_, _36471_);
  or (_36473_, _36461_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  or (_36474_, _36463_, _36386_);
  and (_39171_, _36474_, _36473_);
  or (_36475_, _36461_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  or (_36476_, _36463_, _36400_);
  and (_39175_, _36476_, _36475_);
  or (_36477_, _36461_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  or (_36478_, _36463_, _36290_);
  and (_39178_, _36478_, _36477_);
  and (_36479_, _36460_, _36404_);
  or (_36480_, _36479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  not (_36481_, _36479_);
  or (_36482_, _36481_, _36312_);
  and (_39183_, _36482_, _36480_);
  or (_36483_, _36479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  or (_36484_, _36481_, _36328_);
  and (_39187_, _36484_, _36483_);
  or (_36485_, _36479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  or (_36486_, _36481_, _36343_);
  and (_39191_, _36486_, _36485_);
  or (_36487_, _36479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  or (_36488_, _36481_, _36358_);
  and (_39195_, _36488_, _36487_);
  or (_36489_, _36479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  or (_36490_, _36481_, _36372_);
  and (_39199_, _36490_, _36489_);
  or (_36491_, _36479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  or (_36492_, _36481_, _36386_);
  and (_39203_, _36492_, _36491_);
  or (_36493_, _36479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  or (_36494_, _36481_, _36400_);
  and (_39207_, _36494_, _36493_);
  or (_36495_, _36479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  or (_36496_, _36481_, _36290_);
  and (_39210_, _36496_, _36495_);
  and (_36497_, _36460_, _36423_);
  or (_36498_, _36497_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  not (_36499_, _36497_);
  or (_36500_, _36499_, _36312_);
  and (_39215_, _36500_, _36498_);
  or (_36501_, _36497_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  or (_36502_, _36499_, _36328_);
  and (_39219_, _36502_, _36501_);
  or (_36503_, _36497_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  or (_36504_, _36499_, _36343_);
  and (_39222_, _36504_, _36503_);
  or (_36505_, _36497_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or (_36506_, _36499_, _36358_);
  and (_39226_, _36506_, _36505_);
  or (_36507_, _36497_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  or (_36508_, _36499_, _36372_);
  and (_39230_, _36508_, _36507_);
  or (_36509_, _36497_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  or (_36510_, _36499_, _36386_);
  and (_39234_, _36510_, _36509_);
  or (_36511_, _36497_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  or (_36512_, _36499_, _36400_);
  and (_39238_, _36512_, _36511_);
  or (_36513_, _36497_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  or (_36514_, _36499_, _36290_);
  and (_39241_, _36514_, _36513_);
  and (_36515_, _36460_, _36267_);
  or (_36516_, _36515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  not (_36517_, _36515_);
  or (_36518_, _36517_, _36312_);
  and (_39246_, _36518_, _36516_);
  or (_36519_, _36515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  or (_36520_, _36517_, _36328_);
  and (_39250_, _36520_, _36519_);
  or (_36521_, _36515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  or (_36522_, _36517_, _36343_);
  and (_39254_, _36522_, _36521_);
  or (_36523_, _36515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  or (_36524_, _36517_, _36358_);
  and (_39258_, _36524_, _36523_);
  or (_36525_, _36515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  or (_36526_, _36517_, _36372_);
  and (_39262_, _36526_, _36525_);
  or (_36527_, _36515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  or (_36528_, _36517_, _36386_);
  and (_39266_, _36528_, _36527_);
  or (_36529_, _36515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  or (_36530_, _36517_, _36400_);
  and (_39270_, _36530_, _36529_);
  or (_36531_, _36515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  or (_36532_, _36517_, _36290_);
  and (_39273_, _36532_, _36531_);
  and (_36533_, _36268_, _35989_);
  and (_36534_, _36533_, _36293_);
  or (_36535_, _36534_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  not (_36536_, _36534_);
  or (_36537_, _36536_, _36312_);
  and (_39281_, _36537_, _36535_);
  or (_36538_, _36534_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  or (_36539_, _36536_, _36328_);
  and (_39285_, _36539_, _36538_);
  or (_36540_, _36534_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  or (_36541_, _36536_, _36343_);
  and (_39289_, _36541_, _36540_);
  or (_36542_, _36534_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  or (_36543_, _36536_, _36358_);
  and (_39293_, _36543_, _36542_);
  or (_36544_, _36534_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  or (_36545_, _36536_, _36372_);
  and (_39297_, _36545_, _36544_);
  or (_36546_, _36534_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  or (_36547_, _36536_, _36386_);
  and (_39301_, _36547_, _36546_);
  or (_36548_, _36534_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  or (_36549_, _36536_, _36400_);
  and (_39305_, _36549_, _36548_);
  or (_36550_, _36534_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  or (_36551_, _36536_, _36290_);
  and (_39308_, _36551_, _36550_);
  and (_36552_, _36533_, _36404_);
  or (_36553_, _36552_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  not (_36554_, _36552_);
  or (_36555_, _36554_, _36312_);
  and (_39313_, _36555_, _36553_);
  or (_36556_, _36552_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  or (_36557_, _36554_, _36328_);
  and (_39317_, _36557_, _36556_);
  or (_36558_, _36552_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  or (_36559_, _36554_, _36343_);
  and (_39321_, _36559_, _36558_);
  or (_36560_, _36552_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  or (_36561_, _36554_, _36358_);
  and (_39325_, _36561_, _36560_);
  or (_36562_, _36552_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  or (_36563_, _36554_, _36372_);
  and (_39329_, _36563_, _36562_);
  or (_36564_, _36552_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  or (_36565_, _36554_, _36386_);
  and (_39333_, _36565_, _36564_);
  or (_36566_, _36552_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  or (_36567_, _36554_, _36400_);
  and (_39337_, _36567_, _36566_);
  or (_36568_, _36552_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  or (_36569_, _36554_, _36290_);
  and (_39340_, _36569_, _36568_);
  and (_36570_, _36533_, _36423_);
  or (_36571_, _36570_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  not (_36572_, _36570_);
  or (_36573_, _36572_, _36312_);
  and (_39345_, _36573_, _36571_);
  or (_36574_, _36570_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  or (_36575_, _36572_, _36328_);
  and (_39349_, _36575_, _36574_);
  or (_36576_, _36570_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  or (_36577_, _36572_, _36343_);
  and (_39353_, _36577_, _36576_);
  or (_36578_, _36570_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  or (_36579_, _36572_, _36358_);
  and (_39357_, _36579_, _36578_);
  or (_36580_, _36570_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  or (_36581_, _36572_, _36372_);
  and (_39361_, _36581_, _36580_);
  or (_36582_, _36570_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  or (_36583_, _36572_, _36386_);
  and (_39365_, _36583_, _36582_);
  or (_36584_, _36570_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  or (_36585_, _36572_, _36400_);
  and (_39369_, _36585_, _36584_);
  or (_36586_, _36570_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  or (_36587_, _36572_, _36290_);
  and (_39372_, _36587_, _36586_);
  and (_36588_, _36533_, _36267_);
  or (_36589_, _36588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  not (_36590_, _36588_);
  or (_36591_, _36590_, _36312_);
  and (_39377_, _36591_, _36589_);
  or (_36592_, _36588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  or (_36593_, _36590_, _36328_);
  and (_39381_, _36593_, _36592_);
  or (_36594_, _36588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  or (_36595_, _36590_, _36343_);
  and (_39385_, _36595_, _36594_);
  or (_36596_, _36588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  or (_36597_, _36590_, _36358_);
  and (_39389_, _36597_, _36596_);
  or (_36598_, _36588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  or (_36599_, _36590_, _36372_);
  and (_39393_, _36599_, _36598_);
  or (_36600_, _36588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  or (_36601_, _36590_, _36386_);
  and (_39397_, _36601_, _36600_);
  or (_36602_, _36588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  or (_36603_, _36590_, _36400_);
  and (_39401_, _36603_, _36602_);
  or (_36604_, _36588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  or (_36605_, _36590_, _36290_);
  and (_39404_, _36605_, _36604_);
  and (_36606_, _36293_, _36270_);
  or (_36607_, _36606_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  not (_36608_, _36606_);
  or (_36609_, _36608_, _36312_);
  and (_39410_, _36609_, _36607_);
  or (_36610_, _36606_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  or (_36611_, _36608_, _36328_);
  and (_39414_, _36611_, _36610_);
  or (_36612_, _36606_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  or (_36613_, _36608_, _36343_);
  and (_39418_, _36613_, _36612_);
  or (_36614_, _36606_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  or (_36615_, _36608_, _36358_);
  and (_39422_, _36615_, _36614_);
  or (_36616_, _36606_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  or (_36617_, _36608_, _36372_);
  and (_39426_, _36617_, _36616_);
  or (_36618_, _36606_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  or (_36619_, _36608_, _36386_);
  and (_39430_, _36619_, _36618_);
  or (_36620_, _36606_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  or (_36621_, _36608_, _36400_);
  and (_39434_, _36621_, _36620_);
  or (_36622_, _36606_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  or (_36623_, _36608_, _36290_);
  and (_39437_, _36623_, _36622_);
  and (_36624_, _36404_, _36270_);
  or (_36626_, _36624_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  not (_36627_, _36624_);
  or (_36628_, _36627_, _36312_);
  and (_39442_, _36628_, _36626_);
  or (_36629_, _36624_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  or (_36630_, _36627_, _36328_);
  and (_39446_, _36630_, _36629_);
  or (_36631_, _36624_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  or (_36632_, _36627_, _36343_);
  and (_39450_, _36632_, _36631_);
  or (_36634_, _36624_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  or (_36635_, _36627_, _36358_);
  and (_39454_, _36635_, _36634_);
  or (_36636_, _36624_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  or (_36637_, _36627_, _36372_);
  and (_39458_, _36637_, _36636_);
  or (_36638_, _36624_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  or (_36639_, _36627_, _36386_);
  and (_39462_, _36639_, _36638_);
  or (_36640_, _36624_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  or (_36642_, _36627_, _36400_);
  and (_39466_, _36642_, _36640_);
  or (_36643_, _36624_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  or (_36644_, _36627_, _36290_);
  and (_39469_, _36644_, _36643_);
  and (_36645_, _36423_, _36270_);
  or (_36646_, _36645_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  not (_36647_, _36645_);
  or (_36648_, _36647_, _36312_);
  and (_39474_, _36648_, _36646_);
  or (_36650_, _36645_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  or (_36651_, _36647_, _36328_);
  and (_39478_, _36651_, _36650_);
  or (_36652_, _36645_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  or (_36653_, _36647_, _36343_);
  and (_39482_, _36653_, _36652_);
  or (_36654_, _36645_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  or (_36655_, _36647_, _36358_);
  and (_39486_, _36655_, _36654_);
  or (_36656_, _36645_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  or (_36658_, _36647_, _36372_);
  and (_39490_, _36658_, _36656_);
  or (_36659_, _36645_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  or (_36660_, _36647_, _36386_);
  and (_39494_, _36660_, _36659_);
  or (_36661_, _36645_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  or (_36662_, _36647_, _36400_);
  and (_39498_, _36662_, _36661_);
  or (_36663_, _36645_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  or (_36664_, _36647_, _36290_);
  and (_39501_, _36664_, _36663_);
  or (_36666_, _36271_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  or (_36667_, _36312_, _36273_);
  and (_39506_, _36667_, _36666_);
  or (_36668_, _36271_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  or (_36669_, _36328_, _36273_);
  and (_39510_, _36669_, _36668_);
  or (_36670_, _36271_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  or (_36671_, _36343_, _36273_);
  and (_39514_, _36671_, _36670_);
  or (_36673_, _36271_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  or (_36674_, _36358_, _36273_);
  and (_39518_, _36674_, _36673_);
  or (_36675_, _36271_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  or (_36676_, _36372_, _36273_);
  and (_39522_, _36676_, _36675_);
  or (_36677_, _36271_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  or (_36678_, _36386_, _36273_);
  and (_39526_, _36678_, _36677_);
  or (_36679_, _36271_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  or (_36680_, _36400_, _36273_);
  and (_39530_, _36680_, _36679_);
  and (_36681_, _36066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  and (_36682_, _36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  or (_36683_, _36682_, _36681_);
  and (_36684_, _36683_, _36199_);
  and (_36685_, _36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  and (_36686_, _36066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  or (_36687_, _36686_, _36685_);
  and (_36688_, _36687_, _36218_);
  or (_36689_, _36688_, _36684_);
  or (_36690_, _36689_, _36212_);
  and (_36691_, _36066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  and (_36692_, _36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  or (_36693_, _36692_, _36691_);
  and (_36694_, _36693_, _36199_);
  and (_36695_, _36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  and (_36696_, _36066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  or (_36697_, _36696_, _36695_);
  and (_36698_, _36697_, _36218_);
  or (_36699_, _36698_, _36694_);
  or (_36700_, _36699_, _35985_);
  and (_36701_, _36700_, _36225_);
  and (_36702_, _36701_, _36690_);
  or (_36703_, _36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  or (_36704_, _36066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  and (_36705_, _36704_, _36703_);
  and (_36706_, _36705_, _36199_);
  or (_36707_, _36066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  or (_36708_, _36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  and (_36709_, _36708_, _36707_);
  and (_36710_, _36709_, _36218_);
  or (_36711_, _36710_, _36706_);
  or (_36712_, _36711_, _36212_);
  or (_36713_, _36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  or (_36714_, _36066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  and (_36715_, _36714_, _36713_);
  and (_36716_, _36715_, _36199_);
  or (_36717_, _36066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  or (_36718_, _36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  and (_36719_, _36718_, _36717_);
  and (_36720_, _36719_, _36218_);
  or (_36721_, _36720_, _36716_);
  or (_36722_, _36721_, _35985_);
  and (_36723_, _36722_, _36111_);
  and (_36724_, _36723_, _36712_);
  or (_36725_, _36724_, _36702_);
  or (_36726_, _36725_, _36211_);
  or (_36727_, _36262_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  and (_36728_, _36727_, _37580_);
  and (_00042_, _36728_, _36726_);
  and (_36729_, _36066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  and (_36730_, _36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  or (_36731_, _36730_, _36729_);
  and (_36732_, _36731_, _36199_);
  and (_36733_, _36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  and (_36734_, _36066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  or (_36735_, _36734_, _36733_);
  and (_36736_, _36735_, _36218_);
  or (_36737_, _36736_, _36732_);
  or (_36738_, _36737_, _36212_);
  and (_36739_, _36066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  and (_36740_, _36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  or (_36741_, _36740_, _36739_);
  and (_36742_, _36741_, _36199_);
  and (_36743_, _36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  and (_36744_, _36066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  or (_36745_, _36744_, _36743_);
  and (_36746_, _36745_, _36218_);
  or (_36747_, _36746_, _36742_);
  or (_36748_, _36747_, _35985_);
  and (_36749_, _36748_, _36225_);
  and (_36750_, _36749_, _36738_);
  or (_36751_, _36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  or (_36752_, _36066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  and (_36753_, _36752_, _36751_);
  and (_36754_, _36753_, _36199_);
  or (_36755_, _36066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  or (_36756_, _36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  and (_36757_, _36756_, _36755_);
  and (_36758_, _36757_, _36218_);
  or (_36759_, _36758_, _36754_);
  or (_36760_, _36759_, _36212_);
  or (_36761_, _36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  or (_36762_, _36066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  and (_36763_, _36762_, _36761_);
  and (_36764_, _36763_, _36199_);
  or (_36765_, _36066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  or (_36766_, _36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  and (_36767_, _36766_, _36765_);
  and (_36768_, _36767_, _36218_);
  or (_36769_, _36768_, _36764_);
  or (_36770_, _36769_, _35985_);
  and (_36771_, _36770_, _36111_);
  and (_36772_, _36771_, _36760_);
  or (_36773_, _36772_, _36750_);
  or (_36774_, _36773_, _36211_);
  or (_36775_, _36262_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  and (_36776_, _36775_, _37580_);
  and (_00044_, _36776_, _36774_);
  and (_36777_, _36066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  and (_36778_, _36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  or (_36779_, _36778_, _36777_);
  and (_36780_, _36779_, _36199_);
  and (_36781_, _36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  and (_36782_, _36066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  or (_36783_, _36782_, _36781_);
  and (_36784_, _36783_, _36218_);
  or (_36785_, _36784_, _36780_);
  or (_36786_, _36785_, _36212_);
  and (_36787_, _36066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  and (_36788_, _36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  or (_36789_, _36788_, _36787_);
  and (_36790_, _36789_, _36199_);
  and (_36791_, _36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  and (_36792_, _36066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  or (_36793_, _36792_, _36791_);
  and (_36794_, _36793_, _36218_);
  or (_36795_, _36794_, _36790_);
  or (_36796_, _36795_, _35985_);
  and (_36797_, _36796_, _36225_);
  and (_36798_, _36797_, _36786_);
  or (_36799_, _36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  or (_36800_, _36066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  and (_36801_, _36800_, _36799_);
  and (_36802_, _36801_, _36199_);
  or (_36803_, _36066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  or (_36804_, _36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  and (_36805_, _36804_, _36803_);
  and (_36806_, _36805_, _36218_);
  or (_36807_, _36806_, _36802_);
  or (_36808_, _36807_, _36212_);
  or (_36809_, _36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  or (_36810_, _36066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  and (_36811_, _36810_, _36809_);
  and (_36812_, _36811_, _36199_);
  or (_36813_, _36066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  or (_36814_, _36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  and (_36815_, _36814_, _36813_);
  and (_36816_, _36815_, _36218_);
  or (_36817_, _36816_, _36812_);
  or (_36818_, _36817_, _35985_);
  and (_36819_, _36818_, _36111_);
  and (_36820_, _36819_, _36808_);
  or (_36821_, _36820_, _36798_);
  or (_36822_, _36821_, _36211_);
  or (_36823_, _36262_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  and (_36824_, _36823_, _37580_);
  and (_00046_, _36824_, _36822_);
  and (_36825_, _36066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  and (_36826_, _36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  or (_36827_, _36826_, _36825_);
  and (_36828_, _36827_, _36199_);
  and (_36829_, _36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  and (_36830_, _36066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or (_36831_, _36830_, _36829_);
  and (_36832_, _36831_, _36218_);
  or (_36833_, _36832_, _36828_);
  or (_36834_, _36833_, _36212_);
  and (_36835_, _36066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  and (_36836_, _36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  or (_36837_, _36836_, _36835_);
  and (_36838_, _36837_, _36199_);
  and (_36839_, _36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  and (_36840_, _36066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or (_36841_, _36840_, _36839_);
  and (_36842_, _36841_, _36218_);
  or (_36843_, _36842_, _36838_);
  or (_36844_, _36843_, _35985_);
  and (_36845_, _36844_, _36225_);
  and (_36846_, _36845_, _36834_);
  or (_36847_, _36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  or (_36848_, _36066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  and (_36849_, _36848_, _36847_);
  and (_36850_, _36849_, _36199_);
  or (_36851_, _36066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  or (_36852_, _36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  and (_36853_, _36852_, _36851_);
  and (_36854_, _36853_, _36218_);
  or (_36855_, _36854_, _36850_);
  or (_36856_, _36855_, _36212_);
  or (_36857_, _36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  or (_36858_, _36066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  and (_36860_, _36858_, _36857_);
  and (_36862_, _36860_, _36199_);
  or (_36864_, _36066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  or (_36866_, _36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  and (_36868_, _36866_, _36864_);
  and (_36870_, _36868_, _36218_);
  or (_36872_, _36870_, _36862_);
  or (_36874_, _36872_, _35985_);
  and (_36876_, _36874_, _36111_);
  and (_36878_, _36876_, _36856_);
  or (_36880_, _36878_, _36846_);
  or (_36882_, _36880_, _36211_);
  or (_36884_, _36262_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  and (_36886_, _36884_, _37580_);
  and (_00048_, _36886_, _36882_);
  and (_36889_, _36066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  and (_36891_, _36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  or (_36893_, _36891_, _36889_);
  and (_36895_, _36893_, _36199_);
  and (_36897_, _36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  and (_36899_, _36066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  or (_36901_, _36899_, _36897_);
  and (_36903_, _36901_, _36218_);
  or (_36905_, _36903_, _36895_);
  or (_36907_, _36905_, _36212_);
  and (_36909_, _36066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  and (_36911_, _36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  or (_36913_, _36911_, _36909_);
  and (_36914_, _36913_, _36199_);
  and (_36915_, _36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  and (_36916_, _36066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  or (_36917_, _36916_, _36915_);
  and (_36918_, _36917_, _36218_);
  or (_36919_, _36918_, _36914_);
  or (_36920_, _36919_, _35985_);
  and (_36921_, _36920_, _36225_);
  and (_36922_, _36921_, _36907_);
  or (_36923_, _36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  or (_36924_, _36066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  and (_36925_, _36924_, _36923_);
  and (_36926_, _36925_, _36199_);
  or (_36927_, _36066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  or (_36928_, _36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  and (_36929_, _36928_, _36927_);
  and (_36930_, _36929_, _36218_);
  or (_36931_, _36930_, _36926_);
  or (_36932_, _36931_, _36212_);
  or (_36933_, _36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  or (_36934_, _36066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  and (_36935_, _36934_, _36933_);
  and (_36936_, _36935_, _36199_);
  or (_36937_, _36066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  or (_36938_, _36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  and (_36939_, _36938_, _36937_);
  and (_36940_, _36939_, _36218_);
  or (_36941_, _36940_, _36936_);
  or (_36942_, _36941_, _35985_);
  and (_36943_, _36942_, _36111_);
  and (_36944_, _36943_, _36932_);
  or (_36945_, _36944_, _36922_);
  or (_36946_, _36945_, _36211_);
  or (_36947_, _36262_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  and (_36948_, _36947_, _37580_);
  and (_00050_, _36948_, _36946_);
  and (_36949_, _36066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  and (_36950_, _36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  or (_36951_, _36950_, _36949_);
  and (_36952_, _36951_, _36199_);
  and (_36953_, _36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  and (_36954_, _36066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  or (_36955_, _36954_, _36953_);
  and (_36956_, _36955_, _36218_);
  or (_36957_, _36956_, _36952_);
  or (_36958_, _36957_, _36212_);
  and (_36959_, _36066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  and (_36960_, _36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  or (_36961_, _36960_, _36959_);
  and (_36962_, _36961_, _36199_);
  and (_36963_, _36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  and (_36964_, _36066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  or (_36965_, _36964_, _36963_);
  and (_36966_, _36965_, _36218_);
  or (_36967_, _36966_, _36962_);
  or (_36968_, _36967_, _35985_);
  and (_36969_, _36968_, _36225_);
  and (_36970_, _36969_, _36958_);
  or (_36971_, _36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  or (_36972_, _36066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  and (_36973_, _36972_, _36971_);
  and (_36974_, _36973_, _36199_);
  or (_36975_, _36066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  or (_36976_, _36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  and (_36977_, _36976_, _36975_);
  and (_36978_, _36977_, _36218_);
  or (_36979_, _36978_, _36974_);
  or (_36980_, _36979_, _36212_);
  or (_36981_, _36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  or (_36982_, _36066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  and (_36983_, _36982_, _36981_);
  and (_36984_, _36983_, _36199_);
  or (_36985_, _36066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  or (_36986_, _36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  and (_36987_, _36986_, _36985_);
  and (_36988_, _36987_, _36218_);
  or (_36989_, _36988_, _36984_);
  or (_36990_, _36989_, _35985_);
  and (_36991_, _36990_, _36111_);
  and (_36992_, _36991_, _36980_);
  or (_36993_, _36992_, _36970_);
  or (_36994_, _36993_, _36211_);
  or (_36995_, _36262_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  and (_36996_, _36995_, _37580_);
  and (_00052_, _36996_, _36994_);
  and (_36997_, _36066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  and (_36998_, _36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  or (_36999_, _36998_, _36997_);
  and (_37000_, _36999_, _36199_);
  and (_37001_, _36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  and (_37002_, _36066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  or (_37003_, _37002_, _37001_);
  and (_37004_, _37003_, _36218_);
  or (_37005_, _37004_, _37000_);
  or (_37006_, _37005_, _36212_);
  and (_37007_, _36066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  and (_37008_, _36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  or (_37009_, _37008_, _37007_);
  and (_37010_, _37009_, _36199_);
  and (_37011_, _36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  and (_37012_, _36066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  or (_37013_, _37012_, _37011_);
  and (_37014_, _37013_, _36218_);
  or (_37015_, _37014_, _37010_);
  or (_37016_, _37015_, _35985_);
  and (_37017_, _37016_, _36225_);
  and (_37018_, _37017_, _37006_);
  or (_37019_, _36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  or (_37020_, _36066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  and (_37021_, _37020_, _37019_);
  and (_37022_, _37021_, _36199_);
  or (_37023_, _36066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  or (_37024_, _36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  and (_37025_, _37024_, _37023_);
  and (_37026_, _37025_, _36218_);
  or (_37027_, _37026_, _37022_);
  or (_37028_, _37027_, _36212_);
  or (_37029_, _36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  or (_37030_, _36066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  and (_37031_, _37030_, _37029_);
  and (_37032_, _37031_, _36199_);
  or (_37033_, _36066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  or (_37034_, _36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  and (_37035_, _37034_, _37033_);
  and (_37036_, _37035_, _36218_);
  or (_37037_, _37036_, _37032_);
  or (_37038_, _37037_, _35985_);
  and (_37039_, _37038_, _36111_);
  and (_37040_, _37039_, _37028_);
  or (_37041_, _37040_, _37018_);
  or (_37042_, _37041_, _36211_);
  or (_37043_, _36262_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  and (_37044_, _37043_, _37580_);
  and (_00054_, _37044_, _37042_);
  or (_37045_, \oc8051_gm_cxrom_1.cell0.valid , word_in[7]);
  not (_37046_, \oc8051_gm_cxrom_1.cell0.valid );
  or (_37047_, _37046_, \oc8051_gm_cxrom_1.cell0.data [7]);
  nand (_37048_, _37047_, _37045_);
  nand (_37049_, _37048_, _37580_);
  or (_37050_, \oc8051_gm_cxrom_1.cell0.data [7], _37580_);
  and (_00062_, _37050_, _37049_);
  or (_37051_, word_in[0], \oc8051_gm_cxrom_1.cell0.valid );
  or (_37052_, \oc8051_gm_cxrom_1.cell0.data [0], _37046_);
  nand (_37053_, _37052_, _37051_);
  nand (_37054_, _37053_, _37580_);
  or (_37055_, \oc8051_gm_cxrom_1.cell0.data [0], _37580_);
  and (_00094_, _37055_, _37054_);
  or (_37056_, word_in[1], \oc8051_gm_cxrom_1.cell0.valid );
  or (_37057_, \oc8051_gm_cxrom_1.cell0.data [1], _37046_);
  nand (_37058_, _37057_, _37056_);
  nand (_37059_, _37058_, _37580_);
  or (_37060_, \oc8051_gm_cxrom_1.cell0.data [1], _37580_);
  and (_00096_, _37060_, _37059_);
  or (_37061_, word_in[2], \oc8051_gm_cxrom_1.cell0.valid );
  or (_37062_, \oc8051_gm_cxrom_1.cell0.data [2], _37046_);
  nand (_37063_, _37062_, _37061_);
  nand (_37064_, _37063_, _37580_);
  or (_37065_, \oc8051_gm_cxrom_1.cell0.data [2], _37580_);
  and (_00098_, _37065_, _37064_);
  or (_37066_, word_in[3], \oc8051_gm_cxrom_1.cell0.valid );
  or (_37067_, \oc8051_gm_cxrom_1.cell0.data [3], _37046_);
  nand (_37068_, _37067_, _37066_);
  nand (_37069_, _37068_, _37580_);
  or (_37070_, \oc8051_gm_cxrom_1.cell0.data [3], _37580_);
  and (_00100_, _37070_, _37069_);
  or (_37071_, word_in[4], \oc8051_gm_cxrom_1.cell0.valid );
  or (_37072_, \oc8051_gm_cxrom_1.cell0.data [4], _37046_);
  nand (_37073_, _37072_, _37071_);
  nand (_37074_, _37073_, _37580_);
  or (_37075_, \oc8051_gm_cxrom_1.cell0.data [4], _37580_);
  and (_00102_, _37075_, _37074_);
  or (_37076_, word_in[5], \oc8051_gm_cxrom_1.cell0.valid );
  or (_37077_, \oc8051_gm_cxrom_1.cell0.data [5], _37046_);
  nand (_37078_, _37077_, _37076_);
  nand (_37079_, _37078_, _37580_);
  or (_37080_, \oc8051_gm_cxrom_1.cell0.data [5], _37580_);
  and (_00104_, _37080_, _37079_);
  or (_37081_, word_in[6], \oc8051_gm_cxrom_1.cell0.valid );
  or (_37082_, \oc8051_gm_cxrom_1.cell0.data [6], _37046_);
  nand (_37083_, _37082_, _37081_);
  nand (_37084_, _37083_, _37580_);
  or (_37085_, \oc8051_gm_cxrom_1.cell0.data [6], _37580_);
  and (_00106_, _37085_, _37084_);
  or (_37086_, \oc8051_gm_cxrom_1.cell1.valid , word_in[15]);
  not (_37087_, \oc8051_gm_cxrom_1.cell1.valid );
  or (_37088_, _37087_, \oc8051_gm_cxrom_1.cell1.data [7]);
  nand (_37089_, _37088_, _37086_);
  nand (_37090_, _37089_, _37580_);
  or (_37091_, \oc8051_gm_cxrom_1.cell1.data [7], _37580_);
  and (_00113_, _37091_, _37090_);
  or (_37092_, word_in[8], \oc8051_gm_cxrom_1.cell1.valid );
  or (_37093_, \oc8051_gm_cxrom_1.cell1.data [0], _37087_);
  nand (_37094_, _37093_, _37092_);
  nand (_37095_, _37094_, _37580_);
  or (_37096_, \oc8051_gm_cxrom_1.cell1.data [0], _37580_);
  and (_00145_, _37096_, _37095_);
  or (_37097_, word_in[9], \oc8051_gm_cxrom_1.cell1.valid );
  or (_37098_, \oc8051_gm_cxrom_1.cell1.data [1], _37087_);
  nand (_37099_, _37098_, _37097_);
  nand (_37100_, _37099_, _37580_);
  or (_37101_, \oc8051_gm_cxrom_1.cell1.data [1], _37580_);
  and (_00147_, _37101_, _37100_);
  or (_37102_, word_in[10], \oc8051_gm_cxrom_1.cell1.valid );
  or (_37103_, \oc8051_gm_cxrom_1.cell1.data [2], _37087_);
  nand (_37104_, _37103_, _37102_);
  nand (_37105_, _37104_, _37580_);
  or (_37106_, \oc8051_gm_cxrom_1.cell1.data [2], _37580_);
  and (_00149_, _37106_, _37105_);
  or (_37107_, word_in[11], \oc8051_gm_cxrom_1.cell1.valid );
  or (_37108_, \oc8051_gm_cxrom_1.cell1.data [3], _37087_);
  nand (_37109_, _37108_, _37107_);
  nand (_37110_, _37109_, _37580_);
  or (_37111_, \oc8051_gm_cxrom_1.cell1.data [3], _37580_);
  and (_00151_, _37111_, _37110_);
  or (_37112_, word_in[12], \oc8051_gm_cxrom_1.cell1.valid );
  or (_37113_, \oc8051_gm_cxrom_1.cell1.data [4], _37087_);
  nand (_37114_, _37113_, _37112_);
  nand (_37115_, _37114_, _37580_);
  or (_37116_, \oc8051_gm_cxrom_1.cell1.data [4], _37580_);
  and (_00153_, _37116_, _37115_);
  or (_37117_, word_in[13], \oc8051_gm_cxrom_1.cell1.valid );
  or (_37118_, \oc8051_gm_cxrom_1.cell1.data [5], _37087_);
  nand (_37119_, _37118_, _37117_);
  nand (_37120_, _37119_, _37580_);
  or (_37121_, \oc8051_gm_cxrom_1.cell1.data [5], _37580_);
  and (_00155_, _37121_, _37120_);
  or (_37122_, word_in[14], \oc8051_gm_cxrom_1.cell1.valid );
  or (_37123_, \oc8051_gm_cxrom_1.cell1.data [6], _37087_);
  nand (_37124_, _37123_, _37122_);
  nand (_37125_, _37124_, _37580_);
  or (_37126_, \oc8051_gm_cxrom_1.cell1.data [6], _37580_);
  and (_00157_, _37126_, _37125_);
  or (_37127_, \oc8051_gm_cxrom_1.cell2.valid , word_in[23]);
  not (_37128_, \oc8051_gm_cxrom_1.cell2.valid );
  or (_37129_, _37128_, \oc8051_gm_cxrom_1.cell2.data [7]);
  nand (_37130_, _37129_, _37127_);
  nand (_37131_, _37130_, _37580_);
  or (_37132_, \oc8051_gm_cxrom_1.cell2.data [7], _37580_);
  and (_00165_, _37132_, _37131_);
  or (_37133_, word_in[16], \oc8051_gm_cxrom_1.cell2.valid );
  or (_37134_, \oc8051_gm_cxrom_1.cell2.data [0], _37128_);
  nand (_37135_, _37134_, _37133_);
  nand (_37138_, _37135_, _37580_);
  or (_37144_, \oc8051_gm_cxrom_1.cell2.data [0], _37580_);
  and (_00197_, _37144_, _37138_);
  or (_37155_, word_in[17], \oc8051_gm_cxrom_1.cell2.valid );
  or (_37161_, \oc8051_gm_cxrom_1.cell2.data [1], _37128_);
  nand (_37167_, _37161_, _37155_);
  nand (_37168_, _37167_, _37580_);
  or (_37169_, \oc8051_gm_cxrom_1.cell2.data [1], _37580_);
  and (_00199_, _37169_, _37168_);
  or (_37170_, word_in[18], \oc8051_gm_cxrom_1.cell2.valid );
  or (_37171_, \oc8051_gm_cxrom_1.cell2.data [2], _37128_);
  nand (_37172_, _37171_, _37170_);
  nand (_37173_, _37172_, _37580_);
  or (_37174_, \oc8051_gm_cxrom_1.cell2.data [2], _37580_);
  and (_00201_, _37174_, _37173_);
  or (_37175_, word_in[19], \oc8051_gm_cxrom_1.cell2.valid );
  or (_37176_, \oc8051_gm_cxrom_1.cell2.data [3], _37128_);
  nand (_37177_, _37176_, _37175_);
  nand (_37178_, _37177_, _37580_);
  or (_37179_, \oc8051_gm_cxrom_1.cell2.data [3], _37580_);
  and (_00203_, _37179_, _37178_);
  or (_37180_, word_in[20], \oc8051_gm_cxrom_1.cell2.valid );
  or (_37181_, \oc8051_gm_cxrom_1.cell2.data [4], _37128_);
  nand (_37182_, _37181_, _37180_);
  nand (_37183_, _37182_, _37580_);
  or (_37184_, \oc8051_gm_cxrom_1.cell2.data [4], _37580_);
  and (_00205_, _37184_, _37183_);
  or (_37185_, word_in[21], \oc8051_gm_cxrom_1.cell2.valid );
  or (_37186_, \oc8051_gm_cxrom_1.cell2.data [5], _37128_);
  nand (_37187_, _37186_, _37185_);
  nand (_37188_, _37187_, _37580_);
  or (_37189_, \oc8051_gm_cxrom_1.cell2.data [5], _37580_);
  and (_00207_, _37189_, _37188_);
  or (_37190_, word_in[22], \oc8051_gm_cxrom_1.cell2.valid );
  or (_37191_, \oc8051_gm_cxrom_1.cell2.data [6], _37128_);
  nand (_37192_, _37191_, _37190_);
  nand (_37193_, _37192_, _37580_);
  or (_37194_, \oc8051_gm_cxrom_1.cell2.data [6], _37580_);
  and (_00209_, _37194_, _37193_);
  or (_37195_, \oc8051_gm_cxrom_1.cell3.valid , word_in[31]);
  not (_37196_, \oc8051_gm_cxrom_1.cell3.valid );
  or (_37197_, _37196_, \oc8051_gm_cxrom_1.cell3.data [7]);
  nand (_37198_, _37197_, _37195_);
  nand (_37202_, _37198_, _37580_);
  or (_37205_, \oc8051_gm_cxrom_1.cell3.data [7], _37580_);
  and (_00217_, _37205_, _37202_);
  or (_37209_, word_in[24], \oc8051_gm_cxrom_1.cell3.valid );
  or (_37210_, \oc8051_gm_cxrom_1.cell3.data [0], _37196_);
  nand (_37212_, _37210_, _37209_);
  nand (_37218_, _37212_, _37580_);
  or (_37221_, \oc8051_gm_cxrom_1.cell3.data [0], _37580_);
  and (_00249_, _37221_, _37218_);
  or (_37222_, word_in[25], \oc8051_gm_cxrom_1.cell3.valid );
  or (_37225_, \oc8051_gm_cxrom_1.cell3.data [1], _37196_);
  nand (_37231_, _37225_, _37222_);
  nand (_37233_, _37231_, _37580_);
  or (_37234_, \oc8051_gm_cxrom_1.cell3.data [1], _37580_);
  and (_00251_, _37234_, _37233_);
  or (_37241_, word_in[26], \oc8051_gm_cxrom_1.cell3.valid );
  or (_37244_, \oc8051_gm_cxrom_1.cell3.data [2], _37196_);
  nand (_37245_, _37244_, _37241_);
  nand (_37246_, _37245_, _37580_);
  or (_37249_, \oc8051_gm_cxrom_1.cell3.data [2], _37580_);
  and (_00253_, _37249_, _37246_);
  or (_37256_, word_in[27], \oc8051_gm_cxrom_1.cell3.valid );
  or (_37257_, \oc8051_gm_cxrom_1.cell3.data [3], _37196_);
  nand (_37260_, _37257_, _37256_);
  nand (_37266_, _37260_, _37580_);
  or (_37268_, \oc8051_gm_cxrom_1.cell3.data [3], _37580_);
  and (_00255_, _37268_, _37266_);
  or (_37270_, word_in[28], \oc8051_gm_cxrom_1.cell3.valid );
  or (_37276_, \oc8051_gm_cxrom_1.cell3.data [4], _37196_);
  nand (_37279_, _37276_, _37270_);
  nand (_37280_, _37279_, _37580_);
  or (_37282_, \oc8051_gm_cxrom_1.cell3.data [4], _37580_);
  and (_00257_, _37282_, _37280_);
  or (_37290_, word_in[29], \oc8051_gm_cxrom_1.cell3.valid );
  or (_37291_, \oc8051_gm_cxrom_1.cell3.data [5], _37196_);
  nand (_37292_, _37291_, _37290_);
  nand (_37295_, _37292_, _37580_);
  or (_37301_, \oc8051_gm_cxrom_1.cell3.data [5], _37580_);
  and (_00259_, _37301_, _37295_);
  or (_37303_, word_in[30], \oc8051_gm_cxrom_1.cell3.valid );
  or (_37306_, \oc8051_gm_cxrom_1.cell3.data [6], _37196_);
  nand (_37312_, _37306_, _37303_);
  nand (_37314_, _37312_, _37580_);
  or (_37315_, \oc8051_gm_cxrom_1.cell3.data [6], _37580_);
  and (_00261_, _37315_, _37314_);
  or (_37322_, \oc8051_gm_cxrom_1.cell4.valid , word_in[39]);
  not (_37325_, \oc8051_gm_cxrom_1.cell4.valid );
  or (_37326_, _37325_, \oc8051_gm_cxrom_1.cell4.data [7]);
  nand (_37328_, _37326_, _37322_);
  nand (_37334_, _37328_, _37580_);
  or (_37337_, \oc8051_gm_cxrom_1.cell4.data [7], _37580_);
  and (_00269_, _37337_, _37334_);
  or (_37338_, word_in[32], \oc8051_gm_cxrom_1.cell4.valid );
  or (_37343_, \oc8051_gm_cxrom_1.cell4.data [0], _37325_);
  nand (_37348_, _37343_, _37338_);
  nand (_37349_, _37348_, _37580_);
  or (_37350_, \oc8051_gm_cxrom_1.cell4.data [0], _37580_);
  and (_00302_, _37350_, _37349_);
  or (_37359_, word_in[33], \oc8051_gm_cxrom_1.cell4.valid );
  or (_37360_, \oc8051_gm_cxrom_1.cell4.data [1], _37325_);
  nand (_37361_, _37360_, _37359_);
  nand (_37365_, _37361_, _37580_);
  or (_37371_, \oc8051_gm_cxrom_1.cell4.data [1], _37580_);
  and (_00304_, _37371_, _37365_);
  or (_37372_, word_in[34], \oc8051_gm_cxrom_1.cell4.valid );
  or (_37376_, \oc8051_gm_cxrom_1.cell4.data [2], _37325_);
  nand (_37381_, _37376_, _37372_);
  nand (_37382_, _37381_, _37580_);
  or (_37383_, \oc8051_gm_cxrom_1.cell4.data [2], _37580_);
  and (_00306_, _37383_, _37382_);
  or (_37384_, word_in[35], \oc8051_gm_cxrom_1.cell4.valid );
  or (_37385_, \oc8051_gm_cxrom_1.cell4.data [3], _37325_);
  nand (_37386_, _37385_, _37384_);
  nand (_37387_, _37386_, _37580_);
  or (_37388_, \oc8051_gm_cxrom_1.cell4.data [3], _37580_);
  and (_00307_, _37388_, _37387_);
  or (_37389_, word_in[36], \oc8051_gm_cxrom_1.cell4.valid );
  or (_37390_, \oc8051_gm_cxrom_1.cell4.data [4], _37325_);
  nand (_37391_, _37390_, _37389_);
  nand (_37392_, _37391_, _37580_);
  or (_37393_, \oc8051_gm_cxrom_1.cell4.data [4], _37580_);
  and (_00309_, _37393_, _37392_);
  or (_37394_, word_in[37], \oc8051_gm_cxrom_1.cell4.valid );
  or (_37395_, \oc8051_gm_cxrom_1.cell4.data [5], _37325_);
  nand (_37396_, _37395_, _37394_);
  nand (_37397_, _37396_, _37580_);
  or (_37398_, \oc8051_gm_cxrom_1.cell4.data [5], _37580_);
  and (_00311_, _37398_, _37397_);
  or (_37399_, word_in[38], \oc8051_gm_cxrom_1.cell4.valid );
  or (_37400_, \oc8051_gm_cxrom_1.cell4.data [6], _37325_);
  nand (_37401_, _37400_, _37399_);
  nand (_37402_, _37401_, _37580_);
  or (_37403_, \oc8051_gm_cxrom_1.cell4.data [6], _37580_);
  and (_00313_, _37403_, _37402_);
  or (_37404_, \oc8051_gm_cxrom_1.cell5.valid , word_in[47]);
  not (_37405_, \oc8051_gm_cxrom_1.cell5.valid );
  or (_37406_, _37405_, \oc8051_gm_cxrom_1.cell5.data [7]);
  nand (_37407_, _37406_, _37404_);
  nand (_37408_, _37407_, _37580_);
  or (_37409_, \oc8051_gm_cxrom_1.cell5.data [7], _37580_);
  and (_00321_, _37409_, _37408_);
  or (_37410_, word_in[40], \oc8051_gm_cxrom_1.cell5.valid );
  or (_37411_, \oc8051_gm_cxrom_1.cell5.data [0], _37405_);
  nand (_37412_, _37411_, _37410_);
  nand (_37413_, _37412_, _37580_);
  or (_37414_, \oc8051_gm_cxrom_1.cell5.data [0], _37580_);
  and (_00354_, _37414_, _37413_);
  or (_37415_, word_in[41], \oc8051_gm_cxrom_1.cell5.valid );
  or (_37416_, \oc8051_gm_cxrom_1.cell5.data [1], _37405_);
  nand (_37417_, _37416_, _37415_);
  nand (_37418_, _37417_, _37580_);
  or (_37419_, \oc8051_gm_cxrom_1.cell5.data [1], _37580_);
  and (_00356_, _37419_, _37418_);
  or (_37420_, word_in[42], \oc8051_gm_cxrom_1.cell5.valid );
  or (_37421_, \oc8051_gm_cxrom_1.cell5.data [2], _37405_);
  nand (_37422_, _37421_, _37420_);
  nand (_37423_, _37422_, _37580_);
  or (_37424_, \oc8051_gm_cxrom_1.cell5.data [2], _37580_);
  and (_00358_, _37424_, _37423_);
  or (_37425_, word_in[43], \oc8051_gm_cxrom_1.cell5.valid );
  or (_37426_, \oc8051_gm_cxrom_1.cell5.data [3], _37405_);
  nand (_37427_, _37426_, _37425_);
  nand (_37428_, _37427_, _37580_);
  or (_37429_, \oc8051_gm_cxrom_1.cell5.data [3], _37580_);
  and (_00360_, _37429_, _37428_);
  or (_37430_, word_in[44], \oc8051_gm_cxrom_1.cell5.valid );
  or (_37431_, \oc8051_gm_cxrom_1.cell5.data [4], _37405_);
  nand (_37432_, _37431_, _37430_);
  nand (_37433_, _37432_, _37580_);
  or (_37434_, \oc8051_gm_cxrom_1.cell5.data [4], _37580_);
  and (_00362_, _37434_, _37433_);
  or (_37435_, word_in[45], \oc8051_gm_cxrom_1.cell5.valid );
  or (_37436_, \oc8051_gm_cxrom_1.cell5.data [5], _37405_);
  nand (_37437_, _37436_, _37435_);
  nand (_37438_, _37437_, _37580_);
  or (_37439_, \oc8051_gm_cxrom_1.cell5.data [5], _37580_);
  and (_00364_, _37439_, _37438_);
  or (_37440_, word_in[46], \oc8051_gm_cxrom_1.cell5.valid );
  or (_37441_, \oc8051_gm_cxrom_1.cell5.data [6], _37405_);
  nand (_37442_, _37441_, _37440_);
  nand (_37443_, _37442_, _37580_);
  or (_37444_, \oc8051_gm_cxrom_1.cell5.data [6], _37580_);
  and (_00365_, _37444_, _37443_);
  or (_37445_, \oc8051_gm_cxrom_1.cell6.valid , word_in[55]);
  not (_37446_, \oc8051_gm_cxrom_1.cell6.valid );
  or (_37447_, _37446_, \oc8051_gm_cxrom_1.cell6.data [7]);
  nand (_37448_, _37447_, _37445_);
  nand (_37449_, _37448_, _37580_);
  or (_37450_, \oc8051_gm_cxrom_1.cell6.data [7], _37580_);
  and (_00373_, _37450_, _37449_);
  or (_37451_, word_in[48], \oc8051_gm_cxrom_1.cell6.valid );
  or (_37452_, \oc8051_gm_cxrom_1.cell6.data [0], _37446_);
  nand (_37453_, _37452_, _37451_);
  nand (_37454_, _37453_, _37580_);
  or (_37455_, \oc8051_gm_cxrom_1.cell6.data [0], _37580_);
  and (_00406_, _37455_, _37454_);
  or (_37456_, word_in[49], \oc8051_gm_cxrom_1.cell6.valid );
  or (_37457_, \oc8051_gm_cxrom_1.cell6.data [1], _37446_);
  nand (_37458_, _37457_, _37456_);
  nand (_37459_, _37458_, _37580_);
  or (_37460_, \oc8051_gm_cxrom_1.cell6.data [1], _37580_);
  and (_00408_, _37460_, _37459_);
  or (_37461_, word_in[50], \oc8051_gm_cxrom_1.cell6.valid );
  or (_37462_, \oc8051_gm_cxrom_1.cell6.data [2], _37446_);
  nand (_37463_, _37462_, _37461_);
  nand (_37464_, _37463_, _37580_);
  or (_37465_, \oc8051_gm_cxrom_1.cell6.data [2], _37580_);
  and (_00410_, _37465_, _37464_);
  or (_37466_, word_in[51], \oc8051_gm_cxrom_1.cell6.valid );
  or (_37467_, \oc8051_gm_cxrom_1.cell6.data [3], _37446_);
  nand (_37468_, _37467_, _37466_);
  nand (_37469_, _37468_, _37580_);
  or (_37470_, \oc8051_gm_cxrom_1.cell6.data [3], _37580_);
  and (_00412_, _37470_, _37469_);
  or (_37471_, word_in[52], \oc8051_gm_cxrom_1.cell6.valid );
  or (_37472_, \oc8051_gm_cxrom_1.cell6.data [4], _37446_);
  nand (_37473_, _37472_, _37471_);
  nand (_37474_, _37473_, _37580_);
  or (_37475_, \oc8051_gm_cxrom_1.cell6.data [4], _37580_);
  and (_00414_, _37475_, _37474_);
  or (_37476_, word_in[53], \oc8051_gm_cxrom_1.cell6.valid );
  or (_37477_, \oc8051_gm_cxrom_1.cell6.data [5], _37446_);
  nand (_37478_, _37477_, _37476_);
  nand (_37479_, _37478_, _37580_);
  or (_37480_, \oc8051_gm_cxrom_1.cell6.data [5], _37580_);
  and (_00416_, _37480_, _37479_);
  or (_37481_, word_in[54], \oc8051_gm_cxrom_1.cell6.valid );
  or (_37482_, \oc8051_gm_cxrom_1.cell6.data [6], _37446_);
  nand (_37483_, _37482_, _37481_);
  nand (_37484_, _37483_, _37580_);
  or (_37485_, \oc8051_gm_cxrom_1.cell6.data [6], _37580_);
  and (_00418_, _37485_, _37484_);
  or (_37486_, \oc8051_gm_cxrom_1.cell7.valid , word_in[63]);
  not (_37487_, \oc8051_gm_cxrom_1.cell7.valid );
  or (_37488_, _37487_, \oc8051_gm_cxrom_1.cell7.data [7]);
  nand (_37489_, _37488_, _37486_);
  nand (_37490_, _37489_, _37580_);
  or (_37491_, \oc8051_gm_cxrom_1.cell7.data [7], _37580_);
  and (_00425_, _37491_, _37490_);
  or (_37493_, word_in[56], \oc8051_gm_cxrom_1.cell7.valid );
  or (_37494_, \oc8051_gm_cxrom_1.cell7.data [0], _37487_);
  nand (_37495_, _37494_, _37493_);
  nand (_37496_, _37495_, _37580_);
  or (_37497_, \oc8051_gm_cxrom_1.cell7.data [0], _37580_);
  and (_00458_, _37497_, _37496_);
  or (_37498_, word_in[57], \oc8051_gm_cxrom_1.cell7.valid );
  or (_37499_, \oc8051_gm_cxrom_1.cell7.data [1], _37487_);
  nand (_37500_, _37499_, _37498_);
  nand (_37501_, _37500_, _37580_);
  or (_37502_, \oc8051_gm_cxrom_1.cell7.data [1], _37580_);
  and (_00460_, _37502_, _37501_);
  or (_37503_, word_in[58], \oc8051_gm_cxrom_1.cell7.valid );
  or (_37504_, \oc8051_gm_cxrom_1.cell7.data [2], _37487_);
  nand (_37505_, _37504_, _37503_);
  nand (_37506_, _37505_, _37580_);
  or (_37507_, \oc8051_gm_cxrom_1.cell7.data [2], _37580_);
  and (_00462_, _37507_, _37506_);
  or (_37508_, word_in[59], \oc8051_gm_cxrom_1.cell7.valid );
  or (_37509_, \oc8051_gm_cxrom_1.cell7.data [3], _37487_);
  nand (_37510_, _37509_, _37508_);
  nand (_37511_, _37510_, _37580_);
  or (_37512_, \oc8051_gm_cxrom_1.cell7.data [3], _37580_);
  and (_00464_, _37512_, _37511_);
  or (_37513_, word_in[60], \oc8051_gm_cxrom_1.cell7.valid );
  or (_37514_, \oc8051_gm_cxrom_1.cell7.data [4], _37487_);
  nand (_37515_, _37514_, _37513_);
  nand (_37516_, _37515_, _37580_);
  or (_37517_, \oc8051_gm_cxrom_1.cell7.data [4], _37580_);
  and (_00466_, _37517_, _37516_);
  or (_37518_, word_in[61], \oc8051_gm_cxrom_1.cell7.valid );
  or (_37519_, \oc8051_gm_cxrom_1.cell7.data [5], _37487_);
  nand (_37520_, _37519_, _37518_);
  nand (_37521_, _37520_, _37580_);
  or (_37522_, \oc8051_gm_cxrom_1.cell7.data [5], _37580_);
  and (_00468_, _37522_, _37521_);
  or (_37523_, word_in[62], \oc8051_gm_cxrom_1.cell7.valid );
  or (_37524_, \oc8051_gm_cxrom_1.cell7.data [6], _37487_);
  nand (_37525_, _37524_, _37523_);
  nand (_37526_, _37525_, _37580_);
  or (_37527_, \oc8051_gm_cxrom_1.cell7.data [6], _37580_);
  and (_00470_, _37527_, _37526_);
  or (_37529_, \oc8051_gm_cxrom_1.cell8.valid , word_in[71]);
  not (_37530_, \oc8051_gm_cxrom_1.cell8.valid );
  or (_37531_, _37530_, \oc8051_gm_cxrom_1.cell8.data [7]);
  nand (_37532_, _37531_, _37529_);
  nand (_37533_, _37532_, _37580_);
  or (_37534_, \oc8051_gm_cxrom_1.cell8.data [7], _37580_);
  and (_00477_, _37534_, _37533_);
  or (_37535_, word_in[64], \oc8051_gm_cxrom_1.cell8.valid );
  or (_37536_, \oc8051_gm_cxrom_1.cell8.data [0], _37530_);
  nand (_37537_, _37536_, _37535_);
  nand (_37538_, _37537_, _37580_);
  or (_37539_, \oc8051_gm_cxrom_1.cell8.data [0], _37580_);
  and (_00510_, _37539_, _37538_);
  or (_37540_, word_in[65], \oc8051_gm_cxrom_1.cell8.valid );
  or (_37541_, \oc8051_gm_cxrom_1.cell8.data [1], _37530_);
  nand (_37542_, _37541_, _37540_);
  nand (_37543_, _37542_, _37580_);
  or (_37544_, \oc8051_gm_cxrom_1.cell8.data [1], _37580_);
  and (_00512_, _37544_, _37543_);
  or (_37545_, word_in[66], \oc8051_gm_cxrom_1.cell8.valid );
  or (_37546_, \oc8051_gm_cxrom_1.cell8.data [2], _37530_);
  nand (_37548_, _37546_, _37545_);
  nand (_37550_, _37548_, _37580_);
  or (_37552_, \oc8051_gm_cxrom_1.cell8.data [2], _37580_);
  and (_00514_, _37552_, _37550_);
  or (_37553_, word_in[67], \oc8051_gm_cxrom_1.cell8.valid );
  or (_37554_, \oc8051_gm_cxrom_1.cell8.data [3], _37530_);
  nand (_37555_, _37554_, _37553_);
  nand (_37556_, _37555_, _37580_);
  or (_37557_, \oc8051_gm_cxrom_1.cell8.data [3], _37580_);
  and (_00516_, _37557_, _37556_);
  or (_37558_, word_in[68], \oc8051_gm_cxrom_1.cell8.valid );
  or (_37559_, \oc8051_gm_cxrom_1.cell8.data [4], _37530_);
  nand (_37560_, _37559_, _37558_);
  nand (_37561_, _37560_, _37580_);
  or (_37562_, \oc8051_gm_cxrom_1.cell8.data [4], _37580_);
  and (_00518_, _37562_, _37561_);
  or (_37563_, word_in[69], \oc8051_gm_cxrom_1.cell8.valid );
  or (_37564_, \oc8051_gm_cxrom_1.cell8.data [5], _37530_);
  nand (_37565_, _37564_, _37563_);
  nand (_37566_, _37565_, _37580_);
  or (_37567_, \oc8051_gm_cxrom_1.cell8.data [5], _37580_);
  and (_00520_, _37567_, _37566_);
  or (_37568_, word_in[70], \oc8051_gm_cxrom_1.cell8.valid );
  or (_37569_, \oc8051_gm_cxrom_1.cell8.data [6], _37530_);
  nand (_37570_, _37569_, _37568_);
  nand (_37572_, _37570_, _37580_);
  or (_37574_, \oc8051_gm_cxrom_1.cell8.data [6], _37580_);
  and (_00522_, _37574_, _37572_);
  or (_37577_, \oc8051_gm_cxrom_1.cell9.valid , word_in[79]);
  not (_37579_, \oc8051_gm_cxrom_1.cell9.valid );
  or (_37581_, _37579_, \oc8051_gm_cxrom_1.cell9.data [7]);
  nand (_37583_, _37581_, _37577_);
  nand (_37585_, _37583_, _37580_);
  or (_37587_, \oc8051_gm_cxrom_1.cell9.data [7], _37580_);
  and (_00530_, _37587_, _37585_);
  or (_37589_, word_in[72], \oc8051_gm_cxrom_1.cell9.valid );
  or (_37590_, \oc8051_gm_cxrom_1.cell9.data [0], _37579_);
  nand (_37591_, _37590_, _37589_);
  nand (_37592_, _37591_, _37580_);
  or (_37593_, \oc8051_gm_cxrom_1.cell9.data [0], _37580_);
  and (_00562_, _37593_, _37592_);
  or (_37594_, word_in[73], \oc8051_gm_cxrom_1.cell9.valid );
  or (_37595_, \oc8051_gm_cxrom_1.cell9.data [1], _37579_);
  nand (_37596_, _37595_, _37594_);
  nand (_37597_, _37596_, _37580_);
  or (_37598_, \oc8051_gm_cxrom_1.cell9.data [1], _37580_);
  and (_00564_, _37598_, _37597_);
  or (_37599_, word_in[74], \oc8051_gm_cxrom_1.cell9.valid );
  or (_37600_, \oc8051_gm_cxrom_1.cell9.data [2], _37579_);
  nand (_37601_, _37600_, _37599_);
  nand (_37602_, _37601_, _37580_);
  or (_37603_, \oc8051_gm_cxrom_1.cell9.data [2], _37580_);
  and (_00565_, _37603_, _37602_);
  or (_37604_, word_in[75], \oc8051_gm_cxrom_1.cell9.valid );
  or (_37605_, \oc8051_gm_cxrom_1.cell9.data [3], _37579_);
  nand (_37606_, _37605_, _37604_);
  nand (_37607_, _37606_, _37580_);
  or (_37608_, \oc8051_gm_cxrom_1.cell9.data [3], _37580_);
  and (_00567_, _37608_, _37607_);
  or (_37609_, word_in[76], \oc8051_gm_cxrom_1.cell9.valid );
  or (_37610_, \oc8051_gm_cxrom_1.cell9.data [4], _37579_);
  nand (_37611_, _37610_, _37609_);
  nand (_37612_, _37611_, _37580_);
  or (_37613_, \oc8051_gm_cxrom_1.cell9.data [4], _37580_);
  and (_00569_, _37613_, _37612_);
  or (_37614_, word_in[77], \oc8051_gm_cxrom_1.cell9.valid );
  or (_37615_, \oc8051_gm_cxrom_1.cell9.data [5], _37579_);
  nand (_37616_, _37615_, _37614_);
  nand (_37617_, _37616_, _37580_);
  or (_37618_, \oc8051_gm_cxrom_1.cell9.data [5], _37580_);
  and (_00571_, _37618_, _37617_);
  or (_37619_, word_in[78], \oc8051_gm_cxrom_1.cell9.valid );
  or (_37620_, \oc8051_gm_cxrom_1.cell9.data [6], _37579_);
  nand (_37621_, _37620_, _37619_);
  nand (_37622_, _37621_, _37580_);
  or (_37623_, \oc8051_gm_cxrom_1.cell9.data [6], _37580_);
  and (_00573_, _37623_, _37622_);
  or (_37624_, \oc8051_gm_cxrom_1.cell10.valid , word_in[87]);
  not (_37625_, \oc8051_gm_cxrom_1.cell10.valid );
  or (_37626_, _37625_, \oc8051_gm_cxrom_1.cell10.data [7]);
  nand (_37627_, _37626_, _37624_);
  nand (_37628_, _37627_, _37580_);
  or (_37629_, \oc8051_gm_cxrom_1.cell10.data [7], _37580_);
  and (_00581_, _37629_, _37628_);
  or (_37630_, word_in[80], \oc8051_gm_cxrom_1.cell10.valid );
  or (_37631_, \oc8051_gm_cxrom_1.cell10.data [0], _37625_);
  nand (_37632_, _37631_, _37630_);
  nand (_37633_, _37632_, _37580_);
  or (_37634_, \oc8051_gm_cxrom_1.cell10.data [0], _37580_);
  and (_00613_, _37634_, _37633_);
  or (_37635_, word_in[81], \oc8051_gm_cxrom_1.cell10.valid );
  or (_37636_, \oc8051_gm_cxrom_1.cell10.data [1], _37625_);
  nand (_37637_, _37636_, _37635_);
  nand (_37638_, _37637_, _37580_);
  or (_37639_, \oc8051_gm_cxrom_1.cell10.data [1], _37580_);
  and (_00615_, _37639_, _37638_);
  or (_37640_, word_in[82], \oc8051_gm_cxrom_1.cell10.valid );
  or (_37641_, \oc8051_gm_cxrom_1.cell10.data [2], _37625_);
  nand (_37642_, _37641_, _37640_);
  nand (_37643_, _37642_, _37580_);
  or (_37644_, \oc8051_gm_cxrom_1.cell10.data [2], _37580_);
  and (_00617_, _37644_, _37643_);
  or (_37645_, word_in[83], \oc8051_gm_cxrom_1.cell10.valid );
  or (_37646_, \oc8051_gm_cxrom_1.cell10.data [3], _37625_);
  nand (_37647_, _37646_, _37645_);
  nand (_37648_, _37647_, _37580_);
  or (_37649_, \oc8051_gm_cxrom_1.cell10.data [3], _37580_);
  and (_00619_, _37649_, _37648_);
  or (_37650_, word_in[84], \oc8051_gm_cxrom_1.cell10.valid );
  or (_37651_, \oc8051_gm_cxrom_1.cell10.data [4], _37625_);
  nand (_37652_, _37651_, _37650_);
  nand (_37653_, _37652_, _37580_);
  or (_37654_, \oc8051_gm_cxrom_1.cell10.data [4], _37580_);
  and (_00621_, _37654_, _37653_);
  or (_37655_, word_in[85], \oc8051_gm_cxrom_1.cell10.valid );
  or (_37656_, \oc8051_gm_cxrom_1.cell10.data [5], _37625_);
  nand (_37657_, _37656_, _37655_);
  nand (_37658_, _37657_, _37580_);
  or (_37659_, \oc8051_gm_cxrom_1.cell10.data [5], _37580_);
  and (_00623_, _37659_, _37658_);
  or (_37660_, word_in[86], \oc8051_gm_cxrom_1.cell10.valid );
  or (_37661_, \oc8051_gm_cxrom_1.cell10.data [6], _37625_);
  nand (_37662_, _37661_, _37660_);
  nand (_37663_, _37662_, _37580_);
  or (_37664_, \oc8051_gm_cxrom_1.cell10.data [6], _37580_);
  and (_00625_, _37664_, _37663_);
  or (_37665_, \oc8051_gm_cxrom_1.cell11.valid , word_in[95]);
  not (_37666_, \oc8051_gm_cxrom_1.cell11.valid );
  or (_37667_, _37666_, \oc8051_gm_cxrom_1.cell11.data [7]);
  nand (_37668_, _37667_, _37665_);
  nand (_37669_, _37668_, _37580_);
  or (_37670_, \oc8051_gm_cxrom_1.cell11.data [7], _37580_);
  and (_00633_, _37670_, _37669_);
  or (_37671_, word_in[88], \oc8051_gm_cxrom_1.cell11.valid );
  or (_37672_, \oc8051_gm_cxrom_1.cell11.data [0], _37666_);
  nand (_37673_, _37672_, _37671_);
  nand (_37674_, _37673_, _37580_);
  or (_37675_, \oc8051_gm_cxrom_1.cell11.data [0], _37580_);
  and (_00665_, _37675_, _37674_);
  or (_37676_, word_in[89], \oc8051_gm_cxrom_1.cell11.valid );
  or (_37677_, \oc8051_gm_cxrom_1.cell11.data [1], _37666_);
  nand (_37678_, _37677_, _37676_);
  nand (_37679_, _37678_, _37580_);
  or (_37680_, \oc8051_gm_cxrom_1.cell11.data [1], _37580_);
  and (_00667_, _37680_, _37679_);
  or (_37681_, word_in[90], \oc8051_gm_cxrom_1.cell11.valid );
  or (_37682_, \oc8051_gm_cxrom_1.cell11.data [2], _37666_);
  nand (_37683_, _37682_, _37681_);
  nand (_37684_, _37683_, _37580_);
  or (_37685_, \oc8051_gm_cxrom_1.cell11.data [2], _37580_);
  and (_00669_, _37685_, _37684_);
  or (_37686_, word_in[91], \oc8051_gm_cxrom_1.cell11.valid );
  or (_37687_, \oc8051_gm_cxrom_1.cell11.data [3], _37666_);
  nand (_37688_, _37687_, _37686_);
  nand (_37689_, _37688_, _37580_);
  or (_37690_, \oc8051_gm_cxrom_1.cell11.data [3], _37580_);
  and (_00671_, _37690_, _37689_);
  or (_37691_, word_in[92], \oc8051_gm_cxrom_1.cell11.valid );
  or (_37692_, \oc8051_gm_cxrom_1.cell11.data [4], _37666_);
  nand (_37693_, _37692_, _37691_);
  nand (_37694_, _37693_, _37580_);
  or (_37695_, \oc8051_gm_cxrom_1.cell11.data [4], _37580_);
  and (_00673_, _37695_, _37694_);
  or (_37696_, word_in[93], \oc8051_gm_cxrom_1.cell11.valid );
  or (_37697_, \oc8051_gm_cxrom_1.cell11.data [5], _37666_);
  nand (_37698_, _37697_, _37696_);
  nand (_37699_, _37698_, _37580_);
  or (_37700_, \oc8051_gm_cxrom_1.cell11.data [5], _37580_);
  and (_00675_, _37700_, _37699_);
  or (_37701_, word_in[94], \oc8051_gm_cxrom_1.cell11.valid );
  or (_37702_, \oc8051_gm_cxrom_1.cell11.data [6], _37666_);
  nand (_37703_, _37702_, _37701_);
  nand (_37704_, _37703_, _37580_);
  or (_37705_, \oc8051_gm_cxrom_1.cell11.data [6], _37580_);
  and (_00677_, _37705_, _37704_);
  or (_37706_, \oc8051_gm_cxrom_1.cell12.valid , word_in[103]);
  not (_37707_, \oc8051_gm_cxrom_1.cell12.valid );
  or (_37708_, _37707_, \oc8051_gm_cxrom_1.cell12.data [7]);
  nand (_37709_, _37708_, _37706_);
  nand (_37710_, _37709_, _37580_);
  or (_37711_, \oc8051_gm_cxrom_1.cell12.data [7], _37580_);
  and (_00684_, _37711_, _37710_);
  or (_37712_, word_in[96], \oc8051_gm_cxrom_1.cell12.valid );
  or (_37713_, \oc8051_gm_cxrom_1.cell12.data [0], _37707_);
  nand (_37714_, _37713_, _37712_);
  nand (_37715_, _37714_, _37580_);
  or (_37716_, \oc8051_gm_cxrom_1.cell12.data [0], _37580_);
  and (_00716_, _37716_, _37715_);
  or (_37717_, word_in[97], \oc8051_gm_cxrom_1.cell12.valid );
  or (_37718_, \oc8051_gm_cxrom_1.cell12.data [1], _37707_);
  nand (_37719_, _37718_, _37717_);
  nand (_37720_, _37719_, _37580_);
  or (_37721_, \oc8051_gm_cxrom_1.cell12.data [1], _37580_);
  and (_00718_, _37721_, _37720_);
  or (_37722_, word_in[98], \oc8051_gm_cxrom_1.cell12.valid );
  or (_37723_, \oc8051_gm_cxrom_1.cell12.data [2], _37707_);
  nand (_37724_, _37723_, _37722_);
  nand (_37725_, _37724_, _37580_);
  or (_37726_, \oc8051_gm_cxrom_1.cell12.data [2], _37580_);
  and (_00720_, _37726_, _37725_);
  or (_37727_, word_in[99], \oc8051_gm_cxrom_1.cell12.valid );
  or (_37728_, \oc8051_gm_cxrom_1.cell12.data [3], _37707_);
  nand (_37729_, _37728_, _37727_);
  nand (_37730_, _37729_, _37580_);
  or (_37731_, \oc8051_gm_cxrom_1.cell12.data [3], _37580_);
  and (_00722_, _37731_, _37730_);
  or (_37732_, word_in[100], \oc8051_gm_cxrom_1.cell12.valid );
  or (_37733_, \oc8051_gm_cxrom_1.cell12.data [4], _37707_);
  nand (_37734_, _37733_, _37732_);
  nand (_37735_, _37734_, _37580_);
  or (_37736_, \oc8051_gm_cxrom_1.cell12.data [4], _37580_);
  and (_00724_, _37736_, _37735_);
  or (_37737_, word_in[101], \oc8051_gm_cxrom_1.cell12.valid );
  or (_37738_, \oc8051_gm_cxrom_1.cell12.data [5], _37707_);
  nand (_37739_, _37738_, _37737_);
  nand (_37740_, _37739_, _37580_);
  or (_37741_, \oc8051_gm_cxrom_1.cell12.data [5], _37580_);
  and (_00726_, _37741_, _37740_);
  or (_37742_, word_in[102], \oc8051_gm_cxrom_1.cell12.valid );
  or (_37743_, \oc8051_gm_cxrom_1.cell12.data [6], _37707_);
  nand (_37744_, _37743_, _37742_);
  nand (_37745_, _37744_, _37580_);
  or (_37746_, \oc8051_gm_cxrom_1.cell12.data [6], _37580_);
  and (_00728_, _37746_, _37745_);
  or (_37747_, \oc8051_gm_cxrom_1.cell13.valid , word_in[111]);
  not (_37748_, \oc8051_gm_cxrom_1.cell13.valid );
  or (_37749_, _37748_, \oc8051_gm_cxrom_1.cell13.data [7]);
  nand (_37750_, _37749_, _37747_);
  nand (_37751_, _37750_, _37580_);
  or (_37752_, \oc8051_gm_cxrom_1.cell13.data [7], _37580_);
  and (_00736_, _37752_, _37751_);
  or (_37753_, word_in[104], \oc8051_gm_cxrom_1.cell13.valid );
  or (_37754_, \oc8051_gm_cxrom_1.cell13.data [0], _37748_);
  nand (_37755_, _37754_, _37753_);
  nand (_37756_, _37755_, _37580_);
  or (_37757_, \oc8051_gm_cxrom_1.cell13.data [0], _37580_);
  and (_00768_, _37757_, _37756_);
  or (_37758_, word_in[105], \oc8051_gm_cxrom_1.cell13.valid );
  or (_37759_, \oc8051_gm_cxrom_1.cell13.data [1], _37748_);
  nand (_37760_, _37759_, _37758_);
  nand (_37761_, _37760_, _37580_);
  or (_37762_, \oc8051_gm_cxrom_1.cell13.data [1], _37580_);
  and (_00770_, _37762_, _37761_);
  or (_37763_, word_in[106], \oc8051_gm_cxrom_1.cell13.valid );
  or (_37764_, \oc8051_gm_cxrom_1.cell13.data [2], _37748_);
  nand (_37765_, _37764_, _37763_);
  nand (_37766_, _37765_, _37580_);
  or (_37767_, \oc8051_gm_cxrom_1.cell13.data [2], _37580_);
  and (_00772_, _37767_, _37766_);
  or (_37768_, word_in[107], \oc8051_gm_cxrom_1.cell13.valid );
  or (_37769_, \oc8051_gm_cxrom_1.cell13.data [3], _37748_);
  nand (_37770_, _37769_, _37768_);
  nand (_37771_, _37770_, _37580_);
  or (_37772_, \oc8051_gm_cxrom_1.cell13.data [3], _37580_);
  and (_00774_, _37772_, _37771_);
  or (_37773_, word_in[108], \oc8051_gm_cxrom_1.cell13.valid );
  or (_37774_, \oc8051_gm_cxrom_1.cell13.data [4], _37748_);
  nand (_37775_, _37774_, _37773_);
  nand (_37776_, _37775_, _37580_);
  or (_37777_, \oc8051_gm_cxrom_1.cell13.data [4], _37580_);
  and (_00776_, _37777_, _37776_);
  or (_37778_, word_in[109], \oc8051_gm_cxrom_1.cell13.valid );
  or (_37779_, \oc8051_gm_cxrom_1.cell13.data [5], _37748_);
  nand (_37780_, _37779_, _37778_);
  nand (_37781_, _37780_, _37580_);
  or (_37782_, \oc8051_gm_cxrom_1.cell13.data [5], _37580_);
  and (_00778_, _37782_, _37781_);
  or (_37783_, word_in[110], \oc8051_gm_cxrom_1.cell13.valid );
  or (_37784_, \oc8051_gm_cxrom_1.cell13.data [6], _37748_);
  nand (_37785_, _37784_, _37783_);
  nand (_37786_, _37785_, _37580_);
  or (_37787_, \oc8051_gm_cxrom_1.cell13.data [6], _37580_);
  and (_00780_, _37787_, _37786_);
  or (_37788_, \oc8051_gm_cxrom_1.cell14.valid , word_in[119]);
  not (_37789_, \oc8051_gm_cxrom_1.cell14.valid );
  or (_37790_, _37789_, \oc8051_gm_cxrom_1.cell14.data [7]);
  nand (_37791_, _37790_, _37788_);
  nand (_37792_, _37791_, _37580_);
  or (_37793_, \oc8051_gm_cxrom_1.cell14.data [7], _37580_);
  and (_00787_, _37793_, _37792_);
  or (_37794_, word_in[112], \oc8051_gm_cxrom_1.cell14.valid );
  or (_37795_, \oc8051_gm_cxrom_1.cell14.data [0], _37789_);
  nand (_37796_, _37795_, _37794_);
  nand (_37797_, _37796_, _37580_);
  or (_37798_, \oc8051_gm_cxrom_1.cell14.data [0], _37580_);
  and (_00819_, _37798_, _37797_);
  or (_37799_, word_in[113], \oc8051_gm_cxrom_1.cell14.valid );
  or (_37800_, \oc8051_gm_cxrom_1.cell14.data [1], _37789_);
  nand (_37801_, _37800_, _37799_);
  nand (_37802_, _37801_, _37580_);
  or (_37803_, \oc8051_gm_cxrom_1.cell14.data [1], _37580_);
  and (_00821_, _37803_, _37802_);
  or (_37804_, word_in[114], \oc8051_gm_cxrom_1.cell14.valid );
  or (_37805_, \oc8051_gm_cxrom_1.cell14.data [2], _37789_);
  nand (_37806_, _37805_, _37804_);
  nand (_37807_, _37806_, _37580_);
  or (_37808_, \oc8051_gm_cxrom_1.cell14.data [2], _37580_);
  and (_00823_, _37808_, _37807_);
  or (_37809_, word_in[115], \oc8051_gm_cxrom_1.cell14.valid );
  or (_37810_, \oc8051_gm_cxrom_1.cell14.data [3], _37789_);
  nand (_37811_, _37810_, _37809_);
  nand (_37812_, _37811_, _37580_);
  or (_37813_, \oc8051_gm_cxrom_1.cell14.data [3], _37580_);
  and (_00825_, _37813_, _37812_);
  or (_37814_, word_in[116], \oc8051_gm_cxrom_1.cell14.valid );
  or (_37815_, \oc8051_gm_cxrom_1.cell14.data [4], _37789_);
  nand (_37816_, _37815_, _37814_);
  nand (_37817_, _37816_, _37580_);
  or (_37818_, \oc8051_gm_cxrom_1.cell14.data [4], _37580_);
  and (_00827_, _37818_, _37817_);
  or (_37819_, word_in[117], \oc8051_gm_cxrom_1.cell14.valid );
  or (_37820_, \oc8051_gm_cxrom_1.cell14.data [5], _37789_);
  nand (_37821_, _37820_, _37819_);
  nand (_37822_, _37821_, _37580_);
  or (_37823_, \oc8051_gm_cxrom_1.cell14.data [5], _37580_);
  and (_00829_, _37823_, _37822_);
  or (_37824_, word_in[118], \oc8051_gm_cxrom_1.cell14.valid );
  or (_37825_, \oc8051_gm_cxrom_1.cell14.data [6], _37789_);
  nand (_37826_, _37825_, _37824_);
  nand (_37827_, _37826_, _37580_);
  or (_37828_, \oc8051_gm_cxrom_1.cell14.data [6], _37580_);
  and (_00831_, _37828_, _37827_);
  or (_37829_, \oc8051_gm_cxrom_1.cell15.valid , word_in[127]);
  not (_37830_, \oc8051_gm_cxrom_1.cell15.valid );
  or (_37831_, _37830_, \oc8051_gm_cxrom_1.cell15.data [7]);
  nand (_37832_, _37831_, _37829_);
  nand (_37833_, _37832_, _37580_);
  or (_37834_, \oc8051_gm_cxrom_1.cell15.data [7], _37580_);
  and (_00839_, _37834_, _37833_);
  or (_37835_, word_in[120], \oc8051_gm_cxrom_1.cell15.valid );
  or (_37836_, \oc8051_gm_cxrom_1.cell15.data [0], _37830_);
  nand (_37837_, _37836_, _37835_);
  nand (_37838_, _37837_, _37580_);
  or (_37839_, \oc8051_gm_cxrom_1.cell15.data [0], _37580_);
  and (_00871_, _37839_, _37838_);
  or (_37840_, word_in[121], \oc8051_gm_cxrom_1.cell15.valid );
  or (_37841_, \oc8051_gm_cxrom_1.cell15.data [1], _37830_);
  nand (_37842_, _37841_, _37840_);
  nand (_37843_, _37842_, _37580_);
  or (_37844_, \oc8051_gm_cxrom_1.cell15.data [1], _37580_);
  and (_00873_, _37844_, _37843_);
  or (_37845_, word_in[122], \oc8051_gm_cxrom_1.cell15.valid );
  or (_37846_, \oc8051_gm_cxrom_1.cell15.data [2], _37830_);
  nand (_37847_, _37846_, _37845_);
  nand (_37848_, _37847_, _37580_);
  or (_37849_, \oc8051_gm_cxrom_1.cell15.data [2], _37580_);
  and (_00875_, _37849_, _37848_);
  or (_37850_, word_in[123], \oc8051_gm_cxrom_1.cell15.valid );
  or (_37851_, \oc8051_gm_cxrom_1.cell15.data [3], _37830_);
  nand (_37852_, _37851_, _37850_);
  nand (_37853_, _37852_, _37580_);
  or (_37854_, \oc8051_gm_cxrom_1.cell15.data [3], _37580_);
  and (_00877_, _37854_, _37853_);
  or (_37855_, word_in[124], \oc8051_gm_cxrom_1.cell15.valid );
  or (_37856_, \oc8051_gm_cxrom_1.cell15.data [4], _37830_);
  nand (_37857_, _37856_, _37855_);
  nand (_37858_, _37857_, _37580_);
  or (_37859_, \oc8051_gm_cxrom_1.cell15.data [4], _37580_);
  and (_00879_, _37859_, _37858_);
  or (_37860_, word_in[125], \oc8051_gm_cxrom_1.cell15.valid );
  or (_37861_, \oc8051_gm_cxrom_1.cell15.data [5], _37830_);
  nand (_37862_, _37861_, _37860_);
  nand (_37863_, _37862_, _37580_);
  or (_37864_, \oc8051_gm_cxrom_1.cell15.data [5], _37580_);
  and (_00881_, _37864_, _37863_);
  or (_37865_, word_in[126], \oc8051_gm_cxrom_1.cell15.valid );
  or (_37866_, \oc8051_gm_cxrom_1.cell15.data [6], _37830_);
  nand (_37867_, _37866_, _37865_);
  nand (_37868_, _37867_, _37580_);
  or (_37869_, \oc8051_gm_cxrom_1.cell15.data [6], _37580_);
  and (_00883_, _37869_, _37868_);
  nor (_00914_, _20214_, rst);
  nor (_00918_, _35848_, rst);
  nor (_37870_, _19284_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  and (_37871_, _18640_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_37872_, _18684_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor (_37873_, _37872_, _37871_);
  and (_37874_, _18727_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_37875_, _18771_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor (_37876_, _37875_, _37874_);
  and (_37877_, _37876_, _37873_);
  and (_37878_, _18825_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and (_37879_, _18836_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_37880_, _37879_, _37878_);
  and (_37881_, _37880_, _37877_);
  and (_37882_, _37881_, _19284_);
  nor (_37883_, _37882_, _37870_);
  nor (_37884_, _37883_, _35832_);
  nor (_37885_, _18553_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [7]);
  nor (_37886_, _37885_, _37884_);
  and (_00922_, _37886_, _37580_);
  nor (_01043_, _19702_, rst);
  nor (_01046_, _19462_, rst);
  nor (_01049_, _18935_, rst);
  nor (_01051_, _19186_, rst);
  and (_01054_, _19964_, _37580_);
  nor (_01057_, _20694_, rst);
  nor (_01060_, _20454_, rst);
  nor (_01063_, _36059_, rst);
  nor (_01066_, _36177_, rst);
  nor (_01069_, _35978_, rst);
  nor (_01072_, _36022_, rst);
  nor (_01075_, _36153_, rst);
  nor (_01078_, _35923_, rst);
  nor (_01081_, _36090_, rst);
  nor (_37887_, _19284_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  and (_37888_, _18640_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_37889_, _18684_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor (_37890_, _37889_, _37888_);
  and (_37891_, _18727_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_37892_, _18771_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_37893_, _37892_, _37891_);
  and (_37894_, _37893_, _37890_);
  and (_37895_, _18825_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and (_37896_, _18836_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_37897_, _37896_, _37895_);
  and (_37898_, _37897_, _37894_);
  and (_37899_, _37898_, _19284_);
  nor (_37900_, _37899_, _37887_);
  nor (_37901_, _37900_, _35832_);
  nor (_37902_, _18553_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [0]);
  nor (_37903_, _37902_, _37901_);
  and (_01084_, _37903_, _37580_);
  nor (_37904_, _19284_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  and (_37905_, _18727_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_37906_, _18771_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_37907_, _37906_, _37905_);
  and (_37908_, _18640_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_37909_, _18684_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nor (_37910_, _37909_, _37908_);
  and (_37911_, _18825_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and (_37912_, _18836_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_37913_, _37912_, _37911_);
  and (_37914_, _37913_, _37910_);
  and (_37915_, _37914_, _37907_);
  and (_37916_, _37915_, _19284_);
  nor (_37917_, _37916_, _37904_);
  nor (_37918_, _37917_, _35832_);
  nor (_37919_, _18553_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [1]);
  nor (_37920_, _37919_, _37918_);
  and (_01087_, _37920_, _37580_);
  nor (_37921_, _19284_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  and (_37922_, _18825_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and (_37923_, _18771_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_37924_, _37923_, _37922_);
  and (_37925_, _18640_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_37926_, _18684_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor (_37927_, _37926_, _37925_);
  and (_37928_, _18836_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  and (_37929_, _18727_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  nor (_37930_, _37929_, _37928_);
  and (_37931_, _37930_, _37927_);
  and (_37932_, _37931_, _37924_);
  and (_37933_, _37932_, _19284_);
  nor (_37934_, _37933_, _37921_);
  nor (_37935_, _37934_, _35832_);
  nor (_37936_, _18553_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [2]);
  nor (_37937_, _37936_, _37935_);
  and (_01090_, _37937_, _37580_);
  nor (_37938_, _19284_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  and (_37939_, _18640_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_37940_, _18684_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor (_37941_, _37940_, _37939_);
  and (_37942_, _18727_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_37943_, _18771_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_37944_, _37943_, _37942_);
  and (_37945_, _37944_, _37941_);
  and (_37946_, _18825_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and (_37947_, _18836_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_37948_, _37947_, _37946_);
  and (_37949_, _37948_, _37945_);
  and (_37950_, _37949_, _19284_);
  nor (_37951_, _37950_, _37938_);
  nor (_37952_, _37951_, _35832_);
  nor (_37953_, _18553_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [3]);
  nor (_37954_, _37953_, _37952_);
  and (_01093_, _37954_, _37580_);
  nor (_37955_, _19284_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  and (_37956_, _18836_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  and (_37957_, _18727_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  nor (_37958_, _37957_, _37956_);
  and (_37959_, _18640_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_37960_, _18684_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor (_37961_, _37960_, _37959_);
  and (_37962_, _18825_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and (_37963_, _18771_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_37964_, _37963_, _37962_);
  and (_37965_, _37964_, _37961_);
  and (_37966_, _37965_, _37958_);
  and (_37967_, _37966_, _19284_);
  nor (_37968_, _37967_, _37955_);
  nor (_37969_, _37968_, _35832_);
  nor (_37970_, _18553_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [4]);
  nor (_37971_, _37970_, _37969_);
  and (_01095_, _37971_, _37580_);
  nor (_37972_, _19284_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  and (_37973_, _18836_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  and (_37974_, _18727_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  nor (_37975_, _37974_, _37973_);
  and (_37976_, _18640_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_37977_, _18684_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor (_37978_, _37977_, _37976_);
  and (_37979_, _18825_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and (_37980_, _18771_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_37981_, _37980_, _37979_);
  and (_37982_, _37981_, _37978_);
  and (_37983_, _37982_, _37975_);
  and (_37984_, _37983_, _19284_);
  nor (_37985_, _37984_, _37972_);
  nor (_37986_, _37985_, _35832_);
  nor (_37987_, _18553_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [5]);
  nor (_37988_, _37987_, _37986_);
  and (_01098_, _37988_, _37580_);
  nor (_37989_, _19284_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  and (_37990_, _18836_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  and (_37991_, _18727_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  nor (_37992_, _37991_, _37990_);
  and (_37993_, _18640_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_37994_, _18684_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor (_37995_, _37994_, _37993_);
  and (_37996_, _18825_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and (_37997_, _18771_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor (_37998_, _37997_, _37996_);
  and (_37999_, _37998_, _37995_);
  and (_38000_, _37999_, _37992_);
  and (_38001_, _38000_, _19284_);
  nor (_38002_, _38001_, _37989_);
  nor (_38003_, _38002_, _35832_);
  nor (_38004_, _18553_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [6]);
  nor (_38005_, _38004_, _38003_);
  and (_01101_, _38005_, _37580_);
  not (_38006_, _35889_);
  and (_38007_, _36108_, _38006_);
  nor (_38008_, _36028_, _36158_);
  and (_38009_, _38008_, _35945_);
  and (_38010_, _38009_, _38007_);
  and (_38011_, _36158_, _35946_);
  and (_38012_, _38011_, _38007_);
  and (_38013_, _38012_, _36027_);
  nor (_38014_, _38013_, _38010_);
  nor (_38015_, _36158_, _35945_);
  and (_38016_, _38015_, _38007_);
  and (_38017_, _38016_, _36027_);
  and (_38018_, _36108_, _35945_);
  and (_38019_, _36158_, _38006_);
  and (_38020_, _38019_, _38018_);
  and (_38021_, _38020_, _36027_);
  nor (_38022_, _38021_, _38017_);
  and (_38023_, _38022_, _38014_);
  nor (_38024_, _36108_, _35889_);
  and (_38025_, _38024_, _36027_);
  nor (_38026_, _36158_, _35946_);
  and (_38027_, _38026_, _38025_);
  not (_38028_, _38027_);
  and (_38029_, _38007_, _36028_);
  and (_38030_, _38025_, _35946_);
  nor (_38031_, _38030_, _38029_);
  and (_38032_, _38031_, _38028_);
  and (_38033_, _38032_, _38023_);
  not (_38034_, _38033_);
  and (_38035_, _20923_, _20901_);
  not (_38036_, _38035_);
  nor (_38037_, _22050_, _21984_);
  and (_38038_, _38037_, _38036_);
  and (_38039_, _19996_, _19208_);
  and (_38040_, _38039_, _20934_);
  or (_38041_, _38040_, _21043_);
  nor (_38042_, _19996_, _20869_);
  and (_38043_, _38042_, _20923_);
  or (_38044_, _38043_, _21830_);
  nor (_38045_, _38044_, _38041_);
  and (_38046_, _38045_, _38038_);
  and (_38047_, _21841_, _22160_);
  or (_38048_, _38047_, _22215_);
  nor (_38049_, _38048_, _22204_);
  nor (_38050_, _22270_, _21348_);
  and (_38051_, _38039_, _20749_);
  and (_38052_, _21337_, _19208_);
  or (_38053_, _38052_, _38051_);
  not (_38054_, _38053_);
  and (_38055_, _38054_, _38050_);
  and (_38056_, _38055_, _38049_);
  and (_38057_, _38056_, _38046_);
  and (_38058_, _38057_, _21819_);
  nor (_38059_, _38058_, _18509_);
  nor (_38060_, _38059_, _38023_);
  nor (_38061_, _35889_, _16250_);
  and (_38062_, _35889_, _16250_);
  nor (_38063_, _38062_, _38061_);
  nor (_38064_, _36158_, _16599_);
  and (_38065_, _36158_, _16599_);
  nor (_38066_, _38065_, _38064_);
  nor (_38067_, _38066_, _38063_);
  nor (_38068_, _36108_, _16076_);
  and (_38069_, _36108_, _16076_);
  nor (_38070_, _38069_, _38068_);
  nor (_38071_, _35945_, _15935_);
  and (_38072_, _35945_, _15935_);
  nor (_38073_, _38072_, _38071_);
  nor (_38074_, _38073_, _38070_);
  nor (_38075_, _36027_, _16435_);
  and (_38076_, _36027_, _16435_);
  nor (_38077_, _38076_, _38075_);
  and (_38078_, _38077_, _38074_);
  and (_38079_, _38078_, _38067_);
  and (_38080_, _38079_, _25073_);
  not (_38081_, _38080_);
  nor (_38082_, _38081_, _38060_);
  and (_38083_, _38082_, _38034_);
  and (_38084_, _38025_, _38011_);
  and (_38085_, _38084_, _26068_);
  nor (_38086_, _36064_, _36197_);
  and (_38087_, _18564_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  not (_38088_, _38087_);
  and (_38089_, _38088_, p2in_reg[3]);
  and (_38090_, _38087_, p2_in[3]);
  or (_38091_, _38090_, _38089_);
  or (_38092_, _38091_, _38059_);
  not (_38093_, _38059_);
  or (_38094_, _38093_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_38095_, _38094_, _38092_);
  and (_38096_, _38095_, _38086_);
  not (_38097_, _36197_);
  and (_38098_, _36064_, _38097_);
  and (_38099_, _38088_, p2in_reg[2]);
  and (_38100_, _38087_, p2_in[2]);
  or (_38101_, _38100_, _38099_);
  or (_38102_, _38101_, _38059_);
  or (_38103_, _38093_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_38104_, _38103_, _38102_);
  and (_38105_, _38104_, _38098_);
  or (_38106_, _38105_, _38096_);
  nor (_38107_, _36064_, _38097_);
  and (_38108_, _38088_, p2in_reg[1]);
  and (_38109_, _38087_, p2_in[1]);
  or (_38110_, _38109_, _38108_);
  or (_38111_, _38110_, _38059_);
  or (_38112_, _38093_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_38113_, _38112_, _38111_);
  and (_38114_, _38113_, _38107_);
  and (_38115_, _36064_, _36197_);
  and (_38116_, _38088_, p2in_reg[0]);
  and (_38117_, _38087_, p2_in[0]);
  or (_38118_, _38117_, _38116_);
  or (_38119_, _38118_, _38059_);
  or (_38120_, _38093_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and (_38121_, _38120_, _38119_);
  and (_38122_, _38121_, _38115_);
  or (_38123_, _38122_, _38114_);
  or (_38124_, _38123_, _38106_);
  and (_38125_, _38124_, _38013_);
  and (_38126_, _36108_, _35946_);
  and (_38127_, _38019_, _36028_);
  and (_38128_, _38127_, _38126_);
  and (_38129_, _38086_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_38130_, _38098_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_38131_, _38130_, _38129_);
  and (_38132_, _38115_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_38133_, _38107_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  or (_38134_, _38133_, _38132_);
  or (_38135_, _38134_, _38131_);
  and (_38136_, _38135_, _38128_);
  or (_38137_, _38136_, _38125_);
  and (_38138_, _38088_, p1in_reg[3]);
  and (_38139_, _38087_, p1_in[3]);
  or (_38140_, _38139_, _38138_);
  or (_38141_, _38140_, _38059_);
  or (_38142_, _38093_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_38143_, _38142_, _38141_);
  and (_38144_, _38143_, _38086_);
  and (_38145_, _38088_, p1in_reg[2]);
  and (_38146_, _38087_, p1_in[2]);
  or (_38147_, _38146_, _38145_);
  or (_38148_, _38147_, _38059_);
  or (_38149_, _38093_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_38150_, _38149_, _38148_);
  and (_38151_, _38150_, _38098_);
  or (_38152_, _38151_, _38144_);
  and (_38153_, _38088_, p1in_reg[1]);
  and (_38154_, _38087_, p1_in[1]);
  or (_38155_, _38154_, _38153_);
  or (_38156_, _38155_, _38059_);
  or (_38157_, _38093_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_38158_, _38157_, _38156_);
  and (_38159_, _38158_, _38107_);
  and (_38160_, _38088_, p1in_reg[0]);
  and (_38161_, _38087_, p1_in[0]);
  or (_38162_, _38161_, _38160_);
  or (_38163_, _38162_, _38059_);
  or (_38164_, _38093_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and (_38165_, _38164_, _38163_);
  and (_38166_, _38165_, _38115_);
  or (_38167_, _38166_, _38159_);
  or (_38168_, _38167_, _38152_);
  and (_38169_, _38168_, _38010_);
  and (_38170_, _38115_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and (_38171_, _38086_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_38172_, _38171_, _38170_);
  and (_38173_, _38107_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_38174_, _38098_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_38175_, _38174_, _38173_);
  or (_38176_, _38175_, _38172_);
  and (_38177_, _38176_, _38084_);
  or (_38178_, _38177_, _38169_);
  or (_38179_, _38178_, _38137_);
  and (_38180_, _38179_, _35983_);
  nor (_38181_, _36064_, _17403_);
  and (_38182_, _36064_, _17403_);
  nor (_38183_, _38182_, _38181_);
  nor (_38184_, _36197_, _17598_);
  and (_38185_, _36197_, _17598_);
  nor (_38186_, _38185_, _38184_);
  and (_38187_, _38186_, _38183_);
  and (_38188_, _38187_, _38067_);
  nor (_38189_, _35983_, _16762_);
  and (_38190_, _35983_, _16762_);
  nor (_38191_, _38190_, _38189_);
  and (_38192_, _38191_, _38077_);
  and (_38193_, _38192_, _38074_);
  and (_38194_, _38193_, _38188_);
  nor (_38195_, _38033_, _24920_);
  and (_38196_, _38195_, _38194_);
  not (_38197_, _35983_);
  and (_38198_, _38088_, p2in_reg[7]);
  and (_38199_, _38087_, p2_in[7]);
  or (_38200_, _38199_, _38198_);
  or (_38201_, _38200_, _38059_);
  or (_38202_, _38093_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_38203_, _38202_, _38201_);
  and (_38204_, _38203_, _38086_);
  and (_38205_, _38088_, p2in_reg[6]);
  and (_38206_, _38087_, p2_in[6]);
  or (_38207_, _38206_, _38205_);
  or (_38208_, _38207_, _38059_);
  or (_38209_, _38093_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_38210_, _38209_, _38208_);
  and (_38211_, _38210_, _38098_);
  or (_38212_, _38211_, _38204_);
  and (_38213_, _38088_, p2in_reg[5]);
  and (_38214_, _38087_, p2_in[5]);
  or (_38215_, _38214_, _38213_);
  or (_38216_, _38215_, _38059_);
  or (_38217_, _38093_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_38218_, _38217_, _38216_);
  and (_38219_, _38218_, _38107_);
  and (_38220_, _38088_, p2in_reg[4]);
  and (_38221_, _38087_, p2_in[4]);
  or (_38222_, _38221_, _38220_);
  or (_38223_, _38222_, _38059_);
  or (_38224_, _38093_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_38225_, _38224_, _38223_);
  and (_38226_, _38225_, _38115_);
  or (_38227_, _38226_, _38219_);
  or (_38228_, _38227_, _38212_);
  and (_38229_, _38228_, _38013_);
  and (_38230_, _38086_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_38231_, _38107_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  or (_38232_, _38231_, _38230_);
  and (_38233_, _38115_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  and (_38234_, _38098_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  or (_38235_, _38234_, _38233_);
  or (_38236_, _38235_, _38232_);
  and (_38237_, _38236_, _38128_);
  or (_38238_, _38237_, _38229_);
  and (_38239_, _38088_, p1in_reg[7]);
  and (_38240_, _38087_, p1_in[7]);
  or (_38241_, _38240_, _38239_);
  or (_38242_, _38241_, _38059_);
  or (_38243_, _38093_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_38244_, _38243_, _38242_);
  and (_38245_, _38244_, _38086_);
  and (_38246_, _38088_, p1in_reg[6]);
  and (_38247_, _38087_, p1_in[6]);
  or (_38248_, _38247_, _38246_);
  or (_38249_, _38248_, _38059_);
  or (_38250_, _38093_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_38251_, _38250_, _38249_);
  and (_38252_, _38251_, _38098_);
  or (_38253_, _38252_, _38245_);
  and (_38254_, _38088_, p1in_reg[5]);
  and (_38255_, _38087_, p1_in[5]);
  or (_38256_, _38255_, _38254_);
  or (_38257_, _38256_, _38059_);
  or (_38258_, _38093_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_38259_, _38258_, _38257_);
  and (_38260_, _38259_, _38107_);
  and (_38261_, _38088_, p1in_reg[4]);
  and (_38262_, _38087_, p1_in[4]);
  or (_38263_, _38262_, _38261_);
  or (_38264_, _38263_, _38059_);
  or (_38265_, _38093_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_38266_, _38265_, _38264_);
  and (_38267_, _38266_, _38115_);
  or (_38268_, _38267_, _38260_);
  or (_38269_, _38268_, _38253_);
  and (_38270_, _38269_, _38010_);
  and (_38271_, _38115_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_38272_, _38086_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_38273_, _38272_, _38271_);
  and (_38274_, _38098_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_38275_, _38107_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or (_38276_, _38275_, _38274_);
  or (_38277_, _38276_, _38273_);
  and (_38278_, _38277_, _38084_);
  or (_38279_, _38278_, _38270_);
  or (_38280_, _38279_, _38238_);
  and (_38281_, _38280_, _38197_);
  or (_38282_, _38281_, _38196_);
  or (_38283_, _38282_, _38180_);
  and (_38284_, _38015_, _36027_);
  and (_38285_, _38107_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_38286_, _38098_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or (_38287_, _38286_, _38285_);
  and (_38288_, _38115_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  and (_38289_, _38086_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  or (_38290_, _38289_, _38288_);
  or (_38291_, _38290_, _38287_);
  and (_38292_, _38291_, _35983_);
  and (_38293_, _38107_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_38294_, _38098_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  or (_38295_, _38294_, _38293_);
  and (_38296_, _38115_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_38297_, _38086_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  or (_38298_, _38297_, _38296_);
  or (_38299_, _38298_, _38295_);
  and (_38300_, _38299_, _38197_);
  or (_38301_, _38300_, _38292_);
  and (_38302_, _38301_, _38284_);
  and (_38303_, _38098_, _25420_);
  and (_38304_, _26969_, _26221_);
  nor (_38305_, _26969_, _26221_);
  or (_38306_, _38305_, _38304_);
  and (_38307_, _27250_, _27120_);
  nor (_38308_, _27250_, _27120_);
  nor (_38309_, _38308_, _38307_);
  nor (_38310_, _38309_, _38306_);
  and (_38311_, _38309_, _38306_);
  nor (_38312_, _38311_, _38310_);
  not (_38313_, _26514_);
  and (_38314_, _38313_, _26373_);
  not (_38315_, _26373_);
  and (_38316_, _26514_, _38315_);
  nor (_38317_, _38316_, _38314_);
  and (_38318_, _26817_, _26665_);
  nor (_38319_, _26817_, _26665_);
  or (_38320_, _38319_, _38318_);
  nor (_38321_, _38320_, _38317_);
  and (_38322_, _38320_, _38317_);
  or (_38323_, _38322_, _38321_);
  or (_38324_, _38323_, _38312_);
  nand (_38325_, _38323_, _38312_);
  and (_38326_, _38325_, _38324_);
  and (_38327_, _38326_, _38115_);
  or (_38328_, _38327_, _38303_);
  and (_38329_, _38086_, _25593_);
  and (_38330_, _38107_, _25268_);
  or (_38331_, _38330_, _38329_);
  or (_38332_, _38331_, _38328_);
  and (_38333_, _38332_, _35983_);
  and (_38334_, _38098_, _25928_);
  and (_38335_, _38115_, _25679_);
  or (_38336_, _38335_, _38334_);
  and (_38337_, _38086_, _25138_);
  and (_38338_, _38107_, _25776_);
  or (_38339_, _38338_, _38337_);
  or (_38340_, _38339_, _38336_);
  and (_38341_, _38340_, _38197_);
  or (_38342_, _38341_, _38333_);
  and (_38343_, _38342_, _38009_);
  or (_38344_, _38343_, _38302_);
  and (_38345_, _38344_, _38024_);
  and (_38346_, _38020_, _36028_);
  and (_38347_, _38098_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and (_38348_, _38115_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  or (_38349_, _38348_, _38347_);
  and (_38350_, _38107_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  and (_38351_, _38086_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  or (_38352_, _38351_, _38350_);
  or (_38353_, _38352_, _38349_);
  and (_38354_, _38353_, _35983_);
  and (_38355_, _38086_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and (_38356_, _38107_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or (_38357_, _38356_, _38355_);
  and (_38358_, _38098_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and (_38359_, _38115_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  or (_38360_, _38359_, _38358_);
  or (_38361_, _38360_, _38357_);
  and (_38362_, _38361_, _38197_);
  or (_38363_, _38362_, _38354_);
  and (_38364_, _38363_, _38346_);
  and (_38365_, _38088_, p3in_reg[2]);
  and (_38366_, _38087_, p3_in[2]);
  or (_38367_, _38366_, _38365_);
  or (_38368_, _38367_, _38059_);
  or (_38369_, _38093_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_38370_, _38369_, _38368_);
  and (_38371_, _38370_, _38098_);
  and (_38372_, _38088_, p3in_reg[1]);
  and (_38373_, _38087_, p3_in[1]);
  or (_38374_, _38373_, _38372_);
  or (_38375_, _38374_, _38059_);
  or (_38376_, _38093_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_38377_, _38376_, _38375_);
  and (_38378_, _38377_, _38107_);
  or (_38379_, _38378_, _38371_);
  and (_38380_, _38088_, p3in_reg[0]);
  and (_38381_, _38087_, p3_in[0]);
  or (_38382_, _38381_, _38380_);
  or (_38383_, _38382_, _38059_);
  or (_38384_, _38093_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and (_38385_, _38384_, _38383_);
  and (_38386_, _38385_, _38115_);
  and (_38387_, _38088_, p3in_reg[3]);
  and (_38388_, _38087_, p3_in[3]);
  or (_38389_, _38388_, _38387_);
  or (_38390_, _38389_, _38059_);
  or (_38391_, _38093_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_38392_, _38391_, _38390_);
  and (_38393_, _38392_, _38086_);
  or (_38394_, _38393_, _38386_);
  or (_38395_, _38394_, _38379_);
  and (_38396_, _38395_, _35983_);
  and (_38397_, _38088_, p3in_reg[6]);
  and (_38398_, _38087_, p3_in[6]);
  or (_38399_, _38398_, _38397_);
  or (_38400_, _38399_, _38059_);
  or (_38401_, _38093_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and (_38402_, _38401_, _38400_);
  and (_38403_, _38402_, _38098_);
  and (_38404_, _38088_, p3in_reg[5]);
  and (_38405_, _38087_, p3_in[5]);
  or (_38406_, _38405_, _38404_);
  or (_38407_, _38406_, _38059_);
  or (_38408_, _38093_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_38409_, _38408_, _38407_);
  and (_38410_, _38409_, _38107_);
  or (_38411_, _38410_, _38403_);
  and (_38412_, _38088_, p3in_reg[4]);
  and (_38413_, _38087_, p3_in[4]);
  or (_38414_, _38413_, _38412_);
  or (_38415_, _38414_, _38059_);
  or (_38416_, _38093_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_38417_, _38416_, _38415_);
  and (_38418_, _38417_, _38115_);
  and (_38419_, _38088_, p3in_reg[7]);
  and (_38420_, _38087_, p3_in[7]);
  or (_38421_, _38420_, _38419_);
  or (_38422_, _38421_, _38059_);
  or (_38423_, _38093_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and (_38424_, _38423_, _38422_);
  and (_38425_, _38424_, _38086_);
  or (_38426_, _38425_, _38418_);
  or (_38427_, _38426_, _38411_);
  and (_38428_, _38427_, _38197_);
  or (_38429_, _38428_, _38396_);
  and (_38430_, _38429_, _38017_);
  or (_38431_, _38430_, _38364_);
  and (_38432_, _38088_, p0in_reg[3]);
  and (_38433_, _38087_, p0_in[3]);
  or (_38434_, _38433_, _38432_);
  or (_38435_, _38434_, _38059_);
  or (_38436_, _38093_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_38437_, _38436_, _38435_);
  and (_38438_, _38437_, _38086_);
  and (_38439_, _38088_, p0in_reg[2]);
  and (_38440_, _38087_, p0_in[2]);
  or (_38441_, _38440_, _38439_);
  or (_38442_, _38441_, _38059_);
  nand (_38443_, _38059_, _28309_);
  and (_38444_, _38443_, _38442_);
  and (_38445_, _38444_, _38098_);
  or (_38446_, _38445_, _38438_);
  and (_38447_, _38088_, p0in_reg[1]);
  and (_38448_, _38087_, p0_in[1]);
  or (_38449_, _38448_, _38447_);
  or (_38450_, _38449_, _38059_);
  or (_38451_, _38093_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_38452_, _38451_, _38450_);
  and (_38453_, _38452_, _38107_);
  and (_38454_, _38088_, p0in_reg[0]);
  and (_38455_, _38087_, p0_in[0]);
  or (_38456_, _38455_, _38454_);
  or (_38457_, _38456_, _38059_);
  nand (_38458_, _38059_, _28050_);
  and (_38459_, _38458_, _38457_);
  and (_38460_, _38459_, _38115_);
  or (_38461_, _38460_, _38453_);
  or (_38462_, _38461_, _38446_);
  and (_38463_, _38462_, _35983_);
  and (_38464_, _38088_, p0in_reg[7]);
  and (_38465_, _38087_, p0_in[7]);
  or (_38466_, _38465_, _38464_);
  or (_38467_, _38466_, _38059_);
  or (_38468_, _38093_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_38469_, _38468_, _38467_);
  and (_38470_, _38469_, _38086_);
  and (_38471_, _38088_, p0in_reg[6]);
  and (_38472_, _38087_, p0_in[6]);
  or (_38473_, _38472_, _38471_);
  or (_38474_, _38473_, _38059_);
  or (_38475_, _38093_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_38476_, _38475_, _38474_);
  and (_38477_, _38476_, _38098_);
  or (_38478_, _38477_, _38470_);
  and (_38479_, _38088_, p0in_reg[5]);
  and (_38480_, _38087_, p0_in[5]);
  or (_38481_, _38480_, _38479_);
  or (_38482_, _38481_, _38059_);
  or (_38483_, _38093_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_38484_, _38483_, _38482_);
  and (_38485_, _38484_, _38107_);
  and (_38486_, _38088_, p0in_reg[4]);
  and (_38487_, _38087_, p0_in[4]);
  or (_38488_, _38487_, _38486_);
  or (_38489_, _38488_, _38059_);
  or (_38490_, _38093_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_38491_, _38490_, _38489_);
  and (_38492_, _38491_, _38115_);
  or (_38493_, _38492_, _38485_);
  or (_38494_, _38493_, _38478_);
  and (_38495_, _38494_, _38197_);
  or (_38496_, _38495_, _38463_);
  and (_38497_, _38496_, _38021_);
  and (_38498_, _38086_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and (_38499_, _38107_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  or (_38500_, _38499_, _38498_);
  and (_38501_, _38098_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and (_38502_, _38115_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  or (_38503_, _38502_, _38501_);
  or (_38504_, _38503_, _38500_);
  and (_38505_, _38504_, _38197_);
  and (_38506_, _38086_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_38507_, _38107_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  or (_38508_, _38507_, _38506_);
  and (_38509_, _38098_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and (_38510_, _38115_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  or (_38511_, _38510_, _38509_);
  or (_38512_, _38511_, _38508_);
  and (_38513_, _38512_, _35983_);
  or (_38514_, _38513_, _38505_);
  and (_38515_, _38029_, _38015_);
  and (_38516_, _38515_, _38514_);
  or (_38517_, _38516_, _38497_);
  or (_38518_, _38517_, _38431_);
  or (_38519_, _38518_, _38345_);
  or (_38520_, _38519_, _38283_);
  nand (_38521_, _38196_, _17056_);
  and (_38522_, _38521_, _38520_);
  or (_38523_, _38522_, _38085_);
  not (_38524_, _27250_);
  and (_38525_, _38098_, _38524_);
  or (_38526_, _38525_, _35983_);
  not (_38527_, _26221_);
  and (_38528_, _38086_, _38527_);
  not (_38529_, _26969_);
  and (_38530_, _38115_, _38529_);
  not (_38531_, _27120_);
  and (_38532_, _38107_, _38531_);
  or (_38533_, _38532_, _38530_);
  or (_38534_, _38533_, _38528_);
  or (_38535_, _38534_, _38526_);
  not (_38536_, _26665_);
  and (_38537_, _38098_, _38536_);
  or (_38538_, _38537_, _38197_);
  and (_38539_, _38107_, _38313_);
  and (_38540_, _38115_, _38315_);
  not (_38541_, _26817_);
  and (_38542_, _38086_, _38541_);
  or (_38543_, _38542_, _38540_);
  or (_38544_, _38543_, _38539_);
  or (_38545_, _38544_, _38538_);
  nand (_38546_, _38545_, _38535_);
  nand (_38547_, _38546_, _38085_);
  and (_38548_, _38547_, _38523_);
  or (_38549_, _38548_, _38083_);
  and (_38550_, _38086_, ABINPUT[10]);
  or (_38551_, _38550_, _35983_);
  and (_38552_, _38107_, ABINPUT[8]);
  and (_38553_, _38115_, ABINPUT[7]);
  and (_38554_, _38098_, ABINPUT[9]);
  or (_38555_, _38554_, _38553_);
  or (_38556_, _38555_, _38552_);
  or (_38557_, _38556_, _38551_);
  and (_38558_, _38086_, ABINPUT[6]);
  or (_38559_, _38558_, _38197_);
  and (_38560_, _38107_, ABINPUT[4]);
  and (_38561_, _38115_, ABINPUT[3]);
  and (_38562_, _38098_, ABINPUT[5]);
  or (_38563_, _38562_, _38561_);
  or (_38564_, _38563_, _38560_);
  or (_38565_, _38564_, _38559_);
  nand (_38566_, _38565_, _38557_);
  nand (_38567_, _38566_, _38083_);
  and (_38568_, _38567_, _37580_);
  and (_01521_, _38568_, _38549_);
  not (_38569_, _25007_);
  and (_38570_, _38115_, _35983_);
  and (_38572_, _38570_, _38027_);
  and (_38574_, _38572_, _38569_);
  and (_38576_, _38570_, _38084_);
  and (_38578_, _38576_, _25959_);
  nor (_38580_, _38578_, _38574_);
  and (_38582_, _36027_, _35983_);
  and (_38584_, _38582_, _38086_);
  and (_38586_, _38584_, _38020_);
  nand (_38588_, _38586_, _23784_);
  and (_38590_, _38588_, _38580_);
  nor (_38592_, _38590_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_38594_, _38592_);
  nor (_38596_, _22687_, _16250_);
  and (_38598_, _38596_, _38194_);
  not (_38600_, _38598_);
  and (_38602_, _38570_, _38085_);
  not (_38604_, _24931_);
  and (_38606_, _38086_, _38197_);
  nor (_38608_, _38606_, _38604_);
  and (_38610_, _38608_, _38079_);
  nor (_38612_, _38610_, _38602_);
  and (_38614_, _38612_, _38600_);
  and (_38616_, _38614_, _38594_);
  and (_38618_, _38582_, _38098_);
  and (_38620_, _38618_, _38020_);
  and (_38622_, _38620_, _23784_);
  or (_38624_, _38622_, rst);
  nor (_01523_, _38624_, _38616_);
  or (_38627_, _38616_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  and (_38629_, _38620_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_38631_, _36028_, _35983_);
  and (_38632_, _38631_, _38115_);
  and (_38633_, _38632_, _38016_);
  and (_38634_, _38633_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  or (_38635_, _38634_, _38629_);
  and (_38636_, _38570_, _38346_);
  and (_38637_, _38636_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and (_38638_, _38632_, _38012_);
  and (_38639_, _38638_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  or (_38640_, _38639_, _38637_);
  or (_38641_, _38640_, _38635_);
  and (_38642_, _38582_, _38115_);
  and (_38643_, _38024_, _38015_);
  and (_38644_, _38643_, _38642_);
  and (_38645_, _38644_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_38646_, _38586_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_38647_, _38646_, _38645_);
  and (_38648_, _38582_, _38107_);
  and (_38649_, _38648_, _38020_);
  and (_38650_, _38649_, _35826_);
  and (_38651_, _38642_, _38016_);
  and (_38652_, _38651_, _38424_);
  or (_38653_, _38652_, _38650_);
  or (_38654_, _38653_, _38647_);
  or (_38655_, _38654_, _38641_);
  and (_38656_, _38576_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_38657_, _38642_, _38012_);
  and (_38658_, _38657_, _38203_);
  and (_38659_, _38026_, _38007_);
  and (_38660_, _38659_, _38642_);
  and (_38661_, _38660_, _38244_);
  or (_38662_, _38661_, _38658_);
  and (_38663_, _38572_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  and (_38664_, _38642_, _38020_);
  and (_38665_, _38664_, _38469_);
  or (_38666_, _38665_, _38663_);
  or (_38667_, _38666_, _38662_);
  or (_38668_, _38667_, _38656_);
  nor (_38669_, _38668_, _38655_);
  nand (_38670_, _38669_, _38616_);
  and (_38671_, _38670_, _38627_);
  or (_38672_, _38671_, _38622_);
  nand (_38673_, _38622_, _17122_);
  and (_38674_, _38673_, _37580_);
  and (_01525_, _38674_, _38672_);
  nor (_01528_, _35905_, rst);
  and (_38675_, _38620_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_38676_, _38633_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  or (_38677_, _38676_, _38675_);
  and (_38678_, _38636_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and (_38679_, _38638_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  or (_38680_, _38679_, _38678_);
  or (_38681_, _38680_, _38677_);
  and (_38682_, _38644_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  and (_38683_, _38586_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or (_38684_, _38683_, _38682_);
  and (_38685_, _38649_, _36030_);
  and (_38686_, _38651_, _38385_);
  or (_38687_, _38686_, _38685_);
  or (_38688_, _38687_, _38684_);
  or (_38689_, _38688_, _38681_);
  and (_38690_, _38576_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and (_38691_, _38657_, _38121_);
  and (_38692_, _38660_, _38165_);
  or (_38693_, _38692_, _38691_);
  and (_38694_, _38572_, _38326_);
  and (_38695_, _38664_, _38459_);
  or (_38696_, _38695_, _38694_);
  or (_38697_, _38696_, _38693_);
  or (_38698_, _38697_, _38690_);
  nor (_38699_, _38698_, _38689_);
  nand (_38700_, _38699_, _38616_);
  not (_38701_, _38622_);
  or (_38702_, _38616_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  and (_38703_, _38702_, _38701_);
  and (_38704_, _38703_, _38700_);
  and (_38705_, _38622_, ABINPUT[19]);
  or (_38706_, _38705_, _38704_);
  and (_02204_, _38706_, _37580_);
  and (_38707_, _38620_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_38708_, _38633_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  or (_38709_, _38708_, _38707_);
  and (_38710_, _38570_, _38128_);
  and (_38711_, _38710_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_38713_, _38636_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or (_38714_, _38713_, _38711_);
  or (_38715_, _38714_, _38709_);
  and (_38716_, _38644_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_38717_, _38586_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_38718_, _38717_, _38716_);
  and (_38719_, _38649_, _36182_);
  and (_38720_, _38651_, _38377_);
  or (_38721_, _38720_, _38719_);
  or (_38722_, _38721_, _38718_);
  or (_38723_, _38722_, _38715_);
  and (_38725_, _38576_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_38726_, _38657_, _38113_);
  and (_38727_, _38660_, _38158_);
  or (_38728_, _38727_, _38726_);
  and (_38729_, _38572_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_38730_, _38664_, _38452_);
  or (_38731_, _38730_, _38729_);
  or (_38732_, _38731_, _38728_);
  or (_38733_, _38732_, _38725_);
  nor (_38734_, _38733_, _38723_);
  nand (_38735_, _38734_, _38616_);
  or (_38736_, _38616_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  and (_38737_, _38736_, _38701_);
  and (_38738_, _38737_, _38735_);
  and (_38739_, _38622_, ABINPUT[20]);
  or (_38740_, _38739_, _38738_);
  and (_02206_, _38740_, _37580_);
  or (_38741_, _38616_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  and (_38742_, _38620_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_38743_, _38633_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_38744_, _38743_, _38742_);
  and (_38745_, _38636_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and (_38746_, _38638_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_38747_, _38746_, _38745_);
  or (_38748_, _38747_, _38744_);
  and (_38749_, _38644_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_38750_, _38586_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_38751_, _38750_, _38749_);
  and (_38752_, _38649_, _35963_);
  and (_38753_, _38651_, _38370_);
  or (_38755_, _38753_, _38752_);
  or (_38756_, _38755_, _38751_);
  or (_38757_, _38756_, _38748_);
  and (_38758_, _38576_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_38759_, _38657_, _38104_);
  and (_38760_, _38660_, _38150_);
  or (_38761_, _38760_, _38759_);
  and (_38762_, _38572_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  and (_38763_, _38664_, _38444_);
  or (_38764_, _38763_, _38762_);
  or (_38765_, _38764_, _38761_);
  or (_38766_, _38765_, _38758_);
  nor (_38767_, _38766_, _38757_);
  nand (_38768_, _38767_, _38616_);
  and (_38769_, _38768_, _38741_);
  or (_38770_, _38769_, _38622_);
  nand (_38771_, _38622_, _17707_);
  and (_38772_, _38771_, _37580_);
  and (_02208_, _38772_, _38770_);
  or (_38773_, _38616_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  and (_38775_, _38620_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_38776_, _38633_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  or (_38777_, _38776_, _38775_);
  and (_38778_, _38636_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and (_38779_, _38710_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  or (_38780_, _38779_, _38778_);
  or (_38781_, _38780_, _38777_);
  and (_38782_, _38644_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_38783_, _38586_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_38784_, _38783_, _38782_);
  and (_38785_, _38649_, _35992_);
  and (_38786_, _38651_, _38392_);
  or (_38787_, _38786_, _38785_);
  or (_38788_, _38787_, _38784_);
  or (_38789_, _38788_, _38781_);
  and (_38790_, _38576_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_38791_, _38657_, _38095_);
  and (_38792_, _38660_, _38143_);
  or (_38793_, _38792_, _38791_);
  and (_38794_, _38572_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_38795_, _38664_, _38437_);
  or (_38796_, _38795_, _38794_);
  or (_38797_, _38796_, _38793_);
  or (_38798_, _38797_, _38790_);
  nor (_38799_, _38798_, _38789_);
  nand (_38800_, _38799_, _38616_);
  and (_38801_, _38800_, _38773_);
  or (_38802_, _38801_, _38622_);
  nand (_38803_, _38622_, _17891_);
  and (_38804_, _38803_, _37580_);
  and (_02210_, _38804_, _38802_);
  or (_38805_, _38616_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  and (_38806_, _38620_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_38807_, _38633_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  or (_38808_, _38807_, _38806_);
  and (_38809_, _38636_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and (_38810_, _38710_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  or (_38811_, _38810_, _38809_);
  or (_38812_, _38811_, _38808_);
  and (_38813_, _38644_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_38814_, _38586_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or (_38815_, _38814_, _38813_);
  and (_38816_, _38649_, _36133_);
  and (_38817_, _38651_, _38417_);
  or (_38818_, _38817_, _38816_);
  or (_38819_, _38818_, _38815_);
  or (_38820_, _38819_, _38812_);
  and (_38821_, _38576_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_38822_, _38657_, _38225_);
  and (_38823_, _38660_, _38266_);
  or (_38824_, _38823_, _38822_);
  and (_38825_, _38572_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_38826_, _38664_, _38491_);
  or (_38827_, _38826_, _38825_);
  or (_38828_, _38827_, _38824_);
  or (_38829_, _38828_, _38821_);
  nor (_38830_, _38829_, _38820_);
  nand (_38831_, _38830_, _38616_);
  and (_38832_, _38831_, _38805_);
  or (_38833_, _38832_, _38622_);
  nand (_38834_, _38622_, _18054_);
  and (_38835_, _38834_, _37580_);
  and (_02212_, _38835_, _38833_);
  and (_38836_, _38620_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_38837_, _38633_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  or (_38838_, _38837_, _38836_);
  and (_38839_, _38636_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and (_38840_, _38638_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  or (_38841_, _38840_, _38839_);
  or (_38842_, _38841_, _38838_);
  and (_38843_, _38644_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_38844_, _38586_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or (_38845_, _38844_, _38843_);
  and (_38846_, _38649_, _35908_);
  and (_38847_, _38651_, _38409_);
  or (_38848_, _38847_, _38846_);
  or (_38849_, _38848_, _38845_);
  or (_38850_, _38849_, _38842_);
  and (_38851_, _38576_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_38852_, _38657_, _38218_);
  and (_38853_, _38660_, _38259_);
  or (_38854_, _38853_, _38852_);
  and (_38855_, _38572_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_38856_, _38664_, _38484_);
  or (_38857_, _38856_, _38855_);
  or (_38858_, _38857_, _38854_);
  or (_38859_, _38858_, _38851_);
  nor (_38860_, _38859_, _38850_);
  nand (_38861_, _38860_, _38616_);
  or (_38862_, _38616_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  and (_38863_, _38862_, _38701_);
  and (_38864_, _38863_, _38861_);
  and (_38865_, _38622_, ABINPUT[24]);
  or (_38866_, _38865_, _38864_);
  and (_02214_, _38866_, _37580_);
  and (_38867_, _38620_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_38868_, _38633_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  or (_38869_, _38868_, _38867_);
  and (_38870_, _38636_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and (_38871_, _38638_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  or (_38872_, _38871_, _38870_);
  or (_38873_, _38872_, _38869_);
  and (_38874_, _38644_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_38875_, _38586_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_38876_, _38875_, _38874_);
  and (_38877_, _38649_, _36075_);
  and (_38878_, _38651_, _38402_);
  or (_38879_, _38878_, _38877_);
  or (_38880_, _38879_, _38876_);
  or (_38881_, _38880_, _38873_);
  and (_38882_, _38576_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_38883_, _38657_, _38210_);
  and (_38884_, _38660_, _38251_);
  or (_38885_, _38884_, _38883_);
  and (_38886_, _38572_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_38887_, _38664_, _38476_);
  or (_38888_, _38887_, _38886_);
  or (_38889_, _38888_, _38885_);
  or (_38890_, _38889_, _38882_);
  nor (_38891_, _38890_, _38881_);
  nand (_38892_, _38891_, _38616_);
  or (_38893_, _38616_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  and (_38894_, _38893_, _38701_);
  and (_38895_, _38894_, _38892_);
  and (_38896_, _38622_, ABINPUT[25]);
  or (_38897_, _38896_, _38895_);
  and (_02216_, _38897_, _37580_);
  or (_38898_, _38087_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  not (_38899_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nand (_38900_, _38087_, _38899_);
  and (_38901_, _38900_, _37580_);
  and (_02779_, _38901_, _38898_);
  and (_38902_, _38088_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  and (_38903_, _38087_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  or (_38904_, _38903_, _38902_);
  and (_02783_, _38904_, _37580_);
  nor (_03161_, _35889_, rst);
  nor (_03168_, _36137_, rst);
  nor (_03172_, _35884_, rst);
  and (_38905_, _22435_, _20727_);
  nor (_38906_, _21940_, _35903_);
  not (_38907_, _38906_);
  nor (_38908_, _21940_, _18509_);
  nor (_38909_, _38905_, _38908_);
  and (_38910_, _38909_, _38907_);
  nor (_38911_, _38910_, _38905_);
  nor (_38912_, _22687_, _17023_);
  and (_38913_, _38912_, _38911_);
  and (_38914_, _38913_, _38079_);
  nor (_38915_, ABINPUT[28], ABINPUT[27]);
  nor (_38916_, ABINPUT[30], ABINPUT[29]);
  and (_38917_, _38916_, _38915_);
  nor (_38918_, ABINPUT[32], ABINPUT[31]);
  nor (_38919_, ABINPUT[33], ABINPUT[34]);
  and (_38920_, _38919_, _38918_);
  and (_38921_, _38920_, _38917_);
  not (_38922_, _22435_);
  and (_38923_, _38910_, _38922_);
  and (_38924_, _38923_, _38921_);
  and (_38925_, _38905_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_38926_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_38927_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_38928_, _38927_, _38926_);
  nor (_38929_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor (_38930_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_38931_, _38930_, _38929_);
  and (_38932_, _38931_, _38928_);
  and (_38933_, _38932_, _21501_);
  or (_38934_, _38933_, _38925_);
  nor (_38935_, _38934_, _38924_);
  not (_38936_, \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  and (_38937_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _38936_);
  and (_38938_, _36335_, _36333_);
  and (_38939_, _36378_, _36377_);
  nor (_38940_, _38939_, _38938_);
  and (_38941_, _36364_, _36363_);
  and (_38942_, _36351_, _36350_);
  nor (_38943_, _38942_, _38941_);
  and (_38944_, _38943_, _38940_);
  and (_38945_, _36392_, _36391_);
  and (_38946_, _36320_, _36317_);
  nor (_38947_, _38946_, _38945_);
  and (_38948_, _36309_, _36305_);
  and (_38949_, _36283_, _36282_);
  nor (_38950_, _38949_, _38948_);
  and (_38951_, _38950_, _38947_);
  and (_38952_, _38951_, _38944_);
  nor (_38953_, _38952_, _38937_);
  and (_38954_, _38937_, \oc8051_top_1.oc8051_sfr1.bit_out );
  nor (_38955_, _38954_, _38953_);
  not (_38956_, _38955_);
  and (_38957_, _38956_, _38911_);
  not (_38958_, _38957_);
  and (_38959_, _38958_, _38935_);
  and (_38960_, _22424_, _20858_);
  nor (_38961_, _38960_, _22402_);
  or (_38962_, _38961_, _38959_);
  and (_38963_, _21250_, _21196_);
  and (_38964_, _21141_, _19746_);
  nor (_38965_, _38964_, _38963_);
  not (_38966_, _38965_);
  or (_38967_, _22160_, _21907_);
  or (_38968_, _38967_, _21250_);
  and (_38969_, _38968_, _19746_);
  not (_38970_, _38969_);
  not (_38971_, _38051_);
  and (_38972_, _21687_, _20760_);
  and (_38973_, _21841_, _21305_);
  nor (_38974_, _38973_, _38972_);
  not (_38975_, _38974_);
  and (_38976_, _21305_, _19208_);
  or (_38977_, _38976_, _21316_);
  nor (_38978_, _38977_, _38975_);
  and (_38979_, _38978_, _38971_);
  and (_38980_, _38979_, _38970_);
  not (_38981_, _38980_);
  and (_38982_, _38981_, _38959_);
  nor (_38983_, _38982_, _38966_);
  and (_38984_, _38983_, _38962_);
  nor (_38985_, _38984_, _35903_);
  and (_38986_, _21676_, _19218_);
  and (_38987_, _21337_, _20803_);
  nor (_38988_, _38987_, _38986_);
  nor (_38989_, _38988_, _18509_);
  nor (_38990_, _38989_, _21446_);
  not (_38991_, _38990_);
  nor (_38992_, _38991_, _38985_);
  nor (_38993_, _38569_, _24942_);
  and (_38994_, _38993_, _25105_);
  not (_38995_, _38994_);
  and (_38996_, _38995_, _38905_);
  nor (_38997_, _26242_, _26014_);
  not (_38998_, _38997_);
  and (_38999_, _38998_, _21501_);
  nor (_39000_, _38999_, _38996_);
  not (_39001_, _39000_);
  nor (_39002_, _39001_, _38992_);
  not (_39003_, _39002_);
  nor (_39005_, _39003_, _38914_);
  and (_39006_, _39005_, _38600_);
  nor (_39007_, _21457_, rst);
  and (_03181_, _39007_, _39006_);
  and (_03185_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _37580_);
  and (_03188_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [7], _37580_);
  and (_39009_, _21479_, _38963_);
  nor (_39010_, _39009_, _38989_);
  nor (_39011_, _38978_, _35903_);
  not (_39012_, _39011_);
  not (_39014_, _21457_);
  and (_39015_, _38987_, _22600_);
  and (_39016_, _21885_, _22600_);
  nor (_39017_, _39016_, _39015_);
  and (_39018_, _39017_, _39014_);
  and (_39020_, _39018_, _38907_);
  and (_39021_, _39020_, _39012_);
  and (_39022_, _38965_, _21940_);
  and (_39023_, _39022_, _38979_);
  nor (_39024_, _39023_, _35903_);
  nor (_39026_, _39016_, _22435_);
  not (_39027_, _39026_);
  nor (_39028_, _39027_, _39024_);
  and (_39029_, _39028_, _39021_);
  and (_39030_, _39029_, _39010_);
  and (_39032_, _39030_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  not (_39033_, _39010_);
  and (_39034_, _39033_, _39021_);
  and (_39035_, _20825_, _22600_);
  and (_39036_, _39035_, _19746_);
  not (_39038_, _39036_);
  nor (_39039_, _39024_, _22435_);
  and (_39041_, _39039_, _39038_);
  and (_39042_, _39041_, _39034_);
  and (_39043_, \oc8051_top_1.oc8051_memory_interface1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  not (_39044_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_39045_, \oc8051_top_1.oc8051_memory_interface1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_39046_, _39045_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nand (_39047_, _39046_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nor (_39049_, _39047_, _39044_);
  and (_39050_, _39049_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_39051_, _39050_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_39053_, _39051_, _39043_);
  and (_39054_, _39053_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_39055_, _39054_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_39057_, _39055_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_39058_, _39057_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nand (_39059_, _39058_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand (_39061_, _39059_, _38899_);
  or (_39062_, _39059_, _38899_);
  and (_39063_, _39062_, _39061_);
  and (_39065_, _39063_, _39042_);
  and (_39066_, _39009_, ABINPUT[18]);
  or (_39067_, _39066_, _39065_);
  or (_39069_, _39067_, _39032_);
  and (_39070_, _39021_, _35848_);
  nor (_39071_, _39021_, _37886_);
  nor (_39073_, _39071_, _39070_);
  not (_39074_, _39073_);
  not (_39076_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  not (_39077_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  not (_39078_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  not (_39079_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_39080_, _39073_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor (_39081_, _39073_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_39082_, _39021_, _36090_);
  nor (_39084_, _39021_, _38005_);
  nor (_39085_, _39084_, _39082_);
  and (_39086_, _39085_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_39088_, _39085_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_39089_, _39088_, _39086_);
  and (_39090_, _39021_, _35923_);
  nor (_39092_, _39021_, _37988_);
  nor (_39093_, _39092_, _39090_);
  and (_39094_, _39093_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nor (_39096_, _39093_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_39097_, _39021_, _36153_);
  nor (_39098_, _39021_, _37971_);
  nor (_39100_, _39098_, _39097_);
  nand (_39101_, _39100_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_39102_, _39021_, _36022_);
  nor (_39104_, _39021_, _37954_);
  nor (_39105_, _39104_, _39102_);
  and (_39106_, _39105_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nor (_39108_, _39105_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_39109_, _39021_, _35978_);
  nor (_39111_, _39021_, _37937_);
  nor (_39112_, _39111_, _39109_);
  and (_39113_, _39112_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_39114_, _39021_, _36177_);
  nor (_39115_, _39021_, _37920_);
  nor (_39117_, _39115_, _39114_);
  and (_39118_, _39117_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_39119_, _39021_, _36059_);
  nor (_39121_, _39021_, _37903_);
  nor (_39122_, _39121_, _39119_);
  and (_39123_, _39122_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor (_39125_, _39117_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nor (_39126_, _39125_, _39118_);
  and (_39127_, _39126_, _39123_);
  nor (_39129_, _39127_, _39118_);
  not (_39130_, _39129_);
  nor (_39131_, _39112_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nor (_39133_, _39131_, _39113_);
  and (_39134_, _39133_, _39130_);
  nor (_39135_, _39134_, _39113_);
  nor (_39137_, _39135_, _39108_);
  or (_39138_, _39137_, _39106_);
  or (_39139_, _39100_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_39141_, _39139_, _39101_);
  nand (_39142_, _39141_, _39138_);
  and (_39144_, _39142_, _39101_);
  nor (_39145_, _39144_, _39096_);
  or (_39146_, _39145_, _39094_);
  and (_39147_, _39146_, _39089_);
  nor (_39148_, _39147_, _39086_);
  nor (_39149_, _39148_, _39081_);
  or (_39150_, _39149_, _39080_);
  nor (_39152_, _39150_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_39153_, _39152_, _39079_);
  and (_39154_, _39153_, _39078_);
  and (_39156_, _39154_, _39077_);
  nor (_39157_, \oc8051_top_1.oc8051_memory_interface1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_39158_, _39157_, _39156_);
  and (_39160_, _39158_, _39076_);
  nor (_39161_, _39160_, _39074_);
  and (_39162_, \oc8051_top_1.oc8051_memory_interface1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_39164_, _39162_, _39043_);
  and (_39165_, _39164_, _39150_);
  and (_39166_, _39165_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_39168_, _39166_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_39169_, _39168_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor (_39170_, _39169_, _39073_);
  nor (_39172_, _39170_, _39161_);
  or (_39173_, _39172_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nand (_39174_, _39172_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_39176_, _39174_, _39173_);
  nor (_39177_, _39041_, _39034_);
  and (_39179_, _39177_, _39176_);
  or (_39180_, _39179_, _39069_);
  and (_39181_, _39015_, _35849_);
  and (_39182_, _21435_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and (_39184_, _39182_, _20836_);
  and (_39185_, _39184_, ABINPUT[26]);
  nor (_39186_, _39185_, _39181_);
  nand (_39188_, _39186_, _39006_);
  or (_39189_, _39188_, _39180_);
  and (_39190_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11], \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor (_39192_, _18629_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_39193_, _39192_, _35832_);
  nor (_39194_, _39193_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  not (_39196_, _39194_);
  and (_39197_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4], \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_39198_, _39197_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and (_39200_, _39198_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and (_39201_, _39200_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_39202_, _39201_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and (_39204_, _39202_, _39196_);
  and (_39205_, _39204_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_39206_, _39205_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and (_39208_, _39206_, _39190_);
  and (_39209_, _39208_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and (_39211_, _39209_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and (_39212_, _39211_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or (_39213_, _39212_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nand (_39214_, _39212_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_39216_, _39214_, _39213_);
  or (_39217_, _39216_, _39006_);
  and (_39218_, _39217_, _37580_);
  and (_03191_, _39218_, _39189_);
  not (_39220_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_39221_, _18553_, _39220_);
  not (_39223_, _39221_);
  not (_39224_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  not (_39225_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  not (_39227_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  not (_39228_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  not (_39229_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  not (_39231_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  not (_39232_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  not (_39233_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  not (_39235_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  not (_39236_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_39237_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4], \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_39239_, _39237_, _39236_);
  and (_39240_, _39239_, _39235_);
  and (_39242_, _39240_, _39233_);
  and (_39243_, _39242_, _39232_);
  and (_39244_, _39243_, _39231_);
  and (_39245_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_39247_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_39248_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_39249_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  nor (_39251_, _39249_, _39247_);
  and (_39252_, _39251_, _39248_);
  nor (_39253_, _39252_, _39247_);
  nor (_39255_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_39256_, _39255_, _39245_);
  not (_39257_, _39256_);
  nor (_39259_, _39257_, _39253_);
  nor (_39260_, _39259_, _39245_);
  and (_39261_, _39260_, _39244_);
  and (_39263_, _39261_, _39229_);
  and (_39264_, _39263_, _39228_);
  and (_39265_, _39264_, _39227_);
  and (_39267_, _39265_, _39225_);
  and (_39268_, _39267_, _39224_);
  nor (_39269_, _39267_, _39224_);
  nor (_39271_, _39269_, _39268_);
  not (_39272_, _39271_);
  nor (_39274_, _39265_, _39225_);
  nor (_39275_, _39274_, _39267_);
  not (_39276_, _39275_);
  nor (_39277_, _39264_, _39227_);
  nor (_39278_, _39277_, _39265_);
  not (_39279_, _39278_);
  nor (_39280_, _39263_, _39228_);
  nor (_39282_, _39280_, _39264_);
  not (_39283_, _39282_);
  nor (_39284_, _39261_, _39229_);
  or (_39286_, _39284_, _39263_);
  and (_39287_, _39260_, _39243_);
  nor (_39288_, _39287_, _39231_);
  nor (_39290_, _39288_, _39261_);
  not (_39291_, _39290_);
  and (_39292_, _39260_, _39242_);
  and (_39294_, _39260_, _39240_);
  nor (_39295_, _39294_, _39233_);
  nor (_39296_, _39295_, _39292_);
  not (_39298_, _39296_);
  and (_39299_, _39260_, _39239_);
  nor (_39300_, _39299_, _39235_);
  nor (_39302_, _39300_, _39294_);
  not (_39303_, _39302_);
  and (_39304_, _39260_, _39237_);
  nor (_39306_, _39304_, _39236_);
  nor (_39307_, _39306_, _39299_);
  not (_39309_, _39307_);
  not (_39310_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_39311_, _39260_, _39310_);
  nor (_39312_, _39260_, _39310_);
  nor (_39314_, _39312_, _39311_);
  not (_39315_, _39314_);
  not (_39316_, _19462_);
  and (_39318_, _19186_, _18935_);
  and (_39319_, _39318_, _39316_);
  and (_39320_, _39319_, _19702_);
  not (_39322_, _19186_);
  nor (_39323_, _39322_, _18935_);
  and (_39324_, _39323_, _19462_);
  nor (_39326_, _39324_, _39320_);
  not (_39327_, _20454_);
  and (_39328_, _39327_, _20214_);
  and (_39330_, _20694_, _19975_);
  and (_39331_, _39330_, _39328_);
  not (_39332_, _19702_);
  and (_39334_, _39332_, _19462_);
  and (_39335_, _39334_, _39323_);
  not (_39336_, _20694_);
  nor (_39338_, _20454_, _20214_);
  and (_39339_, _39338_, _39336_);
  and (_39341_, _39339_, _19964_);
  and (_39342_, _39341_, _39335_);
  nor (_39343_, _39342_, _39331_);
  nor (_39344_, _39343_, _39326_);
  not (_39346_, _39344_);
  and (_39347_, _19702_, _19462_);
  and (_39348_, _39347_, _39318_);
  and (_39350_, _20454_, _20214_);
  and (_39351_, _39336_, _19964_);
  nor (_39352_, _39351_, _39330_);
  and (_39354_, _39352_, _39350_);
  and (_39355_, _39354_, _39348_);
  and (_39356_, _20694_, _19964_);
  and (_39358_, _39356_, _39338_);
  and (_39359_, _39358_, _39335_);
  nor (_39360_, _39359_, _39355_);
  and (_39362_, _39350_, _20694_);
  and (_39363_, _39362_, _39320_);
  not (_39364_, _39363_);
  not (_39366_, _20214_);
  and (_39367_, _20454_, _39366_);
  and (_39368_, _39367_, _39330_);
  and (_39370_, _39351_, _39328_);
  or (_39371_, _39370_, _39368_);
  and (_39373_, _39371_, _39335_);
  and (_39374_, _39347_, _39323_);
  and (_39375_, _39367_, _39351_);
  and (_39376_, _39375_, _39374_);
  nor (_39378_, _39376_, _39373_);
  and (_39379_, _39378_, _39364_);
  and (_39380_, _39379_, _39360_);
  and (_39382_, _39319_, _39332_);
  and (_39383_, _39382_, _39331_);
  and (_39384_, _39367_, _39356_);
  and (_39386_, _39384_, _39348_);
  nor (_39387_, _39386_, _39383_);
  not (_39388_, _39387_);
  and (_39390_, _39356_, _39328_);
  not (_39391_, _39390_);
  nor (_39392_, _39391_, _39326_);
  nor (_39394_, _39392_, _39388_);
  nor (_39395_, _20694_, _19964_);
  and (_39396_, _39395_, _39338_);
  and (_39398_, _39396_, _39335_);
  and (_39399_, _39375_, _39335_);
  and (_39400_, _39390_, _39382_);
  or (_39402_, _39400_, _39399_);
  nor (_39403_, _39402_, _39398_);
  and (_39405_, _39403_, _39394_);
  and (_39406_, _39405_, _39380_);
  and (_39407_, _39406_, _39346_);
  not (_39408_, _39350_);
  and (_39409_, _39374_, _39336_);
  nor (_39411_, _39409_, _39335_);
  nor (_39412_, _39411_, _39408_);
  not (_39413_, _39412_);
  not (_39415_, _39320_);
  and (_39416_, _39338_, _39330_);
  not (_39417_, _39416_);
  not (_39419_, _39358_);
  nor (_39420_, _39375_, _39370_);
  and (_39421_, _39420_, _39419_);
  and (_39423_, _39421_, _39417_);
  nor (_39424_, _39423_, _39415_);
  not (_39425_, _39424_);
  and (_39427_, _39367_, _39395_);
  nor (_39428_, _39427_, _39370_);
  nor (_39429_, _39428_, _19186_);
  not (_39431_, _39429_);
  nor (_39432_, _39427_, _39384_);
  nor (_39433_, _39432_, _39415_);
  not (_39435_, _39374_);
  nor (_39436_, _39384_, _39370_);
  nor (_39438_, _39436_, _39435_);
  nor (_39439_, _39438_, _39433_);
  and (_39440_, _39439_, _39431_);
  and (_39441_, _39440_, _39425_);
  and (_39443_, _39441_, _39413_);
  and (_39444_, _39390_, _39348_);
  and (_39445_, _39350_, _39351_);
  and (_39447_, _39445_, _39348_);
  nor (_39448_, _39447_, _39444_);
  and (_39449_, _39348_, _39331_);
  and (_39451_, _39358_, _39322_);
  nor (_39452_, _39451_, _39449_);
  and (_39453_, _39452_, _39448_);
  not (_39455_, _39335_);
  nor (_39456_, _39416_, _39384_);
  nor (_39457_, _39456_, _39455_);
  not (_39459_, _39368_);
  nor (_39460_, _39320_, _39322_);
  nor (_39461_, _39460_, _39459_);
  nor (_39463_, _39461_, _39457_);
  and (_39464_, _39463_, _39453_);
  and (_39465_, _39368_, _39348_);
  and (_39467_, _39375_, _39348_);
  nor (_39468_, _39467_, _39465_);
  and (_39470_, _39395_, _39328_);
  not (_39471_, _39470_);
  nor (_39472_, _39324_, _39319_);
  nor (_39473_, _39472_, _39471_);
  and (_39475_, _39328_, _39336_);
  nor (_39476_, _19462_, _18935_);
  and (_39477_, _39476_, _19186_);
  and (_39479_, _39477_, _19964_);
  and (_39480_, _39479_, _39475_);
  nor (_39481_, _39480_, _39473_);
  and (_39483_, _39481_, _39468_);
  and (_39484_, _39375_, _39322_);
  not (_39485_, _39484_);
  and (_39487_, _39334_, _39318_);
  not (_39488_, _39356_);
  and (_39489_, _39367_, _39488_);
  and (_39491_, _39489_, _39477_);
  nor (_39492_, _39491_, _39487_);
  and (_39493_, _39492_, _39485_);
  not (_39495_, _39348_);
  and (_39496_, _39338_, _20694_);
  nor (_39497_, _39427_, _39496_);
  nor (_39499_, _39497_, _39495_);
  and (_39500_, _39475_, _39348_);
  nor (_39502_, _39500_, _39499_);
  and (_39503_, _39502_, _39493_);
  and (_39504_, _39503_, _39483_);
  and (_39505_, _39504_, _39464_);
  and (_39507_, _39505_, _39443_);
  and (_39508_, _39507_, _39407_);
  nor (_39509_, _39251_, _39248_);
  nor (_39511_, _39509_, _39252_);
  not (_39512_, _39511_);
  nor (_39513_, _39512_, _39508_);
  not (_39515_, _39513_);
  and (_39516_, _39470_, _39382_);
  or (_39517_, _39476_, _39322_);
  and (_39519_, _39517_, _39375_);
  or (_39520_, _39519_, _39447_);
  or (_39521_, _39520_, _39516_);
  or (_39523_, _39402_, _39388_);
  nor (_39524_, _39523_, _39521_);
  nand (_39525_, _39524_, _39380_);
  nor (_39527_, _39525_, _39508_);
  not (_39528_, _39527_);
  nor (_39529_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_39531_, _39529_, _39248_);
  and (_39532_, _39531_, _39528_);
  and (_39533_, _39512_, _39508_);
  nor (_39534_, _39533_, _39513_);
  nand (_39535_, _39534_, _39532_);
  and (_39536_, _39535_, _39515_);
  not (_39537_, _39536_);
  and (_39538_, _39257_, _39253_);
  nor (_39539_, _39538_, _39259_);
  and (_39540_, _39539_, _39537_);
  and (_39541_, _39540_, _39315_);
  not (_39542_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_39543_, _39311_, _39542_);
  or (_39544_, _39543_, _39304_);
  and (_39545_, _39544_, _39541_);
  and (_39546_, _39545_, _39309_);
  and (_39547_, _39546_, _39303_);
  and (_39548_, _39547_, _39298_);
  nor (_39549_, _39292_, _39232_);
  or (_39550_, _39549_, _39287_);
  and (_39551_, _39550_, _39548_);
  and (_39552_, _39551_, _39291_);
  and (_39553_, _39552_, _39286_);
  and (_39554_, _39553_, _39283_);
  and (_39555_, _39554_, _39279_);
  and (_39556_, _39555_, _39276_);
  and (_39557_, _39556_, _39272_);
  nor (_39558_, _39557_, _39223_);
  nor (_39559_, _39221_, _38899_);
  not (_39560_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_39561_, _39268_, _39560_);
  nor (_39562_, _39268_, _39560_);
  nor (_39563_, _39562_, _39561_);
  and (_39564_, _39563_, _39221_);
  or (_39565_, _39564_, _39559_);
  or (_39566_, _39565_, _39558_);
  nand (_39567_, _39563_, _39558_);
  nor (_39568_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , rst);
  and (_39569_, _39568_, _39567_);
  and (_39570_, _39569_, _39566_);
  and (_39571_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _37580_);
  and (_39572_, _39571_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  or (_03194_, _39572_, _39570_);
  nor (_39573_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , rst);
  and (_03199_, _39573_, \oc8051_top_1.oc8051_memory_interface1.int_ack_buff );
  and (_03202_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , _37580_);
  nor (_39574_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  nor (_39575_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_39576_, _39575_, _39574_);
  nor (_39577_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  nor (_39578_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and (_39579_, _39578_, _39577_);
  and (_39580_, _39579_, _39576_);
  nor (_39581_, _39580_, rst);
  and (_39582_, \oc8051_top_1.oc8051_rom1.ea_int , _18520_);
  nand (_39583_, _39582_, _18553_);
  and (_39584_, _39583_, _03202_);
  or (_03205_, _39584_, _39581_);
  and (_39585_, _39580_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  or (_39586_, _39585_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  and (_03208_, _39586_, _37580_);
  nor (_39587_, _39194_, _35832_);
  nor (_39588_, _39508_, _18749_);
  not (_39589_, _39588_);
  nor (_39590_, _39527_, _18662_);
  and (_39591_, _39508_, _18749_);
  nor (_39592_, _39591_, _39588_);
  nand (_39593_, _39592_, _39590_);
  and (_39594_, _39593_, _39589_);
  nor (_39595_, _39594_, _35832_);
  and (_39596_, _39595_, _18618_);
  nor (_39597_, _39595_, _18618_);
  nor (_39598_, _39597_, _39596_);
  nor (_39599_, _39598_, _39587_);
  and (_39600_, _18760_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_39601_, _39600_, _39587_);
  and (_39602_, _39601_, _39525_);
  or (_39603_, _39602_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_39604_, _39603_, _39599_);
  and (_03210_, _39604_, _37580_);
  nor (_39605_, _20411_, _20171_);
  not (_39606_, _19659_);
  and (_39607_, _20651_, _39606_);
  and (_39608_, _39607_, _39605_);
  and (_39609_, _18553_, _37580_);
  and (_39610_, _39609_, _18542_);
  and (_39611_, _39610_, _18869_);
  and (_39612_, _39611_, _19898_);
  nor (_39613_, _19142_, _19419_);
  and (_39614_, _39613_, _39612_);
  and (_03218_, _39614_, _39608_);
  nor (_39615_, \oc8051_top_1.oc8051_memory_interface1.istb_t , rst);
  and (_39616_, _39615_, \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  and (_39617_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [7]);
  and (_03223_, \oc8051_top_1.oc8051_memory_interface1.istb_t , _37580_);
  and (_39618_, _03223_, _39617_);
  or (_03220_, _39618_, _39616_);
  not (_39619_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and (_39620_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_39621_, _39620_, _39619_);
  and (_39622_, _39620_, _39619_);
  nor (_39623_, _39622_, _39621_);
  not (_39624_, _39623_);
  and (_39625_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and (_39626_, _39625_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_39627_, _39625_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_39628_, _39627_, _39626_);
  or (_39629_, _39628_, _39620_);
  and (_39630_, _39629_, _39624_);
  nor (_39631_, _39621_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and (_39632_, _39621_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  or (_39633_, _39632_, _39631_);
  or (_39634_, _39626_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  and (_03229_, _39634_, _37580_);
  and (_39635_, _03229_, _39633_);
  and (_03226_, _39635_, _39630_);
  not (_39636_, \oc8051_top_1.oc8051_rom1.ea_int );
  nor (_39637_, _39194_, _39636_);
  and (_39638_, _39637_, \oc8051_top_1.oc8051_rom1.data_o [31]);
  not (_39639_, _39637_);
  and (_39640_, _39639_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  or (_39641_, _39640_, _39638_);
  and (_03232_, _39641_, _37580_);
  and (_39642_, _39637_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and (_39643_, _39639_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  or (_39644_, _39643_, _39642_);
  and (_03234_, _39644_, _37580_);
  and (_39645_, \oc8051_top_1.oc8051_decoder1.mem_act [2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  not (_39646_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_39647_, \oc8051_top_1.oc8051_decoder1.mem_act [0], _39646_);
  and (_39648_, _39647_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_39649_, _39648_, _39645_);
  and (_03236_, _39649_, _37580_);
  and (_39650_, \oc8051_top_1.oc8051_memory_interface1.dwe_o , \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_39651_, _39650_, _39647_);
  and (_03238_, _39651_, _37580_);
  or (_39652_, _39646_, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  and (_03240_, _39652_, _37580_);
  not (_39653_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  and (_39654_, _39653_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_39655_, _39654_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_39656_, _39646_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  and (_39657_, _39656_, _37580_);
  and (_03242_, _39657_, _39655_);
  or (_39658_, _39646_, \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and (_03244_, _39658_, _37580_);
  nor (_39659_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  and (_39660_, _39659_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_39661_, _39660_, _37580_);
  and (_39662_, _03223_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or (_03246_, _39662_, _39661_);
  and (_39663_, _39636_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or (_39664_, _39663_, _39660_);
  and (_03248_, _39664_, _37580_);
  or (_39665_, _39660_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [15]);
  nand (_39666_, _39660_, _23871_);
  and (_39667_, _39666_, _37580_);
  and (_03250_, _39667_, _39665_);
  and (_03252_, _22666_, _35853_);
  or (_39668_, _38087_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  not (_39669_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nand (_39670_, _38087_, _39669_);
  and (_39671_, _39670_, _37580_);
  and (_03635_, _39671_, _39668_);
  or (_39672_, _38087_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  not (_39673_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nand (_39674_, _38087_, _39673_);
  and (_39675_, _39674_, _37580_);
  and (_03637_, _39675_, _39672_);
  or (_39676_, _38087_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  not (_39677_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nand (_39678_, _38087_, _39677_);
  and (_39679_, _39678_, _37580_);
  and (_03639_, _39679_, _39676_);
  or (_39680_, _38087_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  not (_39681_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nand (_39682_, _38087_, _39681_);
  and (_39683_, _39682_, _37580_);
  and (_03641_, _39683_, _39680_);
  or (_39684_, _38087_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  or (_39685_, _38088_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_39686_, _39685_, _37580_);
  and (_03643_, _39686_, _39684_);
  or (_39687_, _38087_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nand (_39688_, _38087_, _39044_);
  and (_39689_, _39688_, _37580_);
  and (_03645_, _39689_, _39687_);
  or (_39690_, _38087_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  not (_39691_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nand (_39692_, _38087_, _39691_);
  and (_39693_, _39692_, _37580_);
  and (_03647_, _39693_, _39690_);
  or (_39694_, _38087_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  or (_39695_, _38088_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_39696_, _39695_, _37580_);
  and (_03649_, _39696_, _39694_);
  or (_39697_, _38087_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  not (_39698_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nand (_39699_, _38087_, _39698_);
  and (_39700_, _39699_, _37580_);
  and (_03651_, _39700_, _39697_);
  or (_39701_, _38087_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nand (_39702_, _38087_, _39079_);
  and (_39703_, _39702_, _37580_);
  and (_03653_, _39703_, _39701_);
  or (_39704_, _38087_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nand (_39705_, _38087_, _39078_);
  and (_39706_, _39705_, _37580_);
  and (_03655_, _39706_, _39704_);
  or (_39707_, _38087_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nand (_39708_, _38087_, _39077_);
  and (_39709_, _39708_, _37580_);
  and (_03657_, _39709_, _39707_);
  or (_39710_, _38087_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  not (_39711_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nand (_39712_, _38087_, _39711_);
  and (_39713_, _39712_, _37580_);
  and (_03659_, _39713_, _39710_);
  or (_39714_, _38087_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  not (_39715_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nand (_39716_, _38087_, _39715_);
  and (_39717_, _39716_, _37580_);
  and (_03661_, _39717_, _39714_);
  or (_39718_, _38087_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nand (_39719_, _38087_, _39076_);
  and (_39720_, _39719_, _37580_);
  and (_03663_, _39720_, _39718_);
  and (_39721_, _38088_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_39722_, _38087_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  or (_39723_, _39722_, _39721_);
  and (_03695_, _39723_, _37580_);
  and (_39724_, _38088_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and (_39725_, _38087_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  or (_39726_, _39725_, _39724_);
  and (_03697_, _39726_, _37580_);
  and (_39727_, _38088_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and (_39728_, _38087_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or (_39729_, _39728_, _39727_);
  and (_03699_, _39729_, _37580_);
  and (_39730_, _38088_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and (_39731_, _38087_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or (_39732_, _39731_, _39730_);
  and (_03701_, _39732_, _37580_);
  and (_39733_, _38088_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  and (_39734_, _38087_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  or (_39735_, _39734_, _39733_);
  and (_03703_, _39735_, _37580_);
  and (_39736_, _38088_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  and (_39737_, _38087_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  or (_39738_, _39737_, _39736_);
  and (_03705_, _39738_, _37580_);
  and (_39739_, _38088_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  and (_39740_, _38087_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  or (_39741_, _39740_, _39739_);
  and (_03707_, _39741_, _37580_);
  and (_39742_, _38088_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  and (_39743_, _38087_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  or (_39744_, _39743_, _39742_);
  and (_03709_, _39744_, _37580_);
  and (_39745_, _38088_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  and (_39746_, _38087_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  or (_39747_, _39746_, _39745_);
  and (_03711_, _39747_, _37580_);
  and (_39748_, _38088_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  and (_39749_, _38087_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  or (_39750_, _39749_, _39748_);
  and (_03713_, _39750_, _37580_);
  and (_39751_, _38088_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  and (_39752_, _38087_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  or (_39753_, _39752_, _39751_);
  and (_03715_, _39753_, _37580_);
  and (_39754_, _38088_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  and (_39755_, _38087_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  or (_39756_, _39755_, _39754_);
  and (_03717_, _39756_, _37580_);
  and (_39757_, _38088_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  and (_39758_, _38087_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  or (_39760_, _39758_, _39757_);
  and (_03719_, _39760_, _37580_);
  and (_39761_, _38088_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  and (_39762_, _38087_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  or (_39763_, _39762_, _39761_);
  and (_03721_, _39763_, _37580_);
  and (_39764_, _38088_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  and (_39765_, _38087_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  or (_39766_, _39765_, _39764_);
  and (_03723_, _39766_, _37580_);
  and (_39768_, _39639_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_39769_, _39637_, \oc8051_top_1.oc8051_rom1.data_o [0]);
  or (_39770_, _39769_, _39768_);
  and (_05595_, _39770_, _37580_);
  and (_39771_, _39639_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_39772_, _39637_, \oc8051_top_1.oc8051_rom1.data_o [1]);
  or (_39773_, _39772_, _39771_);
  and (_05597_, _39773_, _37580_);
  and (_39774_, _39639_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_39775_, _39637_, \oc8051_top_1.oc8051_rom1.data_o [2]);
  or (_39777_, _39775_, _39774_);
  and (_05599_, _39777_, _37580_);
  and (_39778_, _39639_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_39779_, _39637_, \oc8051_top_1.oc8051_rom1.data_o [3]);
  or (_39780_, _39779_, _39778_);
  and (_05601_, _39780_, _37580_);
  and (_39781_, _39639_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_39782_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [4]);
  and (_39783_, _39782_, _39637_);
  or (_39784_, _39783_, _39781_);
  and (_05603_, _39784_, _37580_);
  and (_39786_, _39639_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_39787_, _39637_, \oc8051_top_1.oc8051_rom1.data_o [5]);
  or (_39788_, _39787_, _39786_);
  and (_05605_, _39788_, _37580_);
  and (_39789_, _39639_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_39790_, _39637_, \oc8051_top_1.oc8051_rom1.data_o [6]);
  or (_39791_, _39790_, _39789_);
  and (_05607_, _39791_, _37580_);
  and (_39792_, _39639_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_39794_, _39637_, \oc8051_top_1.oc8051_rom1.data_o [7]);
  or (_39795_, _39794_, _39792_);
  and (_05609_, _39795_, _37580_);
  and (_39796_, _39637_, \oc8051_top_1.oc8051_rom1.data_o [8]);
  and (_39797_, _39639_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  or (_39798_, _39797_, _39796_);
  and (_05611_, _39798_, _37580_);
  and (_39799_, _39637_, \oc8051_top_1.oc8051_rom1.data_o [9]);
  and (_39800_, _39639_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  or (_39801_, _39800_, _39799_);
  and (_05613_, _39801_, _37580_);
  and (_39803_, _39637_, \oc8051_top_1.oc8051_rom1.data_o [10]);
  and (_39804_, _39639_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  or (_39805_, _39804_, _39803_);
  and (_05615_, _39805_, _37580_);
  and (_39806_, _39637_, \oc8051_top_1.oc8051_rom1.data_o [11]);
  and (_39807_, _39639_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  or (_39808_, _39807_, _39806_);
  and (_05617_, _39808_, _37580_);
  and (_39809_, _39637_, \oc8051_top_1.oc8051_rom1.data_o [12]);
  and (_39811_, _39639_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  or (_39812_, _39811_, _39809_);
  and (_05619_, _39812_, _37580_);
  and (_39813_, _39637_, \oc8051_top_1.oc8051_rom1.data_o [13]);
  and (_39814_, _39639_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  or (_39815_, _39814_, _39813_);
  and (_05621_, _39815_, _37580_);
  and (_39816_, _39637_, \oc8051_top_1.oc8051_rom1.data_o [14]);
  and (_39817_, _39639_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  or (_39818_, _39817_, _39816_);
  and (_05623_, _39818_, _37580_);
  and (_39820_, _39637_, \oc8051_top_1.oc8051_rom1.data_o [15]);
  and (_39821_, _39639_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  or (_39822_, _39821_, _39820_);
  and (_05625_, _39822_, _37580_);
  and (_39823_, _39637_, \oc8051_top_1.oc8051_rom1.data_o [16]);
  and (_39824_, _39639_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  or (_39825_, _39824_, _39823_);
  and (_05627_, _39825_, _37580_);
  and (_39826_, _39637_, \oc8051_top_1.oc8051_rom1.data_o [17]);
  and (_39828_, _39639_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  or (_39829_, _39828_, _39826_);
  and (_05629_, _39829_, _37580_);
  and (_39830_, _39637_, \oc8051_top_1.oc8051_rom1.data_o [18]);
  and (_39831_, _39639_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  or (_39832_, _39831_, _39830_);
  and (_05631_, _39832_, _37580_);
  and (_39833_, _39637_, \oc8051_top_1.oc8051_rom1.data_o [19]);
  and (_39834_, _39639_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  or (_39835_, _39834_, _39833_);
  and (_05633_, _39835_, _37580_);
  and (_39837_, _39637_, \oc8051_top_1.oc8051_rom1.data_o [20]);
  and (_39838_, _39639_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  or (_39839_, _39838_, _39837_);
  and (_05635_, _39839_, _37580_);
  and (_39840_, _39637_, \oc8051_top_1.oc8051_rom1.data_o [21]);
  and (_39841_, _39639_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  or (_39842_, _39841_, _39840_);
  and (_05637_, _39842_, _37580_);
  and (_39843_, _39637_, \oc8051_top_1.oc8051_rom1.data_o [22]);
  and (_39845_, _39639_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  or (_39846_, _39845_, _39843_);
  and (_05639_, _39846_, _37580_);
  and (_39847_, _39637_, \oc8051_top_1.oc8051_rom1.data_o [23]);
  and (_39848_, _39639_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  or (_39849_, _39848_, _39847_);
  and (_05641_, _39849_, _37580_);
  and (_39850_, _39637_, \oc8051_top_1.oc8051_rom1.data_o [24]);
  and (_39851_, _39639_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  or (_39852_, _39851_, _39850_);
  and (_05643_, _39852_, _37580_);
  and (_39854_, _39637_, \oc8051_top_1.oc8051_rom1.data_o [25]);
  and (_39855_, _39639_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  or (_39856_, _39855_, _39854_);
  and (_05645_, _39856_, _37580_);
  and (_39857_, _39637_, \oc8051_top_1.oc8051_rom1.data_o [26]);
  and (_39858_, _39639_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  or (_39859_, _39858_, _39857_);
  and (_05647_, _39859_, _37580_);
  and (_39860_, _39637_, \oc8051_top_1.oc8051_rom1.data_o [27]);
  and (_39862_, _39639_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  or (_39863_, _39862_, _39860_);
  and (_05649_, _39863_, _37580_);
  and (_39864_, _39637_, \oc8051_top_1.oc8051_rom1.data_o [28]);
  and (_39865_, _39639_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  or (_39866_, _39865_, _39864_);
  and (_05651_, _39866_, _37580_);
  and (_39867_, _39637_, \oc8051_top_1.oc8051_rom1.data_o [29]);
  and (_39868_, _39639_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  or (_39869_, _39868_, _39867_);
  and (_05653_, _39869_, _37580_);
  and (_39871_, _39637_, \oc8051_top_1.oc8051_rom1.data_o [30]);
  and (_39872_, _39639_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  or (_39873_, _39872_, _39871_);
  and (_05655_, _39873_, _37580_);
  and (_05658_, _19724_, _37580_);
  and (_05661_, _19484_, _37580_);
  and (_05664_, _18957_, _37580_);
  nor (_05666_, _35856_, rst);
  nor (_05669_, _36043_, rst);
  nor (_05672_, _36193_, rst);
  nor (_05675_, _35957_, rst);
  nor (_05678_, _36006_, rst);
  nor (_05681_, _36129_, rst);
  nor (_05684_, _35941_, rst);
  nor (_05687_, _36104_, rst);
  and (_05717_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], _37580_);
  and (_05719_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _37580_);
  and (_05721_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], _37580_);
  and (_05723_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], _37580_);
  and (_05725_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _37580_);
  and (_05727_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], _37580_);
  and (_05729_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], _37580_);
  or (_39874_, _39030_, _39009_);
  and (_39875_, _39874_, ABINPUT[19]);
  nand (_39876_, _39015_, _37903_);
  or (_39877_, _39122_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nand (_39878_, _39877_, _39177_);
  or (_39879_, _39878_, _39123_);
  and (_39880_, _39042_, _36060_);
  and (_39881_, _39184_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nor (_39882_, _39881_, _39880_);
  and (_39883_, _39882_, _39879_);
  nand (_39884_, _39883_, _39876_);
  nor (_39885_, _39884_, _39875_);
  nand (_39886_, _39885_, _39006_);
  or (_39887_, _39006_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and (_39888_, _39887_, _37580_);
  and (_05731_, _39888_, _39886_);
  and (_39889_, _39874_, ABINPUT[20]);
  and (_39890_, _39042_, _36178_);
  and (_39891_, _39015_, _37920_);
  and (_39892_, _21457_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or (_39893_, _39892_, _39891_);
  or (_39894_, _39893_, _39890_);
  or (_39895_, _39894_, _39889_);
  nor (_39896_, _39126_, _39123_);
  nor (_39897_, _39896_, _39127_);
  and (_39898_, _39897_, _39177_);
  nor (_39899_, _39898_, _39895_);
  nand (_39900_, _39899_, _39006_);
  or (_39901_, _39006_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  and (_39902_, _39901_, _37580_);
  and (_05733_, _39902_, _39900_);
  and (_39903_, _39015_, _37937_);
  and (_39904_, _39874_, ABINPUT[21]);
  and (_39905_, _39042_, _35979_);
  and (_39906_, _39184_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  or (_39907_, _39906_, _39905_);
  or (_39908_, _39907_, _39904_);
  or (_39909_, _39133_, _39130_);
  not (_39910_, _39177_);
  nor (_39911_, _39910_, _39134_);
  and (_39912_, _39911_, _39909_);
  or (_39913_, _39912_, _39908_);
  or (_39914_, _39913_, _39903_);
  and (_39915_, _39914_, _39006_);
  not (_39916_, _39006_);
  not (_39917_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_39918_, _39194_, _39917_);
  and (_39919_, _39194_, _39917_);
  nor (_39920_, _39919_, _39918_);
  and (_39921_, _39920_, _39916_);
  or (_39922_, _39921_, _39915_);
  and (_05735_, _39922_, _37580_);
  and (_39923_, _39874_, ABINPUT[22]);
  and (_39924_, _39042_, _36023_);
  and (_39925_, _39015_, _37954_);
  and (_39926_, _21457_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  or (_39927_, _39926_, _39925_);
  or (_39928_, _39927_, _39924_);
  or (_39929_, _39928_, _39923_);
  or (_39930_, _39108_, _39106_);
  or (_39931_, _39930_, _39135_);
  nand (_39932_, _39930_, _39135_);
  and (_39933_, _39932_, _39931_);
  and (_39934_, _39933_, _39177_);
  or (_39935_, _39934_, _39929_);
  and (_39936_, _39935_, _39006_);
  and (_39937_, _39918_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_39938_, _39918_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_39939_, _39938_, _39937_);
  and (_39940_, _39939_, _39916_);
  or (_39941_, _39940_, _39936_);
  and (_05737_, _39941_, _37580_);
  or (_39942_, _39141_, _39138_);
  nor (_39943_, _39028_, _39034_);
  and (_39944_, _39943_, _39142_);
  and (_39945_, _39944_, _39942_);
  and (_39946_, _39874_, ABINPUT[23]);
  and (_39947_, _39042_, _36154_);
  and (_39948_, _39015_, _37971_);
  and (_39949_, _21457_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or (_39950_, _39949_, _39948_);
  or (_39951_, _39950_, _39947_);
  or (_39952_, _39951_, _39946_);
  or (_39953_, _39952_, _39945_);
  and (_39954_, _39953_, _39006_);
  and (_39955_, _39918_, _39197_);
  nor (_39956_, _39937_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or (_39957_, _39956_, _39955_);
  nor (_39958_, _39957_, _39006_);
  or (_39959_, _39958_, _39954_);
  and (_05739_, _39959_, _37580_);
  and (_39960_, _39874_, ABINPUT[24]);
  and (_39961_, _39042_, _35924_);
  and (_39962_, _39015_, _37988_);
  and (_39963_, _21457_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  or (_39964_, _39963_, _39962_);
  or (_39965_, _39964_, _39961_);
  or (_39966_, _39965_, _39960_);
  or (_39967_, _39096_, _39094_);
  or (_39968_, _39967_, _39144_);
  nand (_39969_, _39967_, _39144_);
  and (_39970_, _39969_, _39968_);
  and (_39971_, _39970_, _39177_);
  or (_39972_, _39971_, _39966_);
  and (_39973_, _39972_, _39006_);
  and (_39974_, _39955_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_39975_, _39955_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  or (_39976_, _39975_, _39974_);
  nor (_39977_, _39976_, _39006_);
  or (_39978_, _39977_, _39973_);
  and (_05741_, _39978_, _37580_);
  and (_39979_, _39015_, _38005_);
  and (_39980_, _39874_, ABINPUT[25]);
  and (_39981_, _39042_, _36091_);
  and (_39982_, _39184_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or (_39983_, _39982_, _39981_);
  or (_39984_, _39983_, _39980_);
  or (_39985_, _39146_, _39089_);
  nor (_39986_, _39910_, _39147_);
  and (_39987_, _39986_, _39985_);
  or (_39988_, _39987_, _39984_);
  or (_39989_, _39988_, _39979_);
  and (_39990_, _39989_, _39006_);
  and (_39991_, _39974_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor (_39992_, _39974_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or (_39993_, _39992_, _39991_);
  nor (_39994_, _39993_, _39006_);
  or (_39995_, _39994_, _39990_);
  and (_05743_, _39995_, _37580_);
  and (_39996_, _39874_, ABINPUT[26]);
  and (_39997_, _39042_, _35849_);
  and (_39998_, _39015_, _37886_);
  and (_39999_, _21457_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  or (_40000_, _39999_, _39998_);
  or (_40001_, _40000_, _39997_);
  or (_40002_, _40001_, _39996_);
  or (_40003_, _39080_, _39081_);
  nand (_40004_, _40003_, _39148_);
  or (_40005_, _40003_, _39148_);
  and (_40006_, _40005_, _40004_);
  and (_40007_, _40006_, _39177_);
  or (_40008_, _40007_, _40002_);
  and (_40009_, _40008_, _39006_);
  nor (_40010_, _39991_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  or (_40011_, _40010_, _39204_);
  nor (_40012_, _40011_, _39006_);
  or (_40013_, _40012_, _40009_);
  and (_05745_, _40013_, _37580_);
  and (_40014_, _39150_, _39698_);
  nor (_40015_, _39150_, _39698_);
  nor (_40016_, _40015_, _40014_);
  or (_40017_, _40016_, _39074_);
  nand (_40018_, _40016_, _39074_);
  and (_40019_, _40018_, _39943_);
  and (_40020_, _40019_, _40017_);
  and (_40021_, _39030_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_40022_, _39042_, _39336_);
  and (_40023_, _39015_, _36060_);
  and (_40024_, _39009_, ABINPUT[11]);
  and (_40025_, _21457_, ABINPUT[19]);
  or (_40026_, _40025_, _40024_);
  or (_40027_, _40026_, _40023_);
  or (_40028_, _40027_, _40022_);
  nor (_40029_, _40028_, _40021_);
  nand (_40030_, _40029_, _39006_);
  or (_40031_, _40030_, _40020_);
  nor (_40032_, _39204_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor (_40033_, _40032_, _39205_);
  or (_40034_, _40033_, _39006_);
  and (_40035_, _40034_, _37580_);
  and (_05747_, _40035_, _40031_);
  and (_40036_, _39150_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_40037_, _40036_, _39074_);
  and (_40038_, _39152_, _39073_);
  nor (_40039_, _40038_, _40037_);
  nand (_40040_, _40039_, _39079_);
  or (_40041_, _40039_, _39079_);
  and (_40042_, _40041_, _39943_);
  and (_40043_, _40042_, _40040_);
  and (_40044_, _39030_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and (_40045_, _39042_, _39327_);
  and (_40046_, _39015_, _36178_);
  and (_40047_, _39009_, ABINPUT[12]);
  and (_40048_, _21457_, ABINPUT[20]);
  or (_40049_, _40048_, _40047_);
  or (_40050_, _40049_, _40046_);
  or (_40051_, _40050_, _40045_);
  nor (_40052_, _40051_, _40044_);
  nand (_40053_, _40052_, _39006_);
  or (_40054_, _40053_, _40043_);
  nor (_40055_, _39205_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  nor (_40056_, _40055_, _39206_);
  or (_40057_, _40056_, _39006_);
  and (_40058_, _40057_, _37580_);
  and (_05749_, _40058_, _40054_);
  and (_40059_, _39153_, _39073_);
  and (_40060_, _40037_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor (_40061_, _40060_, _40059_);
  nand (_40062_, _40061_, _39078_);
  or (_40063_, _40061_, _39078_);
  and (_40064_, _40063_, _39943_);
  and (_40065_, _40064_, _40062_);
  and (_40066_, _39042_, _39366_);
  and (_40067_, _39030_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_40068_, _39015_, _35979_);
  and (_40069_, _39009_, ABINPUT[13]);
  and (_40070_, _21457_, ABINPUT[21]);
  or (_40071_, _40070_, _40069_);
  or (_40072_, _40071_, _40068_);
  or (_40073_, _40072_, _40067_);
  nor (_40074_, _40073_, _40066_);
  nand (_40075_, _40074_, _39006_);
  or (_40076_, _40075_, _40065_);
  nor (_40077_, _39206_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_40078_, _39206_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor (_40079_, _40078_, _40077_);
  or (_40080_, _40079_, _39006_);
  and (_40081_, _40080_, _37580_);
  and (_05751_, _40081_, _40076_);
  and (_40082_, _39043_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_40083_, _40082_, _39150_);
  and (_40084_, _40083_, _39074_);
  and (_40085_, _39154_, _39073_);
  nor (_40086_, _40085_, _40084_);
  nand (_40087_, _40086_, _39077_);
  or (_40088_, _40086_, _39077_);
  and (_40089_, _40088_, _39943_);
  and (_40090_, _40089_, _40087_);
  and (_40091_, _39030_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor (_40092_, _39054_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_40093_, _40092_, _39055_);
  and (_40094_, _40093_, _39042_);
  and (_40095_, _39015_, _36023_);
  and (_40096_, _39009_, ABINPUT[14]);
  and (_40097_, _21457_, ABINPUT[22]);
  or (_40098_, _40097_, _40096_);
  or (_40099_, _40098_, _40095_);
  or (_40100_, _40099_, _40094_);
  nor (_40101_, _40100_, _40091_);
  nand (_40102_, _40101_, _39006_);
  or (_40103_, _40102_, _40090_);
  nor (_40104_, _40078_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor (_40105_, _40104_, _39208_);
  or (_40106_, _40105_, _39006_);
  and (_40107_, _40106_, _37580_);
  and (_05753_, _40107_, _40103_);
  and (_40108_, _39165_, _39074_);
  and (_40109_, _39073_, _39077_);
  and (_40110_, _40109_, _39154_);
  nor (_40111_, _40110_, _40108_);
  nand (_40112_, _40111_, _39711_);
  or (_40113_, _40111_, _39711_);
  and (_40114_, _40113_, _39943_);
  and (_40115_, _40114_, _40112_);
  and (_40116_, _39051_, _39164_);
  and (_40117_, _40116_, _39711_);
  nor (_40118_, _40116_, _39711_);
  or (_40119_, _40118_, _40117_);
  and (_40120_, _40119_, _39042_);
  and (_40121_, _39030_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and (_40122_, _39015_, _36154_);
  and (_40123_, _39009_, ABINPUT[15]);
  and (_40124_, _21457_, ABINPUT[23]);
  or (_40125_, _40124_, _40123_);
  or (_40126_, _40125_, _40122_);
  or (_40127_, _40126_, _40121_);
  nor (_40128_, _40127_, _40120_);
  nand (_40129_, _40128_, _39006_);
  or (_40130_, _40129_, _40115_);
  nor (_40131_, _39208_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor (_40132_, _40131_, _39209_);
  or (_40133_, _40132_, _39006_);
  and (_40134_, _40133_, _37580_);
  and (_05755_, _40134_, _40130_);
  and (_40135_, _39166_, _39074_);
  and (_40136_, _40110_, _39711_);
  nor (_40137_, _40136_, _40135_);
  nor (_40138_, _40137_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_40139_, _40137_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  or (_40140_, _40139_, _40138_);
  and (_40141_, _40140_, _39943_);
  nor (_40142_, _39057_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_40143_, _40142_, _39058_);
  and (_40144_, _40143_, _39042_);
  and (_40145_, _39030_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and (_40146_, _39015_, _35924_);
  and (_40147_, _39009_, ABINPUT[16]);
  and (_40148_, _21457_, ABINPUT[24]);
  or (_40149_, _40148_, _40147_);
  or (_40150_, _40149_, _40146_);
  or (_40151_, _40150_, _40145_);
  or (_40152_, _40151_, _40144_);
  or (_40153_, _40152_, _40141_);
  or (_40154_, _40153_, _39916_);
  nor (_40155_, _39209_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor (_40156_, _40155_, _39211_);
  or (_40157_, _40156_, _39006_);
  and (_40158_, _40157_, _37580_);
  and (_05757_, _40158_, _40154_);
  nand (_40159_, _39015_, _36091_);
  nand (_40160_, _39184_, ABINPUT[25]);
  and (_40161_, _40160_, _40159_);
  nand (_40162_, _39030_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or (_40163_, _39058_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_40164_, _40163_, _39059_);
  nand (_40165_, _40164_, _39042_);
  nand (_40166_, _39009_, ABINPUT[17]);
  and (_40167_, _40166_, _40165_);
  and (_40168_, _40167_, _40162_);
  or (_40169_, _39168_, _39073_);
  or (_40170_, _39158_, _39074_);
  and (_40171_, _40170_, _40169_);
  nor (_40172_, _40171_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_40173_, _40171_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  or (_40174_, _40173_, _40172_);
  or (_40175_, _40174_, _39910_);
  and (_40176_, _40175_, _40168_);
  and (_40177_, _40176_, _40161_);
  nand (_40178_, _40177_, _39006_);
  nor (_40179_, _39211_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor (_40180_, _40179_, _39212_);
  or (_40181_, _40180_, _39006_);
  and (_40182_, _40181_, _37580_);
  and (_05759_, _40182_, _40178_);
  and (_40183_, _39571_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nor (_40191_, _39531_, _39528_);
  nor (_40198_, _40191_, _39532_);
  or (_40202_, _40198_, _39223_);
  or (_40208_, _39221_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_40216_, _40208_, _39568_);
  and (_40221_, _40216_, _40202_);
  or (_05761_, _40221_, _40183_);
  or (_40232_, _39534_, _39532_);
  and (_40239_, _40232_, _39535_);
  or (_40243_, _40239_, _39223_);
  or (_40249_, _39221_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_40257_, _40249_, _39568_);
  and (_40262_, _40257_, _40243_);
  and (_40266_, _39571_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or (_05763_, _40266_, _40262_);
  or (_40280_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _18520_);
  and (_40284_, _40280_, _37580_);
  or (_40290_, _39539_, _39537_);
  nor (_40298_, _39540_, _39223_);
  and (_40303_, _40298_, _40290_);
  nor (_40307_, _39221_, _39677_);
  or (_40315_, _40307_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_40322_, _40315_, _40303_);
  and (_05765_, _40322_, _40284_);
  and (_40331_, _39571_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_40339_, _39540_, _39315_);
  nor (_40344_, _40339_, _39541_);
  or (_40348_, _40344_, _39223_);
  or (_40356_, _39221_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_40357_, _40356_, _39568_);
  and (_40366_, _40357_, _40348_);
  or (_05767_, _40366_, _40331_);
  and (_40380_, _39571_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_40384_, _39544_, _39541_);
  nor (_40390_, _40384_, _39545_);
  or (_40398_, _40390_, _39223_);
  or (_40403_, _39221_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_40407_, _40403_, _39568_);
  and (_40408_, _40407_, _40398_);
  or (_05769_, _40408_, _40380_);
  and (_40409_, _39571_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_40410_, _39545_, _39309_);
  nor (_40411_, _40410_, _39546_);
  or (_40412_, _40411_, _39223_);
  or (_40413_, _39221_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_40414_, _40413_, _39568_);
  and (_40415_, _40414_, _40412_);
  or (_05771_, _40415_, _40409_);
  nor (_40416_, _39546_, _39303_);
  nor (_40417_, _40416_, _39547_);
  or (_40418_, _40417_, _39223_);
  or (_40419_, _39221_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_40420_, _40419_, _39568_);
  and (_40421_, _40420_, _40418_);
  and (_40422_, _39571_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or (_05773_, _40422_, _40421_);
  and (_40423_, _39571_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor (_40424_, _39547_, _39298_);
  nor (_40425_, _40424_, _39548_);
  or (_40426_, _40425_, _39223_);
  or (_40427_, _39221_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_40428_, _40427_, _39568_);
  and (_40429_, _40428_, _40426_);
  or (_05775_, _40429_, _40423_);
  nor (_40430_, _39550_, _39548_);
  nor (_40431_, _40430_, _39551_);
  or (_40432_, _40431_, _39223_);
  or (_40433_, _39221_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_40434_, _40433_, _39568_);
  and (_40435_, _40434_, _40432_);
  and (_40436_, _39571_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  or (_05777_, _40436_, _40435_);
  and (_40437_, _39571_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  nor (_40438_, _39551_, _39291_);
  nor (_40439_, _40438_, _39552_);
  or (_40440_, _40439_, _39223_);
  or (_40441_, _39221_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_40442_, _40441_, _39568_);
  and (_40443_, _40442_, _40440_);
  or (_05779_, _40443_, _40437_);
  nor (_40444_, _39552_, _39286_);
  nor (_40445_, _40444_, _39553_);
  or (_40446_, _40445_, _39223_);
  or (_40447_, _39221_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_40448_, _40447_, _39568_);
  and (_40449_, _40448_, _40446_);
  and (_40450_, _39571_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  or (_05781_, _40450_, _40449_);
  nor (_40451_, _39553_, _39283_);
  nor (_40452_, _40451_, _39554_);
  or (_40453_, _40452_, _39223_);
  or (_40454_, _39221_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_40455_, _40454_, _39568_);
  and (_40456_, _40455_, _40453_);
  and (_40457_, _39571_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  or (_05783_, _40457_, _40456_);
  nor (_40458_, _39554_, _39279_);
  nor (_40459_, _40458_, _39555_);
  or (_40460_, _40459_, _39223_);
  or (_40461_, _39221_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_40462_, _40461_, _39568_);
  and (_40463_, _40462_, _40460_);
  and (_40464_, _39571_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  or (_05785_, _40464_, _40463_);
  nor (_40465_, _39555_, _39276_);
  nor (_40466_, _40465_, _39556_);
  or (_40467_, _40466_, _39223_);
  or (_40468_, _39221_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_40469_, _40468_, _39568_);
  and (_40470_, _40469_, _40467_);
  and (_40471_, _39571_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or (_05787_, _40471_, _40470_);
  or (_40472_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14], _18520_);
  and (_40473_, _40472_, _37580_);
  or (_40474_, _39556_, _39272_);
  and (_40475_, _40474_, _39558_);
  nor (_40476_, _39221_, _39076_);
  or (_40477_, _40476_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_40478_, _40477_, _40475_);
  and (_05789_, _40478_, _40473_);
  and (_40479_, _39580_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  or (_40480_, _40479_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  and (_05791_, _40480_, _37580_);
  and (_40481_, _39580_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  or (_40482_, _40481_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and (_05793_, _40482_, _37580_);
  and (_40483_, _39580_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  or (_40484_, _40483_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  and (_05795_, _40484_, _37580_);
  and (_40485_, _39580_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  or (_40486_, _40485_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_05797_, _40486_, _37580_);
  and (_40487_, _39580_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  or (_40488_, _40487_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and (_05799_, _40488_, _37580_);
  and (_40489_, _39580_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  or (_40490_, _40489_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  and (_05801_, _40490_, _37580_);
  and (_40491_, _39580_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  or (_40492_, _40491_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  and (_05803_, _40492_, _37580_);
  nor (_40493_, _39527_, _35832_);
  or (_40494_, _40493_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nand (_40495_, _40493_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_40496_, _40495_, _39568_);
  and (_05805_, _40496_, _40494_);
  or (_40497_, _39592_, _39590_);
  and (_40498_, _40497_, _39593_);
  or (_40499_, _40498_, _35832_);
  or (_40500_, _18553_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_40501_, _40500_, _39568_);
  and (_05807_, _40501_, _40499_);
  and (_40502_, _39615_, \oc8051_top_1.oc8051_memory_interface1.cdata [0]);
  and (_40503_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [0]);
  and (_40504_, _40503_, _03223_);
  or (_05837_, _40504_, _40502_);
  and (_40505_, _39615_, \oc8051_top_1.oc8051_memory_interface1.cdata [1]);
  and (_40506_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [1]);
  and (_40507_, _40506_, _03223_);
  or (_05839_, _40507_, _40505_);
  and (_40508_, _39615_, \oc8051_top_1.oc8051_memory_interface1.cdata [2]);
  and (_40509_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [2]);
  and (_40510_, _40509_, _03223_);
  or (_05841_, _40510_, _40508_);
  and (_40511_, _39615_, \oc8051_top_1.oc8051_memory_interface1.cdata [3]);
  and (_40512_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [3]);
  and (_40513_, _40512_, _03223_);
  or (_05843_, _40513_, _40511_);
  and (_40514_, _39615_, \oc8051_top_1.oc8051_memory_interface1.cdata [4]);
  and (_40515_, _39782_, _03223_);
  or (_05845_, _40515_, _40514_);
  and (_40516_, _39615_, \oc8051_top_1.oc8051_memory_interface1.cdata [5]);
  and (_40517_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [5]);
  and (_40518_, _40517_, _03223_);
  or (_05847_, _40518_, _40516_);
  and (_40519_, _39615_, \oc8051_top_1.oc8051_memory_interface1.cdata [6]);
  and (_40520_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [6]);
  and (_40521_, _40520_, _03223_);
  or (_05849_, _40521_, _40519_);
  and (_05851_, _39623_, _37580_);
  nor (_05853_, _39633_, rst);
  and (_05855_, _39629_, _37580_);
  and (_40522_, _39637_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_40523_, _39639_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  or (_40524_, _40523_, _40522_);
  and (_05857_, _40524_, _37580_);
  and (_40525_, _39637_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_40526_, _39639_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  or (_40527_, _40526_, _40525_);
  and (_05859_, _40527_, _37580_);
  and (_40528_, _39637_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_40529_, _39639_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  or (_40530_, _40529_, _40528_);
  and (_05861_, _40530_, _37580_);
  and (_40531_, _39637_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_40532_, _39639_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  or (_40533_, _40532_, _40531_);
  and (_05863_, _40533_, _37580_);
  and (_40534_, _39637_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_40535_, _39639_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  or (_40536_, _40535_, _40534_);
  and (_05865_, _40536_, _37580_);
  and (_40537_, _39637_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_40538_, _39639_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  or (_40539_, _40538_, _40537_);
  and (_05867_, _40539_, _37580_);
  and (_40540_, _39637_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_40541_, _39639_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  or (_40542_, _40541_, _40540_);
  and (_05869_, _40542_, _37580_);
  and (_40543_, _39637_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_40544_, _39639_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  or (_40545_, _40544_, _40543_);
  and (_05871_, _40545_, _37580_);
  and (_40546_, _39637_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_40547_, _39639_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  or (_40548_, _40547_, _40546_);
  and (_05873_, _40548_, _37580_);
  and (_40549_, _39637_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_40550_, _39639_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  or (_40551_, _40550_, _40549_);
  and (_05875_, _40551_, _37580_);
  and (_40552_, _39637_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_40553_, _39639_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  or (_40554_, _40553_, _40552_);
  and (_05877_, _40554_, _37580_);
  and (_40555_, _39637_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_40556_, _39639_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  or (_40557_, _40556_, _40555_);
  and (_05879_, _40557_, _37580_);
  and (_40558_, _39637_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_40559_, _39639_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  or (_40560_, _40559_, _40558_);
  and (_05881_, _40560_, _37580_);
  and (_40561_, _39637_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_40562_, _39639_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  or (_40563_, _40562_, _40561_);
  and (_05883_, _40563_, _37580_);
  and (_40564_, _39637_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_40565_, _39639_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  or (_40566_, _40565_, _40564_);
  and (_05885_, _40566_, _37580_);
  and (_40567_, _39637_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_40568_, _39639_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  or (_40569_, _40568_, _40567_);
  and (_05887_, _40569_, _37580_);
  and (_40570_, _39637_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_40571_, _39639_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  or (_40572_, _40571_, _40570_);
  and (_05889_, _40572_, _37580_);
  and (_40573_, _39637_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_40574_, _39639_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  or (_40575_, _40574_, _40573_);
  and (_05891_, _40575_, _37580_);
  and (_40576_, _39637_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_40577_, _39639_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  or (_40578_, _40577_, _40576_);
  and (_05893_, _40578_, _37580_);
  and (_40579_, _39637_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_40580_, _39639_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  or (_40581_, _40580_, _40579_);
  and (_05895_, _40581_, _37580_);
  and (_40582_, _39637_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_40583_, _39639_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  or (_40584_, _40583_, _40582_);
  and (_05897_, _40584_, _37580_);
  and (_40585_, _39637_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_40586_, _39639_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  or (_40587_, _40586_, _40585_);
  and (_05899_, _40587_, _37580_);
  and (_40588_, _39637_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_40589_, _39639_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  or (_40590_, _40589_, _40588_);
  and (_05901_, _40590_, _37580_);
  and (_40591_, _39637_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_40592_, _39639_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  or (_40593_, _40592_, _40591_);
  and (_05903_, _40593_, _37580_);
  and (_40594_, _39637_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and (_40595_, _39639_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  or (_40596_, _40595_, _40594_);
  and (_05905_, _40596_, _37580_);
  and (_40597_, _39637_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and (_40598_, _39639_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  or (_40599_, _40598_, _40597_);
  and (_05907_, _40599_, _37580_);
  and (_40600_, _39637_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and (_40601_, _39639_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  or (_40602_, _40601_, _40600_);
  and (_05909_, _40602_, _37580_);
  and (_40603_, _39637_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and (_40604_, _39639_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  or (_40605_, _40604_, _40603_);
  and (_05911_, _40605_, _37580_);
  and (_40606_, _39637_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and (_40607_, _39639_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  or (_40608_, _40607_, _40606_);
  and (_05913_, _40608_, _37580_);
  and (_40609_, _39637_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and (_40610_, _39639_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  or (_40611_, _40610_, _40609_);
  and (_05915_, _40611_, _37580_);
  and (_40612_, _39637_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and (_40613_, _39639_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  or (_40614_, _40613_, _40612_);
  and (_05917_, _40614_, _37580_);
  and (_40615_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [0], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_40616_, _39647_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_40617_, _40616_, _40615_);
  and (_05919_, _40617_, _37580_);
  and (_40618_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [1], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_40619_, _39647_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_40620_, _40619_, _40618_);
  and (_05921_, _40620_, _37580_);
  and (_40621_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_40622_, _39647_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_40623_, _40622_, _40621_);
  and (_05923_, _40623_, _37580_);
  and (_40624_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [3], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_40625_, _39647_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_40626_, _40625_, _40624_);
  and (_05925_, _40626_, _37580_);
  and (_40627_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [4], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_40628_, _39647_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or (_40629_, _40628_, _40627_);
  and (_05927_, _40629_, _37580_);
  and (_40630_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [5], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_40631_, _39647_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or (_40632_, _40631_, _40630_);
  and (_05929_, _40632_, _37580_);
  and (_40633_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [6], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_40634_, _39647_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_40635_, _40634_, _40633_);
  and (_05931_, _40635_, _37580_);
  and (_40636_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_40637_, _36043_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_40638_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_40639_, _40638_, _39646_);
  and (_40640_, _40639_, _40637_);
  or (_40641_, _40640_, _40636_);
  and (_05933_, _40641_, _37580_);
  and (_40642_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_40643_, _36193_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_40644_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_40645_, _40644_, _39646_);
  and (_40646_, _40645_, _40643_);
  or (_40647_, _40646_, _40642_);
  and (_05935_, _40647_, _37580_);
  and (_40648_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_40649_, _35957_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_40650_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_40651_, _40650_, _39646_);
  and (_40652_, _40651_, _40649_);
  or (_40653_, _40652_, _40648_);
  and (_05937_, _40653_, _37580_);
  and (_40654_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_40655_, _36006_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_40656_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_40657_, _40656_, _39646_);
  and (_40658_, _40657_, _40655_);
  or (_40659_, _40658_, _40654_);
  and (_05939_, _40659_, _37580_);
  and (_40660_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_40661_, _36129_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_40662_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_40663_, _40662_, _39646_);
  and (_40664_, _40663_, _40661_);
  or (_40665_, _40664_, _40660_);
  and (_05941_, _40665_, _37580_);
  and (_40666_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_40667_, _35941_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_40668_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_40669_, _40668_, _39646_);
  and (_40670_, _40669_, _40667_);
  or (_40671_, _40670_, _40666_);
  and (_05943_, _40671_, _37580_);
  and (_40672_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_40673_, _36104_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_40674_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_40675_, _40674_, _39646_);
  and (_40676_, _40675_, _40673_);
  or (_40677_, _40676_, _40672_);
  and (_05945_, _40677_, _37580_);
  and (_40678_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_40679_, _35884_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_40680_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_40681_, _40680_, _39646_);
  and (_40682_, _40681_, _40679_);
  or (_40683_, _40682_, _40678_);
  and (_05947_, _40683_, _37580_);
  and (_40684_, _39653_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or (_40685_, _40684_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_40686_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8], _39646_);
  and (_40687_, _40686_, _37580_);
  and (_05949_, _40687_, _40685_);
  and (_40688_, _39653_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_40689_, _40688_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_40690_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9], _39646_);
  and (_40691_, _40690_, _37580_);
  and (_05951_, _40691_, _40689_);
  and (_40692_, _39653_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_40693_, _40692_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_40694_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10], _39646_);
  and (_40695_, _40694_, _37580_);
  and (_05953_, _40695_, _40693_);
  and (_40696_, _39653_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_40697_, _40696_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_40698_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11], _39646_);
  and (_40699_, _40698_, _37580_);
  and (_05955_, _40699_, _40697_);
  and (_40700_, _39653_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or (_40701_, _40700_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_40702_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12], _39646_);
  and (_40703_, _40702_, _37580_);
  and (_05957_, _40703_, _40701_);
  and (_40704_, _39653_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or (_40705_, _40704_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_40706_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13], _39646_);
  and (_40707_, _40706_, _37580_);
  and (_05959_, _40707_, _40705_);
  and (_40708_, _39653_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_40709_, _40708_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_40710_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14], _39646_);
  and (_40711_, _40710_, _37580_);
  and (_05961_, _40711_, _40709_);
  not (_40712_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  nor (_40713_, _39660_, _40712_);
  and (_40714_, _39660_, ABINPUT[19]);
  or (_40715_, _40714_, _40713_);
  and (_05963_, _40715_, _37580_);
  not (_40716_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1]);
  nor (_40717_, _39660_, _40716_);
  and (_40718_, _39660_, ABINPUT[20]);
  or (_40719_, _40718_, _40717_);
  and (_05965_, _40719_, _37580_);
  not (_40720_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2]);
  nor (_40721_, _39660_, _40720_);
  and (_40722_, _39660_, ABINPUT[21]);
  or (_40723_, _40722_, _40721_);
  and (_05967_, _40723_, _37580_);
  not (_40724_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3]);
  nor (_40725_, _39660_, _40724_);
  and (_40726_, _39660_, ABINPUT[22]);
  or (_40727_, _40726_, _40725_);
  and (_05969_, _40727_, _37580_);
  or (_40728_, _39660_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [4]);
  nand (_40729_, _39660_, _18054_);
  and (_40730_, _40729_, _37580_);
  and (_05971_, _40730_, _40728_);
  or (_40731_, _39660_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [5]);
  nand (_40732_, _39660_, _18228_);
  and (_40733_, _40732_, _37580_);
  and (_05973_, _40733_, _40731_);
  or (_40734_, _39660_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [6]);
  nand (_40735_, _39660_, _18401_);
  and (_40736_, _40735_, _37580_);
  and (_05975_, _40736_, _40734_);
  or (_40737_, _39660_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [7]);
  nand (_40738_, _39660_, _17122_);
  and (_40739_, _40738_, _37580_);
  and (_05977_, _40739_, _40737_);
  or (_40740_, _39660_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [8]);
  nand (_40741_, _39660_, _24043_);
  and (_40742_, _40741_, _37580_);
  and (_05979_, _40742_, _40740_);
  or (_40743_, _39660_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [9]);
  nand (_40744_, _39660_, _24129_);
  and (_40745_, _40744_, _37580_);
  and (_05981_, _40745_, _40743_);
  or (_40746_, _39660_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [10]);
  nand (_40747_, _39660_, _24215_);
  and (_40748_, _40747_, _37580_);
  and (_05983_, _40748_, _40746_);
  or (_40749_, _39660_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [11]);
  nand (_40750_, _39660_, _24301_);
  and (_40751_, _40750_, _37580_);
  and (_05985_, _40751_, _40749_);
  or (_40752_, _39660_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [12]);
  nand (_40753_, _39660_, _24387_);
  and (_40754_, _40753_, _37580_);
  and (_05987_, _40754_, _40752_);
  or (_40755_, _39660_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [13]);
  nand (_40756_, _39660_, _24473_);
  and (_40757_, _40756_, _37580_);
  and (_05989_, _40757_, _40755_);
  or (_40758_, _39660_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [14]);
  nand (_40759_, _39660_, _24559_);
  and (_40760_, _40759_, _37580_);
  and (_05991_, _40760_, _40758_);
  and (_08305_, _36211_, _37580_);
  and (_08308_, _36289_, _37580_);
  nor (_08314_, _35983_, rst);
  and (_08467_, _36311_, _37580_);
  and (_08469_, _36327_, _37580_);
  and (_08471_, _36342_, _37580_);
  and (_08473_, _36357_, _37580_);
  and (_08475_, _36371_, _37580_);
  and (_08477_, _36385_, _37580_);
  and (_08479_, _36399_, _37580_);
  nor (_08481_, _36064_, rst);
  nor (_08483_, _36197_, rst);
  nor (_12267_, _22633_, rst);
  nor (_40761_, _20792_, _19746_);
  nand (_40762_, _39609_, _20967_);
  or (_12269_, _40762_, _40761_);
  and (_40763_, _39367_, _19975_);
  and (_40764_, _40763_, _39374_);
  and (_40765_, _39395_, _39350_);
  and (_40766_, _40765_, _39320_);
  or (_40767_, _40766_, _40764_);
  or (_40768_, _39348_, _39319_);
  nand (_40769_, _40768_, _39339_);
  nand (_40770_, _40769_, _39360_);
  or (_40771_, _40770_, _40767_);
  and (_40772_, _39367_, _20694_);
  and (_40773_, _40772_, _39382_);
  or (_40774_, _40773_, _39465_);
  and (_40775_, _39382_, _39370_);
  and (_40776_, _39445_, _39320_);
  or (_40777_, _40776_, _40775_);
  or (_40778_, _40777_, _40774_);
  or (_40779_, _39500_, _39363_);
  and (_40780_, _39375_, _39324_);
  or (_40781_, _39487_, _40780_);
  or (_40782_, _40781_, _39519_);
  nor (_40783_, _40782_, _40779_);
  nand (_40784_, _40783_, _39453_);
  or (_40785_, _40784_, _40778_);
  or (_40786_, _40785_, _40771_);
  and (_40787_, _40786_, _18564_);
  not (_40788_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_40789_, _18542_, _15565_);
  and (_40790_, _40789_, _21468_);
  nor (_40791_, _40790_, _40788_);
  or (_40792_, _40791_, rst);
  or (_12272_, _40792_, _40787_);
  nand (_40793_, _20214_, _18498_);
  or (_40794_, _18498_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and (_40795_, _40794_, _37580_);
  and (_12275_, _40795_, _40793_);
  and (_40796_, \oc8051_top_1.oc8051_sfr1.wait_data , _37580_);
  and (_40797_, _40796_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  or (_40798_, _22424_, _21610_);
  and (_40799_, _21599_, _21196_);
  and (_40800_, _20792_, _20760_);
  or (_40801_, _40800_, _38964_);
  or (_40802_, _40801_, _40799_);
  or (_40803_, _40802_, _40798_);
  not (_40804_, _21940_);
  and (_40805_, _22523_, _22292_);
  and (_40806_, _21196_, _21130_);
  and (_40807_, _40806_, _20858_);
  or (_40808_, _40807_, _40805_);
  or (_40809_, _40808_, _40804_);
  or (_40810_, _40809_, _40803_);
  and (_40811_, _40810_, _39609_);
  or (_12277_, _40811_, _40797_);
  nor (_40812_, \oc8051_top_1.oc8051_decoder1.state [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_40813_, _40812_, \oc8051_top_1.oc8051_decoder1.state [0]);
  not (_40814_, _22556_);
  and (_40815_, _40814_, _40813_);
  and (_40816_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_40817_, _40816_, _40815_);
  and (_40818_, _21239_, _19746_);
  or (_40819_, _40818_, _21228_);
  and (_40820_, _38042_, _20749_);
  or (_40821_, _40820_, _21326_);
  or (_40822_, _40821_, _21852_);
  or (_40823_, _40822_, _40819_);
  and (_40824_, _40823_, _18553_);
  or (_40825_, _40824_, _40817_);
  and (_12280_, _40825_, _37580_);
  and (_40826_, _40796_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and (_40827_, _22523_, _21973_);
  or (_40828_, _21984_, _38972_);
  or (_40829_, _40828_, _40827_);
  and (_40830_, _21731_, _21841_);
  or (_40831_, _40830_, _40829_);
  or (_40832_, _38976_, _38053_);
  or (_40833_, _40832_, _40831_);
  and (_40834_, _22523_, _22116_);
  and (_40835_, _21294_, _21032_);
  or (_40836_, _40835_, _21348_);
  or (_40837_, _40819_, _40836_);
  or (_40838_, _40837_, _40834_);
  or (_40839_, _40838_, _40833_);
  and (_40840_, _40839_, _39609_);
  or (_12283_, _40840_, _40826_);
  and (_40841_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_40842_, _22094_, _18553_);
  or (_40843_, _40842_, _40841_);
  or (_40844_, _40843_, _40815_);
  and (_12285_, _40844_, _37580_);
  and (_40845_, _38986_, _19996_);
  and (_40846_, _38987_, _19996_);
  or (_40847_, _40846_, _40845_);
  or (_40848_, _40847_, _40807_);
  and (_40849_, _40848_, _22600_);
  not (_40850_, _22292_);
  or (_40851_, _40761_, _40850_);
  not (_40852_, _40806_);
  and (_40853_, _40852_, _40851_);
  not (_40854_, _40853_);
  and (_40855_, _40854_, _40813_);
  or (_40856_, _40855_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_40857_, _40847_, _21479_);
  or (_40858_, _40857_, _40856_);
  or (_40859_, _40858_, _40849_);
  or (_40860_, _15565_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_40861_, _40860_, _37580_);
  and (_12288_, _40861_, _40859_);
  and (_40862_, _40796_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  or (_40863_, _38972_, _21228_);
  and (_40864_, _21294_, _20803_);
  or (_40865_, _40830_, _40800_);
  or (_40866_, _40865_, _40864_);
  or (_40867_, _40866_, _40863_);
  or (_40868_, _40820_, _21863_);
  and (_40869_, _38039_, _21337_);
  or (_40870_, _40869_, _38051_);
  or (_40871_, _21731_, _21599_);
  and (_40872_, _40871_, _20890_);
  or (_40873_, _40872_, _40870_);
  or (_40874_, _40873_, _40868_);
  or (_40875_, _40874_, _40867_);
  and (_40876_, _40875_, _39609_);
  or (_12291_, _40876_, _40862_);
  and (_40877_, _40796_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and (_40878_, _20901_, _20738_);
  or (_40879_, _40878_, _21108_);
  and (_40880_, _20890_, _20760_);
  or (_40881_, _40880_, _40879_);
  and (_40882_, _22523_, _21698_);
  nor (_40883_, _40882_, _21786_);
  nand (_40884_, _40883_, _38055_);
  or (_40885_, _40884_, _40881_);
  and (_40886_, _21841_, _21097_);
  and (_40887_, _21196_, _20814_);
  and (_40888_, _38042_, _20738_);
  and (_40889_, _38043_, _20716_);
  or (_40890_, _40889_, _40888_);
  or (_40891_, _40890_, _40887_);
  or (_40892_, _40891_, _40886_);
  nor (_40893_, _21852_, _21566_);
  nand (_40894_, _40893_, _21720_);
  or (_40895_, _40894_, _40892_);
  or (_40896_, _40895_, _40831_);
  or (_40897_, _40896_, _40885_);
  and (_40898_, _40897_, _39609_);
  or (_12293_, _40898_, _40877_);
  and (_40899_, _21130_, _21032_);
  and (_40900_, _21841_, _20825_);
  or (_40901_, _40900_, _40899_);
  and (_40902_, _38039_, _21130_);
  or (_40903_, _40902_, _21054_);
  and (_40904_, _20825_, _19208_);
  or (_40905_, _40904_, _40903_);
  or (_40906_, _40905_, _40901_);
  and (_40907_, _21841_, _21239_);
  or (_40908_, _40907_, _40906_);
  and (_40909_, _40908_, _18553_);
  nor (_40910_, _22556_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_40911_, \oc8051_top_1.oc8051_sfr1.wait_data , \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or (_40912_, _40911_, _40910_);
  or (_40913_, _40912_, _40909_);
  and (_12296_, _40913_, _37580_);
  and (_40914_, _40830_, _19724_);
  or (_40915_, _40846_, _40828_);
  or (_40916_, _40915_, _40914_);
  or (_40917_, _22050_, _21863_);
  and (_40918_, _20956_, _19996_);
  and (_40919_, _40918_, _21687_);
  nor (_40920_, _40919_, _21775_);
  nand (_40921_, _40920_, _21621_);
  not (_40922_, _22281_);
  or (_40923_, _40922_, _22105_);
  or (_40924_, _40923_, _40921_);
  or (_40925_, _40924_, _40917_);
  or (_40926_, _40925_, _40916_);
  and (_40927_, _38039_, _20956_);
  or (_40928_, _40927_, _21995_);
  and (_40929_, _38042_, _21130_);
  or (_40930_, _40929_, _40845_);
  or (_40931_, _40930_, _40821_);
  or (_40932_, _40931_, _40928_);
  or (_40933_, _22215_, _21152_);
  and (_40934_, _40918_, _20890_);
  or (_40935_, _40934_, _21348_);
  or (_40936_, _40935_, _21951_);
  or (_40937_, _40936_, _38053_);
  or (_40938_, _40937_, _40933_);
  or (_40939_, _40938_, _40932_);
  or (_40940_, _40939_, _40926_);
  and (_40941_, _40940_, _18553_);
  and (_40942_, \oc8051_top_1.oc8051_decoder1.wr , \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_40943_, _22391_, _21479_);
  or (_40944_, _40857_, _40815_);
  or (_40945_, _40944_, _40943_);
  or (_40946_, _40945_, _40942_);
  or (_40947_, _40946_, _40941_);
  and (_12299_, _40947_, _37580_);
  nor (_12341_, _21523_, rst);
  nor (_12343_, _22468_, rst);
  not (_40948_, _39609_);
  or (_12345_, _40853_, _40948_);
  and (_40949_, _20967_, _19746_);
  nor (_40950_, _40949_, _40806_);
  or (_12348_, _40950_, _40948_);
  or (_40951_, _40773_, \oc8051_top_1.oc8051_decoder1.state [1]);
  or (_40952_, _40951_, _40776_);
  or (_40953_, _40952_, _40767_);
  and (_40954_, _40953_, _40790_);
  nor (_40955_, _40789_, _21468_);
  or (_40956_, _40955_, rst);
  or (_12351_, _40956_, _40954_);
  nand (_40957_, _19702_, _18498_);
  or (_40958_, _18498_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and (_40959_, _40958_, _37580_);
  and (_12353_, _40959_, _40957_);
  nand (_40960_, _19462_, _18498_);
  or (_40961_, _18498_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and (_40962_, _40961_, _37580_);
  and (_12356_, _40962_, _40960_);
  nand (_40963_, _18935_, _18498_);
  or (_40964_, _18498_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and (_40965_, _40964_, _37580_);
  and (_12359_, _40965_, _40963_);
  nand (_40966_, _19186_, _18498_);
  or (_40967_, _18498_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and (_40968_, _40967_, _37580_);
  and (_12362_, _40968_, _40966_);
  nand (_40969_, _19975_, _18498_);
  or (_40970_, _18498_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and (_40971_, _40970_, _37580_);
  and (_12365_, _40971_, _40969_);
  nand (_40972_, _20694_, _18498_);
  or (_40973_, _18498_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and (_40974_, _40973_, _37580_);
  and (_12367_, _40974_, _40972_);
  nand (_40975_, _20454_, _18498_);
  or (_40976_, _18498_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and (_40977_, _40976_, _37580_);
  and (_12370_, _40977_, _40975_);
  or (_40978_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], _15565_);
  and (_40979_, _40978_, _40856_);
  and (_40980_, _40979_, _37580_);
  and (_40981_, _22523_, _21742_);
  or (_40982_, _40981_, _40827_);
  and (_40983_, _20967_, _19996_);
  and (_40984_, _40983_, _22523_);
  and (_40985_, _22523_, _21250_);
  or (_40986_, _40985_, _40907_);
  or (_40987_, _40986_, _40984_);
  and (_40988_, _22160_, _20890_);
  or (_40989_, _40805_, _40988_);
  or (_40990_, _40887_, _40886_);
  or (_40991_, _40990_, _40989_);
  or (_40992_, _40991_, _40987_);
  or (_40993_, _40992_, _40982_);
  or (_40994_, _40904_, _38040_);
  and (_40995_, _21698_, _21841_);
  or (_40996_, _40995_, _40818_);
  or (_40997_, _40996_, _40903_);
  or (_40998_, _40997_, _40994_);
  or (_40999_, _21228_, _20988_);
  or (_41000_, _38047_, _22303_);
  or (_41001_, _41000_, _40999_);
  or (_41002_, _40900_, _40889_);
  and (_41003_, _40888_, _20912_);
  and (_41004_, _38042_, _20967_);
  or (_41005_, _41004_, _41003_);
  or (_41006_, _41005_, _41002_);
  or (_41007_, _21370_, _21108_);
  or (_41008_, _41007_, _41006_);
  or (_41009_, _41008_, _41001_);
  or (_41010_, _41009_, _40998_);
  or (_41011_, _41010_, _40993_);
  and (_41012_, _41011_, _39609_);
  or (_35781_, _41012_, _40980_);
  and (_41013_, _40796_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  and (_41014_, _22523_, _21097_);
  and (_41015_, _22523_, _22160_);
  or (_41016_, _40890_, _41015_);
  nor (_41017_, _41016_, _41014_);
  nand (_41018_, _41017_, _21874_);
  or (_41019_, _40881_, _40808_);
  or (_41020_, _41019_, _41018_);
  or (_41021_, _40900_, _21775_);
  or (_41022_, _41021_, _22270_);
  and (_41023_, _41022_, _20781_);
  or (_41024_, _40834_, _38977_);
  or (_41025_, _41024_, _40996_);
  or (_41026_, _41025_, _41023_);
  or (_41027_, _41026_, _41020_);
  and (_41028_, _41027_, _39609_);
  or (_35782_, _41028_, _41013_);
  or (_41029_, _40933_, _40930_);
  or (_41030_, _41029_, _40926_);
  and (_41031_, _41030_, _18553_);
  and (_41032_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_41033_, _41032_, _40945_);
  or (_41034_, _41033_, _41031_);
  and (_35783_, _41034_, _37580_);
  and (_41035_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_41036_, _22259_, _20858_);
  or (_41037_, _41036_, _21326_);
  or (_41038_, _41037_, _40936_);
  or (_41039_, _41038_, _40847_);
  and (_41040_, _41039_, _18553_);
  or (_41041_, _41040_, _41035_);
  or (_41042_, _41041_, _40944_);
  and (_35784_, _41042_, _37580_);
  nor (_41043_, _38988_, _20858_);
  or (_41044_, _41014_, _41043_);
  or (_41045_, _40994_, _40887_);
  and (_41046_, _21032_, _20956_);
  and (_41047_, _40983_, _21687_);
  or (_41048_, _41047_, _40985_);
  or (_41049_, _41048_, _41046_);
  or (_41050_, _41049_, _40882_);
  or (_41051_, _41050_, _41045_);
  or (_41052_, _41051_, _41044_);
  or (_41053_, _40903_, _21043_);
  and (_41054_, _21841_, _35890_);
  or (_41055_, _41054_, _40927_);
  and (_41056_, _22160_, _20803_);
  or (_41057_, _40899_, _38963_);
  or (_41058_, _41057_, _41056_);
  or (_41059_, _41058_, _41055_);
  or (_41060_, _41059_, _41053_);
  or (_41061_, _40984_, _40982_);
  or (_41062_, _40805_, _38973_);
  or (_41063_, _41062_, _22534_);
  or (_41064_, _41063_, _41061_);
  and (_41065_, _38967_, _21841_);
  or (_41066_, _40806_, _22545_);
  or (_41067_, _41066_, _41065_);
  and (_41068_, _22523_, _21599_);
  or (_41069_, _40907_, _41068_);
  or (_41070_, _41069_, _41067_);
  or (_41071_, _41070_, _41064_);
  or (_41072_, _41071_, _41060_);
  or (_41073_, _41072_, _41052_);
  and (_41074_, _41073_, _18553_);
  and (_41075_, \oc8051_top_1.oc8051_sfr1.wait_data , \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  or (_41076_, _40855_, _22611_);
  or (_41077_, _41076_, _41075_);
  or (_41078_, _41077_, _41074_);
  and (_35785_, _41078_, _37580_);
  or (_41079_, _40919_, _22215_);
  and (_41080_, _38039_, _20967_);
  and (_41081_, _40983_, _20890_);
  or (_41082_, _41081_, _41080_);
  or (_41083_, _41082_, _40818_);
  or (_41084_, _41083_, _41079_);
  or (_41085_, _41084_, _21272_);
  and (_41086_, _21698_, _21196_);
  and (_41087_, _21196_, _21097_);
  or (_41088_, _41087_, _41086_);
  or (_41089_, _22545_, _40899_);
  or (_41090_, _41089_, _41088_);
  or (_41091_, _41090_, _41053_);
  or (_41092_, _41069_, _22193_);
  or (_41093_, _41092_, _41045_);
  or (_41094_, _41093_, _41091_);
  or (_41095_, _41094_, _41085_);
  or (_41096_, _41095_, _41064_);
  and (_41097_, _41096_, _18553_);
  and (_41098_, \oc8051_top_1.oc8051_sfr1.wait_data , \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  or (_41099_, _41098_, _41076_);
  or (_41100_, _41099_, _41097_);
  and (_35786_, _41100_, _37580_);
  and (_41101_, _40796_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  and (_41102_, _21742_, _21196_);
  or (_41103_, _41102_, _40907_);
  or (_41104_, _40917_, _40873_);
  or (_41105_, _41104_, _41103_);
  not (_41106_, _35897_);
  or (_41107_, _40863_, _41106_);
  or (_41108_, _40902_, _40820_);
  and (_41109_, _22523_, _20760_);
  or (_41110_, _41109_, _40830_);
  or (_41111_, _41110_, _41108_);
  or (_41112_, _41111_, _41107_);
  and (_41113_, _21032_, _20825_);
  and (_41114_, _21196_, _21907_);
  or (_41115_, _41114_, _41113_);
  and (_41116_, _21305_, _21196_);
  or (_41117_, _21841_, _19208_);
  and (_41118_, _41117_, _21907_);
  or (_41119_, _41118_, _41116_);
  or (_41120_, _41119_, _41115_);
  nor (_41121_, _22083_, _21370_);
  nand (_41122_, _41121_, _35898_);
  or (_41123_, _41122_, _41120_);
  or (_41124_, _41123_, _41112_);
  or (_41125_, _41124_, _41105_);
  and (_41126_, _41125_, _39609_);
  or (_35787_, _41126_, _41101_);
  and (_41127_, _21731_, _21196_);
  and (_41128_, _40900_, _20858_);
  or (_41129_, _41128_, _40880_);
  nor (_41130_, _41129_, _41127_);
  nand (_41131_, _41130_, _40883_);
  or (_41132_, _41131_, _41067_);
  or (_41133_, _41109_, _41114_);
  or (_41134_, _40994_, _22237_);
  or (_41135_, _41134_, _41133_);
  or (_41136_, _21709_, _38963_);
  or (_41137_, _40878_, _21852_);
  or (_41138_, _41137_, _41136_);
  or (_41139_, _40888_, _35832_);
  or (_41140_, _41139_, _21228_);
  or (_41141_, _41140_, _21065_);
  or (_41142_, _41141_, _41138_);
  or (_41143_, _41142_, _41135_);
  or (_41144_, _41143_, _41132_);
  or (_41145_, _22545_, _22600_);
  or (_41146_, \oc8051_top_1.oc8051_decoder1.alu_op [0], _15565_);
  and (_41147_, _41146_, _37580_);
  and (_41148_, _41147_, _41145_);
  and (_35788_, _41148_, _41144_);
  and (_41149_, _21305_, _20792_);
  or (_41150_, _41149_, _40984_);
  or (_41151_, _41108_, _41062_);
  or (_41152_, _41151_, _41150_);
  or (_41153_, _22545_, _21852_);
  and (_41154_, _21196_, _20825_);
  or (_41155_, _41154_, _40907_);
  or (_41156_, _41155_, _41153_);
  or (_41157_, _21643_, \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_41158_, _41157_, _38041_);
  or (_41159_, _41158_, _41156_);
  nand (_41160_, _38049_, _21392_);
  or (_41161_, _41160_, _41159_);
  or (_41162_, _41161_, _41152_);
  or (_41163_, _41162_, _40833_);
  or (_41164_, \oc8051_top_1.oc8051_decoder1.alu_op [1], _15565_);
  and (_41165_, _41164_, _37580_);
  and (_41166_, _41165_, _41145_);
  and (_35789_, _41166_, _41163_);
  or (_41167_, _41110_, _38053_);
  or (_41168_, _41167_, _41150_);
  and (_41169_, _21337_, _21196_);
  nor (_41170_, _41169_, _21359_);
  nand (_41171_, _41170_, _35898_);
  or (_41172_, _38048_, _38041_);
  or (_41173_, _41172_, _41171_);
  or (_41174_, _40868_, _40829_);
  or (_41175_, _41174_, _41173_);
  or (_41176_, _41175_, _41168_);
  and (_41177_, _41176_, _18553_);
  and (_41178_, \oc8051_top_1.oc8051_decoder1.alu_op [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_41179_, _22534_, _15565_);
  or (_41180_, _41179_, _41178_);
  or (_41181_, _41180_, _41177_);
  and (_35790_, _41181_, _37580_);
  and (_41182_, _40796_, \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  nor (_41183_, _41133_, _38977_);
  nand (_41184_, _41183_, _35899_);
  or (_41185_, _38973_, _22061_);
  or (_41186_, _41116_, _40799_);
  or (_41187_, _41186_, _41185_);
  or (_41188_, _41187_, _40906_);
  or (_41189_, _41188_, _41103_);
  or (_41190_, _41189_, _41184_);
  and (_41191_, _41190_, _39609_);
  or (_35792_, _41191_, _41182_);
  not (_41192_, _37750_);
  nor (_41193_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  and (_41194_, _40712_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_41195_, _41194_, _41193_);
  nor (_41196_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  and (_41197_, _40716_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_41198_, _41197_, _41196_);
  nor (_41199_, _41198_, _41195_);
  not (_41200_, _41199_);
  nor (_41201_, _39920_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  and (_41202_, _40720_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_41203_, _41202_, _41201_);
  and (_41204_, _41203_, _41200_);
  nor (_41205_, _39939_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  and (_41206_, _40724_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_41207_, _41206_, _41205_);
  nor (_41208_, _41207_, _41204_);
  not (_41209_, _41198_);
  nor (_41210_, _41209_, _41195_);
  and (_41211_, _41210_, _41208_);
  and (_41212_, _41211_, _41192_);
  not (_41213_, _37832_);
  and (_41214_, _41208_, _41203_);
  and (_41215_, _41214_, _41213_);
  not (_41216_, _37791_);
  and (_41217_, _41198_, _41195_);
  and (_41218_, _41208_, _41217_);
  and (_41219_, _41218_, _41216_);
  or (_41220_, _41219_, _41215_);
  or (_41221_, _41220_, _41212_);
  not (_41222_, _37709_);
  and (_41223_, _41209_, _41195_);
  and (_41224_, _41223_, _41208_);
  and (_41225_, _41224_, _41222_);
  not (_41226_, _37583_);
  nor (_41227_, _41203_, _41200_);
  nor (_41228_, _41227_, _41204_);
  and (_41229_, _41207_, _41204_);
  nor (_41230_, _41229_, _41208_);
  nor (_41231_, _41230_, _41228_);
  and (_41232_, _41210_, _41231_);
  and (_41233_, _41232_, _41226_);
  or (_41234_, _41233_, _41225_);
  or (_41235_, _41234_, _41221_);
  not (_41236_, _37328_);
  and (_41237_, _41207_, _41228_);
  and (_41238_, _41237_, _41223_);
  and (_41239_, _41238_, _41236_);
  not (_41240_, _37448_);
  and (_41241_, _41237_, _41217_);
  and (_41242_, _41241_, _41240_);
  not (_41243_, _37489_);
  and (_41244_, _41237_, _41199_);
  and (_41245_, _41244_, _41243_);
  or (_41246_, _41245_, _41242_);
  or (_41247_, _41246_, _41239_);
  not (_41248_, _37407_);
  and (_41249_, _41237_, _41210_);
  and (_41250_, _41249_, _41248_);
  not (_41251_, _37048_);
  not (_41252_, _41228_);
  and (_41253_, _41230_, _41252_);
  and (_41254_, _41223_, _41253_);
  and (_00004_, _41254_, _41251_);
  or (_00005_, _00004_, _41250_);
  or (_00006_, _00005_, _41247_);
  or (_00007_, _00006_, _41235_);
  not (_00008_, _37089_);
  and (_00009_, _41253_, _41210_);
  and (_00010_, _00009_, _00008_);
  not (_00011_, _37130_);
  and (_00012_, _41253_, _41217_);
  and (_00013_, _00012_, _00011_);
  not (_00014_, _37198_);
  and (_00015_, _41207_, _41227_);
  and (_00016_, _00015_, _00014_);
  or (_00017_, _00016_, _00013_);
  or (_00018_, _00017_, _00010_);
  not (_00019_, _37532_);
  and (_00020_, _41223_, _41231_);
  and (_00021_, _00020_, _00019_);
  not (_00022_, _37627_);
  and (_00023_, _41231_, _41217_);
  and (_00024_, _00023_, _00022_);
  not (_00025_, _37668_);
  and (_00026_, _41231_, _41199_);
  and (_00027_, _00026_, _00025_);
  or (_00028_, _00027_, _00024_);
  or (_00029_, _00028_, _00021_);
  or (_00030_, _00029_, _00018_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [31], _00030_, _00007_);
  and (_00031_, _41224_, _00025_);
  and (_00032_, _00026_, _00022_);
  or (_00033_, _00032_, _00031_);
  and (_00034_, _00023_, _41226_);
  and (_00035_, _41232_, _00019_);
  or (_00036_, _00035_, _00034_);
  or (_00037_, _00036_, _00033_);
  and (_00038_, _41241_, _41248_);
  and (_00039_, _41244_, _41240_);
  and (_00040_, _41249_, _41236_);
  or (_00041_, _00040_, _00039_);
  or (_00043_, _00041_, _00038_);
  and (_00045_, _00020_, _41243_);
  and (_00047_, _00009_, _41251_);
  or (_00049_, _00047_, _00045_);
  or (_00051_, _00049_, _00043_);
  or (_00053_, _00051_, _00037_);
  and (_00055_, _41254_, _41213_);
  and (_00056_, _41214_, _41216_);
  and (_00057_, _41211_, _41222_);
  and (_00058_, _41218_, _41192_);
  or (_00059_, _00058_, _00057_);
  or (_00060_, _00059_, _00056_);
  or (_00061_, _00060_, _00055_);
  and (_00063_, _00012_, _00008_);
  and (_00064_, _41238_, _00014_);
  and (_00066_, _00015_, _00011_);
  or (_00067_, _00066_, _00064_);
  or (_00068_, _00067_, _00063_);
  or (_00069_, _00068_, _00061_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [23], _00069_, _00053_);
  and (_00070_, _00026_, _41226_);
  and (_00071_, _41211_, _00025_);
  and (_00072_, _41224_, _00022_);
  or (_00073_, _00072_, _00071_);
  or (_00074_, _00073_, _00070_);
  and (_00075_, _41218_, _41222_);
  and (_00076_, _00023_, _00019_);
  or (_00077_, _00076_, _00075_);
  or (_00078_, _00077_, _00074_);
  and (_00079_, _00020_, _41240_);
  and (_00080_, _41244_, _41248_);
  and (_00081_, _41241_, _41236_);
  or (_00082_, _00081_, _00080_);
  or (_00083_, _00082_, _00079_);
  and (_00084_, _41232_, _41243_);
  and (_00085_, _00012_, _41251_);
  or (_00086_, _00085_, _00084_);
  or (_00087_, _00086_, _00083_);
  or (_00088_, _00087_, _00078_);
  and (_00089_, _00015_, _00008_);
  and (_00090_, _41249_, _00014_);
  and (_00091_, _41238_, _00011_);
  or (_00092_, _00091_, _00090_);
  or (_00093_, _00092_, _00089_);
  and (_00095_, _41254_, _41216_);
  and (_00097_, _00009_, _41213_);
  and (_00099_, _41214_, _41192_);
  or (_00101_, _00099_, _00097_);
  or (_00103_, _00101_, _00095_);
  or (_00105_, _00103_, _00093_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [15], _00105_, _00088_);
  and (_00107_, _41254_, _41192_);
  and (_00108_, _41244_, _41236_);
  and (_00109_, _41232_, _41240_);
  and (_00110_, _00023_, _41243_);
  or (_00111_, _00110_, _00109_);
  or (_00112_, _00111_, _00108_);
  and (_00114_, _41238_, _00008_);
  and (_00115_, _41249_, _00011_);
  and (_00117_, _41241_, _00014_);
  or (_00118_, _00117_, _00115_);
  or (_00119_, _00118_, _00114_);
  and (_00120_, _00015_, _41251_);
  and (_00121_, _00020_, _41248_);
  or (_00122_, _00121_, _00120_);
  or (_00123_, _00122_, _00119_);
  or (_00124_, _00123_, _00112_);
  or (_00125_, _00124_, _00107_);
  and (_00126_, _00012_, _41213_);
  and (_00127_, _41214_, _41222_);
  or (_00128_, _00127_, _00126_);
  and (_00129_, _00009_, _41216_);
  and (_00130_, _00026_, _00019_);
  and (_00131_, _41224_, _41226_);
  and (_00132_, _41218_, _00025_);
  and (_00133_, _41211_, _00022_);
  or (_00134_, _00133_, _00132_);
  or (_00135_, _00134_, _00131_);
  or (_00136_, _00135_, _00130_);
  or (_00137_, _00136_, _00129_);
  or (_00138_, _00137_, _00128_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [7], _00138_, _00125_);
  not (_00139_, _37796_);
  and (_00140_, _41214_, _00139_);
  not (_00141_, _37755_);
  and (_00142_, _41218_, _00141_);
  not (_00143_, _37714_);
  and (_00144_, _41211_, _00143_);
  or (_00146_, _00144_, _00142_);
  or (_00148_, _00146_, _00140_);
  not (_00150_, _37537_);
  and (_00152_, _41232_, _00150_);
  not (_00154_, _37837_);
  and (_00156_, _41254_, _00154_);
  or (_00158_, _00156_, _00152_);
  or (_00159_, _00158_, _00148_);
  not (_00160_, _37212_);
  and (_00161_, _41238_, _00160_);
  not (_00162_, _37135_);
  and (_00163_, _00015_, _00162_);
  or (_00164_, _00163_, _00161_);
  not (_00166_, _37094_);
  and (_00167_, _00012_, _00166_);
  not (_00169_, _37053_);
  and (_00170_, _00009_, _00169_);
  or (_00171_, _00170_, _00167_);
  or (_00172_, _00171_, _00164_);
  or (_00173_, _00172_, _00159_);
  not (_00174_, _37495_);
  and (_00175_, _00020_, _00174_);
  not (_00176_, _37453_);
  and (_00177_, _41244_, _00176_);
  not (_00178_, _37412_);
  and (_00179_, _41241_, _00178_);
  not (_00180_, _37348_);
  and (_00181_, _41249_, _00180_);
  or (_00182_, _00181_, _00179_);
  or (_00183_, _00182_, _00177_);
  or (_00184_, _00183_, _00175_);
  not (_00185_, _37591_);
  and (_00186_, _00023_, _00185_);
  not (_00187_, _37673_);
  and (_00188_, _41224_, _00187_);
  not (_00189_, _37632_);
  and (_00190_, _00026_, _00189_);
  or (_00191_, _00190_, _00188_);
  or (_00192_, _00191_, _00186_);
  or (_00193_, _00192_, _00184_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [16], _00193_, _00173_);
  not (_00194_, _37801_);
  and (_00195_, _41214_, _00194_);
  not (_00196_, _37760_);
  and (_00198_, _41218_, _00196_);
  not (_00200_, _37719_);
  and (_00202_, _41211_, _00200_);
  or (_00204_, _00202_, _00198_);
  or (_00206_, _00204_, _00195_);
  not (_00208_, _37842_);
  and (_00210_, _41254_, _00208_);
  not (_00211_, _37542_);
  and (_00212_, _41232_, _00211_);
  or (_00213_, _00212_, _00210_);
  or (_00214_, _00213_, _00206_);
  not (_00215_, _37458_);
  and (_00216_, _41244_, _00215_);
  not (_00218_, _37417_);
  and (_00219_, _41241_, _00218_);
  not (_00221_, _37361_);
  and (_00222_, _41249_, _00221_);
  or (_00223_, _00222_, _00219_);
  or (_00224_, _00223_, _00216_);
  not (_00225_, _37099_);
  and (_00226_, _00012_, _00225_);
  not (_00227_, _37500_);
  and (_00228_, _00020_, _00227_);
  or (_00229_, _00228_, _00226_);
  or (_00230_, _00229_, _00224_);
  or (_00231_, _00230_, _00214_);
  not (_00232_, _37058_);
  and (_00233_, _00009_, _00232_);
  not (_00234_, _37231_);
  and (_00235_, _41238_, _00234_);
  not (_00236_, _37167_);
  and (_00237_, _00015_, _00236_);
  or (_00238_, _00237_, _00235_);
  or (_00239_, _00238_, _00233_);
  not (_00240_, _37596_);
  and (_00241_, _00023_, _00240_);
  not (_00242_, _37678_);
  and (_00243_, _41224_, _00242_);
  not (_00244_, _37637_);
  and (_00245_, _00026_, _00244_);
  or (_00246_, _00245_, _00243_);
  or (_00247_, _00246_, _00241_);
  or (_00248_, _00247_, _00239_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [17], _00248_, _00231_);
  not (_00250_, _37806_);
  and (_00252_, _41214_, _00250_);
  not (_00254_, _37765_);
  and (_00256_, _41218_, _00254_);
  not (_00258_, _37724_);
  and (_00260_, _41211_, _00258_);
  or (_00262_, _00260_, _00256_);
  or (_00263_, _00262_, _00252_);
  not (_00264_, _37548_);
  and (_00265_, _41232_, _00264_);
  not (_00266_, _37847_);
  and (_00267_, _41254_, _00266_);
  or (_00268_, _00267_, _00265_);
  or (_00270_, _00268_, _00263_);
  not (_00271_, _37463_);
  and (_00273_, _41244_, _00271_);
  not (_00274_, _37422_);
  and (_00275_, _41241_, _00274_);
  or (_00276_, _00275_, _00273_);
  not (_00277_, _37381_);
  and (_00278_, _41249_, _00277_);
  or (_00279_, _00278_, _00276_);
  not (_00280_, _37505_);
  and (_00281_, _00020_, _00280_);
  not (_00282_, _37104_);
  and (_00283_, _00012_, _00282_);
  or (_00284_, _00283_, _00281_);
  or (_00285_, _00284_, _00279_);
  or (_00286_, _00285_, _00270_);
  not (_00287_, _37063_);
  and (_00288_, _00009_, _00287_);
  not (_00289_, _37245_);
  and (_00290_, _41238_, _00289_);
  not (_00291_, _37172_);
  and (_00292_, _00015_, _00291_);
  or (_00293_, _00292_, _00290_);
  or (_00294_, _00293_, _00288_);
  not (_00295_, _37601_);
  and (_00296_, _00023_, _00295_);
  not (_00297_, _37683_);
  and (_00298_, _41224_, _00297_);
  not (_00299_, _37642_);
  and (_00300_, _00026_, _00299_);
  or (_00301_, _00300_, _00298_);
  or (_00303_, _00301_, _00296_);
  or (_00305_, _00303_, _00294_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [18], _00305_, _00286_);
  not (_00308_, _37811_);
  and (_00310_, _41214_, _00308_);
  not (_00312_, _37770_);
  and (_00314_, _41218_, _00312_);
  not (_00315_, _37729_);
  and (_00316_, _41211_, _00315_);
  or (_00317_, _00316_, _00314_);
  or (_00318_, _00317_, _00310_);
  not (_00319_, _37555_);
  and (_00320_, _41232_, _00319_);
  not (_00322_, _37852_);
  and (_00323_, _41254_, _00322_);
  or (_00325_, _00323_, _00320_);
  or (_00326_, _00325_, _00318_);
  not (_00327_, _37468_);
  and (_00328_, _41244_, _00327_);
  not (_00329_, _37427_);
  and (_00330_, _41241_, _00329_);
  or (_00331_, _00330_, _00328_);
  not (_00332_, _37386_);
  and (_00333_, _41249_, _00332_);
  or (_00334_, _00333_, _00331_);
  not (_00335_, _37510_);
  and (_00336_, _00020_, _00335_);
  not (_00337_, _37109_);
  and (_00338_, _00012_, _00337_);
  or (_00339_, _00338_, _00336_);
  or (_00340_, _00339_, _00334_);
  or (_00341_, _00340_, _00326_);
  not (_00342_, _37068_);
  and (_00343_, _00009_, _00342_);
  not (_00344_, _37260_);
  and (_00345_, _41238_, _00344_);
  not (_00346_, _37177_);
  and (_00347_, _00015_, _00346_);
  or (_00348_, _00347_, _00345_);
  or (_00349_, _00348_, _00343_);
  not (_00350_, _37606_);
  and (_00351_, _00023_, _00350_);
  not (_00352_, _37688_);
  and (_00353_, _41224_, _00352_);
  not (_00355_, _37647_);
  and (_00357_, _00026_, _00355_);
  or (_00359_, _00357_, _00353_);
  or (_00361_, _00359_, _00351_);
  or (_00363_, _00361_, _00349_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [19], _00363_, _00341_);
  not (_00366_, _37611_);
  and (_00367_, _00023_, _00366_);
  not (_00368_, _37560_);
  and (_00369_, _41232_, _00368_);
  or (_00370_, _00369_, _00367_);
  not (_00371_, _37693_);
  and (_00372_, _41224_, _00371_);
  not (_00374_, _37652_);
  and (_00375_, _00026_, _00374_);
  or (_00377_, _00375_, _00372_);
  or (_00378_, _00377_, _00370_);
  not (_00379_, _37473_);
  and (_00380_, _41244_, _00379_);
  not (_00381_, _37432_);
  and (_00382_, _41241_, _00381_);
  not (_00383_, _37391_);
  and (_00384_, _41249_, _00383_);
  or (_00385_, _00384_, _00382_);
  or (_00386_, _00385_, _00380_);
  not (_00387_, _37515_);
  and (_00388_, _00020_, _00387_);
  not (_00389_, _37073_);
  and (_00390_, _00009_, _00389_);
  or (_00391_, _00390_, _00388_);
  or (_00392_, _00391_, _00386_);
  or (_00393_, _00392_, _00378_);
  not (_00394_, _37857_);
  and (_00395_, _41254_, _00394_);
  not (_00396_, _37816_);
  and (_00397_, _41214_, _00396_);
  not (_00398_, _37775_);
  and (_00399_, _41218_, _00398_);
  not (_00400_, _37734_);
  and (_00401_, _41211_, _00400_);
  or (_00402_, _00401_, _00399_);
  or (_00403_, _00402_, _00397_);
  or (_00404_, _00403_, _00395_);
  not (_00405_, _37114_);
  and (_00407_, _00012_, _00405_);
  not (_00409_, _37279_);
  and (_00411_, _41238_, _00409_);
  not (_00413_, _37182_);
  and (_00415_, _00015_, _00413_);
  or (_00417_, _00415_, _00411_);
  or (_00419_, _00417_, _00407_);
  or (_00420_, _00419_, _00404_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [20], _00420_, _00393_);
  not (_00421_, _37821_);
  and (_00422_, _41214_, _00421_);
  not (_00423_, _37780_);
  and (_00424_, _41218_, _00423_);
  not (_00426_, _37739_);
  and (_00427_, _41211_, _00426_);
  or (_00429_, _00427_, _00424_);
  or (_00430_, _00429_, _00422_);
  not (_00431_, _37862_);
  and (_00432_, _41254_, _00431_);
  not (_00433_, _37565_);
  and (_00434_, _41232_, _00433_);
  or (_00435_, _00434_, _00432_);
  or (_00436_, _00435_, _00430_);
  not (_00437_, _37478_);
  and (_00438_, _41244_, _00437_);
  not (_00439_, _37437_);
  and (_00440_, _41241_, _00439_);
  not (_00441_, _37396_);
  and (_00442_, _41249_, _00441_);
  or (_00443_, _00442_, _00440_);
  or (_00444_, _00443_, _00438_);
  not (_00445_, _37119_);
  and (_00446_, _00012_, _00445_);
  not (_00447_, _37520_);
  and (_00448_, _00020_, _00447_);
  or (_00449_, _00448_, _00446_);
  or (_00450_, _00449_, _00444_);
  or (_00451_, _00450_, _00436_);
  not (_00452_, _37078_);
  and (_00453_, _00009_, _00452_);
  not (_00454_, _37292_);
  and (_00455_, _41238_, _00454_);
  not (_00456_, _37187_);
  and (_00457_, _00015_, _00456_);
  or (_00459_, _00457_, _00455_);
  or (_00461_, _00459_, _00453_);
  not (_00463_, _37616_);
  and (_00465_, _00023_, _00463_);
  not (_00467_, _37698_);
  and (_00469_, _41224_, _00467_);
  not (_00471_, _37657_);
  and (_00472_, _00026_, _00471_);
  or (_00473_, _00472_, _00469_);
  or (_00474_, _00473_, _00465_);
  or (_00475_, _00474_, _00461_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [21], _00475_, _00451_);
  not (_00476_, _37826_);
  and (_00478_, _41214_, _00476_);
  not (_00479_, _37785_);
  and (_00481_, _41218_, _00479_);
  not (_00482_, _37744_);
  and (_00483_, _41211_, _00482_);
  or (_00484_, _00483_, _00481_);
  or (_00485_, _00484_, _00478_);
  not (_00486_, _37867_);
  and (_00487_, _41254_, _00486_);
  not (_00488_, _37570_);
  and (_00489_, _41232_, _00488_);
  or (_00490_, _00489_, _00487_);
  or (_00491_, _00490_, _00485_);
  not (_00492_, _37483_);
  and (_00493_, _41244_, _00492_);
  not (_00494_, _37442_);
  and (_00495_, _41241_, _00494_);
  not (_00496_, _37401_);
  and (_00497_, _41249_, _00496_);
  or (_00498_, _00497_, _00495_);
  or (_00499_, _00498_, _00493_);
  not (_00500_, _37124_);
  and (_00501_, _00012_, _00500_);
  not (_00502_, _37525_);
  and (_00503_, _00020_, _00502_);
  or (_00504_, _00503_, _00501_);
  or (_00505_, _00504_, _00499_);
  or (_00506_, _00505_, _00491_);
  not (_00507_, _37083_);
  and (_00508_, _00009_, _00507_);
  not (_00509_, _37312_);
  and (_00511_, _41238_, _00509_);
  not (_00513_, _37192_);
  and (_00515_, _00015_, _00513_);
  or (_00517_, _00515_, _00511_);
  or (_00519_, _00517_, _00508_);
  not (_00521_, _37621_);
  and (_00523_, _00023_, _00521_);
  not (_00524_, _37703_);
  and (_00525_, _41224_, _00524_);
  not (_00526_, _37662_);
  and (_00527_, _00026_, _00526_);
  or (_00528_, _00527_, _00525_);
  or (_00529_, _00528_, _00523_);
  or (_00531_, _00529_, _00519_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [22], _00531_, _00506_);
  and (_00533_, _41214_, _00154_);
  and (_00534_, _41211_, _00141_);
  and (_00535_, _41218_, _00139_);
  or (_00536_, _00535_, _00534_);
  or (_00537_, _00536_, _00533_);
  and (_00538_, _41224_, _00143_);
  and (_00539_, _00020_, _00150_);
  or (_00540_, _00539_, _00538_);
  or (_00541_, _00540_, _00537_);
  and (_00542_, _41249_, _00178_);
  and (_00543_, _41241_, _00176_);
  and (_00544_, _41244_, _00174_);
  or (_00545_, _00544_, _00543_);
  or (_00546_, _00545_, _00542_);
  and (_00547_, _00009_, _00166_);
  and (_00548_, _41238_, _00180_);
  or (_00549_, _00548_, _00547_);
  or (_00550_, _00549_, _00546_);
  or (_00551_, _00550_, _00541_);
  and (_00552_, _41254_, _00169_);
  and (_00553_, _00015_, _00160_);
  and (_00554_, _00012_, _00162_);
  or (_00555_, _00554_, _00553_);
  or (_00556_, _00555_, _00552_);
  and (_00557_, _41232_, _00185_);
  and (_00558_, _00023_, _00189_);
  and (_00559_, _00026_, _00187_);
  or (_00560_, _00559_, _00558_);
  or (_00561_, _00560_, _00557_);
  or (_00563_, _00561_, _00556_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [24], _00563_, _00551_);
  and (_00566_, _41214_, _00208_);
  and (_00568_, _41211_, _00196_);
  and (_00570_, _41218_, _00194_);
  or (_00572_, _00570_, _00568_);
  or (_00574_, _00572_, _00566_);
  and (_00575_, _41224_, _00200_);
  and (_00576_, _00020_, _00211_);
  or (_00577_, _00576_, _00575_);
  or (_00578_, _00577_, _00574_);
  and (_00579_, _41249_, _00218_);
  and (_00580_, _41241_, _00215_);
  and (_00582_, _41244_, _00227_);
  or (_00583_, _00582_, _00580_);
  or (_00585_, _00583_, _00579_);
  and (_00586_, _00009_, _00225_);
  and (_00587_, _41238_, _00221_);
  or (_00588_, _00587_, _00586_);
  or (_00589_, _00588_, _00585_);
  or (_00590_, _00589_, _00578_);
  and (_00591_, _41254_, _00232_);
  and (_00592_, _00015_, _00234_);
  and (_00593_, _00012_, _00236_);
  or (_00594_, _00593_, _00592_);
  or (_00595_, _00594_, _00591_);
  and (_00596_, _41232_, _00240_);
  and (_00597_, _00023_, _00244_);
  and (_00598_, _00026_, _00242_);
  or (_00599_, _00598_, _00597_);
  or (_00600_, _00599_, _00596_);
  or (_00601_, _00600_, _00595_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [25], _00601_, _00590_);
  and (_00602_, _41214_, _00266_);
  and (_00603_, _41211_, _00254_);
  and (_00604_, _41218_, _00250_);
  or (_00605_, _00604_, _00603_);
  or (_00606_, _00605_, _00602_);
  and (_00607_, _41224_, _00258_);
  and (_00608_, _41232_, _00295_);
  or (_00609_, _00608_, _00607_);
  or (_00610_, _00609_, _00606_);
  and (_00611_, _41249_, _00274_);
  and (_00612_, _41241_, _00271_);
  and (_00614_, _41244_, _00280_);
  or (_00616_, _00614_, _00612_);
  or (_00618_, _00616_, _00611_);
  and (_00620_, _00009_, _00282_);
  and (_00622_, _41238_, _00277_);
  or (_00624_, _00622_, _00620_);
  or (_00626_, _00624_, _00618_);
  or (_00627_, _00626_, _00610_);
  and (_00628_, _41254_, _00287_);
  and (_00629_, _00015_, _00289_);
  and (_00630_, _00012_, _00291_);
  or (_00631_, _00630_, _00629_);
  or (_00632_, _00631_, _00628_);
  and (_00634_, _00020_, _00264_);
  and (_00635_, _00023_, _00299_);
  and (_00637_, _00026_, _00297_);
  or (_00638_, _00637_, _00635_);
  or (_00639_, _00638_, _00634_);
  or (_00640_, _00639_, _00632_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [26], _00640_, _00627_);
  and (_00641_, _00023_, _00355_);
  and (_00642_, _00026_, _00352_);
  or (_00643_, _00642_, _00641_);
  and (_00644_, _00020_, _00319_);
  and (_00645_, _41232_, _00350_);
  or (_00646_, _00645_, _00644_);
  or (_00647_, _00646_, _00643_);
  and (_00648_, _00012_, _00346_);
  and (_00649_, _00015_, _00344_);
  or (_00650_, _00649_, _00648_);
  and (_00651_, _41254_, _00342_);
  and (_00652_, _00009_, _00337_);
  or (_00653_, _00652_, _00651_);
  or (_00654_, _00653_, _00650_);
  or (_00655_, _00654_, _00647_);
  and (_00656_, _41238_, _00332_);
  and (_00657_, _41249_, _00329_);
  and (_00658_, _41241_, _00327_);
  and (_00659_, _41244_, _00335_);
  or (_00660_, _00659_, _00658_);
  or (_00661_, _00660_, _00657_);
  or (_00662_, _00661_, _00656_);
  and (_00663_, _41211_, _00312_);
  and (_00664_, _41224_, _00315_);
  and (_00666_, _41214_, _00322_);
  and (_00668_, _41218_, _00308_);
  or (_00670_, _00668_, _00666_);
  or (_00672_, _00670_, _00664_);
  or (_00674_, _00672_, _00663_);
  or (_00676_, _00674_, _00662_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [27], _00676_, _00655_);
  and (_00678_, _00023_, _00374_);
  and (_00679_, _00026_, _00371_);
  or (_00680_, _00679_, _00678_);
  and (_00681_, _00020_, _00368_);
  and (_00682_, _41232_, _00366_);
  or (_00683_, _00682_, _00681_);
  or (_00685_, _00683_, _00680_);
  and (_00686_, _00012_, _00413_);
  and (_00688_, _00015_, _00409_);
  or (_00689_, _00688_, _00686_);
  and (_00690_, _41254_, _00389_);
  and (_00691_, _00009_, _00405_);
  or (_00692_, _00691_, _00690_);
  or (_00693_, _00692_, _00689_);
  or (_00694_, _00693_, _00685_);
  and (_00695_, _41249_, _00381_);
  and (_00696_, _41238_, _00383_);
  and (_00697_, _41241_, _00379_);
  and (_00698_, _41244_, _00387_);
  or (_00699_, _00698_, _00697_);
  or (_00700_, _00699_, _00696_);
  or (_00701_, _00700_, _00695_);
  and (_00702_, _41224_, _00400_);
  and (_00703_, _41211_, _00398_);
  and (_00704_, _41214_, _00394_);
  and (_00705_, _41218_, _00396_);
  or (_00706_, _00705_, _00704_);
  or (_00707_, _00706_, _00703_);
  or (_00708_, _00707_, _00702_);
  or (_00709_, _00708_, _00701_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [28], _00709_, _00694_);
  and (_00710_, _00023_, _00471_);
  and (_00711_, _00026_, _00467_);
  or (_00712_, _00711_, _00710_);
  and (_00713_, _00020_, _00433_);
  and (_00714_, _41232_, _00463_);
  or (_00715_, _00714_, _00713_);
  or (_00717_, _00715_, _00712_);
  and (_00719_, _41238_, _00441_);
  and (_00721_, _41244_, _00447_);
  and (_00723_, _41241_, _00437_);
  or (_00725_, _00723_, _00721_);
  or (_00727_, _00725_, _00719_);
  and (_00729_, _41249_, _00439_);
  and (_00730_, _00009_, _00445_);
  or (_00731_, _00730_, _00729_);
  or (_00732_, _00731_, _00727_);
  or (_00733_, _00732_, _00717_);
  and (_00734_, _41211_, _00423_);
  and (_00735_, _41224_, _00426_);
  and (_00737_, _41214_, _00431_);
  and (_00738_, _41218_, _00421_);
  or (_00740_, _00738_, _00737_);
  or (_00741_, _00740_, _00735_);
  or (_00742_, _00741_, _00734_);
  and (_00743_, _41254_, _00452_);
  and (_00744_, _00012_, _00456_);
  and (_00745_, _00015_, _00454_);
  or (_00746_, _00745_, _00744_);
  or (_00747_, _00746_, _00743_);
  or (_00748_, _00747_, _00742_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [29], _00748_, _00733_);
  and (_00749_, _41224_, _00482_);
  and (_00750_, _41214_, _00486_);
  and (_00751_, _41218_, _00476_);
  or (_00752_, _00751_, _00750_);
  or (_00753_, _00752_, _00749_);
  and (_00754_, _41211_, _00479_);
  and (_00755_, _41232_, _00521_);
  or (_00756_, _00755_, _00754_);
  or (_00757_, _00756_, _00753_);
  and (_00758_, _00015_, _00509_);
  and (_00759_, _00012_, _00513_);
  or (_00760_, _00759_, _00758_);
  and (_00761_, _00009_, _00500_);
  and (_00762_, _41254_, _00507_);
  or (_00763_, _00762_, _00761_);
  or (_00764_, _00763_, _00760_);
  or (_00765_, _00764_, _00757_);
  and (_00766_, _41238_, _00496_);
  and (_00767_, _41249_, _00494_);
  and (_00769_, _41244_, _00502_);
  and (_00771_, _41241_, _00492_);
  or (_00773_, _00771_, _00769_);
  or (_00775_, _00773_, _00767_);
  or (_00777_, _00775_, _00766_);
  and (_00779_, _00020_, _00488_);
  and (_00781_, _00023_, _00526_);
  and (_00782_, _00026_, _00524_);
  or (_00783_, _00782_, _00781_);
  or (_00784_, _00783_, _00779_);
  or (_00785_, _00784_, _00777_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [30], _00785_, _00765_);
  and (_00786_, _41224_, _00185_);
  and (_00788_, _41218_, _00187_);
  and (_00789_, _41211_, _00189_);
  or (_00791_, _00789_, _00788_);
  or (_00792_, _00791_, _00786_);
  and (_00793_, _00026_, _00150_);
  and (_00794_, _41254_, _00141_);
  or (_00795_, _00794_, _00793_);
  or (_00796_, _00795_, _00792_);
  and (_00797_, _00015_, _00169_);
  and (_00798_, _41241_, _00160_);
  and (_00799_, _41249_, _00162_);
  or (_00800_, _00799_, _00798_);
  or (_00801_, _00800_, _00797_);
  and (_00802_, _41244_, _00180_);
  and (_00803_, _41238_, _00166_);
  or (_00804_, _00803_, _00802_);
  or (_00805_, _00804_, _00801_);
  or (_00806_, _00805_, _00796_);
  and (_00807_, _00020_, _00178_);
  and (_00808_, _00023_, _00174_);
  and (_00809_, _41232_, _00176_);
  or (_00810_, _00809_, _00808_);
  or (_00811_, _00810_, _00807_);
  and (_00812_, _00009_, _00139_);
  and (_00813_, _00012_, _00154_);
  and (_00814_, _41214_, _00143_);
  or (_00815_, _00814_, _00813_);
  or (_00816_, _00815_, _00812_);
  or (_00817_, _00816_, _00811_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [0], _00817_, _00806_);
  and (_00818_, _41224_, _00240_);
  and (_00820_, _41218_, _00242_);
  and (_00822_, _41211_, _00244_);
  or (_00824_, _00822_, _00820_);
  or (_00826_, _00824_, _00818_);
  and (_00828_, _00026_, _00211_);
  and (_00830_, _41254_, _00196_);
  or (_00832_, _00830_, _00828_);
  or (_00833_, _00832_, _00826_);
  and (_00834_, _41238_, _00225_);
  and (_00835_, _41249_, _00236_);
  and (_00836_, _41241_, _00234_);
  or (_00837_, _00836_, _00835_);
  or (_00838_, _00837_, _00834_);
  and (_00840_, _00020_, _00218_);
  and (_00841_, _00015_, _00232_);
  or (_00843_, _00841_, _00840_);
  or (_00844_, _00843_, _00838_);
  or (_00845_, _00844_, _00833_);
  and (_00846_, _41244_, _00221_);
  and (_00847_, _00023_, _00227_);
  and (_00848_, _41232_, _00215_);
  or (_00849_, _00848_, _00847_);
  or (_00850_, _00849_, _00846_);
  and (_00851_, _00009_, _00194_);
  and (_00852_, _00012_, _00208_);
  and (_00853_, _41214_, _00200_);
  or (_00854_, _00853_, _00852_);
  or (_00855_, _00854_, _00851_);
  or (_00856_, _00855_, _00850_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [1], _00856_, _00845_);
  and (_00857_, _00009_, _00250_);
  and (_00858_, _00020_, _00274_);
  and (_00859_, _00023_, _00280_);
  and (_00860_, _41232_, _00271_);
  or (_00861_, _00860_, _00859_);
  or (_00862_, _00861_, _00858_);
  and (_00863_, _41238_, _00282_);
  and (_00864_, _41241_, _00289_);
  and (_00865_, _41249_, _00291_);
  or (_00866_, _00865_, _00864_);
  or (_00867_, _00866_, _00863_);
  and (_00868_, _41244_, _00277_);
  and (_00869_, _00015_, _00287_);
  or (_00870_, _00869_, _00868_);
  or (_00872_, _00870_, _00867_);
  or (_00874_, _00872_, _00862_);
  or (_00876_, _00874_, _00857_);
  and (_00878_, _41214_, _00258_);
  and (_00880_, _00012_, _00266_);
  or (_00882_, _00880_, _00878_);
  and (_00884_, _41254_, _00254_);
  and (_00885_, _41224_, _00295_);
  and (_00886_, _00026_, _00264_);
  and (_00887_, _41218_, _00297_);
  and (_00888_, _41211_, _00299_);
  or (_00889_, _00888_, _00887_);
  or (_00890_, _00889_, _00886_);
  or (_00891_, _00890_, _00885_);
  or (_00892_, _00891_, _00884_);
  or (_00893_, _00892_, _00882_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [2], _00893_, _00876_);
  and (_00894_, _41218_, _00352_);
  and (_00895_, _41211_, _00355_);
  or (_00896_, _00895_, _00894_);
  and (_00897_, _00026_, _00319_);
  or (_00898_, _00897_, _00896_);
  and (_00899_, _41224_, _00350_);
  and (_00900_, _00009_, _00308_);
  or (_00901_, _00900_, _00899_);
  or (_00902_, _00901_, _00898_);
  and (_00903_, _00015_, _00342_);
  and (_00904_, _41241_, _00344_);
  and (_00905_, _41249_, _00346_);
  or (_00906_, _00905_, _00904_);
  or (_00907_, _00906_, _00903_);
  and (_00908_, _00020_, _00329_);
  and (_00909_, _41238_, _00337_);
  or (_00910_, _00909_, _00908_);
  or (_00911_, _00910_, _00907_);
  or (_00912_, _00911_, _00902_);
  and (_00913_, _41244_, _00332_);
  and (_00915_, _00023_, _00335_);
  and (_00916_, _41232_, _00327_);
  or (_00917_, _00916_, _00915_);
  or (_00919_, _00917_, _00913_);
  and (_00920_, _41254_, _00312_);
  and (_00921_, _00012_, _00322_);
  and (_00923_, _41214_, _00315_);
  or (_00924_, _00923_, _00921_);
  or (_00925_, _00924_, _00920_);
  or (_00926_, _00925_, _00919_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [3], _00926_, _00912_);
  and (_00927_, _41254_, _00398_);
  and (_00928_, _41244_, _00383_);
  and (_00929_, _41232_, _00379_);
  and (_00930_, _00023_, _00387_);
  or (_00931_, _00930_, _00929_);
  or (_00932_, _00931_, _00928_);
  and (_00933_, _41238_, _00405_);
  and (_00934_, _41249_, _00413_);
  and (_00935_, _41241_, _00409_);
  or (_00936_, _00935_, _00934_);
  or (_00937_, _00936_, _00933_);
  and (_00938_, _00015_, _00389_);
  and (_00939_, _00020_, _00381_);
  or (_00940_, _00939_, _00938_);
  or (_00941_, _00940_, _00937_);
  or (_00942_, _00941_, _00932_);
  or (_00943_, _00942_, _00927_);
  and (_00944_, _41214_, _00400_);
  and (_00945_, _00012_, _00394_);
  or (_00946_, _00945_, _00944_);
  and (_00947_, _00009_, _00396_);
  and (_00948_, _00026_, _00368_);
  and (_00949_, _41224_, _00366_);
  and (_00950_, _41218_, _00371_);
  and (_00951_, _41211_, _00374_);
  or (_00952_, _00951_, _00950_);
  or (_00953_, _00952_, _00949_);
  or (_00954_, _00953_, _00948_);
  or (_00955_, _00954_, _00947_);
  or (_00956_, _00955_, _00946_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [4], _00956_, _00943_);
  and (_00957_, _00009_, _00421_);
  and (_00958_, _41224_, _00463_);
  and (_00959_, _00026_, _00433_);
  and (_00960_, _41218_, _00467_);
  and (_00961_, _41211_, _00471_);
  or (_00962_, _00961_, _00960_);
  or (_00963_, _00962_, _00959_);
  or (_00964_, _00963_, _00958_);
  or (_00965_, _00964_, _00957_);
  and (_00966_, _00020_, _00439_);
  and (_00967_, _41238_, _00445_);
  and (_00968_, _00015_, _00452_);
  and (_00969_, _41249_, _00456_);
  and (_00970_, _41241_, _00454_);
  or (_00971_, _00970_, _00969_);
  or (_00972_, _00971_, _00968_);
  or (_00973_, _00972_, _00967_);
  or (_00974_, _00973_, _00966_);
  or (_00975_, _00974_, _00965_);
  and (_00976_, _41244_, _00441_);
  and (_00977_, _00023_, _00447_);
  and (_00978_, _41232_, _00437_);
  or (_00979_, _00978_, _00977_);
  or (_00980_, _00979_, _00976_);
  and (_00981_, _41254_, _00423_);
  and (_00982_, _00012_, _00431_);
  and (_00983_, _41214_, _00426_);
  or (_00984_, _00983_, _00982_);
  or (_00985_, _00984_, _00981_);
  or (_00986_, _00985_, _00980_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [5], _00986_, _00975_);
  and (_00987_, _41218_, _00524_);
  and (_00988_, _41211_, _00526_);
  or (_00989_, _00988_, _00987_);
  and (_00990_, _00026_, _00488_);
  or (_00991_, _00990_, _00989_);
  and (_00992_, _41224_, _00521_);
  and (_00993_, _00009_, _00476_);
  or (_00994_, _00993_, _00992_);
  or (_00995_, _00994_, _00991_);
  and (_00996_, _00015_, _00507_);
  and (_00997_, _41241_, _00509_);
  and (_00998_, _41249_, _00513_);
  or (_00999_, _00998_, _00997_);
  or (_01000_, _00999_, _00996_);
  and (_01001_, _41244_, _00496_);
  and (_01002_, _41238_, _00500_);
  or (_01003_, _01002_, _01001_);
  or (_01004_, _01003_, _01000_);
  or (_01005_, _01004_, _00995_);
  and (_01006_, _00020_, _00494_);
  and (_01007_, _00023_, _00502_);
  and (_01008_, _41232_, _00492_);
  or (_01009_, _01008_, _01007_);
  or (_01010_, _01009_, _01006_);
  and (_01011_, _41254_, _00479_);
  and (_01012_, _00012_, _00486_);
  and (_01013_, _41214_, _00482_);
  or (_01014_, _01013_, _01012_);
  or (_01015_, _01014_, _01011_);
  or (_01016_, _01015_, _01010_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [6], _01016_, _01005_);
  and (_01017_, _00026_, _00185_);
  and (_01018_, _41211_, _00187_);
  and (_01019_, _41224_, _00189_);
  or (_01020_, _01019_, _01018_);
  or (_01021_, _01020_, _01017_);
  and (_01022_, _41218_, _00143_);
  and (_01023_, _00023_, _00150_);
  or (_01024_, _01023_, _01022_);
  or (_01025_, _01024_, _01021_);
  and (_01026_, _00020_, _00176_);
  and (_01027_, _41244_, _00178_);
  and (_01028_, _41241_, _00180_);
  or (_01029_, _01028_, _01027_);
  or (_01030_, _01029_, _01026_);
  and (_01031_, _41232_, _00174_);
  and (_01032_, _00012_, _00169_);
  or (_01033_, _01032_, _01031_);
  or (_01034_, _01033_, _01030_);
  or (_01035_, _01034_, _01025_);
  and (_01036_, _00015_, _00166_);
  and (_01037_, _41238_, _00162_);
  and (_01038_, _41249_, _00160_);
  or (_01039_, _01038_, _01037_);
  or (_01040_, _01039_, _01036_);
  and (_01041_, _41254_, _00139_);
  and (_01042_, _00009_, _00154_);
  and (_01044_, _41214_, _00141_);
  or (_01045_, _01044_, _01042_);
  or (_01047_, _01045_, _01041_);
  or (_01048_, _01047_, _01040_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [8], _01048_, _01035_);
  and (_01050_, _00026_, _00240_);
  and (_01052_, _41211_, _00242_);
  and (_01053_, _41224_, _00244_);
  or (_01055_, _01053_, _01052_);
  or (_01056_, _01055_, _01050_);
  and (_01058_, _41218_, _00200_);
  and (_01059_, _00023_, _00211_);
  or (_01061_, _01059_, _01058_);
  or (_01062_, _01061_, _01056_);
  and (_01064_, _00020_, _00215_);
  and (_01065_, _41244_, _00218_);
  and (_01067_, _41241_, _00221_);
  or (_01068_, _01067_, _01065_);
  or (_01070_, _01068_, _01064_);
  and (_01071_, _41232_, _00227_);
  and (_01073_, _00012_, _00232_);
  or (_01074_, _01073_, _01071_);
  or (_01076_, _01074_, _01070_);
  or (_01077_, _01076_, _01062_);
  and (_01079_, _00015_, _00225_);
  and (_01080_, _41238_, _00236_);
  and (_01082_, _41249_, _00234_);
  or (_01083_, _01082_, _01080_);
  or (_01085_, _01083_, _01079_);
  and (_01086_, _41254_, _00194_);
  and (_01088_, _00009_, _00208_);
  and (_01089_, _41214_, _00196_);
  or (_01091_, _01089_, _01088_);
  or (_01092_, _01091_, _01086_);
  or (_01094_, _01092_, _01085_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [9], _01094_, _01077_);
  and (_01096_, _41211_, _00297_);
  and (_01097_, _41224_, _00299_);
  or (_01099_, _01097_, _01096_);
  and (_01100_, _00026_, _00295_);
  or (_01102_, _01100_, _01099_);
  and (_01103_, _41218_, _00258_);
  and (_01104_, _00023_, _00264_);
  or (_01105_, _01104_, _01103_);
  or (_01106_, _01105_, _01102_);
  and (_01107_, _41249_, _00289_);
  and (_01108_, _41238_, _00291_);
  or (_01109_, _01108_, _01107_);
  and (_01110_, _00012_, _00287_);
  and (_01111_, _00015_, _00282_);
  or (_01112_, _01111_, _01110_);
  or (_01113_, _01112_, _01109_);
  or (_01114_, _01113_, _01106_);
  and (_01115_, _41232_, _00280_);
  and (_01116_, _00020_, _00271_);
  and (_01117_, _41241_, _00277_);
  and (_01118_, _41244_, _00274_);
  or (_01119_, _01118_, _01117_);
  or (_01120_, _01119_, _01116_);
  or (_01121_, _01120_, _01115_);
  and (_01122_, _41254_, _00250_);
  and (_01123_, _00009_, _00266_);
  and (_01124_, _41214_, _00254_);
  or (_01125_, _01124_, _01123_);
  or (_01126_, _01125_, _01122_);
  or (_01127_, _01126_, _01121_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [10], _01127_, _01114_);
  and (_01128_, _41211_, _00352_);
  and (_01129_, _41224_, _00355_);
  or (_01130_, _01129_, _01128_);
  and (_01131_, _00026_, _00350_);
  or (_01132_, _01131_, _01130_);
  and (_01133_, _41218_, _00315_);
  and (_01134_, _00023_, _00319_);
  or (_01135_, _01134_, _01133_);
  or (_01136_, _01135_, _01132_);
  and (_01137_, _41249_, _00344_);
  and (_01138_, _41238_, _00346_);
  or (_01139_, _01138_, _01137_);
  and (_01140_, _00012_, _00342_);
  and (_01141_, _00015_, _00337_);
  or (_01142_, _01141_, _01140_);
  or (_01143_, _01142_, _01139_);
  or (_01144_, _01143_, _01136_);
  and (_01145_, _41232_, _00335_);
  and (_01146_, _00020_, _00327_);
  and (_01147_, _41241_, _00332_);
  and (_01148_, _41244_, _00329_);
  or (_01149_, _01148_, _01147_);
  or (_01150_, _01149_, _01146_);
  or (_01151_, _01150_, _01145_);
  and (_01152_, _41254_, _00308_);
  and (_01153_, _00009_, _00322_);
  and (_01154_, _41214_, _00312_);
  or (_01155_, _01154_, _01153_);
  or (_01156_, _01155_, _01152_);
  or (_01157_, _01156_, _01151_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [11], _01157_, _01144_);
  and (_01158_, _00026_, _00366_);
  and (_01159_, _41211_, _00371_);
  and (_01160_, _41224_, _00374_);
  or (_01161_, _01160_, _01159_);
  or (_01162_, _01161_, _01158_);
  and (_01163_, _41218_, _00400_);
  and (_01164_, _00023_, _00368_);
  or (_01165_, _01164_, _01163_);
  or (_01166_, _01165_, _01162_);
  and (_01167_, _00020_, _00379_);
  and (_01168_, _41244_, _00381_);
  and (_01169_, _41241_, _00383_);
  or (_01170_, _01169_, _01168_);
  or (_01171_, _01170_, _01167_);
  and (_01172_, _41232_, _00387_);
  and (_01173_, _00012_, _00389_);
  or (_01174_, _01173_, _01172_);
  or (_01175_, _01174_, _01171_);
  or (_01176_, _01175_, _01166_);
  and (_01177_, _00015_, _00405_);
  and (_01178_, _41249_, _00409_);
  and (_01179_, _41238_, _00413_);
  or (_01180_, _01179_, _01178_);
  or (_01181_, _01180_, _01177_);
  and (_01182_, _41254_, _00396_);
  and (_01183_, _00009_, _00394_);
  and (_01184_, _41214_, _00398_);
  or (_01185_, _01184_, _01183_);
  or (_01186_, _01185_, _01182_);
  or (_01187_, _01186_, _01181_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [12], _01187_, _01176_);
  and (_01188_, _41211_, _00467_);
  and (_01189_, _41224_, _00471_);
  or (_01190_, _01189_, _01188_);
  and (_01191_, _00026_, _00463_);
  or (_01192_, _01191_, _01190_);
  and (_01193_, _41218_, _00426_);
  and (_01194_, _00023_, _00433_);
  or (_01195_, _01194_, _01193_);
  or (_01196_, _01195_, _01192_);
  and (_01197_, _41249_, _00454_);
  and (_01198_, _41238_, _00456_);
  or (_01199_, _01198_, _01197_);
  and (_01200_, _00012_, _00452_);
  and (_01201_, _00015_, _00445_);
  or (_01202_, _01201_, _01200_);
  or (_01203_, _01202_, _01199_);
  or (_01204_, _01203_, _01196_);
  and (_01205_, _41232_, _00447_);
  and (_01206_, _00020_, _00437_);
  and (_01207_, _41241_, _00441_);
  and (_01208_, _41244_, _00439_);
  or (_01209_, _01208_, _01207_);
  or (_01210_, _01209_, _01206_);
  or (_01211_, _01210_, _01205_);
  and (_01212_, _41254_, _00421_);
  and (_01213_, _00009_, _00431_);
  and (_01214_, _41214_, _00423_);
  or (_01215_, _01214_, _01213_);
  or (_01216_, _01215_, _01212_);
  or (_01217_, _01216_, _01211_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [13], _01217_, _01204_);
  and (_01218_, _41254_, _00476_);
  and (_01219_, _41232_, _00502_);
  and (_01220_, _00020_, _00492_);
  and (_01221_, _41244_, _00494_);
  and (_01222_, _41241_, _00496_);
  or (_01223_, _01222_, _01221_);
  or (_01224_, _01223_, _01220_);
  or (_01225_, _01224_, _01219_);
  and (_01226_, _41238_, _00513_);
  and (_01227_, _41249_, _00509_);
  or (_01228_, _01227_, _01226_);
  and (_01229_, _00015_, _00500_);
  and (_01230_, _00012_, _00507_);
  or (_01231_, _01230_, _01229_);
  or (_01232_, _01231_, _01228_);
  or (_01233_, _01232_, _01225_);
  or (_01234_, _01233_, _01218_);
  and (_01235_, _41214_, _00479_);
  and (_01236_, _00009_, _00486_);
  or (_01237_, _01236_, _01235_);
  and (_01238_, _41218_, _00482_);
  and (_01239_, _00023_, _00488_);
  and (_01240_, _00026_, _00521_);
  and (_01241_, _41211_, _00524_);
  and (_01242_, _41224_, _00526_);
  or (_01243_, _01242_, _01241_);
  or (_01244_, _01243_, _01240_);
  or (_01245_, _01244_, _01239_);
  or (_01246_, _01245_, _01238_);
  or (_01247_, _01246_, _01237_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [14], _01247_, _01234_);
  nand (_01248_, \oc8051_golden_model_1.PC [1], \oc8051_golden_model_1.PC [0]);
  not (_01249_, \oc8051_golden_model_1.PC [3]);
  or (_01250_, \oc8051_golden_model_1.PC [2], _01249_);
  or (_01251_, _01250_, _01248_);
  or (_01252_, _01251_, _37703_);
  not (_01253_, \oc8051_golden_model_1.PC [1]);
  or (_01254_, _01253_, \oc8051_golden_model_1.PC [0]);
  or (_01255_, _01254_, _01250_);
  or (_01256_, _01255_, _37662_);
  and (_01257_, _01256_, _01252_);
  not (_01258_, \oc8051_golden_model_1.PC [2]);
  or (_01259_, _01258_, \oc8051_golden_model_1.PC [3]);
  or (_01260_, _01259_, _01248_);
  or (_01261_, _01260_, _37525_);
  or (_01262_, _01259_, _01254_);
  or (_01263_, _01262_, _37483_);
  and (_01264_, _01263_, _01261_);
  and (_01265_, _01264_, _01257_);
  nand (_01266_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [3]);
  or (_01267_, _01266_, _01248_);
  or (_01268_, _01267_, _37867_);
  or (_01269_, _01266_, _01254_);
  or (_01270_, _01269_, _37826_);
  and (_01271_, _01270_, _01268_);
  or (_01272_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [3]);
  or (_01273_, _01272_, _01248_);
  or (_01274_, _01273_, _37312_);
  or (_01275_, _01272_, _01254_);
  or (_01276_, _01275_, _37192_);
  and (_01277_, _01276_, _01274_);
  and (_01278_, _01277_, _01271_);
  and (_01279_, _01278_, _01265_);
  not (_01280_, \oc8051_golden_model_1.PC [0]);
  or (_01281_, \oc8051_golden_model_1.PC [1], _01280_);
  or (_01282_, _01281_, _01266_);
  or (_01283_, _01282_, _37785_);
  or (_01284_, \oc8051_golden_model_1.PC [1], \oc8051_golden_model_1.PC [0]);
  or (_01285_, _01284_, _01266_);
  or (_01286_, _01285_, _37744_);
  and (_01287_, _01286_, _01283_);
  or (_01288_, _01272_, _01284_);
  or (_01289_, _01288_, _37083_);
  or (_01290_, _01272_, _01281_);
  or (_01291_, _01290_, _37124_);
  and (_01292_, _01291_, _01289_);
  and (_01293_, _01292_, _01287_);
  or (_01294_, _01281_, _01250_);
  or (_01295_, _01294_, _37621_);
  or (_01296_, _01284_, _01250_);
  or (_01297_, _01296_, _37570_);
  and (_01298_, _01297_, _01295_);
  or (_01299_, _01281_, _01259_);
  or (_01300_, _01299_, _37442_);
  or (_01301_, _01284_, _01259_);
  or (_01302_, _01301_, _37401_);
  and (_01303_, _01302_, _01300_);
  and (_01304_, _01303_, _01298_);
  and (_01305_, _01304_, _01293_);
  and (_01306_, _01305_, _01279_);
  or (_01307_, _01251_, _37668_);
  or (_01308_, _01255_, _37627_);
  and (_01309_, _01308_, _01307_);
  or (_01310_, _01260_, _37489_);
  or (_01311_, _01262_, _37448_);
  and (_01312_, _01311_, _01310_);
  and (_01313_, _01312_, _01309_);
  or (_01314_, _01267_, _37832_);
  or (_01315_, _01269_, _37791_);
  and (_01316_, _01315_, _01314_);
  or (_01317_, _01273_, _37198_);
  or (_01318_, _01275_, _37130_);
  and (_01319_, _01318_, _01317_);
  and (_01320_, _01319_, _01316_);
  and (_01321_, _01320_, _01313_);
  or (_01322_, _01282_, _37750_);
  or (_01323_, _01285_, _37709_);
  and (_01324_, _01323_, _01322_);
  or (_01325_, _01288_, _37048_);
  or (_01326_, _01290_, _37089_);
  and (_01327_, _01326_, _01325_);
  and (_01328_, _01327_, _01324_);
  or (_01329_, _01294_, _37583_);
  or (_01330_, _01296_, _37532_);
  and (_01331_, _01330_, _01329_);
  or (_01332_, _01299_, _37407_);
  or (_01333_, _01301_, _37328_);
  and (_01334_, _01333_, _01332_);
  and (_01335_, _01334_, _01331_);
  and (_01336_, _01335_, _01328_);
  and (_01337_, _01336_, _01321_);
  and (_01338_, _01337_, _01306_);
  or (_01339_, _01251_, _37693_);
  or (_01340_, _01255_, _37652_);
  and (_01341_, _01340_, _01339_);
  or (_01342_, _01260_, _37515_);
  or (_01343_, _01262_, _37473_);
  and (_01344_, _01343_, _01342_);
  and (_01345_, _01344_, _01341_);
  or (_01346_, _01267_, _37857_);
  or (_01347_, _01269_, _37816_);
  and (_01348_, _01347_, _01346_);
  or (_01349_, _01273_, _37279_);
  or (_01350_, _01275_, _37182_);
  and (_01351_, _01350_, _01349_);
  and (_01352_, _01351_, _01348_);
  and (_01353_, _01352_, _01345_);
  or (_01354_, _01282_, _37775_);
  or (_01355_, _01285_, _37734_);
  and (_01356_, _01355_, _01354_);
  or (_01357_, _01288_, _37073_);
  or (_01358_, _01290_, _37114_);
  and (_01359_, _01358_, _01357_);
  and (_01360_, _01359_, _01356_);
  or (_01361_, _01294_, _37611_);
  or (_01362_, _01296_, _37560_);
  and (_01363_, _01362_, _01361_);
  or (_01364_, _01299_, _37432_);
  or (_01365_, _01301_, _37391_);
  and (_01366_, _01365_, _01364_);
  and (_01367_, _01366_, _01363_);
  and (_01368_, _01367_, _01360_);
  nand (_01369_, _01368_, _01353_);
  or (_01370_, _01251_, _37698_);
  or (_01371_, _01255_, _37657_);
  and (_01372_, _01371_, _01370_);
  or (_01373_, _01260_, _37520_);
  or (_01374_, _01262_, _37478_);
  and (_01375_, _01374_, _01373_);
  and (_01376_, _01375_, _01372_);
  or (_01377_, _01267_, _37862_);
  or (_01378_, _01269_, _37821_);
  and (_01379_, _01378_, _01377_);
  or (_01380_, _01273_, _37292_);
  or (_01381_, _01275_, _37187_);
  and (_01382_, _01381_, _01380_);
  and (_01383_, _01382_, _01379_);
  and (_01384_, _01383_, _01376_);
  or (_01385_, _01282_, _37780_);
  or (_01386_, _01285_, _37739_);
  and (_01387_, _01386_, _01385_);
  or (_01388_, _01288_, _37078_);
  or (_01389_, _01290_, _37119_);
  and (_01390_, _01389_, _01388_);
  and (_01391_, _01390_, _01387_);
  or (_01392_, _01294_, _37616_);
  or (_01393_, _01296_, _37565_);
  and (_01394_, _01393_, _01392_);
  or (_01395_, _01299_, _37437_);
  or (_01396_, _01301_, _37396_);
  and (_01397_, _01396_, _01395_);
  and (_01398_, _01397_, _01394_);
  and (_01399_, _01398_, _01391_);
  nand (_01400_, _01399_, _01384_);
  or (_01401_, _01400_, _01369_);
  not (_01402_, _01401_);
  and (_01403_, _01402_, _01338_);
  or (_01404_, _01251_, _37673_);
  or (_01405_, _01255_, _37632_);
  and (_01406_, _01405_, _01404_);
  or (_01407_, _01260_, _37495_);
  or (_01408_, _01262_, _37453_);
  and (_01409_, _01408_, _01407_);
  and (_01410_, _01409_, _01406_);
  or (_01411_, _01267_, _37837_);
  or (_01412_, _01269_, _37796_);
  and (_01413_, _01412_, _01411_);
  or (_01414_, _01273_, _37212_);
  or (_01415_, _01275_, _37135_);
  and (_01416_, _01415_, _01414_);
  and (_01417_, _01416_, _01413_);
  and (_01418_, _01417_, _01410_);
  or (_01419_, _01282_, _37755_);
  or (_01420_, _01285_, _37714_);
  and (_01421_, _01420_, _01419_);
  or (_01422_, _01288_, _37053_);
  or (_01423_, _01290_, _37094_);
  and (_01424_, _01423_, _01422_);
  and (_01425_, _01424_, _01421_);
  or (_01426_, _01294_, _37591_);
  or (_01427_, _01296_, _37537_);
  and (_01428_, _01427_, _01426_);
  or (_01429_, _01299_, _37412_);
  or (_01430_, _01301_, _37348_);
  and (_01431_, _01430_, _01429_);
  and (_01432_, _01431_, _01428_);
  and (_01433_, _01432_, _01425_);
  and (_01434_, _01433_, _01418_);
  or (_01435_, _01251_, _37678_);
  or (_01436_, _01255_, _37637_);
  and (_01437_, _01436_, _01435_);
  or (_01438_, _01260_, _37500_);
  or (_01439_, _01262_, _37458_);
  and (_01440_, _01439_, _01438_);
  and (_01441_, _01440_, _01437_);
  or (_01442_, _01267_, _37842_);
  or (_01443_, _01269_, _37801_);
  and (_01444_, _01443_, _01442_);
  or (_01445_, _01273_, _37231_);
  or (_01446_, _01275_, _37167_);
  and (_01447_, _01446_, _01445_);
  and (_01448_, _01447_, _01444_);
  and (_01449_, _01448_, _01441_);
  or (_01450_, _01282_, _37760_);
  or (_01451_, _01285_, _37719_);
  and (_01452_, _01451_, _01450_);
  or (_01453_, _01288_, _37058_);
  or (_01454_, _01290_, _37099_);
  and (_01455_, _01454_, _01453_);
  and (_01456_, _01455_, _01452_);
  or (_01457_, _01294_, _37596_);
  or (_01458_, _01296_, _37542_);
  and (_01459_, _01458_, _01457_);
  or (_01460_, _01299_, _37417_);
  or (_01461_, _01301_, _37361_);
  and (_01462_, _01461_, _01460_);
  and (_01463_, _01462_, _01459_);
  and (_01464_, _01463_, _01456_);
  nand (_01465_, _01464_, _01449_);
  or (_01466_, _01465_, _01434_);
  not (_01467_, _01466_);
  or (_01468_, _01251_, _37683_);
  or (_01469_, _01255_, _37642_);
  and (_01470_, _01469_, _01468_);
  or (_01471_, _01260_, _37505_);
  or (_01472_, _01262_, _37463_);
  and (_01473_, _01472_, _01471_);
  and (_01474_, _01473_, _01470_);
  or (_01475_, _01267_, _37847_);
  or (_01476_, _01269_, _37806_);
  and (_01477_, _01476_, _01475_);
  or (_01478_, _01273_, _37245_);
  or (_01479_, _01275_, _37172_);
  and (_01480_, _01479_, _01478_);
  and (_01481_, _01480_, _01477_);
  and (_01482_, _01481_, _01474_);
  or (_01483_, _01282_, _37765_);
  or (_01484_, _01285_, _37724_);
  and (_01485_, _01484_, _01483_);
  or (_01486_, _01288_, _37063_);
  or (_01487_, _01290_, _37104_);
  and (_01488_, _01487_, _01486_);
  and (_01489_, _01488_, _01485_);
  or (_01490_, _01294_, _37601_);
  or (_01491_, _01296_, _37548_);
  and (_01492_, _01491_, _01490_);
  or (_01493_, _01299_, _37422_);
  or (_01494_, _01301_, _37381_);
  and (_01495_, _01494_, _01493_);
  and (_01496_, _01495_, _01492_);
  and (_01497_, _01496_, _01489_);
  nand (_01498_, _01497_, _01482_);
  or (_01499_, _01251_, _37688_);
  or (_01500_, _01255_, _37647_);
  and (_01501_, _01500_, _01499_);
  or (_01502_, _01260_, _37510_);
  or (_01503_, _01262_, _37468_);
  and (_01504_, _01503_, _01502_);
  and (_01505_, _01504_, _01501_);
  or (_01506_, _01267_, _37852_);
  or (_01507_, _01269_, _37811_);
  and (_01508_, _01507_, _01506_);
  or (_01509_, _01273_, _37260_);
  or (_01510_, _01275_, _37177_);
  and (_01511_, _01510_, _01509_);
  and (_01512_, _01511_, _01508_);
  and (_01513_, _01512_, _01505_);
  or (_01514_, _01282_, _37770_);
  or (_01515_, _01285_, _37729_);
  and (_01516_, _01515_, _01514_);
  or (_01517_, _01288_, _37068_);
  or (_01518_, _01290_, _37109_);
  and (_01519_, _01518_, _01517_);
  and (_01520_, _01519_, _01516_);
  or (_01522_, _01294_, _37606_);
  or (_01524_, _01296_, _37555_);
  and (_01526_, _01524_, _01522_);
  or (_01527_, _01299_, _37427_);
  or (_01529_, _01301_, _37386_);
  and (_01530_, _01529_, _01527_);
  and (_01531_, _01530_, _01526_);
  and (_01532_, _01531_, _01520_);
  nand (_01533_, _01532_, _01513_);
  not (_01534_, _01533_);
  and (_01535_, _01534_, _01498_);
  and (_01536_, _01535_, _01467_);
  and (_01537_, _01536_, _01403_);
  not (_01538_, _01537_);
  or (_01539_, _01533_, _01498_);
  not (_01540_, _01539_);
  not (_01541_, _01434_);
  and (_01542_, _01465_, _01541_);
  and (_01543_, _01542_, _01540_);
  and (_01544_, _01368_, _01353_);
  or (_01545_, _01400_, _01544_);
  nand (_01546_, _01305_, _01279_);
  or (_01547_, _01337_, _01546_);
  nor (_01548_, _01547_, _01545_);
  and (_01549_, _01548_, _01543_);
  not (_01550_, _01549_);
  and (_01551_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [1]);
  nor (_01552_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [1]);
  nor (_01553_, _01552_, _01551_);
  not (_01554_, _01553_);
  or (_01555_, _01539_, _01466_);
  or (_01556_, _01337_, _01306_);
  or (_01557_, _01556_, _01545_);
  or (_01558_, _01557_, _01555_);
  and (_01559_, _01399_, _01384_);
  or (_01560_, _01559_, _01544_);
  or (_01561_, _01560_, _01556_);
  or (_01562_, _01561_, _01555_);
  and (_01563_, _01562_, _01558_);
  or (_01564_, _01560_, _01547_);
  or (_01565_, _01564_, _01555_);
  or (_01566_, _01559_, _01369_);
  or (_01567_, _01566_, _01556_);
  or (_01568_, _01567_, _01555_);
  and (_01569_, _01568_, _01565_);
  or (_01570_, _01566_, _01547_);
  or (_01572_, _01570_, _01555_);
  or (_01573_, _01556_, _01401_);
  or (_01574_, _01573_, _01555_);
  and (_01575_, _01574_, _01572_);
  and (_01576_, _01575_, _01569_);
  and (_01577_, _01576_, _01563_);
  or (_01578_, _01577_, _01554_);
  nand (_01579_, _01576_, _01563_);
  nor (_01580_, _01248_, _01258_);
  and (_01581_, _01248_, _01258_);
  nor (_01582_, _01581_, _01580_);
  not (_01583_, _01582_);
  or (_01584_, _01583_, _01579_);
  nand (_01585_, _01584_, _01578_);
  nand (_01586_, _01585_, _01550_);
  and (_01587_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.ACC [1]);
  and (_01588_, \oc8051_golden_model_1.DPL [0], \oc8051_golden_model_1.ACC [0]);
  nor (_01589_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.ACC [1]);
  nor (_01590_, _01589_, _01587_);
  and (_01591_, _01590_, _01588_);
  nor (_01592_, _01591_, _01587_);
  and (_01593_, \oc8051_golden_model_1.DPL [2], \oc8051_golden_model_1.ACC [2]);
  nor (_01594_, \oc8051_golden_model_1.DPL [2], \oc8051_golden_model_1.ACC [2]);
  nor (_01595_, _01594_, _01593_);
  not (_01596_, _01595_);
  nor (_01597_, _01596_, _01592_);
  and (_01598_, _01596_, _01592_);
  nor (_01599_, _01598_, _01597_);
  nand (_01600_, _01599_, _01549_);
  nor (_01601_, _01547_, _01401_);
  and (_01602_, _01601_, _01536_);
  not (_01603_, _01555_);
  and (_01604_, _01603_, _01548_);
  nor (_01605_, _01604_, _01602_);
  and (_01606_, _01605_, _01600_);
  nand (_01607_, _01606_, _01586_);
  and (_01608_, _01601_, _01543_);
  not (_01609_, _01608_);
  or (_01610_, _01605_, _01553_);
  and (_01611_, _01610_, _01609_);
  nand (_01612_, _01611_, _01607_);
  not (_01613_, \oc8051_golden_model_1.ACC [1]);
  and (_01614_, _01281_, _01254_);
  nor (_01615_, _01614_, _01613_);
  and (_01616_, \oc8051_golden_model_1.ACC [0], _01280_);
  and (_01617_, _01614_, _01613_);
  nor (_01618_, _01617_, _01615_);
  and (_01619_, _01618_, _01616_);
  nor (_01620_, _01619_, _01615_);
  and (_01621_, _01582_, \oc8051_golden_model_1.ACC [2]);
  nor (_01622_, _01582_, \oc8051_golden_model_1.ACC [2]);
  nor (_01623_, _01622_, _01621_);
  not (_01624_, _01623_);
  and (_01625_, _01624_, _01620_);
  nor (_01626_, _01624_, _01620_);
  nor (_01627_, _01626_, _01625_);
  and (_01628_, _01627_, _01608_);
  not (_01629_, _01545_);
  and (_01630_, _01337_, _01546_);
  and (_01631_, _01630_, _01629_);
  and (_01632_, _01631_, _01603_);
  not (_01633_, _01632_);
  not (_01634_, _01560_);
  and (_01635_, _01634_, _01338_);
  and (_01636_, _01635_, _01603_);
  and (_01637_, _01630_, _01634_);
  and (_01638_, _01637_, _01603_);
  nor (_01639_, _01638_, _01636_);
  and (_01640_, _01639_, _01633_);
  and (_01641_, _01629_, _01338_);
  and (_01642_, _01641_, _01603_);
  not (_01643_, _01566_);
  and (_01644_, _01630_, _01643_);
  and (_01645_, _01644_, _01603_);
  nor (_01646_, _01645_, _01642_);
  and (_01647_, _01630_, _01402_);
  and (_01648_, _01647_, _01603_);
  and (_01649_, _01601_, _01603_);
  nor (_01650_, _01649_, _01648_);
  and (_01651_, _01603_, _01403_);
  and (_01652_, _01643_, _01338_);
  and (_01653_, _01652_, _01603_);
  nor (_01654_, _01653_, _01651_);
  and (_01655_, _01654_, _01650_);
  and (_01656_, _01655_, _01646_);
  and (_01657_, _01656_, _01640_);
  not (_01658_, _01657_);
  nor (_01659_, _01658_, _01628_);
  nand (_01660_, _01659_, _01612_);
  or (_01661_, _01657_, _01553_);
  nand (_01662_, _01661_, _01660_);
  not (_01663_, _01605_);
  nor (_01664_, _01597_, _01593_);
  and (_01665_, \oc8051_golden_model_1.DPL [3], \oc8051_golden_model_1.ACC [3]);
  nor (_01666_, \oc8051_golden_model_1.DPL [3], \oc8051_golden_model_1.ACC [3]);
  nor (_01667_, _01666_, _01665_);
  not (_01668_, _01667_);
  nor (_01669_, _01668_, _01664_);
  and (_01670_, _01668_, _01664_);
  nor (_01671_, _01670_, _01669_);
  nand (_01672_, _01671_, _01549_);
  not (_01673_, _01260_);
  nor (_01674_, _01580_, _01249_);
  nor (_01675_, _01674_, _01673_);
  or (_01676_, _01549_, _01675_);
  or (_01677_, _01676_, _01579_);
  and (_01678_, _01677_, _01672_);
  or (_01679_, _01678_, _01663_);
  nor (_01680_, _01266_, _01253_);
  nor (_01681_, _01551_, \oc8051_golden_model_1.PC [3]);
  nor (_01682_, _01681_, _01680_);
  not (_01683_, _01682_);
  and (_01684_, _01605_, _01577_);
  or (_01685_, _01684_, _01683_);
  and (_01686_, _01685_, _01679_);
  or (_01687_, _01686_, _01608_);
  nor (_01688_, _01626_, _01621_);
  not (_01689_, \oc8051_golden_model_1.ACC [3]);
  nor (_01690_, _01675_, _01689_);
  and (_01691_, _01675_, _01689_);
  nor (_01692_, _01691_, _01690_);
  and (_01693_, _01692_, _01688_);
  nor (_01694_, _01692_, _01688_);
  nor (_01695_, _01694_, _01693_);
  nor (_01696_, _01695_, _01609_);
  nor (_01697_, _01696_, _01658_);
  nand (_01698_, _01697_, _01687_);
  or (_01699_, _01682_, _01657_);
  nand (_01700_, _01699_, _01698_);
  or (_01701_, _01700_, _01662_);
  nor (_01702_, \oc8051_golden_model_1.DPL [0], \oc8051_golden_model_1.ACC [0]);
  nor (_01703_, _01702_, _01588_);
  or (_01704_, _01703_, _01550_);
  or (_01705_, _01549_, _01280_);
  or (_01706_, _01705_, _01579_);
  nand (_01707_, _01706_, _01704_);
  and (_01708_, _01609_, _01605_);
  nand (_01709_, _01708_, _01707_);
  not (_01710_, \oc8051_golden_model_1.ACC [0]);
  and (_01711_, _01710_, \oc8051_golden_model_1.PC [0]);
  or (_01712_, _01711_, _01616_);
  nand (_01713_, _01712_, _01608_);
  and (_01714_, _01713_, _01709_);
  or (_01715_, _01714_, _01658_);
  and (_01716_, _01684_, _01657_);
  or (_01717_, _01716_, \oc8051_golden_model_1.PC [0]);
  and (_01718_, _01717_, _01715_);
  or (_01719_, _01716_, _01253_);
  nor (_01720_, _01590_, _01588_);
  nor (_01721_, _01720_, _01591_);
  or (_01722_, _01721_, _01550_);
  not (_01723_, _01614_);
  nor (_01724_, _01723_, _01549_);
  nand (_01725_, _01724_, _01577_);
  nand (_01726_, _01725_, _01722_);
  and (_01727_, _01726_, _01708_);
  nor (_01728_, _01618_, _01616_);
  nor (_01729_, _01728_, _01619_);
  nor (_01730_, _01729_, _01609_);
  or (_01731_, _01730_, _01727_);
  nand (_01732_, _01731_, _01657_);
  and (_01733_, _01732_, _01719_);
  or (_01734_, _01733_, _01718_);
  or (_01735_, _01734_, _01701_);
  or (_01736_, _01735_, _37709_);
  nand (_01737_, _01733_, _01718_);
  and (_01738_, _01699_, _01698_);
  or (_01739_, _01738_, _01662_);
  or (_01740_, _01739_, _01737_);
  or (_01741_, _01740_, _37489_);
  and (_01742_, _01741_, _01736_);
  nand (_01743_, _01732_, _01719_);
  or (_01744_, _01743_, _01718_);
  or (_01745_, _01744_, _01739_);
  or (_01746_, _01745_, _37448_);
  nand (_01747_, _01743_, _01718_);
  and (_01748_, _01661_, _01660_);
  or (_01749_, _01738_, _01748_);
  or (_01750_, _01749_, _01747_);
  or (_01751_, _01750_, _37089_);
  and (_01752_, _01751_, _01746_);
  and (_01753_, _01752_, _01742_);
  or (_01754_, _01700_, _01748_);
  or (_01755_, _01754_, _01747_);
  or (_01756_, _01755_, _37583_);
  or (_01757_, _01754_, _01744_);
  or (_01758_, _01757_, _37627_);
  and (_01759_, _01758_, _01756_);
  or (_01760_, _01754_, _01737_);
  or (_01761_, _01760_, _37668_);
  or (_01762_, _01749_, _01737_);
  or (_01763_, _01762_, _37198_);
  and (_01764_, _01763_, _01761_);
  and (_01765_, _01764_, _01759_);
  and (_01766_, _01765_, _01753_);
  or (_01767_, _01747_, _01739_);
  or (_01768_, _01767_, _37407_);
  or (_01769_, _01739_, _01734_);
  or (_01770_, _01769_, _37328_);
  and (_01771_, _01770_, _01768_);
  or (_01772_, _01737_, _01701_);
  or (_01773_, _01772_, _37832_);
  or (_01774_, _01749_, _01734_);
  or (_01775_, _01774_, _37048_);
  and (_01776_, _01775_, _01773_);
  and (_01777_, _01776_, _01771_);
  or (_01778_, _01744_, _01701_);
  or (_01779_, _01778_, _37791_);
  or (_01780_, _01749_, _01744_);
  or (_01781_, _01780_, _37130_);
  and (_01782_, _01781_, _01779_);
  or (_01783_, _01747_, _01701_);
  or (_01784_, _01783_, _37750_);
  or (_01785_, _01754_, _01734_);
  or (_01786_, _01785_, _37532_);
  and (_01787_, _01786_, _01784_);
  and (_01788_, _01787_, _01782_);
  and (_01789_, _01788_, _01777_);
  nand (_01790_, _01789_, _01766_);
  nor (_01791_, _01790_, _01538_);
  nor (_01792_, _01783_, _37760_);
  nor (_01793_, _01740_, _37500_);
  nor (_01794_, _01793_, _01792_);
  nor (_01795_, _01745_, _37458_);
  nor (_01796_, _01750_, _37099_);
  nor (_01797_, _01796_, _01795_);
  and (_01798_, _01797_, _01794_);
  nor (_01799_, _01760_, _37678_);
  nor (_01800_, _01762_, _37231_);
  nor (_01801_, _01800_, _01799_);
  nor (_01802_, _01757_, _37637_);
  nor (_01803_, _01785_, _37542_);
  nor (_01804_, _01803_, _01802_);
  and (_01805_, _01804_, _01801_);
  and (_01806_, _01805_, _01798_);
  nor (_01807_, _01767_, _37417_);
  nor (_01808_, _01769_, _37361_);
  nor (_01809_, _01808_, _01807_);
  nor (_01810_, _01778_, _37801_);
  nor (_01811_, _01774_, _37058_);
  nor (_01812_, _01811_, _01810_);
  and (_01813_, _01812_, _01809_);
  nor (_01814_, _01772_, _37842_);
  nor (_01815_, _01780_, _37167_);
  nor (_01816_, _01815_, _01814_);
  nor (_01817_, _01735_, _37719_);
  nor (_01818_, _01755_, _37596_);
  nor (_01819_, _01818_, _01817_);
  and (_01820_, _01819_, _01816_);
  and (_01821_, _01820_, _01813_);
  and (_01822_, _01821_, _01806_);
  not (_01823_, _01822_);
  and (_01824_, _01823_, _01791_);
  nor (_01825_, _01740_, _37515_);
  nor (_01826_, _01774_, _37073_);
  nor (_01827_, _01826_, _01825_);
  nor (_01828_, _01778_, _37816_);
  nor (_01829_, _01762_, _37279_);
  nor (_01830_, _01829_, _01828_);
  and (_01831_, _01830_, _01827_);
  nor (_01832_, _01745_, _37473_);
  nor (_01833_, _01767_, _37432_);
  nor (_01834_, _01833_, _01832_);
  nor (_01835_, _01783_, _37775_);
  nor (_01836_, _01735_, _37734_);
  nor (_01837_, _01836_, _01835_);
  and (_01838_, _01837_, _01834_);
  and (_01839_, _01838_, _01831_);
  nor (_01840_, _01780_, _37182_);
  nor (_01841_, _01750_, _37114_);
  nor (_01842_, _01841_, _01840_);
  nor (_01843_, _01757_, _37652_);
  nor (_01844_, _01785_, _37560_);
  nor (_01845_, _01844_, _01843_);
  and (_01846_, _01845_, _01842_);
  nor (_01847_, _01772_, _37857_);
  nor (_01848_, _01769_, _37391_);
  nor (_01849_, _01848_, _01847_);
  nor (_01850_, _01760_, _37693_);
  nor (_01851_, _01755_, _37611_);
  nor (_01852_, _01851_, _01850_);
  and (_01853_, _01852_, _01849_);
  and (_01854_, _01853_, _01846_);
  and (_01855_, _01854_, _01839_);
  nor (_01856_, _01855_, _01790_);
  not (_01857_, _01465_);
  and (_01858_, _01857_, _01434_);
  and (_01859_, _01858_, _01540_);
  and (_01860_, _01859_, _01641_);
  and (_01861_, _01860_, _01856_);
  not (_01862_, \oc8051_golden_model_1.SP [1]);
  and (_01863_, _01862_, \oc8051_golden_model_1.SP [0]);
  not (_01864_, \oc8051_golden_model_1.SP [0]);
  and (_01865_, \oc8051_golden_model_1.SP [1], _01864_);
  nor (_01866_, _01865_, _01863_);
  not (_01867_, _01866_);
  and (_01868_, _01867_, _01636_);
  and (_01869_, _01637_, _01536_);
  not (_01870_, _01869_);
  nor (_01871_, _01870_, _01790_);
  and (_01872_, _01871_, _01823_);
  and (_01873_, _01465_, _01434_);
  and (_01874_, _01873_, _01540_);
  and (_01875_, _01874_, _01548_);
  and (_01876_, _01856_, _01875_);
  not (_01877_, _01573_);
  and (_01878_, _01859_, _01877_);
  and (_01879_, _01878_, _01867_);
  not (_01880_, _01878_);
  not (_01881_, _01557_);
  and (_01882_, _01535_, _01465_);
  and (_01883_, _01882_, _01881_);
  not (_01884_, _01561_);
  and (_01885_, _01882_, _01884_);
  nor (_01886_, _01885_, _01883_);
  not (_01887_, _01860_);
  and (_01888_, _01874_, _01652_);
  not (_01889_, _01888_);
  and (_01890_, _01652_, _01536_);
  not (_01891_, _01890_);
  nor (_01892_, _01740_, _37525_);
  nor (_01893_, _01762_, _37312_);
  nor (_01894_, _01893_, _01892_);
  nor (_01895_, _01783_, _37785_);
  nor (_01896_, _01785_, _37570_);
  nor (_01897_, _01896_, _01895_);
  and (_01898_, _01897_, _01894_);
  nor (_01899_, _01745_, _37483_);
  nor (_01900_, _01767_, _37442_);
  nor (_01901_, _01900_, _01899_);
  nor (_01902_, _01780_, _37192_);
  nor (_01903_, _01750_, _37124_);
  nor (_01904_, _01903_, _01902_);
  and (_01905_, _01904_, _01901_);
  and (_01906_, _01905_, _01898_);
  nor (_01907_, _01760_, _37703_);
  nor (_01908_, _01757_, _37662_);
  nor (_01909_, _01908_, _01907_);
  nor (_01910_, _01772_, _37867_);
  nor (_01911_, _01755_, _37621_);
  nor (_01912_, _01911_, _01910_);
  and (_01913_, _01912_, _01909_);
  nor (_01914_, _01769_, _37401_);
  nor (_01915_, _01774_, _37083_);
  nor (_01916_, _01915_, _01914_);
  nor (_01917_, _01778_, _37826_);
  nor (_01918_, _01735_, _37744_);
  nor (_01919_, _01918_, _01917_);
  and (_01920_, _01919_, _01916_);
  and (_01921_, _01920_, _01913_);
  and (_01922_, _01921_, _01906_);
  nor (_01923_, _01922_, _01790_);
  or (_01924_, _01760_, _37688_);
  or (_01925_, _01740_, _37510_);
  and (_01926_, _01925_, _01924_);
  or (_01927_, _01745_, _37468_);
  or (_01928_, _01750_, _37109_);
  and (_01929_, _01928_, _01927_);
  and (_01930_, _01929_, _01926_);
  or (_01931_, _01772_, _37852_);
  or (_01932_, _01762_, _37260_);
  and (_01933_, _01932_, _01931_);
  or (_01934_, _01778_, _37811_);
  or (_01935_, _01785_, _37555_);
  and (_01936_, _01935_, _01934_);
  and (_01937_, _01936_, _01933_);
  and (_01938_, _01937_, _01930_);
  or (_01939_, _01767_, _37427_);
  or (_01940_, _01769_, _37386_);
  and (_01941_, _01940_, _01939_);
  or (_01942_, _01757_, _37647_);
  or (_01943_, _01774_, _37068_);
  and (_01944_, _01943_, _01942_);
  and (_01945_, _01944_, _01941_);
  or (_01946_, _01783_, _37770_);
  or (_01947_, _01780_, _37177_);
  and (_01948_, _01947_, _01946_);
  or (_01949_, _01735_, _37729_);
  or (_01950_, _01755_, _37606_);
  and (_01951_, _01950_, _01949_);
  and (_01952_, _01951_, _01948_);
  and (_01953_, _01952_, _01945_);
  and (_01954_, _01953_, _01938_);
  not (_01955_, _01954_);
  and (_01956_, _01955_, _01790_);
  nor (_01957_, _01956_, _01923_);
  and (_01958_, _01874_, _01637_);
  and (_01959_, _01874_, _01601_);
  nor (_01960_, _01959_, _01958_);
  not (_01961_, _01960_);
  and (_01962_, _01961_, _01957_);
  and (_01963_, _01548_, _01536_);
  not (_01964_, _01957_);
  not (_01965_, _01570_);
  and (_01966_, _01859_, _01965_);
  and (_01967_, _01874_, _01965_);
  nor (_01968_, _01967_, _01966_);
  not (_01969_, _01968_);
  not (_01970_, _01498_);
  and (_01971_, _01533_, _01970_);
  and (_01972_, _01971_, _01858_);
  and (_01973_, _01972_, _01965_);
  not (_01974_, _01973_);
  and (_01975_, _01971_, _01873_);
  and (_01976_, _01975_, _01965_);
  and (_01977_, _01533_, _01498_);
  and (_01978_, _01977_, _01858_);
  and (_01979_, _01978_, _01965_);
  or (_01980_, _01979_, _01976_);
  not (_01981_, _01980_);
  not (_01982_, _01977_);
  nor (_01983_, _01982_, _01858_);
  and (_01984_, _01983_, _01965_);
  and (_01985_, _01971_, _01541_);
  and (_01986_, _01985_, _01965_);
  nor (_01987_, _01986_, _01984_);
  and (_01988_, _01987_, _01981_);
  and (_01989_, _01988_, _01974_);
  not (_01990_, _01564_);
  and (_01991_, _01874_, _01990_);
  and (_01992_, _01859_, _01990_);
  nor (_01993_, _01992_, _01991_);
  not (_01994_, _01993_);
  and (_01995_, _01990_, _01536_);
  nor (_01996_, _01995_, _01878_);
  and (_01997_, _01874_, _01877_);
  not (_01998_, \oc8051_golden_model_1.SP [3]);
  and (_01999_, _01859_, _01881_);
  and (_02000_, _01999_, _01998_);
  and (_02001_, _01881_, _01536_);
  not (_02002_, _01567_);
  and (_02003_, _02002_, _01536_);
  nor (_02004_, _02003_, _02001_);
  or (_02005_, _02004_, _01954_);
  and (_02006_, _01877_, _01536_);
  and (_02007_, _01874_, _01881_);
  nor (_02008_, _02007_, _01999_);
  nand (_02009_, _02004_, \oc8051_golden_model_1.PSW [3]);
  and (_02010_, _02009_, _02008_);
  or (_02011_, _02010_, _02006_);
  and (_02012_, _02011_, _02005_);
  nor (_02013_, _02012_, _02000_);
  or (_02014_, _02013_, _01997_);
  and (_02015_, _02014_, _01996_);
  or (_02016_, _02015_, _01994_);
  and (_02017_, _02016_, _01989_);
  or (_02018_, _02017_, _01969_);
  and (_02019_, _02018_, _01964_);
  nor (_02020_, _01989_, _01954_);
  not (_02021_, _02006_);
  and (_02022_, _02021_, _01996_);
  nor (_02023_, _02022_, _01954_);
  not (_02024_, _02007_);
  not (_02025_, _01997_);
  and (_02026_, _02025_, _01996_);
  and (_02027_, _02026_, _02024_);
  and (_02028_, _02027_, _01989_);
  and (_02029_, _02028_, _02013_);
  or (_02030_, _02029_, _02023_);
  and (_02031_, _02030_, _01993_);
  or (_02032_, _02031_, _02020_);
  and (_02033_, _02032_, _01968_);
  nor (_02034_, _02033_, _02019_);
  or (_02035_, _02034_, _01963_);
  not (_02036_, _01963_);
  nor (_02037_, _02036_, _01954_);
  nor (_02038_, _02037_, _01875_);
  nand (_02039_, _02038_, _02035_);
  and (_02040_, _01957_, _01875_);
  nor (_02041_, _02040_, _01602_);
  nand (_02042_, _02041_, _02039_);
  not (_02043_, _01602_);
  and (_02044_, _01858_, _01535_);
  and (_02045_, _02044_, _01990_);
  not (_02046_, _02045_);
  and (_02047_, _01542_, _01535_);
  and (_02048_, _02047_, _01990_);
  and (_02049_, _01971_, _01857_);
  and (_02050_, _02049_, _01990_);
  nor (_02051_, _02050_, _02048_);
  and (_02052_, _02051_, _02046_);
  and (_02053_, _01873_, _01535_);
  and (_02054_, _02053_, _01990_);
  or (_02055_, _02054_, _01995_);
  not (_02056_, _02055_);
  and (_02057_, _01874_, _01403_);
  and (_02058_, _01874_, _01641_);
  nor (_02059_, _02058_, _02057_);
  and (_02060_, _02059_, _02056_);
  and (_02061_, _02060_, _02052_);
  and (_02062_, _01977_, _01542_);
  and (_02063_, _02062_, _01990_);
  nor (_02064_, _02063_, _02001_);
  and (_02065_, _01971_, _01465_);
  and (_02066_, _02065_, _01990_);
  and (_02067_, _01978_, _01990_);
  nor (_02068_, _02067_, _02066_);
  and (_02069_, _02068_, _02064_);
  and (_02070_, _02069_, _02061_);
  and (_02071_, _01647_, _01543_);
  and (_02072_, _01631_, _01543_);
  nor (_02073_, _02072_, _02071_);
  and (_02074_, _01977_, _01467_);
  and (_02075_, _01977_, _01873_);
  nor (_02076_, _02075_, _02074_);
  or (_02077_, _02076_, _01564_);
  and (_02078_, _02077_, _02073_);
  and (_02079_, _01644_, _01543_);
  and (_02080_, _01859_, _01548_);
  nor (_02081_, _02080_, _02079_);
  and (_02082_, _01859_, _01652_);
  and (_02083_, _01859_, _01635_);
  nor (_02084_, _02083_, _02082_);
  nor (_02085_, _01860_, _01869_);
  and (_02086_, _02085_, _02084_);
  and (_02087_, _02086_, _02081_);
  and (_02088_, _02087_, _02078_);
  and (_02089_, _02088_, _02070_);
  nor (_02090_, _02089_, _01280_);
  and (_02091_, _02089_, _01280_);
  or (_02092_, _02091_, _02090_);
  nor (_02093_, _02091_, \oc8051_golden_model_1.PC [1]);
  and (_02094_, _02091_, \oc8051_golden_model_1.PC [1]);
  nor (_02095_, _02094_, _02093_);
  not (_02096_, _02095_);
  and (_02097_, _02096_, _02092_);
  nor (_02098_, _02089_, _01554_);
  and (_02099_, _02089_, _01582_);
  nor (_02100_, _02099_, _02098_);
  not (_02101_, _02100_);
  nor (_02102_, _02089_, _01683_);
  not (_02103_, _01675_);
  and (_02104_, _02089_, _02103_);
  nor (_02105_, _02104_, _02102_);
  and (_02106_, _02105_, _02101_);
  and (_02107_, _02106_, _02097_);
  and (_02108_, _02107_, _00335_);
  and (_02109_, _02105_, _02100_);
  and (_02110_, _02109_, _02097_);
  and (_02111_, _02110_, _00344_);
  nor (_02112_, _02111_, _02108_);
  nor (_02113_, _02095_, _02092_);
  nor (_02114_, _02105_, _02100_);
  and (_02115_, _02114_, _02113_);
  and (_02116_, _02115_, _00308_);
  and (_02117_, _02095_, _02092_);
  nor (_02118_, _02105_, _02101_);
  and (_02119_, _02118_, _02117_);
  and (_02120_, _02119_, _00350_);
  nor (_02121_, _02120_, _02116_);
  and (_02122_, _02121_, _02112_);
  and (_02123_, _02113_, _02106_);
  and (_02124_, _02123_, _00327_);
  and (_02125_, _02117_, _02106_);
  and (_02126_, _02125_, _00329_);
  nor (_02127_, _02126_, _02124_);
  and (_02128_, _02113_, _02109_);
  and (_02129_, _02128_, _00346_);
  and (_02130_, _02117_, _02109_);
  and (_02131_, _02130_, _00337_);
  nor (_02132_, _02131_, _02129_);
  and (_02133_, _02132_, _02127_);
  and (_02134_, _02133_, _02122_);
  and (_02135_, _02117_, _02114_);
  and (_02136_, _02135_, _00312_);
  and (_02137_, _02118_, _02097_);
  and (_02138_, _02137_, _00352_);
  nor (_02139_, _02138_, _02136_);
  and (_02140_, _02114_, _02097_);
  and (_02141_, _02140_, _00322_);
  nor (_02142_, _02096_, _02092_);
  and (_02143_, _02142_, _02114_);
  and (_02144_, _02143_, _00315_);
  nor (_02145_, _02144_, _02141_);
  and (_02146_, _02145_, _02139_);
  and (_02147_, _02142_, _02106_);
  and (_02148_, _02147_, _00332_);
  and (_02149_, _02142_, _02109_);
  and (_02150_, _02149_, _00342_);
  nor (_02151_, _02150_, _02148_);
  and (_02152_, _02118_, _02113_);
  and (_02153_, _02152_, _00355_);
  and (_02154_, _02142_, _02118_);
  and (_02155_, _02154_, _00319_);
  nor (_02156_, _02155_, _02153_);
  and (_02157_, _02156_, _02151_);
  and (_02158_, _02157_, _02146_);
  and (_02159_, _02158_, _02134_);
  nor (_02160_, _02159_, _02043_);
  nor (_02161_, _02160_, _01961_);
  and (_02162_, _02161_, _02042_);
  or (_02163_, _02162_, _01962_);
  and (_02164_, _01635_, _01536_);
  not (_02165_, _02164_);
  not (_02166_, _02079_);
  and (_02167_, _01874_, _01644_);
  and (_02168_, _01644_, _01536_);
  nor (_02169_, _02168_, _02167_);
  and (_02170_, _02169_, _02166_);
  and (_02171_, _01647_, _01536_);
  not (_02172_, _02171_);
  and (_02173_, _01874_, _01647_);
  nor (_02174_, _02173_, _02071_);
  and (_02175_, _02174_, _02172_);
  not (_02176_, _02072_);
  and (_02177_, _01874_, _01631_);
  and (_02178_, _01631_, _01536_);
  nor (_02179_, _02178_, _02177_);
  and (_02180_, _02179_, _02176_);
  and (_02181_, _02180_, _02175_);
  and (_02182_, _02181_, _02170_);
  and (_02183_, _02182_, _02165_);
  nand (_02184_, _02183_, _02163_);
  and (_02185_, _01874_, _01635_);
  nor (_02186_, _02183_, _01955_);
  nor (_02187_, _02186_, _02185_);
  and (_02188_, _02187_, _02184_);
  and (_02189_, _02185_, \oc8051_golden_model_1.SP [3]);
  or (_02190_, _02189_, _02083_);
  nor (_02191_, _02190_, _02188_);
  and (_02192_, _02083_, _01957_);
  or (_02193_, _02192_, _02191_);
  and (_02194_, _02193_, _01891_);
  and (_02195_, _01890_, _01954_);
  or (_02196_, _02195_, _02194_);
  nand (_02197_, _02196_, _01889_);
  and (_02198_, _01888_, _01998_);
  nor (_02199_, _02198_, _02082_);
  and (_02200_, _02199_, _02197_);
  and (_02201_, _01641_, _01536_);
  not (_02202_, _02082_);
  nor (_02203_, _01957_, _02202_);
  or (_02205_, _02203_, _02201_);
  nor (_02207_, _02205_, _02200_);
  and (_02209_, _01954_, _02201_);
  or (_02211_, _02209_, _02207_);
  nand (_02213_, _02211_, _01887_);
  and (_02215_, _01860_, _01957_);
  nor (_02217_, _02215_, _01537_);
  nand (_02218_, _02217_, _02213_);
  nor (_02219_, _01954_, _01538_);
  not (_02220_, _02219_);
  and (_02221_, _02220_, _02218_);
  nor (_02222_, _01774_, _37078_);
  nor (_02223_, _01780_, _37187_);
  nor (_02224_, _02223_, _02222_);
  nor (_02225_, _01735_, _37739_);
  nor (_02226_, _01745_, _37478_);
  nor (_02227_, _02226_, _02225_);
  and (_02228_, _02227_, _02224_);
  nor (_02229_, _01760_, _37698_);
  nor (_02230_, _01755_, _37616_);
  nor (_02231_, _02230_, _02229_);
  nor (_02232_, _01769_, _37396_);
  nor (_02233_, _01750_, _37119_);
  nor (_02234_, _02233_, _02232_);
  and (_02235_, _02234_, _02231_);
  and (_02236_, _02235_, _02228_);
  nor (_02237_, _01772_, _37862_);
  nor (_02238_, _01778_, _37821_);
  nor (_02239_, _02238_, _02237_);
  nor (_02240_, _01783_, _37780_);
  nor (_02241_, _01785_, _37565_);
  nor (_02242_, _02241_, _02240_);
  and (_02243_, _02242_, _02239_);
  nor (_02244_, _01757_, _37657_);
  nor (_02245_, _01762_, _37292_);
  nor (_02246_, _02245_, _02244_);
  nor (_02247_, _01740_, _37520_);
  nor (_02248_, _01767_, _37437_);
  nor (_02249_, _02248_, _02247_);
  and (_02250_, _02249_, _02246_);
  and (_02251_, _02250_, _02243_);
  and (_02252_, _02251_, _02236_);
  nor (_02253_, _02252_, _01790_);
  nor (_02254_, _01860_, _01997_);
  nor (_02255_, _02007_, _01875_);
  and (_02256_, _02255_, _02254_);
  and (_02257_, _02256_, _01960_);
  and (_02258_, _01993_, _01968_);
  and (_02259_, _02258_, _02084_);
  and (_02260_, _02259_, _02257_);
  not (_02261_, _02260_);
  and (_02262_, _02261_, _02253_);
  not (_02263_, _02262_);
  nor (_02264_, _01762_, _37245_);
  nor (_02265_, _01769_, _37381_);
  nor (_02266_, _02265_, _02264_);
  nor (_02267_, _01772_, _37847_);
  nor (_02268_, _01785_, _37548_);
  nor (_02269_, _02268_, _02267_);
  and (_02270_, _02269_, _02266_);
  nor (_02271_, _01778_, _37806_);
  nor (_02272_, _01783_, _37765_);
  nor (_02273_, _02272_, _02271_);
  nor (_02274_, _01740_, _37505_);
  nor (_02275_, _01767_, _37422_);
  nor (_02276_, _02275_, _02274_);
  and (_02277_, _02276_, _02273_);
  and (_02278_, _02277_, _02270_);
  nor (_02279_, _01757_, _37642_);
  nor (_02280_, _01755_, _37601_);
  nor (_02281_, _02280_, _02279_);
  nor (_02282_, _01774_, _37063_);
  nor (_02283_, _01750_, _37104_);
  nor (_02284_, _02283_, _02282_);
  and (_02285_, _02284_, _02281_);
  nor (_02286_, _01735_, _37724_);
  nor (_02287_, _01745_, _37463_);
  nor (_02288_, _02287_, _02286_);
  nor (_02289_, _01760_, _37683_);
  nor (_02290_, _01780_, _37172_);
  nor (_02291_, _02290_, _02289_);
  and (_02292_, _02291_, _02288_);
  and (_02293_, _02292_, _02285_);
  and (_02294_, _02293_, _02278_);
  nor (_02295_, _02294_, _01538_);
  not (_02296_, _02295_);
  nor (_02297_, _01890_, _02006_);
  nor (_02298_, _02164_, _01963_);
  and (_02299_, _02298_, _02297_);
  and (_02300_, _02004_, _01996_);
  and (_02301_, _02300_, _02299_);
  and (_02302_, _02301_, _01989_);
  not (_02303_, _02201_);
  and (_02304_, _02182_, _02303_);
  and (_02305_, _02304_, _02302_);
  nor (_02306_, _02305_, _02294_);
  not (_02307_, _02306_);
  and (_02308_, _02115_, _00250_);
  and (_02309_, _02135_, _00254_);
  nor (_02310_, _02309_, _02308_);
  and (_02311_, _02125_, _00274_);
  and (_02312_, _02110_, _00289_);
  nor (_02313_, _02312_, _02311_);
  and (_02314_, _02313_, _02310_);
  and (_02315_, _02128_, _00291_);
  and (_02316_, _02130_, _00282_);
  nor (_02317_, _02316_, _02315_);
  and (_02318_, _02123_, _00271_);
  and (_02319_, _02147_, _00277_);
  nor (_02320_, _02319_, _02318_);
  and (_02321_, _02320_, _02317_);
  and (_02322_, _02321_, _02314_);
  and (_02323_, _02152_, _00299_);
  and (_02324_, _02154_, _00264_);
  nor (_02325_, _02324_, _02323_);
  and (_02326_, _02140_, _00266_);
  and (_02327_, _02143_, _00258_);
  nor (_02328_, _02327_, _02326_);
  and (_02329_, _02328_, _02325_);
  and (_02330_, _02107_, _00280_);
  and (_02331_, _02149_, _00287_);
  nor (_02332_, _02331_, _02330_);
  and (_02333_, _02137_, _00297_);
  and (_02334_, _02119_, _00295_);
  nor (_02335_, _02334_, _02333_);
  and (_02336_, _02335_, _02332_);
  and (_02337_, _02336_, _02329_);
  and (_02338_, _02337_, _02322_);
  nor (_02339_, _02338_, _02043_);
  and (_02340_, _01977_, _01465_);
  and (_02341_, _02340_, _01641_);
  and (_02342_, _02340_, _01881_);
  nor (_02343_, _02342_, _02341_);
  nand (_02344_, _01977_, _01631_);
  nor (_02345_, _02344_, _01465_);
  not (_02346_, \oc8051_golden_model_1.SP [2]);
  nor (_02347_, _02185_, _01888_);
  nor (_02348_, _02347_, _02346_);
  nor (_02349_, _02348_, _02345_);
  and (_02350_, _02349_, _02343_);
  and (_02351_, _02340_, _01644_);
  not (_02352_, _02351_);
  nor (_02353_, _01982_, _01567_);
  and (_02354_, _02340_, _01601_);
  nor (_02355_, _02354_, _02353_);
  and (_02356_, _02355_, _02352_);
  and (_02357_, _01977_, _01652_);
  and (_02358_, _01977_, _01857_);
  and (_02359_, _02358_, _01635_);
  nor (_02360_, _02359_, _02357_);
  and (_02361_, _02358_, _01647_);
  and (_02362_, _02358_, _01601_);
  nor (_02363_, _02362_, _02361_);
  and (_02364_, _02363_, _02360_);
  and (_02365_, _02364_, _02356_);
  and (_02366_, _02358_, _01881_);
  and (_02367_, _02358_, _01877_);
  nor (_02368_, _02367_, _02366_);
  not (_02369_, _02368_);
  not (_02370_, _02358_);
  not (_02371_, _01644_);
  not (_02372_, _01548_);
  and (_02373_, _01564_, _02372_);
  and (_02374_, _02373_, _02371_);
  nor (_02375_, _02374_, _02370_);
  nor (_02376_, _02375_, _02369_);
  and (_02377_, _02376_, _02365_);
  and (_02378_, _01977_, _01403_);
  and (_02379_, _02378_, _01465_);
  not (_02380_, _02379_);
  and (_02381_, _01999_, \oc8051_golden_model_1.SP [2]);
  not (_02382_, _02340_);
  nor (_02383_, _02373_, _02382_);
  nor (_02384_, _02383_, _02381_);
  and (_02385_, _02384_, _02380_);
  and (_02386_, _02358_, _01403_);
  and (_02387_, _01977_, _01641_);
  and (_02388_, _02387_, _01857_);
  nor (_02389_, _02388_, _02386_);
  and (_02390_, _02340_, _01631_);
  and (_02391_, _02340_, _01635_);
  or (_02392_, _02391_, _02390_);
  not (_02393_, _02392_);
  and (_02394_, _02340_, _01877_);
  and (_02395_, _02340_, _01647_);
  nor (_02396_, _02395_, _02394_);
  and (_02397_, _02396_, _02393_);
  and (_02398_, _02397_, _02389_);
  and (_02399_, _02398_, _02385_);
  and (_02400_, _02399_, _02377_);
  and (_02401_, _02400_, _02350_);
  not (_02402_, _02401_);
  nor (_02403_, _02402_, _02339_);
  and (_02404_, _02403_, _02307_);
  and (_02405_, _02404_, _02296_);
  and (_02406_, _02405_, _02263_);
  not (_02407_, \oc8051_golden_model_1.IRAM[0] [1]);
  not (_02408_, _01875_);
  or (_02409_, _01954_, _01790_);
  nor (_02410_, _02409_, _02408_);
  or (_02411_, _01762_, _37212_);
  or (_02412_, _01750_, _37094_);
  and (_02413_, _02412_, _02411_);
  or (_02414_, _01785_, _37537_);
  or (_02415_, _01780_, _37135_);
  and (_02416_, _02415_, _02414_);
  and (_02417_, _02416_, _02413_);
  or (_02418_, _01740_, _37495_);
  or (_02419_, _01745_, _37453_);
  and (_02420_, _02419_, _02418_);
  or (_02421_, _01772_, _37837_);
  or (_02422_, _01783_, _37755_);
  and (_02423_, _02422_, _02421_);
  and (_02424_, _02423_, _02420_);
  and (_02425_, _02424_, _02417_);
  or (_02426_, _01767_, _37412_);
  or (_02427_, _01774_, _37053_);
  and (_02428_, _02427_, _02426_);
  or (_02429_, _01760_, _37673_);
  or (_02430_, _01757_, _37632_);
  and (_02431_, _02430_, _02429_);
  and (_02432_, _02431_, _02428_);
  or (_02433_, _01778_, _37796_);
  or (_02434_, _01735_, _37714_);
  and (_02435_, _02434_, _02433_);
  or (_02436_, _01755_, _37591_);
  or (_02437_, _01769_, _37348_);
  and (_02438_, _02437_, _02436_);
  and (_02439_, _02438_, _02435_);
  and (_02440_, _02439_, _02432_);
  and (_02441_, _02440_, _02425_);
  nor (_02442_, _02441_, _02036_);
  nor (_02443_, _02409_, _01968_);
  not (_02444_, _01995_);
  nor (_02445_, _02441_, _02444_);
  or (_02446_, _02441_, _02021_);
  nor (_02447_, _02441_, _02004_);
  and (_02448_, _01972_, _02002_);
  and (_02449_, _02053_, _02002_);
  nor (_02450_, _02449_, _02448_);
  and (_02451_, _01874_, _01884_);
  and (_02452_, _01975_, _02002_);
  nor (_02453_, _02452_, _02451_);
  and (_02454_, _02453_, _02450_);
  and (_02455_, _01977_, _01434_);
  and (_02456_, _02455_, _02002_);
  not (_02457_, _02456_);
  and (_02458_, _02053_, _01884_);
  nor (_02459_, _02458_, _02003_);
  and (_02460_, _02459_, _02457_);
  and (_02461_, _02460_, _02454_);
  or (_02462_, _02342_, _01883_);
  and (_02463_, _02462_, _01434_);
  and (_02464_, _01978_, _01881_);
  and (_02465_, _01971_, _01434_);
  and (_02466_, _02465_, _01881_);
  and (_02467_, _01874_, _02002_);
  or (_02468_, _02467_, _02001_);
  or (_02469_, _02468_, _02466_);
  or (_02470_, _02469_, _02464_);
  nor (_02471_, _02470_, _02463_);
  and (_02472_, _02471_, _02461_);
  or (_02473_, _02472_, _02447_);
  nand (_02474_, _02473_, _02024_);
  or (_02475_, _02409_, _02024_);
  nand (_02476_, _02475_, _02474_);
  and (_02477_, _02065_, _01877_);
  nor (_02478_, _02477_, _02394_);
  or (_02479_, _02478_, _01541_);
  and (_02480_, _01999_, _01864_);
  or (_02481_, _02480_, _02006_);
  and (_02482_, _01972_, _01877_);
  or (_02483_, _02053_, _01978_);
  and (_02484_, _02483_, _01877_);
  or (_02485_, _02484_, _02482_);
  nor (_02486_, _02485_, _02481_);
  and (_02487_, _02486_, _02479_);
  nand (_02488_, _02487_, _02476_);
  nand (_02489_, _02488_, _02446_);
  and (_02490_, _02489_, _02025_);
  nor (_02491_, _02409_, _02025_);
  or (_02492_, _02491_, _02490_);
  and (_02493_, _02441_, _01878_);
  and (_02494_, _01533_, _01434_);
  not (_02495_, _02494_);
  nor (_02496_, _02495_, _01564_);
  nor (_02497_, _02496_, _02055_);
  not (_02498_, _02497_);
  nor (_02499_, _02498_, _02493_);
  and (_02500_, _02499_, _02492_);
  or (_02501_, _02500_, _02445_);
  nand (_02502_, _02501_, _01993_);
  not (_02503_, _01989_);
  nor (_02504_, _02409_, _01993_);
  nor (_02505_, _02504_, _02503_);
  nand (_02506_, _02505_, _02502_);
  and (_02507_, _02441_, _02503_);
  and (_02508_, _02053_, _01965_);
  nor (_02509_, _02508_, _01969_);
  not (_02510_, _02509_);
  nor (_02511_, _02510_, _02507_);
  and (_02512_, _02511_, _02506_);
  or (_02513_, _02512_, _02443_);
  and (_02514_, _01978_, _01548_);
  and (_02515_, _01975_, _01548_);
  nor (_02516_, _02515_, _02514_);
  not (_02517_, _02516_);
  nor (_02518_, _02075_, _01536_);
  nor (_02519_, _02053_, _01972_);
  and (_02520_, _02519_, _02518_);
  nor (_02521_, _02520_, _02372_);
  nor (_02522_, _02521_, _02517_);
  and (_02523_, _02522_, _02513_);
  or (_02524_, _02523_, _02442_);
  and (_02525_, _02524_, _02408_);
  or (_02526_, _02525_, _02410_);
  and (_02527_, _02065_, _01601_);
  and (_02528_, _01882_, _01601_);
  nor (_02529_, _02528_, _02527_);
  nor (_02530_, _02529_, _01541_);
  not (_02531_, _01601_);
  not (_02532_, _01972_);
  nor (_02533_, _02455_, _01536_);
  and (_02534_, _02533_, _02532_);
  nor (_02535_, _02534_, _02531_);
  nor (_02536_, _02535_, _02530_);
  and (_02537_, _02536_, _02526_);
  and (_02538_, _02123_, _00176_);
  and (_02539_, _02125_, _00178_);
  nor (_02540_, _02539_, _02538_);
  and (_02541_, _02135_, _00141_);
  and (_02542_, _02137_, _00187_);
  nor (_02543_, _02542_, _02541_);
  and (_02544_, _02543_, _02540_);
  and (_02545_, _02152_, _00189_);
  and (_02546_, _02119_, _00185_);
  nor (_02547_, _02546_, _02545_);
  and (_02548_, _02115_, _00139_);
  and (_02549_, _02143_, _00143_);
  nor (_02550_, _02549_, _02548_);
  and (_02551_, _02550_, _02547_);
  and (_02552_, _02551_, _02544_);
  and (_02553_, _02149_, _00169_);
  and (_02554_, _02128_, _00162_);
  nor (_02555_, _02554_, _02553_);
  and (_02556_, _02107_, _00174_);
  and (_02557_, _02147_, _00180_);
  nor (_02558_, _02557_, _02556_);
  and (_02559_, _02558_, _02555_);
  and (_02560_, _02140_, _00154_);
  and (_02561_, _02154_, _00150_);
  nor (_02562_, _02561_, _02560_);
  and (_02563_, _02110_, _00160_);
  and (_02564_, _02130_, _00166_);
  nor (_02565_, _02564_, _02563_);
  and (_02566_, _02565_, _02562_);
  and (_02567_, _02566_, _02559_);
  and (_02568_, _02567_, _02552_);
  nor (_02569_, _02568_, _02043_);
  or (_02570_, _02569_, _02537_);
  and (_02571_, _02409_, _01959_);
  or (_02572_, _02053_, _01874_);
  and (_02573_, _02572_, _01637_);
  nor (_02574_, _02573_, _02571_);
  and (_02575_, _02574_, _02570_);
  not (_02576_, _01958_);
  nor (_02577_, _02409_, _02576_);
  or (_02578_, _02577_, _02575_);
  and (_02579_, _01882_, _01644_);
  and (_02580_, _02579_, _01434_);
  and (_02581_, _02494_, _01644_);
  nor (_02582_, _02581_, _02580_);
  and (_02583_, _02582_, _02578_);
  not (_02584_, _02441_);
  nor (_02585_, _02584_, _02170_);
  not (_02586_, _01631_);
  nor (_02587_, _02053_, _01975_);
  nor (_02588_, _02455_, _01972_);
  and (_02589_, _02588_, _02587_);
  nor (_02590_, _02589_, _02586_);
  nor (_02591_, _02590_, _02585_);
  and (_02592_, _02591_, _02583_);
  nor (_02593_, _02584_, _02181_);
  and (_02594_, _01975_, _01647_);
  not (_02595_, _01647_);
  not (_02596_, _02455_);
  and (_02597_, _02519_, _02596_);
  nor (_02598_, _02597_, _02595_);
  nor (_02599_, _02598_, _02594_);
  not (_02600_, _01635_);
  and (_02601_, _02587_, _02534_);
  nor (_02602_, _02601_, _02600_);
  not (_02603_, _02602_);
  and (_02604_, _02603_, _02599_);
  not (_02605_, _02604_);
  nor (_02606_, _02605_, _02593_);
  and (_02607_, _02606_, _02592_);
  nor (_02608_, _02441_, _02165_);
  nor (_02609_, _02608_, _02607_);
  and (_02610_, _02185_, _01864_);
  nor (_02611_, _02610_, _02609_);
  not (_02612_, _01652_);
  nor (_02613_, _02601_, _02612_);
  and (_02614_, _02409_, _02083_);
  nor (_02615_, _02614_, _02613_);
  and (_02616_, _02615_, _02611_);
  nor (_02617_, _02441_, _01891_);
  nor (_02618_, _02617_, _02616_);
  and (_02619_, _01888_, _01864_);
  nor (_02620_, _02619_, _02618_);
  and (_02621_, _02075_, _01641_);
  and (_02622_, _02387_, _01858_);
  and (_02623_, _02053_, _01641_);
  and (_02624_, _02465_, _01641_);
  or (_02625_, _02624_, _02201_);
  or (_02626_, _02625_, _02623_);
  or (_02627_, _02626_, _02622_);
  nor (_02628_, _02627_, _02621_);
  not (_02629_, _02628_);
  and (_02630_, _02409_, _02082_);
  nor (_02631_, _02630_, _02629_);
  and (_02632_, _02631_, _02620_);
  nor (_02633_, _02441_, _02303_);
  or (_02634_, _02633_, _02632_);
  and (_02635_, _02634_, _01887_);
  nor (_02636_, _02409_, _01887_);
  or (_02637_, _02636_, _02635_);
  and (_02638_, _01972_, _01403_);
  nor (_02639_, _02638_, _01537_);
  and (_02640_, _01978_, _01403_);
  not (_02641_, _02640_);
  and (_02642_, _01975_, _01403_);
  not (_02643_, _02642_);
  and (_02644_, _02075_, _01403_);
  and (_02645_, _02053_, _01403_);
  nor (_02646_, _02645_, _02644_);
  and (_02647_, _02646_, _02643_);
  and (_02648_, _02647_, _02641_);
  and (_02649_, _02648_, _02639_);
  nand (_02650_, _02649_, _02637_);
  nor (_02651_, _02441_, _01538_);
  not (_02652_, _02651_);
  nand (_02653_, _02652_, _02650_);
  or (_02654_, _02653_, _02407_);
  and (_02655_, _02261_, _01856_);
  not (_02656_, _02655_);
  and (_02657_, _02107_, _00227_);
  and (_02658_, _02130_, _00225_);
  nor (_02659_, _02658_, _02657_);
  and (_02660_, _02119_, _00240_);
  and (_02661_, _02110_, _00234_);
  nor (_02662_, _02661_, _02660_);
  and (_02663_, _02662_, _02659_);
  and (_02664_, _02137_, _00242_);
  and (_02665_, _02149_, _00232_);
  nor (_02666_, _02665_, _02664_);
  and (_02667_, _02135_, _00196_);
  and (_02668_, _02143_, _00200_);
  nor (_02669_, _02668_, _02667_);
  and (_02670_, _02669_, _02666_);
  and (_02671_, _02670_, _02663_);
  and (_02672_, _02115_, _00194_);
  and (_02673_, _02128_, _00236_);
  nor (_02674_, _02673_, _02672_);
  and (_02675_, _02154_, _00211_);
  and (_02676_, _02123_, _00215_);
  nor (_02677_, _02676_, _02675_);
  and (_02678_, _02677_, _02674_);
  and (_02679_, _02152_, _00244_);
  and (_02680_, _02147_, _00221_);
  nor (_02681_, _02680_, _02679_);
  and (_02682_, _02140_, _00208_);
  and (_02683_, _02125_, _00218_);
  nor (_02684_, _02683_, _02682_);
  and (_02685_, _02684_, _02681_);
  and (_02686_, _02685_, _02678_);
  and (_02687_, _02686_, _02671_);
  nor (_02688_, _02687_, _02043_);
  and (_02689_, _01975_, _01631_);
  and (_02690_, _01971_, _01542_);
  and (_02691_, _02690_, _02002_);
  nor (_02692_, _02691_, _02689_);
  and (_02693_, _01975_, _01652_);
  nor (_02694_, _02693_, _02452_);
  and (_02695_, _02694_, _02692_);
  and (_02696_, _02690_, _01631_);
  and (_02697_, _02340_, _02002_);
  nor (_02698_, _02697_, _02696_);
  and (_02699_, _01975_, _01635_);
  nor (_02700_, _02699_, _02515_);
  and (_02701_, _02700_, _02698_);
  nor (_02702_, _02477_, _02341_);
  and (_02703_, _01888_, \oc8051_golden_model_1.SP [1]);
  not (_02704_, _02703_);
  and (_02705_, _02065_, _01403_);
  and (_02706_, _02065_, _01881_);
  nor (_02707_, _02706_, _02705_);
  and (_02708_, _02707_, _02704_);
  and (_02709_, _02708_, _02702_);
  and (_02710_, _02709_, _02701_);
  and (_02711_, _02710_, _02695_);
  not (_02712_, _02690_);
  nor (_02713_, _01635_, _01548_);
  and (_02714_, _02713_, _02612_);
  nor (_02715_, _02714_, _02712_);
  not (_02716_, _02715_);
  and (_02717_, _02340_, _01403_);
  and (_02718_, _02065_, _01641_);
  nor (_02719_, _02718_, _02717_);
  not (_02720_, _02719_);
  nor (_02721_, _01999_, _02185_);
  nor (_02722_, _02721_, _01862_);
  nor (_02723_, _02722_, _02720_);
  and (_02724_, _02723_, _02716_);
  nor (_02725_, _02383_, _02342_);
  and (_02726_, _02725_, _02397_);
  and (_02727_, _02340_, _01652_);
  not (_02728_, _02727_);
  not (_02729_, _02527_);
  nand (_02730_, _02065_, _01647_);
  and (_02731_, _02730_, _02729_);
  and (_02732_, _02731_, _02728_);
  nor (_02733_, _02354_, _02066_);
  and (_02734_, _02065_, _01644_);
  nor (_02735_, _02734_, _02351_);
  and (_02736_, _02735_, _02733_);
  and (_02737_, _02736_, _02732_);
  and (_02738_, _02737_, _02726_);
  and (_02739_, _02738_, _02724_);
  and (_02740_, _02739_, _02711_);
  not (_02741_, _02740_);
  nor (_02742_, _02741_, _02688_);
  nor (_02743_, _02201_, _01537_);
  and (_02744_, _02743_, _02182_);
  and (_02745_, _02744_, _02302_);
  nor (_02746_, _02745_, _01822_);
  not (_02747_, _02746_);
  and (_02748_, _02747_, _02742_);
  and (_02749_, _02748_, _02656_);
  not (_02750_, \oc8051_golden_model_1.IRAM[1] [1]);
  and (_02751_, _02652_, _02650_);
  or (_02752_, _02751_, _02750_);
  and (_02753_, _02752_, _02749_);
  nand (_02754_, _02753_, _02654_);
  not (_02755_, \oc8051_golden_model_1.IRAM[3] [1]);
  or (_02756_, _02751_, _02755_);
  not (_02757_, _02749_);
  not (_02758_, \oc8051_golden_model_1.IRAM[2] [1]);
  or (_02759_, _02653_, _02758_);
  and (_02760_, _02759_, _02757_);
  nand (_02761_, _02760_, _02756_);
  nand (_02762_, _02761_, _02754_);
  nand (_02763_, _02762_, _02406_);
  not (_02764_, _02406_);
  not (_02765_, \oc8051_golden_model_1.IRAM[7] [1]);
  or (_02766_, _02751_, _02765_);
  not (_02767_, \oc8051_golden_model_1.IRAM[6] [1]);
  or (_02768_, _02653_, _02767_);
  and (_02769_, _02768_, _02757_);
  nand (_02770_, _02769_, _02766_);
  not (_02771_, \oc8051_golden_model_1.IRAM[4] [1]);
  or (_02772_, _02653_, _02771_);
  not (_02773_, \oc8051_golden_model_1.IRAM[5] [1]);
  or (_02774_, _02751_, _02773_);
  and (_02775_, _02774_, _02749_);
  nand (_02776_, _02775_, _02772_);
  nand (_02777_, _02776_, _02770_);
  nand (_02778_, _02777_, _02764_);
  nand (_02780_, _02778_, _02763_);
  nand (_02781_, _02780_, _02221_);
  not (_02782_, _02221_);
  nand (_02784_, _02653_, \oc8051_golden_model_1.IRAM[11] [1]);
  nand (_02785_, _02751_, \oc8051_golden_model_1.IRAM[10] [1]);
  and (_02786_, _02785_, _02757_);
  nand (_02787_, _02786_, _02784_);
  not (_02788_, \oc8051_golden_model_1.IRAM[8] [1]);
  or (_02789_, _02653_, _02788_);
  nand (_02790_, _02653_, \oc8051_golden_model_1.IRAM[9] [1]);
  and (_02791_, _02790_, _02749_);
  nand (_02792_, _02791_, _02789_);
  nand (_02793_, _02792_, _02787_);
  nand (_02794_, _02793_, _02406_);
  not (_02795_, \oc8051_golden_model_1.IRAM[15] [1]);
  or (_02796_, _02751_, _02795_);
  not (_02797_, \oc8051_golden_model_1.IRAM[14] [1]);
  or (_02798_, _02653_, _02797_);
  and (_02799_, _02798_, _02757_);
  nand (_02800_, _02799_, _02796_);
  not (_02801_, \oc8051_golden_model_1.IRAM[12] [1]);
  or (_02802_, _02653_, _02801_);
  not (_02803_, \oc8051_golden_model_1.IRAM[13] [1]);
  or (_02804_, _02751_, _02803_);
  and (_02805_, _02804_, _02749_);
  nand (_02806_, _02805_, _02802_);
  nand (_02807_, _02806_, _02800_);
  nand (_02808_, _02807_, _02764_);
  nand (_02809_, _02808_, _02794_);
  nand (_02810_, _02809_, _02782_);
  nand (_02811_, _02810_, _02781_);
  not (_02812_, _02811_);
  or (_02813_, _02812_, _01886_);
  not (_02814_, _02001_);
  nor (_02815_, _02814_, _01790_);
  not (_02816_, _02815_);
  and (_02817_, _01884_, _01536_);
  not (_02818_, _02817_);
  nor (_02819_, _02818_, _01790_);
  and (_02820_, _01533_, _01857_);
  and (_02821_, _02820_, _01884_);
  nor (_02822_, _02821_, _02819_);
  not (_02823_, _01562_);
  and (_02824_, _02819_, _01823_);
  or (_02825_, _02824_, _02823_);
  or (_02826_, _02825_, _02822_);
  nor (_02827_, _01867_, _01562_);
  not (_02828_, _02827_);
  and (_02829_, _02049_, _01881_);
  nor (_02830_, _02829_, _02366_);
  and (_02831_, _02830_, _02828_);
  and (_02832_, _02831_, _02826_);
  and (_02833_, _02832_, _02816_);
  and (_02834_, _02833_, _02813_);
  and (_02835_, _02815_, _01823_);
  nor (_02836_, _02835_, _02834_);
  nor (_02837_, _02024_, _01790_);
  and (_02838_, _02837_, _01855_);
  nor (_02839_, _02838_, _02836_);
  not (_02840_, _01999_);
  nor (_02841_, _02840_, _01790_);
  nor (_02842_, _01867_, _01558_);
  nor (_02843_, _02842_, _02841_);
  and (_02844_, _02843_, _02839_);
  and (_02845_, _02841_, _01823_);
  nor (_02846_, _02845_, _02844_);
  and (_02847_, _02820_, _01877_);
  nor (_02848_, _02847_, _02846_);
  nor (_02849_, _02021_, _01790_);
  and (_02850_, _01882_, _01877_);
  and (_02851_, _02850_, _02811_);
  nor (_02852_, _02851_, _02849_);
  and (_02853_, _02852_, _02848_);
  and (_02854_, _02849_, _01823_);
  nor (_02855_, _02854_, _02853_);
  nor (_02856_, _02025_, _01790_);
  and (_02857_, _02856_, _01855_);
  nor (_02858_, _02857_, _02855_);
  and (_02859_, _02858_, _01880_);
  nor (_02860_, _02859_, _01879_);
  not (_02861_, _01991_);
  nor (_02862_, _02861_, _01790_);
  and (_02863_, _02862_, _01855_);
  or (_02864_, _02863_, _02860_);
  nor (_02865_, _01867_, _01565_);
  and (_02866_, _02820_, _01965_);
  nor (_02867_, _02866_, _02865_);
  not (_02868_, _02867_);
  nor (_02869_, _02868_, _02864_);
  nor (_02870_, _02408_, _01790_);
  and (_02871_, _01882_, _01965_);
  and (_02872_, _02811_, _02871_);
  nor (_02873_, _02872_, _02870_);
  and (_02874_, _02873_, _02869_);
  nor (_02875_, _02874_, _01876_);
  nor (_02876_, _02875_, _01604_);
  and (_02877_, _01867_, _01604_);
  nor (_02878_, _02877_, _02876_);
  nor (_02879_, _01790_, _02043_);
  not (_02880_, _02879_);
  nor (_02881_, _01790_, _02531_);
  or (_02882_, _02049_, _01978_);
  and (_02883_, _02882_, _02881_);
  nor (_02884_, _01983_, _02065_);
  not (_02885_, _02884_);
  and (_02886_, _02885_, _02881_);
  nor (_02887_, _02886_, _02883_);
  not (_02888_, _02528_);
  nor (_02889_, _02888_, _01790_);
  not (_02890_, _02889_);
  and (_02891_, _02890_, _02887_);
  and (_02892_, _02891_, _02880_);
  nor (_02893_, _02892_, _01823_);
  and (_02894_, _02358_, _01637_);
  and (_02895_, _02049_, _01637_);
  or (_02896_, _02895_, _02894_);
  or (_02897_, _02896_, _02893_);
  nor (_02898_, _02897_, _02878_);
  and (_02899_, _01882_, _01637_);
  and (_02900_, _02899_, _02811_);
  nor (_02901_, _02900_, _01871_);
  and (_02902_, _02901_, _02898_);
  nor (_02903_, _02902_, _01872_);
  nor (_02904_, _02903_, _01638_);
  and (_02905_, _01867_, _01638_);
  nor (_02906_, _02905_, _02904_);
  not (_02907_, _02177_);
  nor (_02908_, _02907_, _01790_);
  not (_02909_, _02908_);
  nor (_02910_, _02176_, _01790_);
  not (_02911_, _02910_);
  not (_02912_, _02167_);
  nor (_02913_, _02912_, _01790_);
  nor (_02914_, _02166_, _01790_);
  nor (_02915_, _02914_, _02913_);
  and (_02916_, _02915_, _02911_);
  and (_02917_, _02916_, _02909_);
  nor (_02918_, _02917_, _01823_);
  nor (_02919_, _02918_, _01632_);
  not (_02920_, _02919_);
  nor (_02921_, _02920_, _02906_);
  and (_02922_, _01867_, _01632_);
  nor (_02923_, _02922_, _02921_);
  nor (_02924_, _02174_, _01790_);
  and (_02925_, _02924_, _01822_);
  nor (_02926_, _02925_, _01636_);
  not (_02927_, _02926_);
  nor (_02928_, _02927_, _02923_);
  nor (_02929_, _02928_, _01868_);
  and (_02930_, _02049_, _01641_);
  nor (_02931_, _02930_, _02388_);
  not (_02932_, _02931_);
  nor (_02933_, _02932_, _02929_);
  nor (_02934_, _02303_, _01790_);
  and (_02935_, _01882_, _01641_);
  and (_02936_, _02811_, _02935_);
  nor (_02937_, _02936_, _02934_);
  and (_02938_, _02937_, _02933_);
  and (_02939_, _02934_, _01823_);
  nor (_02940_, _02939_, _02938_);
  nor (_02941_, _01887_, _01790_);
  nor (_02942_, _02058_, _01642_);
  nor (_02943_, _02942_, _01867_);
  nor (_02944_, _02943_, _02941_);
  not (_02945_, _02944_);
  nor (_02946_, _02945_, _02940_);
  nor (_02947_, _02946_, _01861_);
  and (_02948_, _02049_, _01403_);
  nor (_02949_, _02948_, _02386_);
  not (_02950_, _02949_);
  nor (_02951_, _02950_, _02947_);
  and (_02952_, _01882_, _01403_);
  and (_02953_, _02811_, _02952_);
  nor (_02954_, _02953_, _01791_);
  and (_02955_, _02954_, _02951_);
  nor (_02956_, _02955_, _01824_);
  not (_02957_, _02956_);
  not (_02958_, _02941_);
  and (_02959_, _02584_, _01871_);
  nor (_02960_, _01565_, _01864_);
  nor (_02961_, _02409_, _02861_);
  not (_02962_, _02862_);
  and (_02963_, _02819_, _02584_);
  nor (_02964_, _02963_, _02823_);
  nor (_02965_, _02495_, _01561_);
  nor (_02966_, _02965_, _02819_);
  not (_02967_, _02966_);
  and (_02968_, _02967_, _02964_);
  nor (_02969_, _01562_, _01864_);
  nor (_02970_, _02495_, _01557_);
  nor (_02971_, _02970_, _02969_);
  not (_02972_, _02971_);
  nor (_02973_, _02972_, _02968_);
  not (_02974_, _02973_);
  not (_02975_, \oc8051_golden_model_1.IRAM[0] [0]);
  or (_02976_, _02653_, _02975_);
  not (_02977_, \oc8051_golden_model_1.IRAM[1] [0]);
  or (_02978_, _02751_, _02977_);
  and (_02979_, _02978_, _02749_);
  nand (_02980_, _02979_, _02976_);
  not (_02981_, \oc8051_golden_model_1.IRAM[3] [0]);
  or (_02982_, _02751_, _02981_);
  not (_02983_, \oc8051_golden_model_1.IRAM[2] [0]);
  or (_02984_, _02653_, _02983_);
  and (_02985_, _02984_, _02757_);
  nand (_02986_, _02985_, _02982_);
  nand (_02987_, _02986_, _02980_);
  nand (_02988_, _02987_, _02406_);
  not (_02989_, \oc8051_golden_model_1.IRAM[7] [0]);
  or (_02990_, _02751_, _02989_);
  not (_02991_, \oc8051_golden_model_1.IRAM[6] [0]);
  or (_02992_, _02653_, _02991_);
  and (_02993_, _02992_, _02757_);
  nand (_02994_, _02993_, _02990_);
  not (_02995_, \oc8051_golden_model_1.IRAM[4] [0]);
  or (_02996_, _02653_, _02995_);
  not (_02997_, \oc8051_golden_model_1.IRAM[5] [0]);
  or (_02998_, _02751_, _02997_);
  and (_02999_, _02998_, _02749_);
  nand (_03000_, _02999_, _02996_);
  nand (_03001_, _03000_, _02994_);
  nand (_03002_, _03001_, _02764_);
  nand (_03003_, _03002_, _02988_);
  nand (_03004_, _03003_, _02221_);
  nand (_03005_, _02653_, \oc8051_golden_model_1.IRAM[11] [0]);
  nand (_03006_, _02751_, \oc8051_golden_model_1.IRAM[10] [0]);
  and (_03007_, _03006_, _02757_);
  nand (_03008_, _03007_, _03005_);
  not (_03009_, \oc8051_golden_model_1.IRAM[8] [0]);
  or (_03010_, _02653_, _03009_);
  nand (_03011_, _02653_, \oc8051_golden_model_1.IRAM[9] [0]);
  and (_03012_, _03011_, _02749_);
  nand (_03013_, _03012_, _03010_);
  nand (_03014_, _03013_, _03008_);
  nand (_03015_, _03014_, _02406_);
  nand (_03016_, _02653_, \oc8051_golden_model_1.IRAM[15] [0]);
  nand (_03017_, _02751_, \oc8051_golden_model_1.IRAM[14] [0]);
  and (_03018_, _03017_, _02757_);
  nand (_03019_, _03018_, _03016_);
  nand (_03020_, _02751_, \oc8051_golden_model_1.IRAM[12] [0]);
  nand (_03021_, _02653_, \oc8051_golden_model_1.IRAM[13] [0]);
  and (_03022_, _03021_, _02749_);
  nand (_03023_, _03022_, _03020_);
  nand (_03024_, _03023_, _03019_);
  nand (_03025_, _03024_, _02764_);
  nand (_03026_, _03025_, _03015_);
  nand (_03027_, _03026_, _02782_);
  and (_03028_, _03027_, _03004_);
  nor (_03029_, _03028_, _01886_);
  nor (_03030_, _03029_, _02974_);
  and (_03031_, _02815_, _02441_);
  nor (_03032_, _03031_, _02837_);
  and (_03033_, _03032_, _03030_);
  not (_03034_, _03033_);
  and (_03035_, _03034_, _02475_);
  nor (_03036_, _01558_, _01864_);
  nor (_03037_, _03036_, _03035_);
  and (_03038_, _02841_, _02441_);
  nor (_03039_, _02495_, _01573_);
  nor (_03040_, _03039_, _03038_);
  and (_03041_, _03040_, _03037_);
  nand (_03042_, _03027_, _03004_);
  and (_03043_, _03042_, _02850_);
  not (_03044_, _03043_);
  and (_03045_, _03044_, _03041_);
  and (_03046_, _02849_, _02441_);
  nor (_03047_, _03046_, _02856_);
  and (_03048_, _03047_, _03045_);
  nor (_03049_, _03048_, _02491_);
  or (_03050_, _03049_, _01878_);
  nand (_03051_, _01878_, _01864_);
  nand (_03052_, _03051_, _03050_);
  and (_03053_, _03052_, _02962_);
  nor (_03054_, _03053_, _02961_);
  nor (_03055_, _02495_, _01570_);
  or (_03056_, _03055_, _03054_);
  nor (_03057_, _03056_, _02960_);
  and (_03058_, _03042_, _02871_);
  nor (_03059_, _03058_, _02870_);
  and (_03060_, _03059_, _03057_);
  nor (_03061_, _03060_, _02410_);
  nor (_03062_, _03061_, _01604_);
  and (_03063_, _01604_, _01864_);
  nor (_03064_, _03063_, _03062_);
  nor (_03065_, _02892_, _02584_);
  and (_03066_, _02494_, _01637_);
  nor (_03067_, _03066_, _03065_);
  not (_03068_, _03067_);
  nor (_03069_, _03068_, _03064_);
  and (_03070_, _03042_, _02899_);
  nor (_03071_, _03070_, _01871_);
  and (_03072_, _03071_, _03069_);
  nor (_03073_, _03072_, _02959_);
  nor (_03074_, _03073_, _01638_);
  and (_03075_, _01638_, _01864_);
  nor (_03076_, _03075_, _03074_);
  nor (_03077_, _02917_, _02584_);
  nor (_03078_, _03077_, _01632_);
  not (_03079_, _03078_);
  nor (_03080_, _03079_, _03076_);
  and (_03081_, _01632_, _01864_);
  nor (_03082_, _03081_, _03080_);
  and (_03083_, _02924_, _02441_);
  nor (_03084_, _03083_, _01636_);
  not (_03085_, _03084_);
  nor (_03086_, _03085_, _03082_);
  and (_03087_, _01636_, _01864_);
  nor (_03088_, _03087_, _03086_);
  and (_03089_, _03042_, _02935_);
  and (_03090_, _02494_, _01641_);
  or (_03091_, _03090_, _02934_);
  or (_03092_, _03091_, _03089_);
  nor (_03093_, _03092_, _03088_);
  and (_03094_, _02934_, _02584_);
  nor (_03095_, _03094_, _03093_);
  nor (_03096_, _02942_, _01864_);
  nor (_03097_, _03096_, _03095_);
  and (_03098_, _03097_, _02958_);
  nor (_03099_, _03098_, _02636_);
  and (_03100_, _03042_, _02952_);
  and (_03101_, _02494_, _01403_);
  or (_03102_, _03101_, _01791_);
  or (_03103_, _03102_, _03100_);
  nor (_03104_, _03103_, _03099_);
  and (_03105_, _02584_, _01791_);
  nor (_03106_, _03105_, _03104_);
  nor (_03107_, _02879_, _02870_);
  nor (_03108_, _02934_, _02908_);
  and (_03109_, _03108_, _03107_);
  nor (_03110_, _02815_, _02837_);
  nor (_03111_, _02841_, _02819_);
  and (_03112_, _03111_, _03110_);
  and (_03113_, _03112_, _03109_);
  and (_03114_, _03113_, _02916_);
  nor (_03115_, _02862_, _01871_);
  nor (_03116_, _02849_, _02856_);
  and (_03117_, _03116_, _03115_);
  not (_03118_, _01791_);
  and (_03119_, _02690_, _01965_);
  not (_03120_, _03119_);
  and (_03121_, _02952_, _01434_);
  nor (_03122_, _01985_, _02065_);
  nor (_03123_, _03122_, _01573_);
  nor (_03124_, _03123_, _03121_);
  and (_03125_, _03124_, _03120_);
  not (_03126_, _02482_);
  and (_03127_, _02707_, _03126_);
  and (_03128_, _03127_, _02389_);
  nor (_03129_, _02899_, _02935_);
  and (_03130_, _03129_, _01563_);
  not (_03131_, _01565_);
  or (_03132_, _01604_, _03131_);
  not (_03133_, _03132_);
  and (_03134_, _03133_, _02942_);
  and (_03135_, _03134_, _03130_);
  and (_03136_, _03135_, _03128_);
  and (_03137_, _03136_, _03125_);
  not (_03138_, _02894_);
  not (_03139_, _01858_);
  and (_03140_, _01971_, _01637_);
  nand (_03141_, _03140_, _03139_);
  and (_03142_, _03141_, _03138_);
  and (_03143_, _02047_, _01403_);
  nor (_03144_, _03143_, _02948_);
  and (_03145_, _01972_, _01637_);
  and (_03146_, _02340_, _01637_);
  nor (_03147_, _03146_, _03145_);
  and (_03148_, _03147_, _03144_);
  and (_03149_, _03148_, _03142_);
  and (_03150_, _02368_, _01981_);
  and (_03151_, _02719_, _02343_);
  and (_03152_, _03151_, _03150_);
  nor (_03153_, _02394_, _01883_);
  nor (_03154_, _02829_, _01885_);
  and (_03155_, _03154_, _03153_);
  nor (_03156_, _02871_, _01878_);
  nor (_03157_, _02850_, _01984_);
  and (_03158_, _03157_, _03156_);
  and (_03159_, _03158_, _03155_);
  and (_03160_, _02049_, _01965_);
  nor (_03162_, _02930_, _03160_);
  nor (_03163_, _01982_, _01561_);
  and (_03164_, _01971_, _01884_);
  nor (_03165_, _03164_, _03163_);
  and (_03166_, _03165_, _03162_);
  and (_03167_, _03166_, _01640_);
  and (_03169_, _03167_, _03159_);
  and (_03170_, _03169_, _03152_);
  and (_03171_, _03170_, _03149_);
  and (_03173_, _03171_, _03137_);
  and (_03174_, _03173_, _03118_);
  nor (_03176_, _02924_, _02941_);
  and (_03177_, _03176_, _03174_);
  and (_03179_, _03177_, _03117_);
  and (_03180_, _03179_, _02891_);
  and (_03182_, _03180_, _03114_);
  and (_03183_, _38087_, _37580_);
  not (_03184_, _03183_);
  nor (_03186_, _03184_, _03182_);
  not (_03187_, _03186_);
  nor (_03189_, _03187_, _03106_);
  and (_03190_, _03189_, _02957_);
  not (_03192_, \oc8051_golden_model_1.IRAM[0] [3]);
  or (_03193_, _02653_, _03192_);
  not (_03195_, \oc8051_golden_model_1.IRAM[1] [3]);
  or (_03196_, _02751_, _03195_);
  and (_03197_, _03196_, _02749_);
  nand (_03198_, _03197_, _03193_);
  not (_03200_, \oc8051_golden_model_1.IRAM[3] [3]);
  or (_03201_, _02751_, _03200_);
  not (_03203_, \oc8051_golden_model_1.IRAM[2] [3]);
  or (_03204_, _02653_, _03203_);
  and (_03206_, _03204_, _02757_);
  nand (_03207_, _03206_, _03201_);
  nand (_03209_, _03207_, _03198_);
  nand (_03211_, _03209_, _02406_);
  not (_03213_, \oc8051_golden_model_1.IRAM[7] [3]);
  or (_03214_, _02751_, _03213_);
  not (_03216_, \oc8051_golden_model_1.IRAM[6] [3]);
  or (_03217_, _02653_, _03216_);
  and (_03219_, _03217_, _02757_);
  nand (_03221_, _03219_, _03214_);
  not (_03222_, \oc8051_golden_model_1.IRAM[4] [3]);
  or (_03224_, _02653_, _03222_);
  not (_03225_, \oc8051_golden_model_1.IRAM[5] [3]);
  or (_03227_, _02751_, _03225_);
  and (_03228_, _03227_, _02749_);
  nand (_03230_, _03228_, _03224_);
  nand (_03231_, _03230_, _03221_);
  nand (_03233_, _03231_, _02764_);
  nand (_03235_, _03233_, _03211_);
  nand (_03237_, _03235_, _02221_);
  nand (_03239_, _02653_, \oc8051_golden_model_1.IRAM[11] [3]);
  nand (_03241_, _02751_, \oc8051_golden_model_1.IRAM[10] [3]);
  and (_03243_, _03241_, _02757_);
  nand (_03245_, _03243_, _03239_);
  nand (_03247_, _02751_, \oc8051_golden_model_1.IRAM[8] [3]);
  nand (_03249_, _02653_, \oc8051_golden_model_1.IRAM[9] [3]);
  and (_03251_, _03249_, _02749_);
  nand (_03253_, _03251_, _03247_);
  nand (_03254_, _03253_, _03245_);
  nand (_03255_, _03254_, _02406_);
  nand (_03256_, _02653_, \oc8051_golden_model_1.IRAM[15] [3]);
  nand (_03257_, _02751_, \oc8051_golden_model_1.IRAM[14] [3]);
  and (_03258_, _03257_, _02757_);
  nand (_03259_, _03258_, _03256_);
  nand (_03260_, _02751_, \oc8051_golden_model_1.IRAM[12] [3]);
  nand (_03261_, _02653_, \oc8051_golden_model_1.IRAM[13] [3]);
  and (_03262_, _03261_, _02749_);
  nand (_03263_, _03262_, _03260_);
  nand (_03264_, _03263_, _03259_);
  nand (_03265_, _03264_, _02764_);
  nand (_03266_, _03265_, _03255_);
  nand (_03267_, _03266_, _02782_);
  nand (_03268_, _03267_, _03237_);
  and (_03269_, _03268_, _02952_);
  and (_03270_, _03268_, _02935_);
  and (_03271_, _03268_, _02899_);
  and (_03272_, \oc8051_golden_model_1.SP [1], \oc8051_golden_model_1.SP [0]);
  and (_03273_, _03272_, \oc8051_golden_model_1.SP [2]);
  nor (_03274_, _03273_, \oc8051_golden_model_1.SP [3]);
  and (_03275_, _03273_, \oc8051_golden_model_1.SP [3]);
  nor (_03276_, _03275_, _03274_);
  not (_03277_, _03276_);
  nor (_03278_, _03277_, _01565_);
  not (_03279_, _01558_);
  and (_03280_, _02837_, _01922_);
  nor (_03281_, _03277_, _01562_);
  nor (_03282_, _01885_, \oc8051_golden_model_1.PSW [3]);
  and (_03283_, _03268_, _01885_);
  nor (_03284_, _03283_, _03282_);
  nor (_03285_, _03284_, _02819_);
  and (_03286_, _02819_, _01954_);
  nor (_03287_, _03286_, _02823_);
  not (_03288_, _03287_);
  nor (_03289_, _03288_, _03285_);
  or (_03290_, _03289_, _01883_);
  nor (_03291_, _03290_, _03281_);
  and (_03292_, _03268_, _01883_);
  nor (_03293_, _03292_, _02815_);
  not (_03294_, _03293_);
  nor (_03295_, _03294_, _03291_);
  nor (_03296_, _02409_, _02814_);
  or (_03297_, _03296_, _02837_);
  nor (_03298_, _03297_, _03295_);
  nor (_03299_, _03298_, _03280_);
  nor (_03300_, _03299_, _03279_);
  nor (_03301_, _03276_, _01558_);
  nor (_03302_, _03301_, _02841_);
  not (_03303_, _03302_);
  nor (_03304_, _03303_, _03300_);
  and (_03305_, _02841_, _01955_);
  nor (_03306_, _03305_, _02850_);
  not (_03307_, _03306_);
  nor (_03308_, _03307_, _03304_);
  and (_03309_, _03268_, _02850_);
  nor (_03310_, _03309_, _02849_);
  not (_03311_, _03310_);
  nor (_03312_, _03311_, _03308_);
  and (_03313_, _02849_, _01955_);
  or (_03314_, _03313_, _02856_);
  nor (_03315_, _03314_, _03312_);
  and (_03316_, _02856_, _01922_);
  nor (_03317_, _03316_, _03315_);
  and (_03318_, _03317_, _01880_);
  and (_03319_, _03276_, _01878_);
  nor (_03320_, _03319_, _03318_);
  nor (_03321_, _03320_, _02862_);
  nor (_03322_, _01957_, _02962_);
  or (_03323_, _03322_, _03321_);
  and (_03324_, _03323_, _01565_);
  or (_03325_, _03324_, _02871_);
  nor (_03326_, _03325_, _03278_);
  and (_03327_, _03268_, _02871_);
  nor (_03328_, _03327_, _02870_);
  not (_03329_, _03328_);
  nor (_03330_, _03329_, _03326_);
  and (_03331_, _01923_, _01875_);
  nor (_03332_, _03331_, _03330_);
  nor (_03333_, _03332_, _01604_);
  and (_03334_, _03276_, _01604_);
  not (_03335_, _03334_);
  and (_03336_, _03335_, _02892_);
  not (_03337_, _03336_);
  nor (_03338_, _03337_, _03333_);
  nor (_03339_, _02892_, _01955_);
  nor (_03340_, _03339_, _03338_);
  nor (_03341_, _03340_, _02899_);
  or (_03342_, _03341_, _01871_);
  nor (_03343_, _03342_, _03271_);
  and (_03344_, _01955_, _01871_);
  nor (_03345_, _03344_, _03343_);
  nor (_03346_, _03345_, _01638_);
  and (_03347_, _03276_, _01638_);
  not (_03348_, _03347_);
  and (_03349_, _03348_, _02917_);
  not (_03350_, _03349_);
  nor (_03351_, _03350_, _03346_);
  nor (_03352_, _02917_, _01955_);
  nor (_03353_, _03352_, _01632_);
  not (_03354_, _03353_);
  nor (_03355_, _03354_, _03351_);
  and (_03356_, _03276_, _01632_);
  nor (_03357_, _03356_, _02924_);
  not (_03358_, _03357_);
  nor (_03359_, _03358_, _03355_);
  and (_03360_, _02924_, _01954_);
  nor (_03361_, _03360_, _01636_);
  not (_03362_, _03361_);
  nor (_03363_, _03362_, _03359_);
  and (_03364_, _03276_, _01636_);
  nor (_03365_, _03364_, _02935_);
  not (_03366_, _03365_);
  nor (_03367_, _03366_, _03363_);
  or (_03368_, _03367_, _02934_);
  nor (_03369_, _03368_, _03270_);
  not (_03370_, _02942_);
  and (_03371_, _02934_, _01955_);
  nor (_03372_, _03371_, _03370_);
  not (_03373_, _03372_);
  nor (_03374_, _03373_, _03369_);
  nor (_03375_, _03276_, _02942_);
  nor (_03376_, _03375_, _02941_);
  not (_03377_, _03376_);
  nor (_03378_, _03377_, _03374_);
  not (_03379_, _01922_);
  and (_03380_, _02941_, _03379_);
  or (_03381_, _03380_, _02952_);
  nor (_03382_, _03381_, _03378_);
  or (_03383_, _03382_, _01791_);
  nor (_03384_, _03383_, _03269_);
  and (_03385_, _01955_, _01791_);
  nor (_03386_, _03385_, _03384_);
  and (_03387_, _02253_, _01860_);
  nor (_03388_, _03272_, \oc8051_golden_model_1.SP [2]);
  nor (_03389_, _03388_, _03273_);
  and (_03390_, _03389_, _01636_);
  not (_03391_, _02294_);
  and (_03392_, _03391_, _01871_);
  nor (_03393_, _02892_, _03391_);
  and (_03394_, _02253_, _01875_);
  and (_03395_, _03389_, _01878_);
  and (_03396_, _01971_, _01877_);
  not (_03397_, \oc8051_golden_model_1.IRAM[0] [2]);
  or (_03398_, _02653_, _03397_);
  not (_03399_, \oc8051_golden_model_1.IRAM[1] [2]);
  or (_03400_, _02751_, _03399_);
  and (_03401_, _03400_, _02749_);
  nand (_03402_, _03401_, _03398_);
  not (_03403_, \oc8051_golden_model_1.IRAM[3] [2]);
  or (_03404_, _02751_, _03403_);
  not (_03405_, \oc8051_golden_model_1.IRAM[2] [2]);
  or (_03406_, _02653_, _03405_);
  and (_03407_, _03406_, _02757_);
  nand (_03408_, _03407_, _03404_);
  nand (_03409_, _03408_, _03402_);
  nand (_03410_, _03409_, _02406_);
  not (_03411_, \oc8051_golden_model_1.IRAM[7] [2]);
  or (_03412_, _02751_, _03411_);
  not (_03413_, \oc8051_golden_model_1.IRAM[6] [2]);
  or (_03414_, _02653_, _03413_);
  and (_03415_, _03414_, _02757_);
  nand (_03416_, _03415_, _03412_);
  not (_03417_, \oc8051_golden_model_1.IRAM[4] [2]);
  or (_03418_, _02653_, _03417_);
  not (_03419_, \oc8051_golden_model_1.IRAM[5] [2]);
  or (_03420_, _02751_, _03419_);
  and (_03421_, _03420_, _02749_);
  nand (_03422_, _03421_, _03418_);
  nand (_03423_, _03422_, _03416_);
  nand (_03424_, _03423_, _02764_);
  nand (_03425_, _03424_, _03410_);
  nand (_03426_, _03425_, _02221_);
  nand (_03427_, _02653_, \oc8051_golden_model_1.IRAM[11] [2]);
  not (_03428_, \oc8051_golden_model_1.IRAM[10] [2]);
  or (_03429_, _02653_, _03428_);
  and (_03430_, _03429_, _02757_);
  nand (_03431_, _03430_, _03427_);
  not (_03432_, \oc8051_golden_model_1.IRAM[8] [2]);
  or (_03433_, _02653_, _03432_);
  nand (_03434_, _02653_, \oc8051_golden_model_1.IRAM[9] [2]);
  and (_03435_, _03434_, _02749_);
  nand (_03436_, _03435_, _03433_);
  nand (_03437_, _03436_, _03431_);
  nand (_03438_, _03437_, _02406_);
  not (_03439_, \oc8051_golden_model_1.IRAM[15] [2]);
  or (_03440_, _02751_, _03439_);
  not (_03441_, \oc8051_golden_model_1.IRAM[14] [2]);
  or (_03442_, _02653_, _03441_);
  and (_03443_, _03442_, _02757_);
  nand (_03444_, _03443_, _03440_);
  not (_03445_, \oc8051_golden_model_1.IRAM[12] [2]);
  or (_03446_, _02653_, _03445_);
  not (_03447_, \oc8051_golden_model_1.IRAM[13] [2]);
  or (_03448_, _02751_, _03447_);
  and (_03449_, _03448_, _02749_);
  nand (_03450_, _03449_, _03446_);
  nand (_03451_, _03450_, _03444_);
  nand (_03452_, _03451_, _02764_);
  nand (_03453_, _03452_, _03438_);
  nand (_03454_, _03453_, _02782_);
  nand (_03455_, _03454_, _03426_);
  not (_03456_, _03455_);
  or (_03457_, _03456_, _01886_);
  nor (_03458_, _03164_, _02819_);
  and (_03459_, _02819_, _03391_);
  or (_03460_, _03459_, _02823_);
  or (_03461_, _03460_, _03458_);
  nor (_03462_, _03389_, _01562_);
  and (_03463_, _01971_, _01881_);
  nor (_03464_, _03463_, _03462_);
  and (_03465_, _03464_, _03461_);
  and (_03466_, _03465_, _02816_);
  and (_03467_, _03466_, _03457_);
  and (_03468_, _02815_, _03391_);
  nor (_03469_, _03468_, _03467_);
  and (_03470_, _02837_, _02252_);
  nor (_03471_, _03470_, _03469_);
  nor (_03472_, _03389_, _01558_);
  nor (_03473_, _03472_, _02841_);
  and (_03474_, _03473_, _03471_);
  and (_03475_, _02841_, _03391_);
  nor (_03476_, _03475_, _03474_);
  nor (_03477_, _03476_, _03396_);
  and (_03478_, _03455_, _02850_);
  nor (_03479_, _03478_, _02849_);
  and (_03480_, _03479_, _03477_);
  and (_03481_, _02849_, _03391_);
  nor (_03482_, _03481_, _03480_);
  and (_03483_, _02856_, _02252_);
  nor (_03484_, _03483_, _03482_);
  and (_03485_, _03484_, _01880_);
  nor (_03486_, _03485_, _03395_);
  and (_03487_, _02252_, _02862_);
  or (_03488_, _03487_, _03486_);
  and (_03489_, _01971_, _01965_);
  nor (_03490_, _03389_, _01565_);
  nor (_03491_, _03490_, _03489_);
  not (_03492_, _03491_);
  nor (_03493_, _03492_, _03488_);
  and (_03494_, _03455_, _02871_);
  nor (_03495_, _03494_, _02870_);
  and (_03496_, _03495_, _03493_);
  nor (_03497_, _03496_, _03394_);
  nor (_03498_, _03497_, _01604_);
  and (_03499_, _03389_, _01604_);
  nor (_03500_, _03499_, _03498_);
  or (_03501_, _03500_, _03140_);
  nor (_03502_, _03501_, _03393_);
  and (_03503_, _03455_, _02899_);
  nor (_03504_, _03503_, _01871_);
  and (_03505_, _03504_, _03502_);
  nor (_03506_, _03505_, _03392_);
  nor (_03507_, _03506_, _01638_);
  and (_03508_, _03389_, _01638_);
  nor (_03509_, _03508_, _03507_);
  nor (_03510_, _02917_, _03391_);
  nor (_03511_, _03510_, _01632_);
  not (_03512_, _03511_);
  nor (_03513_, _03512_, _03509_);
  and (_03514_, _03389_, _01632_);
  nor (_03515_, _03514_, _03513_);
  and (_03516_, _02924_, _02294_);
  nor (_03517_, _03516_, _01636_);
  not (_03518_, _03517_);
  nor (_03519_, _03518_, _03515_);
  nor (_03520_, _03519_, _03390_);
  and (_03521_, _01971_, _01641_);
  nor (_03522_, _03521_, _03520_);
  and (_03523_, _03455_, _02935_);
  nor (_03524_, _03523_, _02934_);
  and (_03525_, _03524_, _03522_);
  and (_03526_, _02934_, _03391_);
  nor (_03527_, _03526_, _03525_);
  nor (_03528_, _03389_, _02942_);
  nor (_03529_, _03528_, _02941_);
  not (_03530_, _03529_);
  nor (_03531_, _03530_, _03527_);
  nor (_03532_, _03531_, _03387_);
  and (_03533_, _01971_, _01403_);
  nor (_03534_, _03533_, _03532_);
  and (_03535_, _03455_, _02952_);
  nor (_03536_, _03535_, _01791_);
  and (_03537_, _03536_, _03534_);
  and (_03538_, _03391_, _01791_);
  nor (_03539_, _03538_, _03537_);
  nor (_03540_, _03539_, _03187_);
  not (_03541_, _03540_);
  nor (_03542_, _03541_, _03386_);
  and (_03543_, _03542_, _03190_);
  or (_03544_, _03543_, \oc8051_golden_model_1.IRAM[15] [7]);
  and (_03545_, \oc8051_golden_model_1.SP [2], \oc8051_golden_model_1.SP [1]);
  and (_03546_, _03545_, _01864_);
  nor (_03547_, _03389_, _01865_);
  nor (_03548_, _03547_, _03546_);
  and (_03549_, _03545_, \oc8051_golden_model_1.SP [3]);
  and (_03550_, _03549_, _01864_);
  nor (_03551_, _03546_, _03276_);
  nor (_03552_, _03551_, _03550_);
  and (_03553_, _02942_, _01563_);
  and (_03554_, _03553_, _03133_);
  and (_03555_, _03554_, _01640_);
  nor (_03556_, _03555_, _03184_);
  and (_03557_, _03556_, _03552_);
  and (_03558_, _03557_, _03548_);
  and (_03559_, _03558_, _01863_);
  not (_03560_, _03559_);
  and (_03561_, _03560_, _03544_);
  not (_03562_, _03543_);
  not (_03563_, \oc8051_golden_model_1.IRAM[0] [7]);
  or (_03564_, _02653_, _03563_);
  not (_03565_, \oc8051_golden_model_1.IRAM[1] [7]);
  or (_03566_, _02751_, _03565_);
  and (_03567_, _03566_, _02749_);
  nand (_03568_, _03567_, _03564_);
  not (_03569_, \oc8051_golden_model_1.IRAM[3] [7]);
  or (_03570_, _02751_, _03569_);
  not (_03571_, \oc8051_golden_model_1.IRAM[2] [7]);
  or (_03572_, _02653_, _03571_);
  and (_03573_, _03572_, _02757_);
  nand (_03574_, _03573_, _03570_);
  nand (_03575_, _03574_, _03568_);
  nand (_03576_, _03575_, _02406_);
  not (_03577_, \oc8051_golden_model_1.IRAM[7] [7]);
  or (_03578_, _02751_, _03577_);
  not (_03579_, \oc8051_golden_model_1.IRAM[6] [7]);
  or (_03580_, _02653_, _03579_);
  and (_03581_, _03580_, _02757_);
  nand (_03582_, _03581_, _03578_);
  not (_03583_, \oc8051_golden_model_1.IRAM[4] [7]);
  or (_03584_, _02653_, _03583_);
  not (_03585_, \oc8051_golden_model_1.IRAM[5] [7]);
  or (_03586_, _02751_, _03585_);
  and (_03587_, _03586_, _02749_);
  nand (_03588_, _03587_, _03584_);
  nand (_03589_, _03588_, _03582_);
  nand (_03590_, _03589_, _02764_);
  nand (_03591_, _03590_, _03576_);
  nand (_03592_, _03591_, _02221_);
  nand (_03593_, _02653_, \oc8051_golden_model_1.IRAM[11] [7]);
  not (_03594_, \oc8051_golden_model_1.IRAM[10] [7]);
  or (_03595_, _02653_, _03594_);
  and (_03596_, _03595_, _02757_);
  nand (_03597_, _03596_, _03593_);
  nand (_03598_, _02751_, \oc8051_golden_model_1.IRAM[8] [7]);
  nand (_03599_, _02653_, \oc8051_golden_model_1.IRAM[9] [7]);
  and (_03600_, _03599_, _02749_);
  nand (_03601_, _03600_, _03598_);
  nand (_03602_, _03601_, _03597_);
  nand (_03603_, _03602_, _02406_);
  nand (_03604_, _02653_, \oc8051_golden_model_1.IRAM[15] [7]);
  nand (_03605_, _02751_, \oc8051_golden_model_1.IRAM[14] [7]);
  and (_03606_, _03605_, _02757_);
  nand (_03607_, _03606_, _03604_);
  nand (_03608_, _02751_, \oc8051_golden_model_1.IRAM[12] [7]);
  nand (_03609_, _02653_, \oc8051_golden_model_1.IRAM[13] [7]);
  and (_03610_, _03609_, _02749_);
  nand (_03611_, _03610_, _03608_);
  nand (_03612_, _03611_, _03607_);
  nand (_03613_, _03612_, _02764_);
  nand (_03614_, _03613_, _03603_);
  nand (_03615_, _03614_, _02782_);
  nand (_03616_, _03615_, _03592_);
  or (_03617_, _03616_, _01790_);
  and (_03618_, _02584_, _01822_);
  and (_03619_, _03618_, _02294_);
  and (_03620_, _03619_, _01955_);
  and (_03621_, _01922_, _01790_);
  not (_03622_, _01855_);
  and (_03623_, _02252_, _03622_);
  and (_03624_, _03623_, _03621_);
  and (_03625_, _03624_, _03620_);
  and (_03626_, _03625_, \oc8051_golden_model_1.SBUF [7]);
  and (_03627_, _02441_, _01822_);
  and (_03628_, _03627_, _02294_);
  and (_03629_, _03628_, _01955_);
  not (_03630_, _02252_);
  and (_03631_, _03630_, _01855_);
  and (_03632_, _03631_, _03621_);
  and (_03633_, _03632_, _03629_);
  and (_03634_, _03633_, \oc8051_golden_model_1.IE [7]);
  nor (_03636_, _03634_, _03626_);
  nor (_03638_, _02252_, _01855_);
  and (_03640_, _03638_, _03621_);
  and (_03642_, _02294_, _01954_);
  and (_03644_, _03642_, _03627_);
  and (_03646_, _03644_, _03640_);
  and (_03648_, _03646_, \oc8051_golden_model_1.P3 [7]);
  not (_03650_, _03648_);
  and (_03652_, _03621_, _02252_);
  and (_03654_, _03652_, _01855_);
  and (_03656_, _03654_, _01954_);
  nor (_03658_, _02441_, _01822_);
  and (_03660_, _03658_, _03391_);
  and (_03662_, _03660_, _03656_);
  and (_03664_, _03662_, \oc8051_golden_model_1.PCON [7]);
  and (_03665_, _03644_, _03632_);
  and (_03666_, _03665_, \oc8051_golden_model_1.P2 [7]);
  nor (_03667_, _03666_, _03664_);
  and (_03668_, _03667_, _03650_);
  and (_03669_, _03668_, _03636_);
  and (_03670_, _03640_, _03629_);
  and (_03671_, _03670_, \oc8051_golden_model_1.IP [7]);
  not (_03672_, _03671_);
  not (_03673_, _01790_);
  nor (_03674_, _01922_, _03673_);
  and (_03675_, _03674_, _03623_);
  and (_03676_, _03675_, _03644_);
  and (_03677_, _03676_, \oc8051_golden_model_1.PSW [7]);
  not (_03678_, _03677_);
  and (_03679_, _03674_, _03631_);
  and (_03680_, _03679_, _03644_);
  and (_03681_, _03680_, \oc8051_golden_model_1.ACC [7]);
  and (_03682_, _03674_, _03638_);
  and (_03683_, _03682_, _03644_);
  and (_03684_, _03683_, \oc8051_golden_model_1.B [7]);
  nor (_03685_, _03684_, _03681_);
  and (_03686_, _03685_, _03678_);
  and (_03687_, _03686_, _03672_);
  not (_03688_, _03654_);
  nor (_03689_, _02294_, _01954_);
  nand (_03690_, _03689_, _03627_);
  nor (_03691_, _03690_, _03688_);
  and (_03692_, _03691_, \oc8051_golden_model_1.TH0 [7]);
  and (_03693_, _03629_, _03654_);
  and (_03694_, _03693_, \oc8051_golden_model_1.TCON [7]);
  nor (_03696_, _03694_, _03692_);
  and (_03698_, _03644_, _03624_);
  and (_03700_, _03698_, \oc8051_golden_model_1.P1 [7]);
  not (_03702_, _03658_);
  nand (_03704_, _02294_, _01955_);
  or (_03706_, _03704_, _03702_);
  nor (_03708_, _03706_, _03688_);
  and (_03710_, _03708_, \oc8051_golden_model_1.TL1 [7]);
  nor (_03712_, _03710_, _03700_);
  and (_03714_, _03712_, _03696_);
  and (_03716_, _03624_, _03629_);
  and (_03718_, _03716_, \oc8051_golden_model_1.SCON [7]);
  nand (_03720_, _03689_, _03618_);
  nor (_03722_, _03720_, _03688_);
  and (_03724_, _03722_, \oc8051_golden_model_1.TH1 [7]);
  nor (_03725_, _03724_, _03718_);
  and (_03726_, _03620_, _03654_);
  and (_03727_, _03726_, \oc8051_golden_model_1.TMOD [7]);
  nor (_03728_, _02584_, _01822_);
  nor (_03729_, _03704_, _03688_);
  and (_03730_, _03729_, _03728_);
  and (_03731_, _03730_, \oc8051_golden_model_1.TL0 [7]);
  nor (_03732_, _03731_, _03727_);
  and (_03733_, _03732_, _03725_);
  and (_03734_, _03733_, _03714_);
  and (_03735_, _03734_, _03687_);
  and (_03736_, _03735_, _03669_);
  and (_03737_, _03644_, _03654_);
  and (_03738_, _03737_, \oc8051_golden_model_1.P0 [7]);
  not (_03739_, _03738_);
  nand (_03740_, _03642_, _03658_);
  nor (_03741_, _03740_, _03688_);
  and (_03742_, _03741_, \oc8051_golden_model_1.DPH [7]);
  not (_03743_, _03742_);
  and (_03744_, _03642_, _03618_);
  and (_03745_, _03744_, _03654_);
  and (_03746_, _03745_, \oc8051_golden_model_1.SP [7]);
  nand (_03747_, _03642_, _03728_);
  nor (_03748_, _03747_, _03688_);
  and (_03749_, _03748_, \oc8051_golden_model_1.DPL [7]);
  nor (_03750_, _03749_, _03746_);
  and (_03751_, _03750_, _03743_);
  and (_03752_, _03751_, _03739_);
  and (_03753_, _03752_, _03736_);
  and (_03754_, _03753_, _03617_);
  not (_03755_, _03754_);
  not (_03756_, \oc8051_golden_model_1.IRAM[0] [6]);
  or (_03757_, _02653_, _03756_);
  not (_03758_, \oc8051_golden_model_1.IRAM[1] [6]);
  or (_03759_, _02751_, _03758_);
  and (_03760_, _03759_, _02749_);
  nand (_03761_, _03760_, _03757_);
  not (_03762_, \oc8051_golden_model_1.IRAM[3] [6]);
  or (_03763_, _02751_, _03762_);
  not (_03764_, \oc8051_golden_model_1.IRAM[2] [6]);
  or (_03765_, _02653_, _03764_);
  and (_03766_, _03765_, _02757_);
  nand (_03767_, _03766_, _03763_);
  nand (_03768_, _03767_, _03761_);
  nand (_03769_, _03768_, _02406_);
  not (_03770_, \oc8051_golden_model_1.IRAM[7] [6]);
  or (_03771_, _02751_, _03770_);
  not (_03772_, \oc8051_golden_model_1.IRAM[6] [6]);
  or (_03773_, _02653_, _03772_);
  and (_03774_, _03773_, _02757_);
  nand (_03775_, _03774_, _03771_);
  not (_03776_, \oc8051_golden_model_1.IRAM[4] [6]);
  or (_03777_, _02653_, _03776_);
  not (_03778_, \oc8051_golden_model_1.IRAM[5] [6]);
  or (_03779_, _02751_, _03778_);
  and (_03780_, _03779_, _02749_);
  nand (_03781_, _03780_, _03777_);
  nand (_03782_, _03781_, _03775_);
  nand (_03783_, _03782_, _02764_);
  nand (_03784_, _03783_, _03769_);
  nand (_03785_, _03784_, _02221_);
  nand (_03786_, _02653_, \oc8051_golden_model_1.IRAM[11] [6]);
  nand (_03787_, _02751_, \oc8051_golden_model_1.IRAM[10] [6]);
  and (_03788_, _03787_, _02757_);
  nand (_03789_, _03788_, _03786_);
  nand (_03790_, _02751_, \oc8051_golden_model_1.IRAM[8] [6]);
  nand (_03791_, _02653_, \oc8051_golden_model_1.IRAM[9] [6]);
  and (_03792_, _03791_, _02749_);
  nand (_03793_, _03792_, _03790_);
  nand (_03794_, _03793_, _03789_);
  nand (_03795_, _03794_, _02406_);
  nand (_03796_, _02653_, \oc8051_golden_model_1.IRAM[15] [6]);
  nand (_03797_, _02751_, \oc8051_golden_model_1.IRAM[14] [6]);
  and (_03798_, _03797_, _02757_);
  nand (_03799_, _03798_, _03796_);
  nand (_03800_, _02751_, \oc8051_golden_model_1.IRAM[12] [6]);
  nand (_03801_, _02653_, \oc8051_golden_model_1.IRAM[13] [6]);
  and (_03802_, _03801_, _02749_);
  nand (_03803_, _03802_, _03800_);
  nand (_03804_, _03803_, _03799_);
  nand (_03805_, _03804_, _02764_);
  nand (_03806_, _03805_, _03795_);
  nand (_03807_, _03806_, _02782_);
  nand (_03808_, _03807_, _03785_);
  or (_03809_, _03808_, _01790_);
  and (_03810_, _03662_, \oc8051_golden_model_1.PCON [6]);
  not (_03811_, _03810_);
  and (_03812_, _03625_, \oc8051_golden_model_1.SBUF [6]);
  and (_03813_, _03633_, \oc8051_golden_model_1.IE [6]);
  nor (_03814_, _03813_, _03812_);
  and (_03815_, _03814_, _03811_);
  and (_03816_, _03693_, \oc8051_golden_model_1.TCON [6]);
  not (_03817_, _03816_);
  and (_03818_, _03698_, \oc8051_golden_model_1.P1 [6]);
  not (_03819_, _03818_);
  and (_03820_, _03665_, \oc8051_golden_model_1.P2 [6]);
  and (_03821_, _03646_, \oc8051_golden_model_1.P3 [6]);
  nor (_03822_, _03821_, _03820_);
  and (_03823_, _03822_, _03819_);
  and (_03824_, _03823_, _03817_);
  and (_03825_, _03670_, \oc8051_golden_model_1.IP [6]);
  and (_03826_, _03683_, \oc8051_golden_model_1.B [6]);
  nor (_03827_, _03826_, _03825_);
  and (_03828_, _03676_, \oc8051_golden_model_1.PSW [6]);
  and (_03829_, _03680_, \oc8051_golden_model_1.ACC [6]);
  nor (_03830_, _03829_, _03828_);
  and (_03831_, _03830_, _03827_);
  and (_03832_, _03628_, _03656_);
  nand (_03833_, _03832_, \oc8051_golden_model_1.P0 [6]);
  and (_03834_, _03833_, _03831_);
  and (_03835_, _03834_, _03824_);
  and (_03836_, _03835_, _03815_);
  and (_03837_, _03726_, \oc8051_golden_model_1.TMOD [6]);
  and (_03838_, _03716_, \oc8051_golden_model_1.SCON [6]);
  nor (_03839_, _03838_, _03837_);
  and (_03840_, _03691_, \oc8051_golden_model_1.TH0 [6]);
  and (_03841_, _03722_, \oc8051_golden_model_1.TH1 [6]);
  nor (_03842_, _03841_, _03840_);
  and (_03843_, _03842_, _03839_);
  and (_03844_, _03730_, \oc8051_golden_model_1.TL0 [6]);
  and (_03845_, _03729_, _03658_);
  and (_03846_, _03845_, \oc8051_golden_model_1.TL1 [6]);
  nor (_03847_, _03846_, _03844_);
  and (_03848_, _03847_, _03843_);
  and (_03849_, _03658_, _02294_);
  and (_03850_, _03849_, _03656_);
  and (_03851_, _03850_, \oc8051_golden_model_1.DPH [6]);
  not (_03852_, _03851_);
  and (_03853_, _03619_, _03656_);
  and (_03854_, _03853_, \oc8051_golden_model_1.SP [6]);
  and (_03855_, _03728_, _02294_);
  and (_03856_, _03855_, _03656_);
  and (_03857_, _03856_, \oc8051_golden_model_1.DPL [6]);
  nor (_03858_, _03857_, _03854_);
  and (_03859_, _03858_, _03852_);
  and (_03860_, _03859_, _03848_);
  and (_03861_, _03860_, _03836_);
  and (_03862_, _03861_, _03809_);
  not (_03863_, _03862_);
  not (_03864_, \oc8051_golden_model_1.IRAM[0] [5]);
  or (_03865_, _02653_, _03864_);
  not (_03866_, \oc8051_golden_model_1.IRAM[1] [5]);
  or (_03867_, _02751_, _03866_);
  and (_03868_, _03867_, _02749_);
  nand (_03869_, _03868_, _03865_);
  not (_03870_, \oc8051_golden_model_1.IRAM[3] [5]);
  or (_03871_, _02751_, _03870_);
  not (_03872_, \oc8051_golden_model_1.IRAM[2] [5]);
  or (_03873_, _02653_, _03872_);
  and (_03874_, _03873_, _02757_);
  nand (_03875_, _03874_, _03871_);
  nand (_03876_, _03875_, _03869_);
  nand (_03877_, _03876_, _02406_);
  not (_03878_, \oc8051_golden_model_1.IRAM[7] [5]);
  or (_03879_, _02751_, _03878_);
  not (_03880_, \oc8051_golden_model_1.IRAM[6] [5]);
  or (_03881_, _02653_, _03880_);
  and (_03882_, _03881_, _02757_);
  nand (_03883_, _03882_, _03879_);
  not (_03884_, \oc8051_golden_model_1.IRAM[4] [5]);
  or (_03885_, _02653_, _03884_);
  not (_03886_, \oc8051_golden_model_1.IRAM[5] [5]);
  or (_03887_, _02751_, _03886_);
  and (_03888_, _03887_, _02749_);
  nand (_03889_, _03888_, _03885_);
  nand (_03890_, _03889_, _03883_);
  nand (_03891_, _03890_, _02764_);
  nand (_03892_, _03891_, _03877_);
  nand (_03893_, _03892_, _02221_);
  nand (_03894_, _02653_, \oc8051_golden_model_1.IRAM[11] [5]);
  nand (_03895_, _02751_, \oc8051_golden_model_1.IRAM[10] [5]);
  and (_03896_, _03895_, _02757_);
  nand (_03897_, _03896_, _03894_);
  nand (_03898_, _02751_, \oc8051_golden_model_1.IRAM[8] [5]);
  nand (_03899_, _02653_, \oc8051_golden_model_1.IRAM[9] [5]);
  and (_03900_, _03899_, _02749_);
  nand (_03901_, _03900_, _03898_);
  nand (_03902_, _03901_, _03897_);
  nand (_03903_, _03902_, _02406_);
  nand (_03904_, _02653_, \oc8051_golden_model_1.IRAM[15] [5]);
  nand (_03905_, _02751_, \oc8051_golden_model_1.IRAM[14] [5]);
  and (_03906_, _03905_, _02757_);
  nand (_03907_, _03906_, _03904_);
  nand (_03908_, _02751_, \oc8051_golden_model_1.IRAM[12] [5]);
  nand (_03909_, _02653_, \oc8051_golden_model_1.IRAM[13] [5]);
  and (_03910_, _03909_, _02749_);
  nand (_03911_, _03910_, _03908_);
  nand (_03912_, _03911_, _03907_);
  nand (_03913_, _03912_, _02764_);
  nand (_03914_, _03913_, _03903_);
  nand (_03915_, _03914_, _02782_);
  nand (_03916_, _03915_, _03893_);
  or (_03917_, _03916_, _01790_);
  and (_03918_, _03850_, \oc8051_golden_model_1.DPH [5]);
  not (_03919_, _03918_);
  and (_03920_, _03853_, \oc8051_golden_model_1.SP [5]);
  and (_03921_, _03856_, \oc8051_golden_model_1.DPL [5]);
  nor (_03922_, _03921_, _03920_);
  and (_03923_, _03922_, _03919_);
  and (_03924_, _03625_, \oc8051_golden_model_1.SBUF [5]);
  not (_03925_, _03924_);
  and (_03926_, _03726_, \oc8051_golden_model_1.TMOD [5]);
  and (_03927_, _03716_, \oc8051_golden_model_1.SCON [5]);
  nor (_03928_, _03927_, _03926_);
  and (_03929_, _03928_, _03925_);
  and (_03930_, _03730_, \oc8051_golden_model_1.TL0 [5]);
  not (_03931_, _03930_);
  and (_03932_, _03722_, \oc8051_golden_model_1.TH1 [5]);
  and (_03933_, _03633_, \oc8051_golden_model_1.IE [5]);
  nor (_03934_, _03933_, _03932_);
  and (_03935_, _03934_, _03931_);
  and (_03936_, _03935_, _03929_);
  and (_03937_, _03936_, _03923_);
  and (_03938_, _03693_, \oc8051_golden_model_1.TCON [5]);
  and (_03939_, _03691_, \oc8051_golden_model_1.TH0 [5]);
  nor (_03940_, _03939_, _03938_);
  and (_03941_, _03845_, \oc8051_golden_model_1.TL1 [5]);
  not (_03942_, _03941_);
  and (_03943_, _03942_, _03940_);
  and (_03944_, _03676_, \oc8051_golden_model_1.PSW [5]);
  and (_03945_, _03680_, \oc8051_golden_model_1.ACC [5]);
  nor (_03946_, _03945_, _03944_);
  and (_03947_, _03670_, \oc8051_golden_model_1.IP [5]);
  and (_03948_, _03683_, \oc8051_golden_model_1.B [5]);
  nor (_03949_, _03948_, _03947_);
  and (_03950_, _03949_, _03946_);
  and (_03951_, _03698_, \oc8051_golden_model_1.P1 [5]);
  not (_03952_, _03951_);
  and (_03953_, _03665_, \oc8051_golden_model_1.P2 [5]);
  and (_03954_, _03646_, \oc8051_golden_model_1.P3 [5]);
  nor (_03955_, _03954_, _03953_);
  and (_03956_, _03955_, _03952_);
  and (_03957_, _03956_, _03950_);
  and (_03958_, _03662_, \oc8051_golden_model_1.PCON [5]);
  and (_03959_, _03832_, \oc8051_golden_model_1.P0 [5]);
  nor (_03960_, _03959_, _03958_);
  and (_03961_, _03960_, _03957_);
  and (_03962_, _03961_, _03943_);
  and (_03963_, _03962_, _03937_);
  and (_03964_, _03963_, _03917_);
  not (_03965_, _03964_);
  or (_03966_, _03268_, _01790_);
  and (_03967_, _03670_, \oc8051_golden_model_1.IP [3]);
  and (_03968_, _03680_, \oc8051_golden_model_1.ACC [3]);
  nor (_03969_, _03968_, _03967_);
  and (_03970_, _03676_, \oc8051_golden_model_1.PSW [3]);
  and (_03971_, _03683_, \oc8051_golden_model_1.B [3]);
  nor (_03972_, _03971_, _03970_);
  and (_03973_, _03972_, _03969_);
  and (_03974_, _03832_, \oc8051_golden_model_1.P0 [3]);
  not (_03975_, _03974_);
  and (_03976_, _03698_, \oc8051_golden_model_1.P1 [3]);
  not (_03977_, _03976_);
  and (_03978_, _03665_, \oc8051_golden_model_1.P2 [3]);
  and (_03979_, _03646_, \oc8051_golden_model_1.P3 [3]);
  nor (_03980_, _03979_, _03978_);
  and (_03981_, _03980_, _03977_);
  and (_03982_, _03981_, _03975_);
  and (_03983_, _03982_, _03973_);
  and (_03984_, _03662_, \oc8051_golden_model_1.PCON [3]);
  not (_03985_, _03984_);
  and (_03986_, _03625_, \oc8051_golden_model_1.SBUF [3]);
  and (_03987_, _03633_, \oc8051_golden_model_1.IE [3]);
  nor (_03988_, _03987_, _03986_);
  and (_03989_, _03988_, _03985_);
  and (_03990_, _03856_, \oc8051_golden_model_1.DPL [3]);
  and (_03991_, _03853_, \oc8051_golden_model_1.SP [3]);
  nor (_03992_, _03991_, _03990_);
  and (_03993_, _03992_, _03989_);
  and (_03994_, _03993_, _03983_);
  and (_03995_, _03730_, \oc8051_golden_model_1.TL0 [3]);
  not (_03996_, _03995_);
  and (_03997_, _03726_, \oc8051_golden_model_1.TMOD [3]);
  and (_03998_, _03716_, \oc8051_golden_model_1.SCON [3]);
  nor (_03999_, _03998_, _03997_);
  and (_04000_, _03693_, \oc8051_golden_model_1.TCON [3]);
  and (_04001_, _03722_, \oc8051_golden_model_1.TH1 [3]);
  nor (_04002_, _04001_, _04000_);
  and (_04003_, _04002_, _03999_);
  and (_04004_, _04003_, _03996_);
  and (_04005_, _03845_, \oc8051_golden_model_1.TL1 [3]);
  not (_04006_, _04005_);
  and (_04007_, _03691_, \oc8051_golden_model_1.TH0 [3]);
  and (_04008_, _03850_, \oc8051_golden_model_1.DPH [3]);
  nor (_04009_, _04008_, _04007_);
  and (_04010_, _04009_, _04006_);
  and (_04011_, _04010_, _04004_);
  and (_04012_, _04011_, _03994_);
  and (_04013_, _04012_, _03966_);
  not (_04014_, _04013_);
  or (_04015_, _02811_, _01790_);
  and (_04016_, _03676_, \oc8051_golden_model_1.PSW [1]);
  and (_04017_, _03680_, \oc8051_golden_model_1.ACC [1]);
  nor (_04018_, _04017_, _04016_);
  and (_04019_, _03670_, \oc8051_golden_model_1.IP [1]);
  and (_04020_, _03683_, \oc8051_golden_model_1.B [1]);
  nor (_04021_, _04020_, _04019_);
  and (_04022_, _04021_, _04018_);
  and (_04023_, _03737_, \oc8051_golden_model_1.P0 [1]);
  and (_04024_, _03741_, \oc8051_golden_model_1.DPH [1]);
  nor (_04025_, _04024_, _04023_);
  and (_04026_, _03625_, \oc8051_golden_model_1.SBUF [1]);
  and (_04027_, _03633_, \oc8051_golden_model_1.IE [1]);
  nor (_04028_, _04027_, _04026_);
  and (_04029_, _03646_, \oc8051_golden_model_1.P3 [1]);
  and (_04030_, _03662_, \oc8051_golden_model_1.PCON [1]);
  and (_04031_, _03665_, \oc8051_golden_model_1.P2 [1]);
  or (_04032_, _04031_, _04030_);
  nor (_04033_, _04032_, _04029_);
  and (_04034_, _04033_, _04028_);
  and (_04035_, _03691_, \oc8051_golden_model_1.TH0 [1]);
  and (_04036_, _03693_, \oc8051_golden_model_1.TCON [1]);
  nor (_04037_, _04036_, _04035_);
  and (_04038_, _03698_, \oc8051_golden_model_1.P1 [1]);
  and (_04039_, _03708_, \oc8051_golden_model_1.TL1 [1]);
  nor (_04040_, _04039_, _04038_);
  and (_04041_, _04040_, _04037_);
  and (_04042_, _03722_, \oc8051_golden_model_1.TH1 [1]);
  and (_04043_, _03716_, \oc8051_golden_model_1.SCON [1]);
  nor (_04044_, _04043_, _04042_);
  and (_04045_, _03726_, \oc8051_golden_model_1.TMOD [1]);
  and (_04046_, _03730_, \oc8051_golden_model_1.TL0 [1]);
  nor (_04047_, _04046_, _04045_);
  and (_04048_, _04047_, _04044_);
  and (_04049_, _04048_, _04041_);
  and (_04050_, _03745_, \oc8051_golden_model_1.SP [1]);
  and (_04051_, _03748_, \oc8051_golden_model_1.DPL [1]);
  nor (_04052_, _04051_, _04050_);
  and (_04053_, _04052_, _04049_);
  and (_04054_, _04053_, _04034_);
  and (_04055_, _04054_, _04025_);
  and (_04056_, _04055_, _04022_);
  and (_04057_, _04056_, _04015_);
  not (_04058_, _04057_);
  or (_04059_, _03042_, _01790_);
  and (_04060_, _03722_, \oc8051_golden_model_1.TH1 [0]);
  and (_04061_, _03625_, \oc8051_golden_model_1.SBUF [0]);
  nor (_04062_, _04061_, _04060_);
  and (_04063_, _03691_, \oc8051_golden_model_1.TH0 [0]);
  and (_04064_, _03716_, \oc8051_golden_model_1.SCON [0]);
  nor (_04065_, _04064_, _04063_);
  and (_04066_, _04065_, _04062_);
  and (_04067_, _03850_, \oc8051_golden_model_1.DPH [0]);
  not (_04068_, _04067_);
  and (_04069_, _03726_, \oc8051_golden_model_1.TMOD [0]);
  and (_04070_, _03633_, \oc8051_golden_model_1.IE [0]);
  nor (_04071_, _04070_, _04069_);
  and (_04072_, _04071_, _04068_);
  and (_04073_, _03730_, \oc8051_golden_model_1.TL0 [0]);
  and (_04074_, _03845_, \oc8051_golden_model_1.TL1 [0]);
  nor (_04075_, _04074_, _04073_);
  and (_04076_, _04075_, _04072_);
  and (_04077_, _04076_, _04066_);
  and (_04078_, _03662_, \oc8051_golden_model_1.PCON [0]);
  not (_04079_, _04078_);
  and (_04080_, _03693_, \oc8051_golden_model_1.TCON [0]);
  not (_04081_, _04080_);
  and (_04082_, _03670_, \oc8051_golden_model_1.IP [0]);
  and (_04083_, _03683_, \oc8051_golden_model_1.B [0]);
  nor (_04084_, _04083_, _04082_);
  and (_04085_, _03676_, \oc8051_golden_model_1.PSW [0]);
  and (_04086_, _03680_, \oc8051_golden_model_1.ACC [0]);
  nor (_04087_, _04086_, _04085_);
  and (_04088_, _04087_, _04084_);
  and (_04089_, _04088_, _04081_);
  and (_04090_, _04089_, _04079_);
  and (_04091_, _03856_, \oc8051_golden_model_1.DPL [0]);
  and (_04092_, _03853_, \oc8051_golden_model_1.SP [0]);
  nor (_04093_, _04092_, _04091_);
  and (_04094_, _03832_, \oc8051_golden_model_1.P0 [0]);
  not (_04095_, _04094_);
  and (_04096_, _03698_, \oc8051_golden_model_1.P1 [0]);
  not (_04097_, _04096_);
  and (_04098_, _03665_, \oc8051_golden_model_1.P2 [0]);
  and (_04099_, _03646_, \oc8051_golden_model_1.P3 [0]);
  nor (_04100_, _04099_, _04098_);
  and (_04101_, _04100_, _04097_);
  and (_04102_, _04101_, _04095_);
  and (_04103_, _04102_, _04093_);
  and (_04104_, _04103_, _04090_);
  and (_04105_, _04104_, _04077_);
  nand (_04106_, _04105_, _04059_);
  and (_04107_, _04106_, _04058_);
  or (_04108_, _03455_, _01790_);
  and (_04109_, _03853_, \oc8051_golden_model_1.SP [2]);
  and (_04110_, _03850_, \oc8051_golden_model_1.DPH [2]);
  nor (_04111_, _04110_, _04109_);
  and (_04112_, _03730_, \oc8051_golden_model_1.TL0 [2]);
  and (_04113_, _03845_, \oc8051_golden_model_1.TL1 [2]);
  nor (_04114_, _04113_, _04112_);
  and (_04115_, _04114_, _04111_);
  and (_04116_, _03693_, \oc8051_golden_model_1.TCON [2]);
  not (_04117_, _04116_);
  and (_04118_, _03726_, \oc8051_golden_model_1.TMOD [2]);
  and (_04119_, _03716_, \oc8051_golden_model_1.SCON [2]);
  nor (_04120_, _04119_, _04118_);
  and (_04121_, _04120_, _04117_);
  and (_04122_, _03856_, \oc8051_golden_model_1.DPL [2]);
  not (_04123_, _04122_);
  and (_04124_, _03691_, \oc8051_golden_model_1.TH0 [2]);
  and (_04125_, _03722_, \oc8051_golden_model_1.TH1 [2]);
  nor (_04126_, _04125_, _04124_);
  and (_04127_, _04126_, _04123_);
  and (_04128_, _04127_, _04121_);
  and (_04129_, _04128_, _04115_);
  and (_04130_, _03662_, \oc8051_golden_model_1.PCON [2]);
  not (_04131_, _04130_);
  and (_04132_, _03625_, \oc8051_golden_model_1.SBUF [2]);
  and (_04133_, _03633_, \oc8051_golden_model_1.IE [2]);
  nor (_04134_, _04133_, _04132_);
  and (_04135_, _04134_, _04131_);
  and (_04136_, _03832_, \oc8051_golden_model_1.P0 [2]);
  not (_04137_, _04136_);
  and (_04138_, _03670_, \oc8051_golden_model_1.IP [2]);
  and (_04139_, _03680_, \oc8051_golden_model_1.ACC [2]);
  nor (_04140_, _04139_, _04138_);
  and (_04141_, _03676_, \oc8051_golden_model_1.PSW [2]);
  and (_04142_, _03683_, \oc8051_golden_model_1.B [2]);
  nor (_04143_, _04142_, _04141_);
  and (_04144_, _04143_, _04140_);
  and (_04145_, _03698_, \oc8051_golden_model_1.P1 [2]);
  not (_04146_, _04145_);
  and (_04147_, _03665_, \oc8051_golden_model_1.P2 [2]);
  and (_04148_, _03646_, \oc8051_golden_model_1.P3 [2]);
  nor (_04149_, _04148_, _04147_);
  and (_04150_, _04149_, _04146_);
  and (_04151_, _04150_, _04144_);
  and (_04152_, _04151_, _04137_);
  and (_04153_, _04152_, _04135_);
  and (_04154_, _04153_, _04129_);
  and (_04155_, _04154_, _04108_);
  not (_04156_, _04155_);
  and (_04157_, _04156_, _04107_);
  and (_04158_, _04157_, _04014_);
  not (_04159_, \oc8051_golden_model_1.IRAM[0] [4]);
  or (_04160_, _02653_, _04159_);
  not (_04161_, \oc8051_golden_model_1.IRAM[1] [4]);
  or (_04162_, _02751_, _04161_);
  and (_04163_, _04162_, _02749_);
  nand (_04164_, _04163_, _04160_);
  not (_04165_, \oc8051_golden_model_1.IRAM[3] [4]);
  or (_04166_, _02751_, _04165_);
  not (_04167_, \oc8051_golden_model_1.IRAM[2] [4]);
  or (_04168_, _02653_, _04167_);
  and (_04169_, _04168_, _02757_);
  nand (_04170_, _04169_, _04166_);
  nand (_04171_, _04170_, _04164_);
  nand (_04172_, _04171_, _02406_);
  not (_04173_, \oc8051_golden_model_1.IRAM[7] [4]);
  or (_04174_, _02751_, _04173_);
  not (_04175_, \oc8051_golden_model_1.IRAM[6] [4]);
  or (_04176_, _02653_, _04175_);
  and (_04177_, _04176_, _02757_);
  nand (_04178_, _04177_, _04174_);
  not (_04179_, \oc8051_golden_model_1.IRAM[4] [4]);
  or (_04180_, _02653_, _04179_);
  not (_04181_, \oc8051_golden_model_1.IRAM[5] [4]);
  or (_04182_, _02751_, _04181_);
  and (_04183_, _04182_, _02749_);
  nand (_04184_, _04183_, _04180_);
  nand (_04185_, _04184_, _04178_);
  nand (_04186_, _04185_, _02764_);
  nand (_04187_, _04186_, _04172_);
  nand (_04188_, _04187_, _02221_);
  nand (_04189_, _02653_, \oc8051_golden_model_1.IRAM[11] [4]);
  nand (_04190_, _02751_, \oc8051_golden_model_1.IRAM[10] [4]);
  and (_04191_, _04190_, _02757_);
  nand (_04192_, _04191_, _04189_);
  nand (_04193_, _02751_, \oc8051_golden_model_1.IRAM[8] [4]);
  nand (_04194_, _02653_, \oc8051_golden_model_1.IRAM[9] [4]);
  and (_04195_, _04194_, _02749_);
  nand (_04196_, _04195_, _04193_);
  nand (_04197_, _04196_, _04192_);
  nand (_04198_, _04197_, _02406_);
  nand (_04199_, _02653_, \oc8051_golden_model_1.IRAM[15] [4]);
  nand (_04200_, _02751_, \oc8051_golden_model_1.IRAM[14] [4]);
  and (_04201_, _04200_, _02757_);
  nand (_04202_, _04201_, _04199_);
  nand (_04203_, _02751_, \oc8051_golden_model_1.IRAM[12] [4]);
  nand (_04204_, _02653_, \oc8051_golden_model_1.IRAM[13] [4]);
  and (_04205_, _04204_, _02749_);
  nand (_04206_, _04205_, _04203_);
  nand (_04207_, _04206_, _04202_);
  nand (_04208_, _04207_, _02764_);
  nand (_04209_, _04208_, _04198_);
  nand (_04210_, _04209_, _02782_);
  nand (_04211_, _04210_, _04188_);
  or (_04212_, _04211_, _01790_);
  and (_04213_, _03662_, \oc8051_golden_model_1.PCON [4]);
  not (_04214_, _04213_);
  and (_04215_, _03625_, \oc8051_golden_model_1.SBUF [4]);
  and (_04216_, _03633_, \oc8051_golden_model_1.IE [4]);
  nor (_04217_, _04216_, _04215_);
  and (_04218_, _04217_, _04214_);
  and (_04219_, _03665_, \oc8051_golden_model_1.P2 [4]);
  and (_04220_, _03646_, \oc8051_golden_model_1.P3 [4]);
  nor (_04221_, _04220_, _04219_);
  and (_04222_, _04221_, _04218_);
  and (_04223_, _03676_, \oc8051_golden_model_1.PSW [4]);
  and (_04224_, _03683_, \oc8051_golden_model_1.B [4]);
  nor (_04225_, _04224_, _04223_);
  and (_04226_, _03670_, \oc8051_golden_model_1.IP [4]);
  and (_04227_, _03680_, \oc8051_golden_model_1.ACC [4]);
  nor (_04228_, _04227_, _04226_);
  and (_04229_, _04228_, _04225_);
  and (_04230_, _03693_, \oc8051_golden_model_1.TCON [4]);
  and (_04231_, _03691_, \oc8051_golden_model_1.TH0 [4]);
  nor (_04232_, _04231_, _04230_);
  and (_04233_, _03698_, \oc8051_golden_model_1.P1 [4]);
  and (_04234_, _03708_, \oc8051_golden_model_1.TL1 [4]);
  nor (_04235_, _04234_, _04233_);
  and (_04236_, _04235_, _04232_);
  and (_04237_, _03716_, \oc8051_golden_model_1.SCON [4]);
  and (_04238_, _03722_, \oc8051_golden_model_1.TH1 [4]);
  nor (_04239_, _04238_, _04237_);
  and (_04240_, _03726_, \oc8051_golden_model_1.TMOD [4]);
  and (_04241_, _03730_, \oc8051_golden_model_1.TL0 [4]);
  nor (_04242_, _04241_, _04240_);
  and (_04243_, _04242_, _04239_);
  and (_04244_, _04243_, _04236_);
  and (_04245_, _04244_, _04229_);
  and (_04246_, _04245_, _04222_);
  and (_04247_, _03737_, \oc8051_golden_model_1.P0 [4]);
  not (_04248_, _04247_);
  and (_04249_, _03741_, \oc8051_golden_model_1.DPH [4]);
  not (_04250_, _04249_);
  and (_04251_, _03745_, \oc8051_golden_model_1.SP [4]);
  and (_04252_, _03748_, \oc8051_golden_model_1.DPL [4]);
  nor (_04253_, _04252_, _04251_);
  and (_04254_, _04253_, _04250_);
  and (_04255_, _04254_, _04248_);
  and (_04256_, _04255_, _04246_);
  and (_04257_, _04256_, _04212_);
  not (_04258_, _04257_);
  and (_04259_, _04258_, _04158_);
  and (_04260_, _04259_, _03965_);
  and (_04261_, _04260_, _03863_);
  nor (_04262_, _04261_, _03755_);
  and (_04263_, _04261_, _03755_);
  nor (_04264_, _04263_, _04262_);
  and (_04265_, _04264_, _01791_);
  and (_04266_, _01284_, \oc8051_golden_model_1.PC [2]);
  and (_04267_, _04266_, \oc8051_golden_model_1.PC [3]);
  and (_04268_, \oc8051_golden_model_1.PC [5], \oc8051_golden_model_1.PC [4]);
  and (_04269_, _04268_, \oc8051_golden_model_1.PC [6]);
  and (_04270_, _04269_, \oc8051_golden_model_1.PC [7]);
  and (_04271_, _04270_, _04267_);
  and (_04272_, _04267_, _04269_);
  nor (_04273_, _04272_, \oc8051_golden_model_1.PC [7]);
  nor (_04274_, _04273_, _04271_);
  not (_04275_, _04274_);
  nand (_04276_, _04275_, _02058_);
  and (_04277_, _02107_, _41243_);
  and (_04278_, _02110_, _00014_);
  nor (_04279_, _04278_, _04277_);
  and (_04280_, _02135_, _41192_);
  and (_04281_, _02152_, _00022_);
  nor (_04282_, _04281_, _04280_);
  and (_04283_, _04282_, _04279_);
  and (_04284_, _02128_, _00011_);
  and (_04285_, _02130_, _00008_);
  nor (_04286_, _04285_, _04284_);
  and (_04287_, _02123_, _41240_);
  and (_04288_, _02147_, _41236_);
  nor (_04289_, _04288_, _04287_);
  and (_04290_, _04289_, _04286_);
  and (_04291_, _04290_, _04283_);
  and (_04292_, _02143_, _41222_);
  and (_04293_, _02137_, _00025_);
  nor (_04294_, _04293_, _04292_);
  and (_04295_, _02140_, _41213_);
  and (_04296_, _02154_, _00019_);
  nor (_04297_, _04296_, _04295_);
  and (_04298_, _04297_, _04294_);
  and (_04299_, _02125_, _41248_);
  and (_04300_, _02149_, _41251_);
  nor (_04301_, _04300_, _04299_);
  and (_04302_, _02115_, _41216_);
  and (_04303_, _02119_, _41226_);
  nor (_04304_, _04303_, _04302_);
  and (_04305_, _04304_, _04301_);
  and (_04306_, _04305_, _04298_);
  and (_04307_, _04306_, _04291_);
  nor (_04308_, _04307_, _03754_);
  and (_04309_, _04308_, _02910_);
  not (_04310_, _01604_);
  not (_04311_, _02870_);
  nor (_04312_, _02253_, _01856_);
  and (_04313_, _04312_, _02409_);
  and (_04314_, _04313_, _01964_);
  and (_04315_, _04314_, _03654_);
  and (_04316_, _04315_, \oc8051_golden_model_1.TCON [7]);
  and (_04317_, _04313_, _01957_);
  and (_04318_, _03682_, _04317_);
  and (_04319_, _04318_, \oc8051_golden_model_1.B [7]);
  nor (_04320_, _04319_, _04316_);
  and (_04321_, _03675_, _04317_);
  and (_04322_, _04321_, \oc8051_golden_model_1.PSW [7]);
  not (_04323_, _04322_);
  and (_04324_, _04314_, _03640_);
  and (_04325_, _04324_, \oc8051_golden_model_1.IP [7]);
  and (_04326_, _03679_, _04317_);
  and (_04327_, _04326_, \oc8051_golden_model_1.ACC [7]);
  nor (_04328_, _04327_, _04325_);
  and (_04329_, _04328_, _04323_);
  and (_04330_, _04329_, _04320_);
  and (_04331_, _04314_, _03624_);
  and (_04332_, _04331_, \oc8051_golden_model_1.SCON [7]);
  and (_04333_, _04314_, _03632_);
  and (_04334_, _04333_, \oc8051_golden_model_1.IE [7]);
  nor (_04335_, _04334_, _04332_);
  and (_04336_, _03624_, _04317_);
  and (_04337_, _04336_, \oc8051_golden_model_1.P1INREG [7]);
  and (_04338_, _03640_, _04317_);
  and (_04339_, _04338_, \oc8051_golden_model_1.P3INREG [7]);
  nor (_04340_, _04339_, _04337_);
  and (_04341_, _03656_, \oc8051_golden_model_1.P0INREG [7]);
  and (_04342_, _03632_, _04317_);
  and (_04343_, _04342_, \oc8051_golden_model_1.P2INREG [7]);
  nor (_04344_, _04343_, _04341_);
  and (_04345_, _04344_, _04340_);
  and (_04346_, _04345_, _04335_);
  and (_04347_, _04346_, _04330_);
  and (_04348_, _04347_, _03617_);
  nor (_04349_, _04348_, _03660_);
  and (_04350_, _03660_, \oc8051_golden_model_1.PSW [7]);
  nor (_04351_, _04350_, _04349_);
  nor (_04352_, _04351_, _04311_);
  not (_04353_, _02856_);
  and (_04354_, _03656_, \oc8051_golden_model_1.P0 [7]);
  and (_04355_, _04336_, \oc8051_golden_model_1.P1 [7]);
  nor (_04356_, _04355_, _04354_);
  and (_04357_, _04342_, \oc8051_golden_model_1.P2 [7]);
  and (_04358_, _04338_, \oc8051_golden_model_1.P3 [7]);
  nor (_04359_, _04358_, _04357_);
  and (_04360_, _04359_, _04356_);
  and (_04361_, _04360_, _04335_);
  and (_04362_, _04361_, _04330_);
  and (_04363_, _04362_, _03617_);
  nor (_04364_, _04363_, _03660_);
  or (_04365_, _04364_, _04353_);
  not (_04366_, _02837_);
  not (_04367_, _03660_);
  nand (_04368_, _04363_, _04367_);
  or (_04369_, _04368_, _04366_);
  not (_04370_, _03616_);
  and (_04371_, _04211_, _03916_);
  and (_04372_, _03042_, _02811_);
  and (_04373_, _03455_, _03268_);
  and (_04374_, _04373_, _04372_);
  and (_04375_, _04374_, _04371_);
  and (_04376_, _04375_, _03808_);
  or (_04377_, _04376_, _04370_);
  nand (_04378_, _04376_, _04370_);
  and (_04379_, _04378_, _04377_);
  nor (_04380_, _01557_, _01534_);
  not (_04381_, _04380_);
  or (_04382_, _04381_, _04379_);
  and (_04383_, _01562_, \oc8051_golden_model_1.ACC [7]);
  and (_04384_, _04269_, _01680_);
  and (_04385_, _04384_, \oc8051_golden_model_1.PC [7]);
  nor (_04386_, _04384_, \oc8051_golden_model_1.PC [7]);
  nor (_04387_, _04386_, _04385_);
  not (_04388_, _04387_);
  nor (_04389_, _04388_, _01562_);
  or (_04390_, _04389_, _04383_);
  or (_04391_, _04390_, _04380_);
  and (_04392_, _04391_, _04382_);
  or (_04393_, _04392_, _01883_);
  not (_04394_, _01883_);
  nor (_04395_, \oc8051_golden_model_1.SP [1], \oc8051_golden_model_1.SP [0]);
  and (_04396_, _04395_, _02346_);
  nor (_04397_, _04396_, _01998_);
  nor (_04398_, \oc8051_golden_model_1.SP [2], \oc8051_golden_model_1.SP [1]);
  and (_04399_, _04398_, _01998_);
  and (_04400_, _04399_, _01864_);
  nor (_04401_, _04400_, _04397_);
  nor (_04402_, _04401_, _02347_);
  not (_04403_, _02871_);
  and (_04404_, _03268_, _04403_);
  and (_04405_, _02871_, _01954_);
  not (_04406_, _04405_);
  nand (_04407_, _04406_, _02347_);
  nor (_04408_, _04407_, _04404_);
  nor (_04409_, _04408_, _04402_);
  not (_04410_, _04409_);
  nor (_04411_, _04395_, _02346_);
  nor (_04412_, _04411_, _04396_);
  nor (_04413_, _04412_, _02347_);
  not (_04414_, _04413_);
  nand (_04415_, _03455_, _04403_);
  and (_04416_, _02871_, _02294_);
  not (_04417_, _04416_);
  and (_04418_, _04417_, _02347_);
  nand (_04419_, _04418_, _04415_);
  and (_04420_, _04419_, _04414_);
  or (_04421_, _03028_, _02871_);
  not (_04422_, _02347_);
  and (_04423_, _02871_, _02441_);
  nor (_04424_, _04423_, _04422_);
  nand (_04425_, _04424_, _04421_);
  nor (_04426_, _02347_, \oc8051_golden_model_1.SP [0]);
  not (_04427_, _04426_);
  and (_04428_, _04427_, _04425_);
  or (_04429_, _04428_, \oc8051_golden_model_1.IRAM[9] [7]);
  nor (_04430_, _02347_, _01866_);
  not (_04431_, _04430_);
  or (_04432_, _02811_, _02871_);
  or (_04433_, _04403_, _01822_);
  and (_04434_, _04433_, _02347_);
  nand (_04435_, _04434_, _04432_);
  and (_04436_, _04435_, _04431_);
  not (_04437_, _04436_);
  not (_04438_, _04428_);
  or (_04439_, _04438_, \oc8051_golden_model_1.IRAM[8] [7]);
  and (_04440_, _04439_, _04437_);
  and (_04441_, _04440_, _04429_);
  nand (_04442_, _04428_, _03594_);
  or (_04443_, _04428_, \oc8051_golden_model_1.IRAM[11] [7]);
  and (_04444_, _04443_, _04436_);
  and (_04445_, _04444_, _04442_);
  nor (_04446_, _04445_, _04441_);
  nand (_04447_, _04446_, _04420_);
  not (_04448_, _04420_);
  or (_04449_, _04428_, \oc8051_golden_model_1.IRAM[13] [7]);
  or (_04450_, _04438_, \oc8051_golden_model_1.IRAM[12] [7]);
  and (_04451_, _04450_, _04437_);
  and (_04452_, _04451_, _04449_);
  or (_04453_, _04438_, \oc8051_golden_model_1.IRAM[14] [7]);
  or (_04454_, _04428_, \oc8051_golden_model_1.IRAM[15] [7]);
  and (_04455_, _04454_, _04436_);
  and (_04456_, _04455_, _04453_);
  nor (_04457_, _04456_, _04452_);
  nand (_04458_, _04457_, _04448_);
  nand (_04459_, _04458_, _04447_);
  nand (_04460_, _04459_, _04410_);
  or (_04461_, _04428_, _03565_);
  nand (_04462_, _04428_, \oc8051_golden_model_1.IRAM[0] [7]);
  and (_04463_, _04462_, _04437_);
  nand (_04464_, _04463_, _04461_);
  nand (_04465_, _04428_, \oc8051_golden_model_1.IRAM[2] [7]);
  or (_04466_, _04428_, _03569_);
  and (_04467_, _04466_, _04436_);
  nand (_04468_, _04467_, _04465_);
  nand (_04469_, _04468_, _04464_);
  nand (_04470_, _04469_, _04420_);
  nand (_04471_, _04428_, \oc8051_golden_model_1.IRAM[4] [7]);
  or (_04472_, _04428_, _03585_);
  and (_04473_, _04472_, _04437_);
  nand (_04474_, _04473_, _04471_);
  nand (_04475_, _04428_, \oc8051_golden_model_1.IRAM[6] [7]);
  or (_04476_, _04428_, _03577_);
  and (_04477_, _04476_, _04436_);
  nand (_04478_, _04477_, _04475_);
  nand (_04479_, _04478_, _04474_);
  nand (_04480_, _04479_, _04448_);
  nand (_04481_, _04480_, _04470_);
  nand (_04482_, _04481_, _04409_);
  and (_04483_, _04482_, _04460_);
  or (_04484_, _04483_, _04394_);
  and (_04485_, _04484_, _04393_);
  or (_04486_, _04485_, _02815_);
  and (_04487_, _04257_, _03964_);
  not (_04488_, _04106_);
  and (_04489_, _04488_, _04057_);
  and (_04490_, _04155_, _04013_);
  and (_04491_, _04490_, _04489_);
  and (_04492_, _04491_, _04487_);
  and (_04493_, _04492_, _03862_);
  nor (_04494_, _04493_, _03755_);
  and (_04495_, _04493_, _03755_);
  nor (_04496_, _04495_, _04494_);
  or (_04497_, _04496_, _02816_);
  and (_04498_, _04497_, _04486_);
  or (_04499_, _04498_, _02837_);
  and (_04500_, _04499_, _04369_);
  or (_04501_, _04500_, _03279_);
  nor (_04502_, _04387_, _01558_);
  nor (_04503_, _04502_, _02841_);
  and (_04504_, _04503_, _04501_);
  and (_04505_, _04370_, _02841_);
  or (_04506_, _04505_, _02856_);
  or (_04507_, _04506_, _04504_);
  and (_04508_, _04507_, _04365_);
  or (_04509_, _04508_, _01878_);
  not (_04510_, _03692_);
  and (_04511_, _03732_, _04510_);
  nor (_04512_, _03710_, _03694_);
  and (_04513_, _04512_, _04511_);
  and (_04514_, _03665_, \oc8051_golden_model_1.P2INREG [7]);
  and (_04515_, _03646_, \oc8051_golden_model_1.P3INREG [7]);
  nor (_04516_, _04515_, _04514_);
  and (_04517_, _03698_, \oc8051_golden_model_1.P1INREG [7]);
  and (_04518_, _03737_, \oc8051_golden_model_1.P0INREG [7]);
  nor (_04519_, _04518_, _04517_);
  and (_04520_, _04519_, _04516_);
  and (_04521_, _04520_, _04513_);
  not (_04522_, _03664_);
  and (_04523_, _03636_, _04522_);
  and (_04524_, _04523_, _03725_);
  and (_04525_, _03751_, _03687_);
  and (_04526_, _04525_, _04524_);
  and (_04527_, _04526_, _04521_);
  and (_04528_, _04527_, _03617_);
  nand (_04529_, _04528_, _01878_);
  and (_04530_, _04529_, _02962_);
  and (_04531_, _04530_, _04509_);
  nor (_04532_, _04363_, _04367_);
  not (_04533_, _04532_);
  and (_04534_, _04533_, _04368_);
  and (_04535_, _04534_, _02862_);
  or (_04536_, _04535_, _04531_);
  and (_04537_, _04536_, _01565_);
  or (_04538_, _04388_, _01565_);
  nand (_04539_, _04538_, _01989_);
  or (_04540_, _04539_, _04537_);
  nand (_04541_, _04528_, _02503_);
  and (_04542_, _04541_, _04540_);
  or (_04543_, _04542_, _02871_);
  nand (_04544_, _04483_, _03673_);
  and (_04545_, _04527_, _02871_);
  nand (_04546_, _04545_, _04544_);
  and (_04547_, _04546_, _04311_);
  and (_04548_, _04547_, _04543_);
  or (_04549_, _04548_, _04352_);
  and (_04550_, _04549_, _04310_);
  nand (_04551_, _04387_, _01604_);
  nand (_04552_, _04551_, _02887_);
  or (_04553_, _04552_, _04550_);
  or (_04554_, _04370_, _02887_);
  and (_04555_, _04554_, _04553_);
  or (_04556_, _04555_, _02889_);
  or (_04557_, _04483_, _02890_);
  and (_04558_, _04557_, _02880_);
  and (_04559_, _04558_, _04556_);
  not (_04560_, _04307_);
  nor (_04561_, _04560_, _03616_);
  not (_04562_, _02568_);
  and (_04563_, _02687_, _04562_);
  and (_04564_, _02140_, _00486_);
  and (_04565_, _02137_, _00524_);
  nor (_04566_, _04565_, _04564_);
  and (_04567_, _02123_, _00492_);
  and (_04568_, _02149_, _00507_);
  nor (_04569_, _04568_, _04567_);
  and (_04570_, _04569_, _04566_);
  and (_04571_, _02152_, _00526_);
  and (_04572_, _02119_, _00521_);
  nor (_04573_, _04572_, _04571_);
  and (_04574_, _02115_, _00476_);
  and (_04575_, _02143_, _00482_);
  nor (_04576_, _04575_, _04574_);
  and (_04577_, _04576_, _04573_);
  and (_04578_, _04577_, _04570_);
  and (_04579_, _02147_, _00496_);
  and (_04580_, _02110_, _00509_);
  nor (_04581_, _04580_, _04579_);
  and (_04582_, _02107_, _00502_);
  and (_04583_, _02125_, _00494_);
  nor (_04584_, _04583_, _04582_);
  and (_04585_, _04584_, _04581_);
  and (_04586_, _02128_, _00513_);
  and (_04587_, _02130_, _00500_);
  nor (_04588_, _04587_, _04586_);
  and (_04589_, _02135_, _00479_);
  and (_04590_, _02154_, _00488_);
  nor (_04591_, _04590_, _04589_);
  and (_04592_, _04591_, _04588_);
  and (_04593_, _04592_, _04585_);
  and (_04594_, _04593_, _04578_);
  and (_04595_, _04594_, _04560_);
  and (_04596_, _02140_, _00431_);
  and (_04597_, _02110_, _00454_);
  nor (_04598_, _04597_, _04596_);
  and (_04599_, _02115_, _00421_);
  and (_04600_, _02154_, _00433_);
  nor (_04601_, _04600_, _04599_);
  and (_04602_, _04601_, _04598_);
  and (_04603_, _02125_, _00439_);
  and (_04604_, _02123_, _00437_);
  nor (_04605_, _04604_, _04603_);
  and (_04606_, _02137_, _00467_);
  and (_04607_, _02107_, _00447_);
  nor (_04608_, _04607_, _04606_);
  and (_04609_, _04608_, _04605_);
  and (_04610_, _04609_, _04602_);
  and (_04611_, _02135_, _00423_);
  and (_04612_, _02143_, _00426_);
  nor (_04613_, _04612_, _04611_);
  and (_04614_, _02119_, _00463_);
  and (_04615_, _02128_, _00456_);
  nor (_04616_, _04615_, _04614_);
  and (_04617_, _04616_, _04613_);
  and (_04618_, _02152_, _00471_);
  and (_04619_, _02147_, _00441_);
  nor (_04620_, _04619_, _04618_);
  and (_04621_, _02149_, _00452_);
  and (_04622_, _02130_, _00445_);
  nor (_04623_, _04622_, _04621_);
  and (_04624_, _04623_, _04620_);
  and (_04625_, _04624_, _04617_);
  and (_04626_, _04625_, _04610_);
  and (_04627_, _02140_, _00394_);
  and (_04628_, _02154_, _00368_);
  nor (_04629_, _04628_, _04627_);
  and (_04630_, _02125_, _00381_);
  and (_04631_, _02130_, _00405_);
  nor (_04632_, _04631_, _04630_);
  and (_04633_, _04632_, _04629_);
  and (_04634_, _02115_, _00396_);
  and (_04635_, _02135_, _00398_);
  nor (_04636_, _04635_, _04634_);
  and (_04637_, _02107_, _00387_);
  and (_04638_, _02147_, _00383_);
  nor (_04639_, _04638_, _04637_);
  and (_04640_, _04639_, _04636_);
  and (_04641_, _04640_, _04633_);
  and (_04642_, _02152_, _00374_);
  and (_04643_, _02119_, _00366_);
  nor (_04644_, _04643_, _04642_);
  and (_04645_, _02110_, _00409_);
  and (_04646_, _02149_, _00389_);
  nor (_04647_, _04646_, _04645_);
  and (_04648_, _04647_, _04644_);
  and (_04649_, _02143_, _00400_);
  and (_04650_, _02123_, _00379_);
  nor (_04651_, _04650_, _04649_);
  and (_04652_, _02137_, _00371_);
  and (_04653_, _02128_, _00413_);
  nor (_04654_, _04653_, _04652_);
  and (_04655_, _04654_, _04651_);
  and (_04656_, _04655_, _04648_);
  and (_04657_, _04656_, _04641_);
  and (_04658_, _04657_, _04626_);
  and (_04659_, _04658_, _04595_);
  nor (_04660_, _02338_, _02159_);
  and (_04661_, _04660_, _04659_);
  and (_04662_, _04661_, _04563_);
  and (_04663_, _04662_, \oc8051_golden_model_1.TH1 [7]);
  and (_04664_, _02338_, _02159_);
  nor (_04665_, _02687_, _02568_);
  and (_04666_, _04665_, _04659_);
  and (_04667_, _04666_, _04664_);
  and (_04668_, _04667_, \oc8051_golden_model_1.DPH [7]);
  nor (_04669_, _04668_, _04663_);
  and (_04670_, _02687_, _02568_);
  and (_04671_, _04670_, _04664_);
  not (_04672_, _04626_);
  and (_04673_, _04657_, _04672_);
  and (_04674_, _04673_, _04595_);
  and (_04675_, _04674_, _04671_);
  and (_04676_, _04675_, \oc8051_golden_model_1.P2INREG [7]);
  not (_04677_, _04676_);
  not (_04678_, _02159_);
  and (_04679_, _02338_, _04678_);
  and (_04680_, _04679_, _04563_);
  and (_04681_, _04680_, _04659_);
  and (_04682_, _04681_, \oc8051_golden_model_1.TMOD [7]);
  not (_04683_, _02687_);
  and (_04684_, _04683_, _02568_);
  and (_04685_, _04684_, _04679_);
  and (_04686_, _04685_, _04659_);
  and (_04687_, _04686_, \oc8051_golden_model_1.TL0 [7]);
  nor (_04688_, _04687_, _04682_);
  and (_04689_, _04688_, _04677_);
  and (_04690_, _04679_, _04670_);
  and (_04691_, _04690_, _04674_);
  and (_04692_, _04691_, \oc8051_golden_model_1.IE [7]);
  not (_04693_, _04692_);
  not (_04694_, _04657_);
  and (_04695_, _04694_, _04626_);
  and (_04696_, _04695_, _04595_);
  and (_04697_, _04696_, _04690_);
  and (_04698_, _04697_, \oc8051_golden_model_1.SCON [7]);
  and (_04699_, _04696_, _04680_);
  and (_04700_, _04699_, \oc8051_golden_model_1.SBUF [7]);
  nor (_04701_, _04700_, _04698_);
  and (_04702_, _04701_, _04693_);
  and (_04703_, _04671_, _04659_);
  and (_04704_, _04703_, \oc8051_golden_model_1.P0INREG [7]);
  not (_04705_, _04704_);
  and (_04706_, _04696_, _04671_);
  and (_04707_, _04706_, \oc8051_golden_model_1.P1INREG [7]);
  nor (_04708_, _04657_, _04626_);
  and (_04709_, _04708_, _04595_);
  and (_04710_, _04709_, _04671_);
  and (_04711_, _04710_, \oc8051_golden_model_1.P3INREG [7]);
  nor (_04712_, _04711_, _04707_);
  and (_04713_, _04712_, _04705_);
  and (_04714_, _04713_, _04702_);
  and (_04715_, _04714_, _04689_);
  and (_04716_, _04715_, _04669_);
  and (_04717_, _04670_, _04661_);
  and (_04718_, _04717_, \oc8051_golden_model_1.TH0 [7]);
  and (_04719_, _04679_, _04666_);
  and (_04720_, _04719_, \oc8051_golden_model_1.TL1 [7]);
  nor (_04721_, _04720_, _04718_);
  and (_04722_, _04690_, _04659_);
  and (_04723_, _04722_, \oc8051_golden_model_1.TCON [7]);
  not (_04724_, _02338_);
  and (_04725_, _04724_, _02159_);
  and (_04726_, _04725_, _04666_);
  and (_04727_, _04726_, \oc8051_golden_model_1.PCON [7]);
  nor (_04728_, _04727_, _04723_);
  and (_04729_, _04728_, _04721_);
  and (_04730_, _04709_, _04690_);
  and (_04731_, _04730_, \oc8051_golden_model_1.IP [7]);
  nor (_04732_, _04594_, _04307_);
  and (_04733_, _04732_, _04671_);
  and (_04734_, _04733_, _04673_);
  and (_04735_, _04734_, \oc8051_golden_model_1.ACC [7]);
  nor (_04736_, _04735_, _04731_);
  and (_04737_, _04733_, _04695_);
  and (_04738_, _04737_, \oc8051_golden_model_1.PSW [7]);
  and (_04739_, _04733_, _04708_);
  and (_04740_, _04739_, \oc8051_golden_model_1.B [7]);
  nor (_04741_, _04740_, _04738_);
  and (_04742_, _04741_, _04736_);
  and (_04743_, _04664_, _04659_);
  and (_04744_, _04743_, _04684_);
  and (_04745_, _04744_, \oc8051_golden_model_1.DPL [7]);
  and (_04746_, _04743_, _04563_);
  and (_04747_, _04746_, \oc8051_golden_model_1.SP [7]);
  nor (_04748_, _04747_, _04745_);
  and (_04749_, _04748_, _04742_);
  and (_04750_, _04749_, _04729_);
  and (_04751_, _04750_, _04716_);
  not (_04752_, _04751_);
  nor (_04753_, _04752_, _04561_);
  nor (_04754_, _04753_, _02880_);
  not (_04755_, _02899_);
  and (_04756_, _03142_, _04755_);
  and (_04757_, _04756_, _03147_);
  not (_04758_, _04757_);
  or (_04759_, _04758_, _04754_);
  or (_04760_, _04759_, _04559_);
  nor (_04761_, _04757_, _01790_);
  nor (_04762_, _04761_, _01871_);
  and (_04763_, _04762_, _04760_);
  and (_04764_, _04560_, _01871_);
  or (_04765_, _04764_, _01638_);
  or (_04766_, _04765_, _04763_);
  and (_04767_, _04388_, _01638_);
  nor (_04768_, _04767_, _02914_);
  and (_04769_, _04768_, _04766_);
  and (_04770_, _04307_, _03754_);
  nor (_04771_, _04770_, _04308_);
  nor (_04772_, _04771_, _02913_);
  nor (_04773_, _04772_, _02915_);
  or (_04774_, _04773_, _04769_);
  not (_04775_, _02913_);
  not (_04776_, \oc8051_golden_model_1.ACC [7]);
  nor (_04777_, _03754_, _04776_);
  and (_04778_, _03754_, _04776_);
  nor (_04779_, _04778_, _04777_);
  or (_04780_, _04779_, _04775_);
  and (_04781_, _04780_, _02911_);
  and (_04782_, _04781_, _04774_);
  or (_04783_, _04782_, _04309_);
  and (_04784_, _04783_, _02909_);
  and (_04785_, _04777_, _02908_);
  or (_04786_, _04785_, _01632_);
  or (_04787_, _04786_, _04784_);
  not (_04788_, _02071_);
  nor (_04789_, _04788_, _01790_);
  and (_04790_, _04388_, _01632_);
  nor (_04791_, _04790_, _04789_);
  and (_04792_, _04791_, _04787_);
  not (_04793_, _02173_);
  nor (_04794_, _04793_, _01790_);
  not (_04795_, _04789_);
  nor (_04796_, _04770_, _04795_);
  or (_04797_, _04796_, _04794_);
  or (_04798_, _04797_, _04792_);
  not (_04799_, _01636_);
  nand (_04800_, _04778_, _04794_);
  and (_04801_, _04800_, _04799_);
  and (_04802_, _04801_, _04798_);
  nand (_04803_, _04387_, _01636_);
  nor (_04804_, _02718_, _02387_);
  nand (_04805_, _04804_, _04803_);
  or (_04806_, _04805_, _04802_);
  not (_04807_, _02930_);
  or (_04808_, _04804_, _04379_);
  and (_04809_, _04808_, _04807_);
  and (_04810_, _04809_, _04806_);
  and (_04811_, _04379_, _02930_);
  or (_04812_, _04811_, _02935_);
  or (_04813_, _04812_, _04810_);
  not (_04814_, _02934_);
  not (_04815_, _02935_);
  not (_04816_, _04483_);
  or (_04817_, _04428_, \oc8051_golden_model_1.IRAM[9] [6]);
  or (_04818_, _04438_, \oc8051_golden_model_1.IRAM[8] [6]);
  and (_04819_, _04818_, _04437_);
  and (_04820_, _04819_, _04817_);
  or (_04821_, _04438_, \oc8051_golden_model_1.IRAM[10] [6]);
  or (_04822_, _04428_, \oc8051_golden_model_1.IRAM[11] [6]);
  and (_04823_, _04822_, _04436_);
  and (_04824_, _04823_, _04821_);
  nor (_04825_, _04824_, _04820_);
  nand (_04826_, _04825_, _04420_);
  or (_04827_, _04428_, \oc8051_golden_model_1.IRAM[13] [6]);
  or (_04828_, _04438_, \oc8051_golden_model_1.IRAM[12] [6]);
  and (_04829_, _04828_, _04437_);
  and (_04830_, _04829_, _04827_);
  or (_04831_, _04438_, \oc8051_golden_model_1.IRAM[14] [6]);
  or (_04832_, _04428_, \oc8051_golden_model_1.IRAM[15] [6]);
  and (_04833_, _04832_, _04436_);
  and (_04834_, _04833_, _04831_);
  nor (_04835_, _04834_, _04830_);
  nand (_04836_, _04835_, _04448_);
  nand (_04837_, _04836_, _04826_);
  nand (_04838_, _04837_, _04410_);
  or (_04839_, _04428_, _03758_);
  nand (_04840_, _04428_, \oc8051_golden_model_1.IRAM[0] [6]);
  and (_04841_, _04840_, _04437_);
  nand (_04842_, _04841_, _04839_);
  nand (_04843_, _04428_, \oc8051_golden_model_1.IRAM[2] [6]);
  or (_04844_, _04428_, _03762_);
  and (_04845_, _04844_, _04436_);
  nand (_04846_, _04845_, _04843_);
  nand (_04847_, _04846_, _04842_);
  nand (_04848_, _04847_, _04420_);
  nand (_04849_, _04428_, \oc8051_golden_model_1.IRAM[4] [6]);
  or (_04850_, _04428_, _03778_);
  and (_04851_, _04850_, _04437_);
  nand (_04852_, _04851_, _04849_);
  nand (_04853_, _04428_, \oc8051_golden_model_1.IRAM[6] [6]);
  or (_04854_, _04428_, _03770_);
  and (_04855_, _04854_, _04436_);
  nand (_04856_, _04855_, _04853_);
  nand (_04857_, _04856_, _04852_);
  nand (_04858_, _04857_, _04448_);
  nand (_04859_, _04858_, _04848_);
  nand (_04860_, _04859_, _04409_);
  and (_04861_, _04860_, _04838_);
  not (_04862_, _04861_);
  or (_04863_, _04428_, \oc8051_golden_model_1.IRAM[9] [1]);
  nand (_04864_, _04428_, _02788_);
  and (_04865_, _04864_, _04437_);
  and (_04866_, _04865_, _04863_);
  or (_04867_, _04438_, \oc8051_golden_model_1.IRAM[10] [1]);
  or (_04868_, _04428_, \oc8051_golden_model_1.IRAM[11] [1]);
  and (_04869_, _04868_, _04436_);
  and (_04870_, _04869_, _04867_);
  nor (_04871_, _04870_, _04866_);
  nand (_04872_, _04871_, _04420_);
  or (_04873_, _04428_, \oc8051_golden_model_1.IRAM[13] [1]);
  nand (_04874_, _04428_, _02801_);
  and (_04875_, _04874_, _04437_);
  and (_04876_, _04875_, _04873_);
  nand (_04877_, _04428_, _02797_);
  or (_04878_, _04428_, \oc8051_golden_model_1.IRAM[15] [1]);
  and (_04879_, _04878_, _04436_);
  and (_04880_, _04879_, _04877_);
  nor (_04881_, _04880_, _04876_);
  nand (_04882_, _04881_, _04448_);
  nand (_04883_, _04882_, _04872_);
  nand (_04884_, _04883_, _04410_);
  or (_04885_, _04428_, _02750_);
  nand (_04886_, _04428_, \oc8051_golden_model_1.IRAM[0] [1]);
  and (_04887_, _04886_, _04437_);
  nand (_04888_, _04887_, _04885_);
  nand (_04889_, _04428_, \oc8051_golden_model_1.IRAM[2] [1]);
  or (_04890_, _04428_, _02755_);
  and (_04891_, _04890_, _04436_);
  nand (_04892_, _04891_, _04889_);
  nand (_04893_, _04892_, _04888_);
  nand (_04894_, _04893_, _04420_);
  nand (_04895_, _04428_, \oc8051_golden_model_1.IRAM[4] [1]);
  or (_04896_, _04428_, _02773_);
  and (_04897_, _04896_, _04437_);
  nand (_04898_, _04897_, _04895_);
  nand (_04899_, _04428_, \oc8051_golden_model_1.IRAM[6] [1]);
  or (_04900_, _04428_, _02765_);
  and (_04901_, _04900_, _04436_);
  nand (_04902_, _04901_, _04899_);
  nand (_04903_, _04902_, _04898_);
  nand (_04904_, _04903_, _04448_);
  nand (_04905_, _04904_, _04894_);
  nand (_04906_, _04905_, _04409_);
  and (_04907_, _04906_, _04884_);
  or (_04908_, _04428_, \oc8051_golden_model_1.IRAM[9] [0]);
  nand (_04909_, _04428_, _03009_);
  and (_04910_, _04909_, _04437_);
  and (_04911_, _04910_, _04908_);
  or (_04912_, _04438_, \oc8051_golden_model_1.IRAM[10] [0]);
  or (_04913_, _04428_, \oc8051_golden_model_1.IRAM[11] [0]);
  and (_04914_, _04913_, _04436_);
  and (_04915_, _04914_, _04912_);
  nor (_04916_, _04915_, _04911_);
  nand (_04917_, _04916_, _04420_);
  or (_04918_, _04428_, \oc8051_golden_model_1.IRAM[13] [0]);
  or (_04919_, _04438_, \oc8051_golden_model_1.IRAM[12] [0]);
  and (_04920_, _04919_, _04437_);
  and (_04921_, _04920_, _04918_);
  or (_04922_, _04438_, \oc8051_golden_model_1.IRAM[14] [0]);
  or (_04923_, _04428_, \oc8051_golden_model_1.IRAM[15] [0]);
  and (_04924_, _04923_, _04436_);
  and (_04925_, _04924_, _04922_);
  nor (_04926_, _04925_, _04921_);
  nand (_04927_, _04926_, _04448_);
  nand (_04928_, _04927_, _04917_);
  nand (_04929_, _04928_, _04410_);
  or (_04930_, _04428_, _02977_);
  nand (_04931_, _04428_, \oc8051_golden_model_1.IRAM[0] [0]);
  and (_04932_, _04931_, _04437_);
  nand (_04933_, _04932_, _04930_);
  nand (_04934_, _04428_, \oc8051_golden_model_1.IRAM[2] [0]);
  or (_04935_, _04428_, _02981_);
  and (_04936_, _04935_, _04436_);
  nand (_04937_, _04936_, _04934_);
  nand (_04938_, _04937_, _04933_);
  nand (_04939_, _04938_, _04420_);
  nand (_04940_, _04428_, \oc8051_golden_model_1.IRAM[4] [0]);
  or (_04941_, _04428_, _02997_);
  and (_04942_, _04941_, _04437_);
  nand (_04943_, _04942_, _04940_);
  nand (_04944_, _04428_, \oc8051_golden_model_1.IRAM[6] [0]);
  or (_04945_, _04428_, _02989_);
  and (_04946_, _04945_, _04436_);
  nand (_04947_, _04946_, _04944_);
  nand (_04948_, _04947_, _04943_);
  nand (_04949_, _04948_, _04448_);
  nand (_04950_, _04949_, _04939_);
  nand (_04951_, _04950_, _04409_);
  and (_04952_, _04951_, _04929_);
  nor (_04953_, _04952_, _04907_);
  or (_04954_, _04428_, \oc8051_golden_model_1.IRAM[9] [3]);
  or (_04955_, _04438_, \oc8051_golden_model_1.IRAM[8] [3]);
  and (_04956_, _04955_, _04437_);
  and (_04957_, _04956_, _04954_);
  or (_04958_, _04438_, \oc8051_golden_model_1.IRAM[10] [3]);
  or (_04959_, _04428_, \oc8051_golden_model_1.IRAM[11] [3]);
  and (_04960_, _04959_, _04436_);
  and (_04961_, _04960_, _04958_);
  nor (_04962_, _04961_, _04957_);
  nand (_04963_, _04962_, _04420_);
  or (_04964_, _04428_, \oc8051_golden_model_1.IRAM[13] [3]);
  or (_04965_, _04438_, \oc8051_golden_model_1.IRAM[12] [3]);
  and (_04966_, _04965_, _04437_);
  and (_04967_, _04966_, _04964_);
  or (_04968_, _04438_, \oc8051_golden_model_1.IRAM[14] [3]);
  or (_04969_, _04428_, \oc8051_golden_model_1.IRAM[15] [3]);
  and (_04970_, _04969_, _04436_);
  and (_04971_, _04970_, _04968_);
  nor (_04972_, _04971_, _04967_);
  nand (_04973_, _04972_, _04448_);
  nand (_04974_, _04973_, _04963_);
  nand (_04975_, _04974_, _04410_);
  or (_04976_, _04428_, _03195_);
  nand (_04977_, _04428_, \oc8051_golden_model_1.IRAM[0] [3]);
  and (_04978_, _04977_, _04437_);
  nand (_04979_, _04978_, _04976_);
  nand (_04980_, _04428_, \oc8051_golden_model_1.IRAM[2] [3]);
  or (_04981_, _04428_, _03200_);
  and (_04982_, _04981_, _04436_);
  nand (_04983_, _04982_, _04980_);
  nand (_04984_, _04983_, _04979_);
  nand (_04985_, _04984_, _04420_);
  nand (_04986_, _04428_, \oc8051_golden_model_1.IRAM[4] [3]);
  or (_04987_, _04428_, _03225_);
  and (_04988_, _04987_, _04437_);
  nand (_04989_, _04988_, _04986_);
  nand (_04990_, _04428_, \oc8051_golden_model_1.IRAM[6] [3]);
  or (_04991_, _04428_, _03213_);
  and (_04992_, _04991_, _04436_);
  nand (_04993_, _04992_, _04990_);
  nand (_04994_, _04993_, _04989_);
  nand (_04995_, _04994_, _04448_);
  nand (_04996_, _04995_, _04985_);
  nand (_04997_, _04996_, _04409_);
  and (_04998_, _04997_, _04975_);
  or (_04999_, _04428_, \oc8051_golden_model_1.IRAM[9] [2]);
  nand (_05000_, _04428_, _03432_);
  and (_05001_, _05000_, _04437_);
  and (_05002_, _05001_, _04999_);
  nand (_05003_, _04428_, _03428_);
  or (_05004_, _04428_, \oc8051_golden_model_1.IRAM[11] [2]);
  and (_05005_, _05004_, _04436_);
  and (_05006_, _05005_, _05003_);
  nor (_05007_, _05006_, _05002_);
  nand (_05008_, _05007_, _04420_);
  or (_05009_, _04428_, \oc8051_golden_model_1.IRAM[13] [2]);
  nand (_05010_, _04428_, _03445_);
  and (_05011_, _05010_, _04437_);
  and (_05012_, _05011_, _05009_);
  nand (_05013_, _04428_, _03441_);
  or (_05014_, _04428_, \oc8051_golden_model_1.IRAM[15] [2]);
  and (_05015_, _05014_, _04436_);
  and (_05016_, _05015_, _05013_);
  nor (_05017_, _05016_, _05012_);
  nand (_05018_, _05017_, _04448_);
  nand (_05019_, _05018_, _05008_);
  nand (_05020_, _05019_, _04410_);
  or (_05021_, _04428_, _03399_);
  nand (_05022_, _04428_, \oc8051_golden_model_1.IRAM[0] [2]);
  and (_05023_, _05022_, _04437_);
  nand (_05024_, _05023_, _05021_);
  nand (_05025_, _04428_, \oc8051_golden_model_1.IRAM[2] [2]);
  or (_05026_, _04428_, _03403_);
  and (_05027_, _05026_, _04436_);
  nand (_05028_, _05027_, _05025_);
  nand (_05029_, _05028_, _05024_);
  nand (_05030_, _05029_, _04420_);
  nand (_05031_, _04428_, \oc8051_golden_model_1.IRAM[4] [2]);
  or (_05032_, _04428_, _03419_);
  and (_05033_, _05032_, _04437_);
  nand (_05034_, _05033_, _05031_);
  nand (_05035_, _04428_, \oc8051_golden_model_1.IRAM[6] [2]);
  or (_05036_, _04428_, _03411_);
  and (_05037_, _05036_, _04436_);
  nand (_05038_, _05037_, _05035_);
  nand (_05039_, _05038_, _05034_);
  nand (_05040_, _05039_, _04448_);
  nand (_05041_, _05040_, _05030_);
  nand (_05042_, _05041_, _04409_);
  and (_05043_, _05042_, _05020_);
  nor (_05044_, _05043_, _04998_);
  and (_05045_, _05044_, _04953_);
  or (_05046_, _04428_, \oc8051_golden_model_1.IRAM[9] [5]);
  or (_05047_, _04438_, \oc8051_golden_model_1.IRAM[8] [5]);
  and (_05048_, _05047_, _04437_);
  and (_05049_, _05048_, _05046_);
  or (_05050_, _04438_, \oc8051_golden_model_1.IRAM[10] [5]);
  or (_05051_, _04428_, \oc8051_golden_model_1.IRAM[11] [5]);
  and (_05052_, _05051_, _04436_);
  and (_05053_, _05052_, _05050_);
  nor (_05054_, _05053_, _05049_);
  nand (_05055_, _05054_, _04420_);
  or (_05056_, _04428_, \oc8051_golden_model_1.IRAM[13] [5]);
  or (_05057_, _04438_, \oc8051_golden_model_1.IRAM[12] [5]);
  and (_05058_, _05057_, _04437_);
  and (_05059_, _05058_, _05056_);
  or (_05060_, _04438_, \oc8051_golden_model_1.IRAM[14] [5]);
  or (_05061_, _04428_, \oc8051_golden_model_1.IRAM[15] [5]);
  and (_05062_, _05061_, _04436_);
  and (_05063_, _05062_, _05060_);
  nor (_05064_, _05063_, _05059_);
  nand (_05065_, _05064_, _04448_);
  nand (_05066_, _05065_, _05055_);
  nand (_05067_, _05066_, _04410_);
  or (_05068_, _04428_, _03866_);
  nand (_05069_, _04428_, \oc8051_golden_model_1.IRAM[0] [5]);
  and (_05070_, _05069_, _04437_);
  nand (_05071_, _05070_, _05068_);
  nand (_05072_, _04428_, \oc8051_golden_model_1.IRAM[2] [5]);
  or (_05073_, _04428_, _03870_);
  and (_05074_, _05073_, _04436_);
  nand (_05075_, _05074_, _05072_);
  nand (_05076_, _05075_, _05071_);
  nand (_05077_, _05076_, _04420_);
  nand (_05078_, _04428_, \oc8051_golden_model_1.IRAM[4] [5]);
  or (_05079_, _04428_, _03886_);
  and (_05080_, _05079_, _04437_);
  nand (_05081_, _05080_, _05078_);
  nand (_05082_, _04428_, \oc8051_golden_model_1.IRAM[6] [5]);
  or (_05083_, _04428_, _03878_);
  and (_05084_, _05083_, _04436_);
  nand (_05085_, _05084_, _05082_);
  nand (_05086_, _05085_, _05081_);
  nand (_05087_, _05086_, _04448_);
  nand (_05088_, _05087_, _05077_);
  nand (_05089_, _05088_, _04409_);
  and (_05090_, _05089_, _05067_);
  or (_05091_, _04428_, \oc8051_golden_model_1.IRAM[9] [4]);
  or (_05092_, _04438_, \oc8051_golden_model_1.IRAM[8] [4]);
  and (_05093_, _05092_, _04437_);
  and (_05094_, _05093_, _05091_);
  or (_05095_, _04438_, \oc8051_golden_model_1.IRAM[10] [4]);
  or (_05096_, _04428_, \oc8051_golden_model_1.IRAM[11] [4]);
  and (_05097_, _05096_, _04436_);
  and (_05098_, _05097_, _05095_);
  nor (_05099_, _05098_, _05094_);
  nand (_05100_, _05099_, _04420_);
  or (_05101_, _04428_, \oc8051_golden_model_1.IRAM[13] [4]);
  or (_05102_, _04438_, \oc8051_golden_model_1.IRAM[12] [4]);
  and (_05103_, _05102_, _04437_);
  and (_05104_, _05103_, _05101_);
  or (_05105_, _04438_, \oc8051_golden_model_1.IRAM[14] [4]);
  or (_05106_, _04428_, \oc8051_golden_model_1.IRAM[15] [4]);
  and (_05107_, _05106_, _04436_);
  and (_05108_, _05107_, _05105_);
  nor (_05109_, _05108_, _05104_);
  nand (_05110_, _05109_, _04448_);
  nand (_05111_, _05110_, _05100_);
  nand (_05112_, _05111_, _04410_);
  or (_05113_, _04428_, _04161_);
  nand (_05114_, _04428_, \oc8051_golden_model_1.IRAM[0] [4]);
  and (_05115_, _05114_, _04437_);
  nand (_05116_, _05115_, _05113_);
  nand (_05117_, _04428_, \oc8051_golden_model_1.IRAM[2] [4]);
  or (_05118_, _04428_, _04165_);
  and (_05119_, _05118_, _04436_);
  nand (_05120_, _05119_, _05117_);
  nand (_05121_, _05120_, _05116_);
  nand (_05122_, _05121_, _04420_);
  nand (_05123_, _04428_, \oc8051_golden_model_1.IRAM[4] [4]);
  or (_05124_, _04428_, _04181_);
  and (_05125_, _05124_, _04437_);
  nand (_05126_, _05125_, _05123_);
  nand (_05127_, _04428_, \oc8051_golden_model_1.IRAM[6] [4]);
  or (_05128_, _04428_, _04173_);
  and (_05129_, _05128_, _04436_);
  nand (_05130_, _05129_, _05127_);
  nand (_05131_, _05130_, _05126_);
  nand (_05132_, _05131_, _04448_);
  nand (_05133_, _05132_, _05122_);
  nand (_05134_, _05133_, _04409_);
  and (_05135_, _05134_, _05112_);
  nor (_05136_, _05135_, _05090_);
  and (_05137_, _05136_, _05045_);
  and (_05138_, _05137_, _04862_);
  nor (_05139_, _05138_, _04816_);
  and (_05140_, _05138_, _04816_);
  or (_05141_, _05140_, _05139_);
  or (_05142_, _05141_, _04815_);
  and (_05143_, _05142_, _04814_);
  and (_05144_, _05143_, _04813_);
  and (_05145_, _04496_, _02934_);
  or (_05146_, _05145_, _02058_);
  or (_05147_, _05146_, _05144_);
  and (_05148_, _05147_, _04276_);
  or (_05149_, _05148_, _01642_);
  and (_05150_, _04388_, _01642_);
  nor (_05151_, _05150_, _02941_);
  and (_05152_, _05151_, _05149_);
  nand (_05153_, _04349_, _02941_);
  nor (_05154_, _02705_, _02378_);
  nand (_05155_, _05154_, _05153_);
  or (_05156_, _05155_, _05152_);
  not (_05157_, _02948_);
  not (_05158_, _03808_);
  not (_05159_, _03916_);
  not (_05160_, _04211_);
  nor (_05161_, _03042_, _02811_);
  nor (_05162_, _03455_, _03268_);
  and (_05163_, _05162_, _05161_);
  and (_05164_, _05163_, _05160_);
  and (_05165_, _05164_, _05159_);
  nand (_05166_, _05165_, _05158_);
  nor (_05167_, _05166_, _04370_);
  and (_05168_, _05166_, _04370_);
  or (_05169_, _05168_, _05167_);
  and (_05170_, _05169_, _05157_);
  and (_05171_, _01533_, _01403_);
  not (_05172_, _05171_);
  or (_05173_, _05172_, _05170_);
  and (_05174_, _05173_, _05156_);
  and (_05175_, _05169_, _02948_);
  or (_05176_, _05175_, _02952_);
  or (_05177_, _05176_, _05174_);
  not (_05178_, _02952_);
  and (_05179_, _04952_, _04907_);
  and (_05180_, _05043_, _04998_);
  and (_05181_, _05180_, _05179_);
  and (_05182_, _05135_, _05090_);
  and (_05183_, _05182_, _05181_);
  and (_05184_, _05183_, _04861_);
  nand (_05185_, _05184_, _04483_);
  or (_05186_, _05184_, _04483_);
  and (_05187_, _05186_, _05185_);
  or (_05188_, _05187_, _05178_);
  and (_05189_, _05188_, _03118_);
  and (_05190_, _05189_, _05177_);
  or (_05191_, _05190_, _04265_);
  and (_05192_, _05191_, _03186_);
  or (_05193_, _05192_, _03562_);
  and (_05194_, _05193_, _03561_);
  not (_05195_, _02058_);
  and (_05196_, \oc8051_golden_model_1.PC [9], \oc8051_golden_model_1.PC [8]);
  and (_05197_, _05196_, \oc8051_golden_model_1.PC [10]);
  and (_05198_, _05197_, _04385_);
  and (_05199_, _05198_, \oc8051_golden_model_1.PC [11]);
  and (_05200_, _05199_, \oc8051_golden_model_1.PC [12]);
  and (_05201_, _05200_, \oc8051_golden_model_1.PC [13]);
  and (_05202_, _05201_, \oc8051_golden_model_1.PC [14]);
  nor (_05203_, _05202_, \oc8051_golden_model_1.PC [15]);
  and (_05204_, _04385_, \oc8051_golden_model_1.PC [8]);
  and (_05205_, _05204_, \oc8051_golden_model_1.PC [9]);
  and (_05206_, _05205_, \oc8051_golden_model_1.PC [10]);
  and (_05207_, _05206_, \oc8051_golden_model_1.PC [11]);
  and (_05208_, _05207_, \oc8051_golden_model_1.PC [12]);
  and (_05209_, _05208_, \oc8051_golden_model_1.PC [13]);
  and (_05210_, _05209_, \oc8051_golden_model_1.PC [14]);
  and (_05211_, _05210_, \oc8051_golden_model_1.PC [15]);
  nor (_05212_, _05211_, _05203_);
  and (_05213_, _05212_, _05195_);
  and (_05214_, _05197_, _04271_);
  and (_05215_, _05214_, \oc8051_golden_model_1.PC [11]);
  and (_05216_, _05215_, \oc8051_golden_model_1.PC [12]);
  and (_05217_, _05216_, \oc8051_golden_model_1.PC [13]);
  and (_05218_, _05217_, \oc8051_golden_model_1.PC [14]);
  nor (_05219_, _05218_, \oc8051_golden_model_1.PC [15]);
  and (_05220_, _04271_, \oc8051_golden_model_1.PC [8]);
  and (_05221_, _05220_, \oc8051_golden_model_1.PC [9]);
  and (_05222_, _05221_, \oc8051_golden_model_1.PC [10]);
  and (_05223_, _05222_, \oc8051_golden_model_1.PC [11]);
  and (_05224_, _05223_, \oc8051_golden_model_1.PC [12]);
  and (_05225_, _05224_, \oc8051_golden_model_1.PC [13]);
  and (_05226_, _05225_, \oc8051_golden_model_1.PC [14]);
  and (_05227_, _05226_, \oc8051_golden_model_1.PC [15]);
  nor (_05228_, _05227_, _05219_);
  and (_05229_, _05228_, _02058_);
  or (_05230_, _05229_, _05213_);
  and (_05231_, _05230_, _03556_);
  and (_05232_, _05231_, _03559_);
  or (_37136_, _05232_, _05194_);
  not (_05233_, \oc8051_golden_model_1.B [7]);
  nor (_05234_, _38087_, _05233_);
  nor (_05235_, _03683_, _05233_);
  and (_05236_, _04779_, _03683_);
  or (_05237_, _05236_, _05235_);
  and (_05238_, _05237_, _02167_);
  not (_05239_, _03683_);
  nor (_05240_, _05239_, _03616_);
  or (_05241_, _05240_, _05235_);
  nor (_05242_, _02465_, _02049_);
  nor (_05243_, _05242_, _02531_);
  not (_05244_, _05243_);
  not (_05245_, _02354_);
  and (_05246_, _02690_, _01601_);
  nor (_05247_, _05246_, _02362_);
  and (_05248_, _05247_, _05245_);
  and (_05249_, _05248_, _05244_);
  or (_05250_, _05249_, _05241_);
  nor (_05251_, _04318_, _05233_);
  and (_05252_, _04364_, _04318_);
  or (_05253_, _05252_, _05251_);
  and (_05254_, _05253_, _01997_);
  and (_05255_, _04496_, _03683_);
  or (_05256_, _05255_, _05235_);
  or (_05257_, _05256_, _02814_);
  and (_05258_, _03683_, \oc8051_golden_model_1.ACC [7]);
  or (_05259_, _05258_, _05235_);
  and (_05260_, _05259_, _02817_);
  nor (_05261_, _02817_, _05233_);
  or (_05262_, _05261_, _02001_);
  or (_05263_, _05262_, _05260_);
  and (_05264_, _05263_, _02024_);
  and (_05265_, _05264_, _05257_);
  and (_05266_, _04368_, _04318_);
  or (_05267_, _05266_, _05251_);
  and (_05268_, _05267_, _02007_);
  or (_05269_, _05268_, _01999_);
  or (_05270_, _05269_, _05265_);
  or (_05271_, _05241_, _02840_);
  and (_05272_, _05271_, _05270_);
  or (_05273_, _05272_, _02006_);
  or (_05274_, _05259_, _02021_);
  and (_05275_, _05274_, _02025_);
  and (_05276_, _05275_, _05273_);
  or (_05277_, _05276_, _05254_);
  and (_05278_, _05277_, _02861_);
  and (_05279_, _02044_, _01965_);
  or (_05280_, _05251_, _04533_);
  and (_05281_, _05280_, _01991_);
  and (_05282_, _05281_, _05267_);
  or (_05283_, _05282_, _05279_);
  or (_05284_, _05283_, _05278_);
  not (_05285_, _05279_);
  and (_05286_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [7]);
  and (_05287_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [6]);
  and (_05288_, _05287_, _05286_);
  and (_05289_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [7]);
  and (_05290_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [6]);
  nor (_05291_, _05290_, _05289_);
  nor (_05292_, _05291_, _05288_);
  and (_05293_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [4]);
  and (_05294_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [3]);
  and (_05295_, _05294_, _05293_);
  and (_05296_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [7]);
  and (_05297_, _05296_, _05287_);
  and (_05298_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [5]);
  nor (_05299_, _05296_, _05287_);
  nor (_05300_, _05299_, _05297_);
  and (_05301_, _05300_, _05298_);
  nor (_05302_, _05301_, _05297_);
  and (_05303_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [4]);
  and (_05304_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [5]);
  and (_05305_, _05304_, _05303_);
  nor (_05306_, _05304_, _05303_);
  nor (_05307_, _05306_, _05305_);
  not (_05308_, _05307_);
  nor (_05309_, _05308_, _05302_);
  and (_05310_, _05308_, _05302_);
  nor (_05311_, _05310_, _05309_);
  and (_05312_, _05311_, _05295_);
  nor (_05313_, _05311_, _05295_);
  nor (_05314_, _05313_, _05312_);
  and (_05315_, _05314_, _05292_);
  and (_05316_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [5]);
  and (_05317_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [6]);
  and (_05318_, _05317_, _05316_);
  nor (_05319_, _05317_, _05316_);
  nor (_05320_, _05319_, _05318_);
  and (_05321_, _05320_, _05288_);
  nor (_05322_, _05320_, _05288_);
  nor (_05324_, _05322_, _05321_);
  and (_05325_, _05324_, _05305_);
  nor (_05326_, _05324_, _05305_);
  nor (_05327_, _05326_, _05325_);
  and (_05328_, _05327_, _05286_);
  nor (_05329_, _05327_, _05286_);
  nor (_05330_, _05329_, _05328_);
  and (_05331_, _05330_, _05315_);
  nor (_05332_, _05312_, _05309_);
  not (_05333_, _05332_);
  nor (_05334_, _05330_, _05315_);
  nor (_05335_, _05334_, _05331_);
  and (_05336_, _05335_, _05333_);
  nor (_05337_, _05336_, _05331_);
  nor (_05338_, _05325_, _05321_);
  not (_05339_, _05338_);
  and (_05340_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [6]);
  and (_05341_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [7]);
  and (_05342_, _05341_, _05340_);
  nor (_05343_, _05341_, _05340_);
  nor (_05344_, _05343_, _05342_);
  and (_05345_, _05344_, _05318_);
  nor (_05346_, _05344_, _05318_);
  nor (_05347_, _05346_, _05345_);
  and (_05348_, _05347_, _05328_);
  nor (_05349_, _05347_, _05328_);
  nor (_05350_, _05349_, _05348_);
  and (_05351_, _05350_, _05339_);
  nor (_05352_, _05350_, _05339_);
  nor (_05353_, _05352_, _05351_);
  not (_05354_, _05353_);
  nor (_05355_, _05354_, _05337_);
  and (_05356_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [7]);
  not (_05357_, _05356_);
  nor (_05358_, _05357_, _05317_);
  nor (_05359_, _05358_, _05345_);
  nor (_05360_, _05351_, _05348_);
  nor (_05361_, _05360_, _05359_);
  and (_05362_, _05360_, _05359_);
  nor (_05363_, _05362_, _05361_);
  and (_05364_, _05363_, _05355_);
  or (_05365_, _05361_, _05342_);
  or (_05366_, _05365_, _05364_);
  and (_05367_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [6]);
  and (_05368_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [7]);
  and (_05369_, _05368_, _05367_);
  not (_05370_, _05367_);
  and (_05371_, _05368_, _05370_);
  and (_05372_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [4]);
  and (_05373_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [5]);
  and (_05374_, _05373_, _05287_);
  and (_05375_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [6]);
  and (_05376_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [5]);
  nor (_05377_, _05376_, _05375_);
  nor (_05378_, _05377_, _05374_);
  and (_05379_, _05378_, _05372_);
  nor (_05380_, _05378_, _05372_);
  nor (_05381_, _05380_, _05379_);
  and (_05382_, _05381_, _05371_);
  nor (_05383_, _05382_, _05369_);
  nor (_05384_, _05300_, _05298_);
  nor (_05385_, _05384_, _05301_);
  not (_05386_, _05385_);
  nor (_05387_, _05386_, _05383_);
  and (_05388_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [3]);
  and (_05389_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [2]);
  and (_05390_, _05389_, _05388_);
  nor (_05391_, _05379_, _05374_);
  nor (_05392_, _05294_, _05293_);
  nor (_05393_, _05392_, _05295_);
  not (_05394_, _05393_);
  nor (_05395_, _05394_, _05391_);
  and (_05396_, _05394_, _05391_);
  nor (_05397_, _05396_, _05395_);
  and (_05398_, _05397_, _05390_);
  nor (_05399_, _05397_, _05390_);
  nor (_05400_, _05399_, _05398_);
  and (_05401_, _05386_, _05383_);
  nor (_05402_, _05401_, _05387_);
  and (_05403_, _05402_, _05400_);
  nor (_05404_, _05403_, _05387_);
  not (_05405_, _05404_);
  nor (_05406_, _05314_, _05292_);
  nor (_05407_, _05406_, _05315_);
  and (_05408_, _05407_, _05405_);
  nor (_05409_, _05398_, _05395_);
  not (_05410_, _05409_);
  nor (_05411_, _05407_, _05405_);
  nor (_05412_, _05411_, _05408_);
  and (_05413_, _05412_, _05410_);
  nor (_05414_, _05413_, _05408_);
  nor (_05415_, _05335_, _05333_);
  nor (_05416_, _05415_, _05336_);
  not (_05417_, _05416_);
  nor (_05418_, _05417_, _05414_);
  and (_05419_, _05354_, _05337_);
  nor (_05420_, _05419_, _05355_);
  and (_05421_, _05420_, _05418_);
  and (_05422_, _05421_, _05363_);
  and (_05423_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [7]);
  and (_05424_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [6]);
  and (_05425_, _05424_, _05423_);
  and (_05426_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [5]);
  and (_05427_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [7]);
  nor (_05428_, _05427_, _05367_);
  nor (_05429_, _05428_, _05425_);
  and (_05430_, _05429_, _05426_);
  nor (_05431_, _05430_, _05425_);
  and (_05432_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [6]);
  nor (_05433_, _05432_, _05423_);
  nor (_05434_, _05433_, _05369_);
  not (_05435_, _05434_);
  nor (_05436_, _05435_, _05431_);
  and (_05437_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [3]);
  and (_05438_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [4]);
  and (_05439_, _05438_, _05373_);
  nor (_05440_, _05438_, _05373_);
  nor (_05441_, _05440_, _05439_);
  and (_05442_, _05441_, _05437_);
  nor (_05443_, _05441_, _05437_);
  nor (_05444_, _05443_, _05442_);
  and (_05445_, _05435_, _05431_);
  nor (_05446_, _05445_, _05436_);
  and (_05447_, _05446_, _05444_);
  nor (_05448_, _05447_, _05436_);
  nor (_05449_, _05381_, _05371_);
  nor (_05450_, _05449_, _05382_);
  not (_05451_, _05450_);
  nor (_05452_, _05451_, _05448_);
  and (_05453_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [2]);
  and (_05454_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [1]);
  and (_05455_, _05454_, _05453_);
  nor (_05456_, _05442_, _05439_);
  nor (_05457_, _05389_, _05388_);
  nor (_05458_, _05457_, _05390_);
  not (_05459_, _05458_);
  nor (_05460_, _05459_, _05456_);
  and (_05461_, _05459_, _05456_);
  nor (_05462_, _05461_, _05460_);
  and (_05463_, _05462_, _05455_);
  nor (_05464_, _05462_, _05455_);
  nor (_05465_, _05464_, _05463_);
  and (_05466_, _05451_, _05448_);
  nor (_05467_, _05466_, _05452_);
  and (_05468_, _05467_, _05465_);
  nor (_05469_, _05468_, _05452_);
  nor (_05470_, _05402_, _05400_);
  nor (_05471_, _05470_, _05403_);
  not (_05472_, _05471_);
  nor (_05473_, _05472_, _05469_);
  nor (_05474_, _05463_, _05460_);
  not (_05475_, _05474_);
  and (_05476_, _05472_, _05469_);
  nor (_05477_, _05476_, _05473_);
  and (_05478_, _05477_, _05475_);
  nor (_05479_, _05478_, _05473_);
  nor (_05480_, _05412_, _05410_);
  nor (_05481_, _05480_, _05413_);
  not (_05482_, _05481_);
  nor (_05483_, _05482_, _05479_);
  and (_05484_, _05417_, _05414_);
  nor (_05485_, _05484_, _05418_);
  and (_05486_, _05485_, _05483_);
  nor (_05487_, _05420_, _05418_);
  nor (_05488_, _05487_, _05421_);
  and (_05489_, _05488_, _05486_);
  nor (_05490_, _05488_, _05486_);
  and (_05491_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [5]);
  and (_05492_, _05491_, _05367_);
  and (_05493_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [4]);
  and (_05494_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [5]);
  nor (_05495_, _05494_, _05424_);
  nor (_05496_, _05495_, _05492_);
  and (_05497_, _05496_, _05493_);
  nor (_05498_, _05497_, _05492_);
  not (_05499_, _05498_);
  nor (_05500_, _05429_, _05426_);
  nor (_05501_, _05500_, _05430_);
  and (_05502_, _05501_, _05499_);
  and (_05503_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [2]);
  and (_05504_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [4]);
  and (_05505_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [3]);
  and (_05506_, _05505_, _05504_);
  nor (_05507_, _05505_, _05504_);
  nor (_05508_, _05507_, _05506_);
  and (_05509_, _05508_, _05503_);
  nor (_05510_, _05508_, _05503_);
  nor (_05511_, _05510_, _05509_);
  nor (_05512_, _05501_, _05499_);
  nor (_05513_, _05512_, _05502_);
  and (_05514_, _05513_, _05511_);
  nor (_05515_, _05514_, _05502_);
  nor (_05516_, _05446_, _05444_);
  nor (_05517_, _05516_, _05447_);
  not (_05518_, _05517_);
  nor (_05519_, _05518_, _05515_);
  and (_05520_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [0]);
  and (_05521_, _05520_, _05454_);
  nor (_05522_, _05509_, _05506_);
  nor (_05523_, _05454_, _05453_);
  nor (_05524_, _05523_, _05455_);
  not (_05525_, _05524_);
  nor (_05526_, _05525_, _05522_);
  and (_05527_, _05525_, _05522_);
  nor (_05528_, _05527_, _05526_);
  and (_05529_, _05528_, _05521_);
  nor (_05530_, _05528_, _05521_);
  nor (_05531_, _05530_, _05529_);
  and (_05532_, _05518_, _05515_);
  nor (_05533_, _05532_, _05519_);
  and (_05534_, _05533_, _05531_);
  nor (_05535_, _05534_, _05519_);
  nor (_05536_, _05467_, _05465_);
  nor (_05537_, _05536_, _05468_);
  not (_05538_, _05537_);
  nor (_05539_, _05538_, _05535_);
  nor (_05540_, _05529_, _05526_);
  not (_05541_, _05540_);
  and (_05542_, _05538_, _05535_);
  nor (_05543_, _05542_, _05539_);
  and (_05544_, _05543_, _05541_);
  nor (_05545_, _05544_, _05539_);
  nor (_05546_, _05477_, _05475_);
  nor (_05547_, _05546_, _05478_);
  not (_05548_, _05547_);
  nor (_05549_, _05548_, _05545_);
  and (_05550_, _05482_, _05479_);
  nor (_05551_, _05550_, _05483_);
  and (_05552_, _05551_, _05549_);
  nor (_05553_, _05485_, _05483_);
  nor (_05554_, _05553_, _05486_);
  nand (_05555_, _05554_, _05552_);
  and (_05556_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [4]);
  and (_05557_, _05556_, _05491_);
  and (_05558_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [3]);
  nor (_05559_, _05556_, _05491_);
  nor (_05560_, _05559_, _05557_);
  and (_05561_, _05560_, _05558_);
  nor (_05562_, _05561_, _05557_);
  not (_05563_, _05562_);
  nor (_05564_, _05496_, _05493_);
  nor (_05565_, _05564_, _05497_);
  and (_05566_, _05565_, _05563_);
  and (_05567_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [1]);
  and (_05568_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [3]);
  and (_05569_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [2]);
  and (_05570_, _05569_, _05568_);
  nor (_05571_, _05569_, _05568_);
  nor (_05572_, _05571_, _05570_);
  and (_05573_, _05572_, _05567_);
  nor (_05574_, _05572_, _05567_);
  nor (_05575_, _05574_, _05573_);
  nor (_05576_, _05565_, _05563_);
  nor (_05577_, _05576_, _05566_);
  and (_05578_, _05577_, _05575_);
  nor (_05579_, _05578_, _05566_);
  not (_05580_, _05579_);
  nor (_05581_, _05513_, _05511_);
  nor (_05582_, _05581_, _05514_);
  and (_05583_, _05582_, _05580_);
  nor (_05584_, _05573_, _05570_);
  and (_05585_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [1]);
  and (_05586_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [0]);
  nor (_05587_, _05586_, _05585_);
  nor (_05588_, _05587_, _05521_);
  not (_05589_, _05588_);
  nor (_05590_, _05589_, _05584_);
  and (_05591_, _05589_, _05584_);
  nor (_05592_, _05591_, _05590_);
  nor (_05593_, _05582_, _05580_);
  nor (_05594_, _05593_, _05583_);
  and (_05596_, _05594_, _05592_);
  nor (_05598_, _05596_, _05583_);
  nor (_05600_, _05533_, _05531_);
  nor (_05602_, _05600_, _05534_);
  not (_05604_, _05602_);
  nor (_05606_, _05604_, _05598_);
  and (_05608_, _05604_, _05598_);
  nor (_05610_, _05608_, _05606_);
  and (_05612_, _05610_, _05590_);
  nor (_05614_, _05612_, _05606_);
  nor (_05616_, _05543_, _05541_);
  nor (_05618_, _05616_, _05544_);
  not (_05620_, _05618_);
  nor (_05622_, _05620_, _05614_);
  and (_05624_, _05548_, _05545_);
  nor (_05626_, _05624_, _05549_);
  and (_05628_, _05626_, _05622_);
  nor (_05630_, _05551_, _05549_);
  nor (_05632_, _05630_, _05552_);
  and (_05634_, _05632_, _05628_);
  nor (_05636_, _05632_, _05628_);
  nor (_05638_, _05636_, _05634_);
  and (_05640_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [4]);
  and (_05642_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [3]);
  and (_05644_, _05642_, _05640_);
  and (_05646_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [2]);
  nor (_05648_, _05642_, _05640_);
  nor (_05650_, _05648_, _05644_);
  and (_05652_, _05650_, _05646_);
  nor (_05654_, _05652_, _05644_);
  not (_05656_, _05654_);
  nor (_05657_, _05560_, _05558_);
  nor (_05659_, _05657_, _05561_);
  and (_05660_, _05659_, _05656_);
  and (_05662_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [0]);
  and (_05663_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [2]);
  and (_05665_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [1]);
  and (_05667_, _05665_, _05663_);
  nor (_05668_, _05665_, _05663_);
  nor (_05670_, _05668_, _05667_);
  and (_05671_, _05670_, _05662_);
  nor (_05673_, _05670_, _05662_);
  nor (_05674_, _05673_, _05671_);
  nor (_05676_, _05659_, _05656_);
  nor (_05677_, _05676_, _05660_);
  and (_05679_, _05677_, _05674_);
  nor (_05680_, _05679_, _05660_);
  not (_05682_, _05680_);
  nor (_05683_, _05577_, _05575_);
  nor (_05685_, _05683_, _05578_);
  and (_05686_, _05685_, _05682_);
  not (_05688_, _05520_);
  nor (_05690_, _05671_, _05667_);
  nor (_05692_, _05690_, _05688_);
  and (_05694_, _05690_, _05688_);
  nor (_05696_, _05694_, _05692_);
  nor (_05698_, _05685_, _05682_);
  nor (_05700_, _05698_, _05686_);
  and (_05702_, _05700_, _05696_);
  nor (_05704_, _05702_, _05686_);
  not (_05706_, _05704_);
  nor (_05708_, _05594_, _05592_);
  nor (_05710_, _05708_, _05596_);
  and (_05712_, _05710_, _05706_);
  nor (_05714_, _05710_, _05706_);
  nor (_05716_, _05714_, _05712_);
  and (_05718_, _05716_, _05692_);
  nor (_05720_, _05718_, _05712_);
  nor (_05722_, _05610_, _05590_);
  nor (_05724_, _05722_, _05612_);
  not (_05726_, _05724_);
  nor (_05728_, _05726_, _05720_);
  and (_05730_, _05620_, _05614_);
  nor (_05732_, _05730_, _05622_);
  and (_05734_, _05732_, _05728_);
  nor (_05736_, _05626_, _05622_);
  nor (_05738_, _05736_, _05628_);
  nand (_05740_, _05738_, _05734_);
  or (_05742_, _05738_, _05734_);
  and (_05744_, _05742_, _05740_);
  and (_05746_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [3]);
  and (_05748_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [2]);
  and (_05750_, _05748_, _05746_);
  and (_05752_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [1]);
  nor (_05754_, _05748_, _05746_);
  nor (_05756_, _05754_, _05750_);
  and (_05758_, _05756_, _05752_);
  nor (_05760_, _05758_, _05750_);
  not (_05762_, _05760_);
  nor (_05764_, _05650_, _05646_);
  nor (_05766_, _05764_, _05652_);
  and (_05768_, _05766_, _05762_);
  and (_05770_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [0]);
  and (_05772_, _05770_, _05665_);
  and (_05774_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [1]);
  and (_05776_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [0]);
  nor (_05778_, _05776_, _05774_);
  nor (_05780_, _05778_, _05772_);
  nor (_05782_, _05766_, _05762_);
  nor (_05784_, _05782_, _05768_);
  and (_05786_, _05784_, _05780_);
  nor (_05788_, _05786_, _05768_);
  not (_05790_, _05788_);
  nor (_05792_, _05677_, _05674_);
  nor (_05794_, _05792_, _05679_);
  and (_05796_, _05794_, _05790_);
  nor (_05798_, _05794_, _05790_);
  nor (_05800_, _05798_, _05796_);
  and (_05802_, _05800_, _05772_);
  nor (_05804_, _05802_, _05796_);
  not (_05806_, _05804_);
  nor (_05808_, _05700_, _05696_);
  nor (_05810_, _05808_, _05702_);
  and (_05812_, _05810_, _05806_);
  nor (_05814_, _05716_, _05692_);
  nor (_05816_, _05814_, _05718_);
  and (_05818_, _05816_, _05812_);
  and (_05820_, _05726_, _05720_);
  nor (_05822_, _05820_, _05728_);
  and (_05824_, _05822_, _05818_);
  nor (_05826_, _05732_, _05728_);
  nor (_05828_, _05826_, _05734_);
  and (_05830_, _05828_, _05824_);
  nor (_05832_, _05828_, _05824_);
  nor (_05834_, _05832_, _05830_);
  and (_05836_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [2]);
  and (_05838_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [1]);
  and (_05840_, _05838_, _05836_);
  and (_05842_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [0]);
  nor (_05844_, _05838_, _05836_);
  nor (_05846_, _05844_, _05840_);
  and (_05848_, _05846_, _05842_);
  nor (_05850_, _05848_, _05840_);
  not (_05852_, _05850_);
  nor (_05854_, _05756_, _05752_);
  nor (_05856_, _05854_, _05758_);
  and (_05858_, _05856_, _05852_);
  nor (_05860_, _05856_, _05852_);
  nor (_05862_, _05860_, _05858_);
  and (_05864_, _05862_, _05770_);
  nor (_05866_, _05864_, _05858_);
  not (_05868_, _05866_);
  nor (_05870_, _05784_, _05780_);
  nor (_05872_, _05870_, _05786_);
  and (_05874_, _05872_, _05868_);
  nor (_05876_, _05800_, _05772_);
  nor (_05878_, _05876_, _05802_);
  and (_05880_, _05878_, _05874_);
  nor (_05882_, _05810_, _05806_);
  nor (_05884_, _05882_, _05812_);
  and (_05886_, _05884_, _05880_);
  nor (_05888_, _05816_, _05812_);
  nor (_05890_, _05888_, _05818_);
  and (_05892_, _05890_, _05886_);
  nor (_05894_, _05822_, _05818_);
  nor (_05896_, _05894_, _05824_);
  and (_05898_, _05896_, _05892_);
  and (_05900_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [0]);
  and (_05902_, _05900_, _05838_);
  nor (_05904_, _05846_, _05842_);
  nor (_05906_, _05904_, _05848_);
  and (_05908_, _05906_, _05902_);
  nor (_05910_, _05862_, _05770_);
  nor (_05912_, _05910_, _05864_);
  and (_05914_, _05912_, _05908_);
  nor (_05916_, _05872_, _05868_);
  nor (_05918_, _05916_, _05874_);
  and (_05920_, _05918_, _05914_);
  nor (_05922_, _05878_, _05874_);
  nor (_05924_, _05922_, _05880_);
  and (_05926_, _05924_, _05920_);
  nor (_05928_, _05884_, _05880_);
  nor (_05930_, _05928_, _05886_);
  and (_05932_, _05930_, _05926_);
  nor (_05934_, _05890_, _05886_);
  nor (_05936_, _05934_, _05892_);
  and (_05938_, _05936_, _05932_);
  nor (_05940_, _05896_, _05892_);
  nor (_05942_, _05940_, _05898_);
  and (_05944_, _05942_, _05938_);
  nor (_05946_, _05944_, _05898_);
  not (_05948_, _05946_);
  and (_05950_, _05948_, _05834_);
  or (_05952_, _05950_, _05830_);
  nand (_05954_, _05952_, _05744_);
  and (_05956_, _05954_, _05740_);
  not (_05958_, _05956_);
  and (_05960_, _05958_, _05638_);
  or (_05962_, _05960_, _05634_);
  or (_05964_, _05554_, _05552_);
  and (_05966_, _05964_, _05555_);
  nand (_05968_, _05966_, _05962_);
  and (_05970_, _05968_, _05555_);
  nor (_05972_, _05970_, _05490_);
  or (_05974_, _05972_, _05489_);
  nor (_05976_, _05421_, _05355_);
  and (_05978_, _05976_, _05363_);
  nor (_05980_, _05976_, _05363_);
  or (_05982_, _05980_, _05978_);
  and (_05984_, _05982_, _05974_);
  or (_05986_, _05984_, _05422_);
  or (_05988_, _05986_, _05366_);
  or (_05990_, _05988_, _05285_);
  and (_05992_, _05990_, _02408_);
  and (_05993_, _05992_, _05284_);
  not (_05994_, _05249_);
  not (_05995_, _04318_);
  nor (_05996_, _04351_, _05995_);
  or (_05997_, _05996_, _05251_);
  and (_05998_, _05997_, _01875_);
  or (_05999_, _05998_, _05994_);
  or (_06000_, _05999_, _05993_);
  and (_06001_, _06000_, _05250_);
  or (_06002_, _06001_, _02528_);
  and (_06003_, _04483_, _03683_);
  or (_06004_, _05235_, _02888_);
  or (_06005_, _06004_, _06003_);
  and (_06006_, _06005_, _02043_);
  and (_06007_, _06006_, _06002_);
  and (_06008_, _02044_, _01601_);
  nor (_06009_, _04753_, _05239_);
  or (_06010_, _06009_, _05235_);
  and (_06011_, _06010_, _01602_);
  or (_06012_, _06011_, _06008_);
  or (_06013_, _06012_, _06007_);
  not (_06014_, \oc8051_golden_model_1.B [1]);
  nor (_06015_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.B [5]);
  nor (_06016_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.B [3]);
  and (_06017_, _06016_, _06015_);
  and (_06018_, _06017_, _06014_);
  nor (_06019_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.B [7]);
  not (_06020_, \oc8051_golden_model_1.B [0]);
  and (_06021_, _06020_, \oc8051_golden_model_1.ACC [7]);
  and (_06022_, _06021_, _06019_);
  and (_06023_, _06022_, _06018_);
  and (_06024_, _06019_, _06018_);
  or (_06025_, _06024_, _04776_);
  not (_06026_, \oc8051_golden_model_1.ACC [6]);
  and (_06027_, \oc8051_golden_model_1.B [0], _06026_);
  nor (_06028_, _06027_, _04776_);
  nor (_06029_, _06028_, _06014_);
  and (_06030_, _06019_, _06017_);
  not (_06031_, _06030_);
  nor (_06032_, _06031_, _06029_);
  nor (_06033_, _06032_, _06025_);
  nor (_06034_, _06033_, _06023_);
  and (_06035_, _06032_, \oc8051_golden_model_1.B [0]);
  nor (_06036_, _06035_, _06026_);
  and (_06037_, _06036_, _06014_);
  nor (_06038_, _06036_, _06014_);
  nor (_06039_, _06038_, _06037_);
  nor (_06040_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [5]);
  nor (_06041_, _06040_, _05491_);
  nor (_06042_, _06041_, \oc8051_golden_model_1.ACC [4]);
  nor (_06043_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.ACC [4]);
  and (_06044_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.ACC [4]);
  nor (_06045_, _06044_, _06020_);
  nor (_06046_, _06045_, _06043_);
  nor (_06047_, _06046_, _06042_);
  not (_06048_, _06047_);
  and (_06049_, _06048_, _06039_);
  nor (_06050_, _06034_, \oc8051_golden_model_1.B [2]);
  nor (_06051_, _06050_, _06037_);
  not (_06052_, _06051_);
  nor (_06053_, _06052_, _06049_);
  and (_06054_, _06017_, _05233_);
  and (_06055_, \oc8051_golden_model_1.B [2], _04776_);
  not (_06056_, _06055_);
  and (_06057_, _06056_, _06054_);
  not (_06058_, _06057_);
  nor (_06059_, _06058_, _06053_);
  nor (_06060_, _06059_, _06034_);
  nor (_06061_, _06060_, _06023_);
  nor (_06062_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.B [4]);
  nor (_06063_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.B [7]);
  and (_06064_, _06063_, \oc8051_golden_model_1.ACC [7]);
  and (_06065_, _06064_, _06062_);
  nor (_06066_, _06065_, _06054_);
  nor (_06067_, _06061_, \oc8051_golden_model_1.B [3]);
  not (_06068_, \oc8051_golden_model_1.B [2]);
  nor (_06069_, _06048_, _06039_);
  nor (_06070_, _06069_, _06049_);
  not (_06071_, _06070_);
  and (_06072_, _06071_, _06059_);
  nor (_06073_, _06059_, _06036_);
  nor (_06074_, _06073_, _06072_);
  and (_06075_, _06074_, _06068_);
  nor (_06076_, _06074_, _06068_);
  nor (_06077_, _06076_, _06075_);
  not (_06078_, _06077_);
  not (_06079_, \oc8051_golden_model_1.ACC [5]);
  nor (_06080_, _06059_, _06079_);
  and (_06081_, _06059_, _06041_);
  or (_06082_, _06081_, _06080_);
  and (_06083_, _06082_, _06014_);
  nor (_06084_, _06082_, _06014_);
  not (_06085_, \oc8051_golden_model_1.ACC [4]);
  and (_06086_, \oc8051_golden_model_1.B [0], _06085_);
  nor (_06087_, _06086_, _06084_);
  nor (_06088_, _06087_, _06083_);
  nor (_06089_, _06088_, _06078_);
  or (_06090_, _06089_, _06075_);
  nor (_06091_, _06090_, _06067_);
  nor (_06092_, _06091_, _06066_);
  nor (_06093_, _06092_, _06061_);
  nor (_06094_, _06093_, _06023_);
  nor (_06095_, _06094_, \oc8051_golden_model_1.B [4]);
  not (_06096_, \oc8051_golden_model_1.B [3]);
  not (_06097_, _06092_);
  and (_06098_, _06088_, _06078_);
  nor (_06099_, _06098_, _06089_);
  nor (_06100_, _06099_, _06097_);
  nor (_06101_, _06092_, _06074_);
  nor (_06102_, _06101_, _06100_);
  and (_06103_, _06102_, _06096_);
  nor (_06104_, _06102_, _06096_);
  nor (_06105_, _06104_, _06103_);
  not (_06106_, _06105_);
  nor (_06107_, _06092_, _06082_);
  nor (_06108_, _06084_, _06083_);
  and (_06109_, _06108_, _06086_);
  nor (_06110_, _06108_, _06086_);
  nor (_06111_, _06110_, _06109_);
  and (_06112_, _06111_, _06092_);
  or (_06113_, _06112_, _06107_);
  nor (_06114_, _06113_, \oc8051_golden_model_1.B [2]);
  and (_06115_, _06113_, \oc8051_golden_model_1.B [2]);
  nor (_06116_, _06092_, _06085_);
  nor (_06117_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [4]);
  nor (_06118_, _06117_, _05640_);
  and (_06119_, _06092_, _06118_);
  or (_06120_, _06119_, _06116_);
  and (_06121_, _06120_, _06014_);
  nor (_06122_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [3]);
  nor (_06123_, _06122_, _05746_);
  nor (_06124_, _06123_, \oc8051_golden_model_1.ACC [2]);
  nor (_06125_, \oc8051_golden_model_1.ACC [3], \oc8051_golden_model_1.ACC [2]);
  and (_06126_, \oc8051_golden_model_1.ACC [3], \oc8051_golden_model_1.ACC [2]);
  nor (_06127_, _06126_, _06020_);
  nor (_06128_, _06127_, _06125_);
  nor (_06129_, _06128_, _06124_);
  not (_06130_, _06129_);
  nor (_06131_, _06120_, _06014_);
  nor (_06132_, _06131_, _06121_);
  and (_06133_, _06132_, _06130_);
  nor (_06134_, _06133_, _06121_);
  nor (_06135_, _06134_, _06115_);
  nor (_06136_, _06135_, _06114_);
  nor (_06137_, _06136_, _06106_);
  or (_06138_, _06137_, _06103_);
  nor (_06139_, _06138_, _06095_);
  not (_06140_, \oc8051_golden_model_1.B [5]);
  and (_06141_, _06063_, _06140_);
  not (_06142_, _06141_);
  and (_06143_, \oc8051_golden_model_1.B [4], _04776_);
  nor (_06144_, _06143_, _06142_);
  not (_06145_, _06144_);
  nor (_06146_, _06145_, _06139_);
  nor (_06147_, _06146_, _06094_);
  nor (_06148_, _06147_, _06023_);
  nor (_06149_, _06064_, _06141_);
  nor (_06150_, _06148_, \oc8051_golden_model_1.B [5]);
  not (_06151_, \oc8051_golden_model_1.B [4]);
  and (_06152_, _06136_, _06106_);
  nor (_06153_, _06152_, _06137_);
  not (_06154_, _06153_);
  and (_06155_, _06154_, _06146_);
  nor (_06156_, _06146_, _06102_);
  nor (_06157_, _06156_, _06155_);
  and (_06158_, _06157_, _06151_);
  nor (_06159_, _06157_, _06151_);
  nor (_06160_, _06159_, _06158_);
  not (_06161_, _06160_);
  nor (_06162_, _06146_, _06113_);
  nor (_06163_, _06115_, _06114_);
  and (_06164_, _06163_, _06134_);
  nor (_06165_, _06163_, _06134_);
  nor (_06166_, _06165_, _06164_);
  not (_06167_, _06166_);
  and (_06168_, _06167_, _06146_);
  nor (_06169_, _06168_, _06162_);
  nor (_06170_, _06169_, \oc8051_golden_model_1.B [3]);
  and (_06171_, _06169_, \oc8051_golden_model_1.B [3]);
  nor (_06172_, _06132_, _06130_);
  nor (_06173_, _06172_, _06133_);
  not (_06174_, _06173_);
  and (_06175_, _06174_, _06146_);
  nor (_06176_, _06146_, _06120_);
  nor (_06177_, _06176_, _06175_);
  and (_06178_, _06177_, _06068_);
  nor (_06179_, _06146_, _01689_);
  and (_06180_, _06146_, _06123_);
  or (_06181_, _06180_, _06179_);
  and (_06182_, _06181_, _06014_);
  nor (_06183_, _06181_, _06014_);
  not (_06184_, \oc8051_golden_model_1.ACC [2]);
  and (_06185_, \oc8051_golden_model_1.B [0], _06184_);
  nor (_06186_, _06185_, _06183_);
  nor (_06187_, _06186_, _06182_);
  nor (_06188_, _06177_, _06068_);
  nor (_06189_, _06188_, _06178_);
  not (_06190_, _06189_);
  nor (_06191_, _06190_, _06187_);
  nor (_06192_, _06191_, _06178_);
  nor (_06193_, _06192_, _06171_);
  nor (_06194_, _06193_, _06170_);
  nor (_06195_, _06194_, _06161_);
  or (_06196_, _06195_, _06158_);
  nor (_06197_, _06196_, _06150_);
  nor (_06198_, _06197_, _06149_);
  nor (_06199_, _06198_, _06148_);
  not (_06200_, _06198_);
  and (_06201_, _06194_, _06161_);
  nor (_06202_, _06201_, _06195_);
  nor (_06203_, _06202_, _06200_);
  nor (_06204_, _06198_, _06157_);
  nor (_06205_, _06204_, _06203_);
  and (_06206_, _06205_, _06140_);
  nor (_06207_, _06205_, _06140_);
  nor (_06208_, _06207_, _06206_);
  not (_06209_, _06208_);
  nor (_06210_, _06198_, _06169_);
  nor (_06211_, _06171_, _06170_);
  nor (_06212_, _06211_, _06192_);
  and (_06213_, _06211_, _06192_);
  or (_06214_, _06213_, _06212_);
  and (_06215_, _06214_, _06198_);
  or (_06216_, _06215_, _06210_);
  and (_06217_, _06216_, _06151_);
  nor (_06218_, _06216_, _06151_);
  and (_06219_, _06190_, _06187_);
  nor (_06220_, _06219_, _06191_);
  nor (_06221_, _06220_, _06200_);
  nor (_06222_, _06198_, _06177_);
  nor (_06223_, _06222_, _06221_);
  and (_06224_, _06223_, _06096_);
  nor (_06225_, _06183_, _06182_);
  nor (_06226_, _06225_, _06185_);
  and (_06227_, _06225_, _06185_);
  or (_06228_, _06227_, _06226_);
  nor (_06229_, _06228_, _06200_);
  nor (_06230_, _06198_, _06181_);
  nor (_06231_, _06230_, _06229_);
  and (_06232_, _06231_, _06068_);
  nor (_06233_, _06231_, _06068_);
  nor (_06234_, _06198_, _06184_);
  nor (_06235_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [2]);
  nor (_06236_, _06235_, _05836_);
  and (_06237_, _06198_, _06236_);
  or (_06238_, _06237_, _06234_);
  and (_06239_, _06238_, _06014_);
  and (_06240_, \oc8051_golden_model_1.B [0], _01613_);
  not (_06241_, _06240_);
  nor (_06242_, _06238_, _06014_);
  nor (_06243_, _06242_, _06239_);
  and (_06244_, _06243_, _06241_);
  nor (_06245_, _06244_, _06239_);
  nor (_06246_, _06245_, _06233_);
  nor (_06247_, _06246_, _06232_);
  nor (_06248_, _06223_, _06096_);
  nor (_06249_, _06248_, _06224_);
  not (_06250_, _06249_);
  nor (_06251_, _06250_, _06247_);
  nor (_06252_, _06251_, _06224_);
  nor (_06253_, _06252_, _06218_);
  nor (_06254_, _06253_, _06217_);
  nor (_06255_, _06254_, _06209_);
  nor (_06256_, _06255_, _06206_);
  and (_06257_, _05233_, \oc8051_golden_model_1.ACC [7]);
  nor (_06258_, _06257_, _06063_);
  nor (_06259_, _06258_, _06256_);
  not (_06260_, _06063_);
  nor (_06261_, _06199_, _06023_);
  nor (_06262_, _06261_, _06260_);
  nor (_06263_, _06262_, _06259_);
  and (_06264_, _06263_, _06199_);
  nor (_06265_, _06264_, _06023_);
  and (_06266_, _06265_, \oc8051_golden_model_1.B [7]);
  and (_06267_, _06265_, _05233_);
  nor (_06268_, _06267_, _05356_);
  not (_06269_, _06268_);
  not (_06270_, \oc8051_golden_model_1.B [6]);
  and (_06271_, _06254_, _06209_);
  nor (_06272_, _06271_, _06255_);
  nor (_06273_, _06272_, _06263_);
  not (_06274_, _06263_);
  nor (_06275_, _06274_, _06205_);
  nor (_06276_, _06275_, _06273_);
  nor (_06277_, _06276_, _06270_);
  and (_06278_, _06276_, _06270_);
  nor (_06279_, _06218_, _06217_);
  nor (_06280_, _06279_, _06252_);
  and (_06281_, _06279_, _06252_);
  or (_06282_, _06281_, _06280_);
  nor (_06283_, _06282_, _06263_);
  nor (_06284_, _06274_, _06216_);
  nor (_06285_, _06284_, _06283_);
  nor (_06286_, _06285_, _06140_);
  and (_06287_, _06285_, _06140_);
  not (_06288_, _06287_);
  and (_06289_, _06250_, _06247_);
  nor (_06290_, _06289_, _06251_);
  nor (_06291_, _06290_, _06263_);
  nor (_06292_, _06274_, _06223_);
  nor (_06293_, _06292_, _06291_);
  nor (_06294_, _06293_, _06151_);
  and (_06295_, _06263_, _06231_);
  nor (_06296_, _06233_, _06232_);
  and (_06297_, _06296_, _06245_);
  nor (_06298_, _06296_, _06245_);
  nor (_06299_, _06298_, _06297_);
  nor (_06300_, _06299_, _06263_);
  or (_06301_, _06300_, _06295_);
  nor (_06302_, _06301_, _06096_);
  and (_06303_, _06301_, _06096_);
  nor (_06304_, _06303_, _06302_);
  nor (_06305_, _06243_, _06241_);
  or (_06306_, _06305_, _06244_);
  nor (_06307_, _06306_, _06263_);
  and (_06308_, _06263_, _06238_);
  nor (_06309_, _06308_, _06307_);
  and (_06310_, _06309_, \oc8051_golden_model_1.B [2]);
  nor (_06311_, _06309_, \oc8051_golden_model_1.B [2]);
  nor (_06312_, _06311_, _06310_);
  and (_06313_, _06312_, _06304_);
  and (_06314_, _06263_, _01613_);
  and (_06315_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [1]);
  nor (_06316_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [1]);
  nor (_06317_, _06316_, _06315_);
  nor (_06318_, _06263_, _06317_);
  nor (_06319_, _06318_, _06314_);
  and (_06320_, _06319_, _06014_);
  nor (_06321_, _06319_, _06014_);
  and (_06322_, _06020_, \oc8051_golden_model_1.ACC [0]);
  not (_06323_, _06322_);
  nor (_06324_, _06323_, _06321_);
  nor (_06325_, _06324_, _06320_);
  and (_06326_, _06325_, _06313_);
  not (_06327_, _06326_);
  and (_06328_, _06310_, _06304_);
  nor (_06329_, _06328_, _06302_);
  and (_06330_, _06329_, _06327_);
  and (_06331_, _06293_, _06151_);
  nor (_06332_, _06331_, _06330_);
  or (_06333_, _06332_, _06294_);
  and (_06334_, _06333_, _06288_);
  nor (_06335_, _06334_, _06286_);
  nor (_06336_, _06335_, _06278_);
  or (_06337_, _06336_, _06277_);
  and (_06338_, _06337_, _06269_);
  nor (_06339_, _06338_, _06266_);
  nor (_06340_, _06331_, _06294_);
  nor (_06341_, _06287_, _06286_);
  and (_06342_, _06341_, _06340_);
  nor (_06343_, _06278_, _06277_);
  and (_06344_, _06343_, _06269_);
  and (_06345_, _06344_, _06342_);
  nor (_06346_, _06321_, _06320_);
  and (_06347_, \oc8051_golden_model_1.B [0], _01710_);
  not (_06348_, _06347_);
  and (_06349_, _06348_, _06346_);
  and (_06350_, _06349_, _06323_);
  and (_06351_, _06350_, _06313_);
  and (_06352_, _06351_, _06345_);
  nor (_06353_, _06352_, _06339_);
  and (_06354_, _06353_, _06264_);
  not (_06355_, _06008_);
  or (_06356_, _06023_, _06355_);
  or (_06357_, _06356_, _06354_);
  and (_06358_, _06357_, _01870_);
  and (_06359_, _06358_, _06013_);
  and (_06360_, _04560_, _03683_);
  or (_06361_, _06360_, _05235_);
  and (_06362_, _06361_, _01869_);
  or (_06363_, _06362_, _02079_);
  or (_06364_, _06363_, _06359_);
  and (_06365_, _04771_, _03683_);
  or (_06366_, _05235_, _02166_);
  or (_06367_, _06366_, _06365_);
  and (_06368_, _06367_, _02912_);
  and (_06369_, _06368_, _06364_);
  or (_06370_, _06369_, _05238_);
  and (_06371_, _06370_, _02176_);
  or (_06372_, _05235_, _03755_);
  and (_06373_, _06361_, _02072_);
  and (_06374_, _06373_, _06372_);
  or (_06375_, _06374_, _06371_);
  and (_06376_, _06375_, _02907_);
  and (_06377_, _05259_, _02177_);
  and (_06378_, _06377_, _06372_);
  or (_06379_, _06378_, _02071_);
  or (_06380_, _06379_, _06376_);
  nor (_06381_, _04770_, _05239_);
  or (_06382_, _05235_, _04788_);
  or (_06383_, _06382_, _06381_);
  and (_06384_, _06383_, _04793_);
  and (_06385_, _06384_, _06380_);
  nor (_06386_, _04778_, _05239_);
  or (_06387_, _06386_, _05235_);
  and (_06389_, _06387_, _02173_);
  or (_06390_, _06389_, _02201_);
  or (_06391_, _06390_, _06385_);
  or (_06392_, _05256_, _02303_);
  and (_06393_, _06392_, _01887_);
  and (_06394_, _06393_, _06391_);
  and (_06395_, _05253_, _01860_);
  or (_06396_, _06395_, _01537_);
  or (_06397_, _06396_, _06394_);
  and (_06398_, _04264_, _03683_);
  or (_06400_, _05235_, _01538_);
  or (_06401_, _06400_, _06398_);
  and (_06402_, _06401_, _38087_);
  and (_06403_, _06402_, _06397_);
  or (_06404_, _06403_, _05234_);
  and (_37137_, _06404_, _37580_);
  nor (_06405_, _38087_, _04776_);
  and (_06406_, _03616_, _04776_);
  nor (_06407_, _03616_, _04776_);
  nor (_06408_, _06407_, _06406_);
  nor (_06410_, _03808_, _06026_);
  and (_06411_, _03808_, _06026_);
  nor (_06412_, _06411_, _06410_);
  nor (_06413_, _03916_, _06079_);
  and (_06414_, _03916_, _06079_);
  nor (_06415_, _06414_, _06413_);
  not (_06416_, _06415_);
  nor (_06417_, _04211_, _06085_);
  and (_06418_, _04211_, _06085_);
  nor (_06419_, _06418_, _06417_);
  and (_06421_, _03268_, _01689_);
  not (_06422_, _06421_);
  nor (_06423_, _03268_, _01689_);
  not (_06424_, _06423_);
  nor (_06425_, _03455_, _06184_);
  and (_06426_, _03455_, _06184_);
  nor (_06427_, _06426_, _06425_);
  not (_06428_, _06427_);
  nor (_06429_, _02811_, _01613_);
  and (_06430_, _02811_, _01613_);
  nor (_06432_, _06430_, _06429_);
  and (_06433_, _03028_, \oc8051_golden_model_1.ACC [0]);
  and (_06434_, _06433_, _06432_);
  nor (_06435_, _06434_, _06429_);
  nor (_06436_, _06435_, _06428_);
  nor (_06437_, _06436_, _06425_);
  nand (_06438_, _06437_, _06424_);
  and (_06439_, _06438_, _06422_);
  and (_06440_, _06439_, _06419_);
  nor (_06441_, _06440_, _06417_);
  nor (_06443_, _06441_, _06416_);
  or (_06444_, _06443_, _06413_);
  and (_06445_, _06444_, _06412_);
  nor (_06446_, _06445_, _06410_);
  nor (_06447_, _06446_, _06408_);
  and (_06448_, _06446_, _06408_);
  nor (_06449_, _06448_, _06447_);
  and (_06450_, _01972_, _01652_);
  not (_06451_, _06450_);
  nor (_06452_, _02690_, _01977_);
  nor (_06453_, _06452_, _02612_);
  and (_06454_, _01971_, _01467_);
  and (_06455_, _06454_, _01652_);
  or (_06456_, _06455_, _02693_);
  nor (_06457_, _06456_, _06453_);
  and (_06458_, _06457_, _06451_);
  not (_06459_, _06458_);
  nand (_06460_, _06459_, _06449_);
  nor (_06461_, _04483_, \oc8051_golden_model_1.ACC [7]);
  and (_06462_, _01882_, _01647_);
  nand (_06463_, _06462_, _06461_);
  nor (_06464_, _03680_, _04776_);
  and (_06465_, _04560_, _03680_);
  nor (_06466_, _06465_, _06464_);
  or (_06467_, _06466_, _04778_);
  nor (_06468_, _06467_, _02176_);
  and (_06469_, _04771_, _03680_);
  nor (_06470_, _06469_, _06464_);
  nand (_06471_, _06470_, _02079_);
  not (_06472_, _03680_);
  nor (_06473_, _06472_, _03616_);
  nor (_06474_, _06473_, _06464_);
  nand (_06475_, _06474_, _05994_);
  and (_06476_, _02044_, _01548_);
  and (_06477_, _03658_, \oc8051_golden_model_1.PSW [7]);
  and (_06478_, _06477_, _03689_);
  and (_06479_, _06478_, _03638_);
  and (_06480_, _06479_, _03379_);
  nor (_06481_, _06480_, _03673_);
  and (_06482_, _06479_, _01923_);
  or (_06483_, _06482_, _06481_);
  nor (_06484_, _06483_, _04776_);
  and (_06485_, _06483_, _04776_);
  nor (_06486_, _06485_, _06484_);
  not (_06487_, _06486_);
  nor (_06488_, _06479_, _03379_);
  nor (_06489_, _06488_, _06480_);
  nor (_06490_, _06489_, _06026_);
  and (_06491_, _06489_, _06026_);
  and (_06492_, _06478_, _03622_);
  nor (_06493_, _06492_, _03630_);
  nor (_06494_, _06493_, _06479_);
  and (_06495_, _06494_, _06079_);
  nor (_06496_, _06494_, _06079_);
  nor (_06497_, _06478_, _03622_);
  nor (_06498_, _06497_, _06492_);
  nor (_06499_, _06498_, _06085_);
  nor (_06500_, _06499_, _06496_);
  nor (_06501_, _06500_, _06495_);
  nor (_06502_, _06496_, _06495_);
  not (_06503_, _06502_);
  and (_06504_, _06498_, _06085_);
  or (_06505_, _06504_, _06499_);
  or (_06506_, _06505_, _06503_);
  nor (_06507_, _04350_, _01955_);
  nor (_06508_, _06507_, _06478_);
  nor (_06509_, _06508_, _01689_);
  and (_06510_, _06508_, _01689_);
  nor (_06511_, _06510_, _06509_);
  nor (_06512_, _06477_, _03391_);
  nor (_06513_, _06512_, _04350_);
  nor (_06514_, _06513_, _06184_);
  and (_06515_, _06513_, _06184_);
  nor (_06516_, _06515_, _06514_);
  and (_06517_, _06516_, _06511_);
  not (_06518_, \oc8051_golden_model_1.PSW [7]);
  nor (_06519_, _02441_, _06518_);
  nor (_06520_, _06519_, _01823_);
  nor (_06521_, _06520_, _06477_);
  and (_06522_, _06521_, _01613_);
  nor (_06523_, _06521_, _01613_);
  nor (_06524_, _02441_, \oc8051_golden_model_1.PSW [7]);
  and (_06525_, _02441_, \oc8051_golden_model_1.PSW [7]);
  nor (_06526_, _06525_, _06524_);
  or (_06527_, _06526_, \oc8051_golden_model_1.ACC [0]);
  nor (_06528_, _06527_, _06523_);
  nor (_06529_, _06528_, _06522_);
  nand (_06530_, _06529_, _06517_);
  and (_06531_, _06514_, _06511_);
  nor (_06532_, _06531_, _06509_);
  and (_06533_, _06532_, _06530_);
  nor (_06534_, _06533_, _06506_);
  nor (_06535_, _06534_, _06501_);
  nor (_06536_, _06535_, _06491_);
  or (_06537_, _06536_, _06490_);
  and (_06538_, _06537_, _06487_);
  nor (_06539_, _06537_, _06487_);
  nor (_06540_, _06539_, _06538_);
  nand (_06541_, _06540_, _06476_);
  and (_06542_, _05184_, \oc8051_golden_model_1.PSW [7]);
  and (_06543_, _06542_, _04816_);
  nor (_06544_, _06542_, _04816_);
  or (_06545_, _06544_, _06543_);
  nor (_06546_, _06545_, _04776_);
  and (_06547_, _06545_, _04776_);
  nor (_06548_, _06547_, _06546_);
  not (_06549_, _06548_);
  and (_06550_, _05183_, \oc8051_golden_model_1.PSW [7]);
  nor (_06551_, _06550_, _04861_);
  nor (_06552_, _06551_, _06542_);
  nor (_06553_, _06552_, _06026_);
  and (_06554_, _05181_, _05135_);
  and (_06555_, _06554_, \oc8051_golden_model_1.PSW [7]);
  nor (_06556_, _06555_, _05090_);
  nor (_06557_, _06556_, _06550_);
  and (_06558_, _06557_, _06079_);
  nor (_06559_, _06557_, _06079_);
  and (_06560_, _05179_, \oc8051_golden_model_1.PSW [7]);
  and (_06561_, _06560_, _05180_);
  nor (_06562_, _06561_, _05135_);
  nor (_06563_, _06562_, _06555_);
  nor (_06564_, _06563_, _06085_);
  nor (_06565_, _06564_, _06559_);
  nor (_06566_, _06565_, _06558_);
  nor (_06567_, _06559_, _06558_);
  not (_06568_, _06567_);
  and (_06569_, _06563_, _06085_);
  or (_06570_, _06569_, _06564_);
  or (_06571_, _06570_, _06568_);
  and (_06572_, _05179_, _05043_);
  and (_06573_, _06572_, \oc8051_golden_model_1.PSW [7]);
  nor (_06574_, _06573_, _04998_);
  nor (_06575_, _06574_, _06561_);
  nor (_06576_, _06575_, _01689_);
  and (_06577_, _06575_, _01689_);
  nor (_06578_, _06577_, _06576_);
  nor (_06579_, _06560_, _05043_);
  nor (_06580_, _06579_, _06573_);
  nor (_06581_, _06580_, _06184_);
  and (_06582_, _06580_, _06184_);
  nor (_06583_, _06582_, _06581_);
  and (_06584_, _06583_, _06578_);
  and (_06585_, _04952_, \oc8051_golden_model_1.PSW [7]);
  nor (_06586_, _06585_, _04907_);
  nor (_06587_, _06586_, _06560_);
  nor (_06588_, _06587_, _01613_);
  and (_06589_, _06587_, _01613_);
  nor (_06590_, _04952_, \oc8051_golden_model_1.PSW [7]);
  nor (_06591_, _06590_, _06585_);
  and (_06592_, _06591_, _01710_);
  nor (_06593_, _06592_, _06589_);
  or (_06594_, _06593_, _06588_);
  nand (_06595_, _06594_, _06584_);
  and (_06596_, _06581_, _06578_);
  nor (_06597_, _06596_, _06576_);
  and (_06598_, _06597_, _06595_);
  nor (_06599_, _06598_, _06571_);
  nor (_06600_, _06599_, _06566_);
  and (_06601_, _06552_, _06026_);
  nor (_06602_, _06553_, _06601_);
  not (_06603_, _06602_);
  nor (_06604_, _06603_, _06600_);
  or (_06605_, _06604_, _06553_);
  and (_06606_, _06605_, _06549_);
  nor (_06607_, _06605_, _06549_);
  nor (_06608_, _06607_, _06606_);
  and (_06609_, _01882_, _01548_);
  nand (_06610_, _06609_, _06608_);
  nor (_06611_, _02482_, _02367_);
  nor (_06612_, _03123_, _02394_);
  and (_06613_, _06612_, _06611_);
  not (_06614_, _06613_);
  nand (_06615_, _06614_, _03616_);
  and (_06616_, _02044_, _02002_);
  nor (_06617_, _06616_, _02001_);
  not (_06618_, _02003_);
  nor (_06619_, _04528_, _06618_);
  and (_06620_, _01882_, _02002_);
  not (_06621_, _06620_);
  or (_06622_, _04483_, _06621_);
  nor (_06623_, _01567_, _01534_);
  nand (_06624_, _06623_, _03616_);
  and (_06625_, _02044_, _01884_);
  or (_06626_, _06625_, \oc8051_golden_model_1.ACC [7]);
  nand (_06627_, _06625_, \oc8051_golden_model_1.ACC [7]);
  and (_06628_, _06627_, _06626_);
  or (_06629_, _06623_, _06620_);
  or (_06630_, _06629_, _06628_);
  and (_06631_, _06630_, _06624_);
  and (_06632_, _06631_, _06618_);
  and (_06633_, _06632_, _06622_);
  or (_06634_, _06633_, _06619_);
  and (_06635_, _06634_, _06617_);
  and (_06636_, _02044_, _01881_);
  and (_06637_, _04496_, _03680_);
  nor (_06638_, _06637_, _06464_);
  nor (_06639_, _06638_, _02814_);
  or (_06640_, _06639_, _06636_);
  or (_06641_, _06640_, _06635_);
  not (_06642_, _06636_);
  nor (_06643_, \oc8051_golden_model_1.ACC [2], \oc8051_golden_model_1.ACC [1]);
  nor (_06644_, _06643_, _01689_);
  and (_06645_, _06644_, _06044_);
  and (_06646_, _06645_, \oc8051_golden_model_1.ACC [6]);
  and (_06647_, _06646_, \oc8051_golden_model_1.ACC [7]);
  nor (_06648_, _06646_, \oc8051_golden_model_1.ACC [7]);
  nor (_06649_, _06648_, _06647_);
  and (_06650_, _06644_, \oc8051_golden_model_1.ACC [4]);
  nor (_06651_, _06650_, \oc8051_golden_model_1.ACC [5]);
  nor (_06652_, _06651_, _06645_);
  nor (_06653_, _06645_, \oc8051_golden_model_1.ACC [6]);
  nor (_06654_, _06653_, _06646_);
  nor (_06655_, _06654_, _06652_);
  not (_06656_, _06655_);
  and (_06657_, _06656_, _06649_);
  nor (_06658_, \oc8051_golden_model_1.PSW [7], \oc8051_golden_model_1.ACC [7]);
  nor (_06659_, _06658_, _06655_);
  nor (_06660_, _06659_, _06649_);
  nor (_06661_, _06660_, _06657_);
  or (_06662_, _06661_, _06642_);
  and (_06663_, _06662_, _02008_);
  and (_06664_, _06663_, _06641_);
  nor (_06665_, _04326_, _04776_);
  and (_06666_, _04368_, _04326_);
  nor (_06667_, _06666_, _06665_);
  nor (_06668_, _06667_, _02024_);
  nor (_06669_, _06474_, _02840_);
  or (_06670_, _06669_, _06614_);
  or (_06671_, _06670_, _06668_);
  or (_06672_, _06671_, _06664_);
  and (_06673_, _06672_, _06615_);
  or (_06674_, _06673_, _02850_);
  not (_06675_, _02850_);
  or (_06676_, _04483_, _06675_);
  and (_06677_, _06676_, _02021_);
  and (_06678_, _06677_, _06674_);
  and (_06679_, _02044_, _01877_);
  nor (_06680_, _04528_, _02021_);
  or (_06681_, _06680_, _06679_);
  or (_06682_, _06681_, _06678_);
  nand (_06683_, _06679_, _01689_);
  and (_06684_, _06683_, _06682_);
  or (_06685_, _06684_, _01997_);
  and (_06686_, _04364_, _04326_);
  nor (_06687_, _06686_, _06665_);
  nand (_06688_, _06687_, _01997_);
  and (_06689_, _06688_, _02861_);
  and (_06690_, _06689_, _06685_);
  and (_06691_, _06666_, _04533_);
  nor (_06692_, _06691_, _06665_);
  nor (_06693_, _06692_, _02861_);
  or (_06694_, _06693_, _05279_);
  or (_06695_, _06694_, _06690_);
  nor (_06696_, _05936_, _05932_);
  nor (_06697_, _06696_, _05938_);
  or (_06698_, _06697_, _05285_);
  and (_06699_, _01548_, _01533_);
  not (_06700_, _06699_);
  and (_06701_, _06700_, _06698_);
  and (_06702_, _06701_, _06695_);
  and (_06703_, _05165_, \oc8051_golden_model_1.PSW [7]);
  and (_06704_, _06703_, _05158_);
  nor (_06705_, _06704_, _03616_);
  and (_06706_, _06704_, _03616_);
  nor (_06707_, _06706_, _06705_);
  and (_06708_, _06707_, \oc8051_golden_model_1.ACC [7]);
  nor (_06709_, _06707_, \oc8051_golden_model_1.ACC [7]);
  nor (_06710_, _06709_, _06708_);
  not (_06711_, _06710_);
  nor (_06712_, _06703_, _05158_);
  nor (_06713_, _06712_, _06704_);
  nor (_06714_, _06713_, _06026_);
  and (_06715_, _05164_, \oc8051_golden_model_1.PSW [7]);
  nor (_06716_, _06715_, _05159_);
  nor (_06717_, _06716_, _06703_);
  and (_06718_, _06717_, _06079_);
  nor (_06719_, _06717_, _06079_);
  and (_06720_, _05161_, \oc8051_golden_model_1.PSW [7]);
  and (_06721_, _06720_, _05162_);
  nor (_06722_, _06721_, _05160_);
  nor (_06723_, _06722_, _06715_);
  nor (_06724_, _06723_, _06085_);
  nor (_06725_, _06724_, _06719_);
  nor (_06726_, _06725_, _06718_);
  nor (_06727_, _06719_, _06718_);
  not (_06728_, _06727_);
  and (_06729_, _06723_, _06085_);
  or (_06730_, _06729_, _06724_);
  or (_06731_, _06730_, _06728_);
  not (_06732_, _03268_);
  and (_06733_, _05161_, _03456_);
  and (_06734_, _06733_, \oc8051_golden_model_1.PSW [7]);
  nor (_06735_, _06734_, _06732_);
  nor (_06736_, _06735_, _06721_);
  nor (_06737_, _06736_, _01689_);
  and (_06738_, _06736_, _01689_);
  nor (_06739_, _06738_, _06737_);
  nor (_06740_, _06720_, _03456_);
  nor (_06741_, _06740_, _06734_);
  nor (_06742_, _06741_, _06184_);
  and (_06743_, _06741_, _06184_);
  nor (_06744_, _06743_, _06742_);
  and (_06745_, _06744_, _06739_);
  and (_06746_, _03028_, \oc8051_golden_model_1.PSW [7]);
  nor (_06747_, _06746_, _02812_);
  nor (_06748_, _06747_, _06720_);
  nor (_06749_, _06748_, _01613_);
  and (_06750_, _06748_, _01613_);
  and (_06751_, _03042_, _06518_);
  nor (_06752_, _06751_, _06746_);
  and (_06753_, _06752_, _01710_);
  nor (_06754_, _06753_, _06750_);
  or (_06755_, _06754_, _06749_);
  nand (_06756_, _06755_, _06745_);
  and (_06757_, _06742_, _06739_);
  nor (_06758_, _06757_, _06737_);
  and (_06759_, _06758_, _06756_);
  nor (_06760_, _06759_, _06731_);
  nor (_06761_, _06760_, _06726_);
  and (_06762_, _06713_, _06026_);
  nor (_06763_, _06714_, _06762_);
  not (_06764_, _06763_);
  nor (_06765_, _06764_, _06761_);
  or (_06766_, _06765_, _06714_);
  and (_06767_, _06766_, _06711_);
  nor (_06768_, _06766_, _06711_);
  nor (_06769_, _06768_, _06767_);
  nor (_06770_, _06769_, _06700_);
  or (_06771_, _06770_, _06609_);
  or (_06772_, _06771_, _06702_);
  and (_06773_, _06772_, _02036_);
  and (_06774_, _06773_, _06610_);
  nor (_06775_, _06476_, _01963_);
  not (_06776_, _06775_);
  not (_06777_, _06476_);
  and (_06778_, _03698_, \oc8051_golden_model_1.P1INREG [6]);
  not (_06779_, _06778_);
  and (_06780_, _03665_, \oc8051_golden_model_1.P2INREG [6]);
  and (_06781_, _03646_, \oc8051_golden_model_1.P3INREG [6]);
  nor (_06782_, _06781_, _06780_);
  and (_06783_, _06782_, _03817_);
  and (_06784_, _06783_, _06779_);
  and (_06785_, _03832_, \oc8051_golden_model_1.P0INREG [6]);
  not (_06786_, _06785_);
  and (_06787_, _06786_, _03831_);
  and (_06788_, _06787_, _06784_);
  and (_06789_, _06788_, _03815_);
  and (_06790_, _06789_, _03860_);
  and (_06791_, _06790_, _03809_);
  not (_06792_, _06791_);
  nand (_06793_, _03832_, \oc8051_golden_model_1.P0INREG [3]);
  and (_06794_, _03698_, \oc8051_golden_model_1.P1INREG [3]);
  not (_06795_, _06794_);
  and (_06796_, _03665_, \oc8051_golden_model_1.P2INREG [3]);
  and (_06797_, _03646_, \oc8051_golden_model_1.P3INREG [3]);
  nor (_06798_, _06797_, _06796_);
  and (_06799_, _06798_, _06795_);
  and (_06800_, _06799_, _03973_);
  and (_06801_, _06800_, _06793_);
  and (_06802_, _06801_, _03993_);
  and (_06803_, _06802_, _04011_);
  and (_06804_, _06803_, _03966_);
  not (_06805_, _06804_);
  and (_06806_, _03665_, \oc8051_golden_model_1.P2INREG [2]);
  and (_06807_, _03646_, \oc8051_golden_model_1.P3INREG [2]);
  nor (_06808_, _06807_, _06806_);
  and (_06809_, _03698_, \oc8051_golden_model_1.P1INREG [2]);
  and (_06810_, _03737_, \oc8051_golden_model_1.P0INREG [2]);
  nor (_06811_, _06810_, _06809_);
  and (_06812_, _06811_, _06808_);
  and (_06813_, _06812_, _04144_);
  and (_06814_, _06813_, _04135_);
  and (_06815_, _06814_, _04129_);
  and (_06816_, _06815_, _04108_);
  not (_06817_, _06816_);
  and (_06818_, _03665_, \oc8051_golden_model_1.P2INREG [1]);
  and (_06819_, _03646_, \oc8051_golden_model_1.P3INREG [1]);
  nor (_06820_, _06819_, _06818_);
  and (_06821_, _03698_, \oc8051_golden_model_1.P1INREG [1]);
  and (_06822_, _03737_, \oc8051_golden_model_1.P0INREG [1]);
  nor (_06823_, _06822_, _06821_);
  and (_06824_, _06823_, _06820_);
  not (_06825_, _04035_);
  and (_06826_, _04047_, _06825_);
  nor (_06827_, _04039_, _04036_);
  and (_06828_, _06827_, _06826_);
  and (_06829_, _06828_, _06824_);
  not (_06830_, _04030_);
  and (_06831_, _04044_, _06830_);
  and (_06832_, _06831_, _04028_);
  not (_06833_, _04024_);
  and (_06834_, _04052_, _06833_);
  and (_06835_, _06834_, _04022_);
  and (_06836_, _06835_, _06832_);
  and (_06837_, _06836_, _06829_);
  and (_06838_, _06837_, _04015_);
  not (_06839_, _06838_);
  and (_06840_, _03665_, \oc8051_golden_model_1.P2INREG [0]);
  and (_06841_, _03646_, \oc8051_golden_model_1.P3INREG [0]);
  nor (_06842_, _06841_, _06840_);
  and (_06843_, _03698_, \oc8051_golden_model_1.P1INREG [0]);
  and (_06844_, _03737_, \oc8051_golden_model_1.P0INREG [0]);
  nor (_06845_, _06844_, _06843_);
  and (_06846_, _06845_, _06842_);
  and (_06847_, _06846_, _04093_);
  and (_06848_, _06847_, _04090_);
  and (_06849_, _06848_, _04077_);
  and (_06850_, _06849_, _04059_);
  nor (_06851_, _06850_, _06518_);
  and (_06852_, _06851_, _06839_);
  and (_06853_, _06852_, _06817_);
  and (_06854_, _06853_, _06805_);
  and (_06855_, _03698_, \oc8051_golden_model_1.P1INREG [5]);
  not (_06856_, _06855_);
  and (_06857_, _03665_, \oc8051_golden_model_1.P2INREG [5]);
  and (_06858_, _03646_, \oc8051_golden_model_1.P3INREG [5]);
  nor (_06859_, _06858_, _06857_);
  and (_06860_, _06859_, _06856_);
  and (_06861_, _06860_, _03950_);
  and (_06862_, _03832_, \oc8051_golden_model_1.P0INREG [5]);
  nor (_06863_, _06862_, _03958_);
  and (_06864_, _06863_, _06861_);
  and (_06865_, _06864_, _03943_);
  and (_06866_, _06865_, _03937_);
  and (_06867_, _06866_, _03917_);
  not (_06868_, _04231_);
  and (_06869_, _04242_, _06868_);
  nor (_06870_, _04234_, _04230_);
  and (_06871_, _06870_, _06869_);
  and (_06872_, _03665_, \oc8051_golden_model_1.P2INREG [4]);
  and (_06873_, _03646_, \oc8051_golden_model_1.P3INREG [4]);
  nor (_06874_, _06873_, _06872_);
  and (_06875_, _03698_, \oc8051_golden_model_1.P1INREG [4]);
  and (_06876_, _03737_, \oc8051_golden_model_1.P0INREG [4]);
  nor (_06877_, _06876_, _06875_);
  and (_06878_, _06877_, _06874_);
  and (_06879_, _06878_, _06871_);
  and (_06880_, _04239_, _04218_);
  and (_06881_, _04254_, _04229_);
  and (_06882_, _06881_, _06880_);
  and (_06883_, _06882_, _06879_);
  and (_06884_, _06883_, _04212_);
  nor (_06885_, _06884_, _06867_);
  and (_06886_, _06885_, _06854_);
  and (_06887_, _06886_, _06792_);
  nor (_06888_, _06887_, _04528_);
  and (_06889_, _06887_, _04528_);
  nor (_06890_, _06889_, _06888_);
  and (_06891_, _06890_, \oc8051_golden_model_1.ACC [7]);
  nor (_06892_, _06890_, \oc8051_golden_model_1.ACC [7]);
  nor (_06893_, _06892_, _06891_);
  not (_06894_, _06893_);
  nor (_06895_, _06886_, _06792_);
  nor (_06896_, _06895_, _06887_);
  nor (_06897_, _06896_, _06026_);
  not (_06898_, _06867_);
  not (_06899_, _06884_);
  and (_06900_, _06854_, _06899_);
  nor (_06901_, _06900_, _06898_);
  nor (_06902_, _06901_, _06886_);
  nor (_06903_, _06902_, _06079_);
  and (_06904_, _06902_, _06079_);
  nor (_06905_, _06904_, _06903_);
  not (_06906_, _06905_);
  nor (_06907_, _06854_, _06899_);
  nor (_06908_, _06907_, _06900_);
  nor (_06909_, _06908_, _06085_);
  and (_06910_, _06908_, _06085_);
  or (_06911_, _06910_, _06909_);
  or (_06912_, _06911_, _06906_);
  nor (_06913_, _06853_, _06805_);
  nor (_06914_, _06913_, _06854_);
  and (_06915_, _06914_, _01689_);
  nor (_06916_, _06914_, _01689_);
  nor (_06917_, _06852_, _06817_);
  nor (_06918_, _06917_, _06853_);
  nor (_06919_, _06918_, _06184_);
  nor (_06920_, _06919_, _06916_);
  or (_06921_, _06920_, _06915_);
  nor (_06922_, _06916_, _06915_);
  and (_06923_, _06918_, _06184_);
  nor (_06924_, _06923_, _06919_);
  and (_06925_, _06924_, _06922_);
  nor (_06926_, _06851_, _06839_);
  nor (_06927_, _06926_, _06852_);
  nor (_06928_, _06927_, _01613_);
  and (_06929_, _06927_, _01613_);
  and (_06930_, _06850_, _06518_);
  nor (_06931_, _06930_, _06851_);
  and (_06932_, _06931_, _01710_);
  nor (_06933_, _06932_, _06929_);
  or (_06934_, _06933_, _06928_);
  nand (_06935_, _06934_, _06925_);
  and (_06936_, _06935_, _06921_);
  nor (_06937_, _06936_, _06912_);
  nor (_06938_, _06909_, _06903_);
  or (_06939_, _06938_, _06904_);
  not (_06940_, _06939_);
  nor (_06941_, _06940_, _06937_);
  and (_06942_, _06896_, _06026_);
  nor (_06943_, _06897_, _06942_);
  not (_06944_, _06943_);
  nor (_06945_, _06944_, _06941_);
  or (_06946_, _06945_, _06897_);
  and (_06947_, _06946_, _06894_);
  nor (_06948_, _06946_, _06894_);
  nor (_06949_, _06948_, _06947_);
  nand (_06950_, _06949_, _06777_);
  and (_06951_, _06950_, _06776_);
  or (_06952_, _06951_, _06774_);
  and (_06953_, _06952_, _06541_);
  or (_06954_, _06953_, _01549_);
  or (_06955_, _01790_, _01550_);
  and (_06956_, _06955_, _02408_);
  and (_06957_, _06956_, _06954_);
  not (_06958_, _04326_);
  nor (_06959_, _04351_, _06958_);
  nor (_06960_, _06959_, _06665_);
  nor (_06961_, _06960_, _02408_);
  or (_06962_, _06961_, _05994_);
  or (_06963_, _06962_, _06957_);
  and (_06964_, _06963_, _06475_);
  or (_06965_, _06964_, _02528_);
  and (_06966_, _04483_, _03680_);
  or (_06967_, _06966_, _06464_);
  or (_06968_, _06967_, _02888_);
  and (_06969_, _06968_, _02043_);
  and (_06970_, _06969_, _06965_);
  nor (_06971_, _04753_, _06472_);
  nor (_06972_, _06971_, _06464_);
  nor (_06973_, _06972_, _02043_);
  or (_06974_, _06973_, _06008_);
  or (_06975_, _06974_, _06970_);
  or (_06976_, _06020_, \oc8051_golden_model_1.ACC [7]);
  and (_06977_, _06976_, _06024_);
  or (_06978_, _06977_, _06355_);
  and (_06979_, _06978_, _06975_);
  or (_06980_, _06979_, _01608_);
  or (_06981_, _01790_, _01609_);
  and (_06982_, _06981_, _06980_);
  or (_06983_, _06982_, _01869_);
  and (_06984_, _02044_, _01637_);
  not (_06985_, _06984_);
  nand (_06986_, _06466_, _01869_);
  and (_06987_, _06986_, _06985_);
  and (_06988_, _06987_, _06983_);
  and (_06989_, _06984_, _01790_);
  and (_06990_, _01983_, _01644_);
  or (_06991_, _06990_, _06989_);
  or (_06992_, _06991_, _06988_);
  and (_06993_, _01978_, _01644_);
  nor (_06994_, _02734_, _06993_);
  not (_06995_, _06994_);
  or (_06996_, _06995_, _06990_);
  nand (_06997_, _06994_, _06408_);
  and (_06998_, _06997_, _06996_);
  and (_06999_, _02049_, _01644_);
  nor (_07000_, _06999_, _06998_);
  and (_07001_, _07000_, _06992_);
  or (_07002_, _06999_, _06995_);
  and (_07003_, _07002_, _06408_);
  or (_07004_, _07003_, _02579_);
  or (_07005_, _07004_, _07001_);
  not (_07006_, _02579_);
  and (_07007_, _04483_, \oc8051_golden_model_1.ACC [7]);
  nor (_07008_, _07007_, _06461_);
  or (_07009_, _07008_, _07006_);
  and (_07010_, _07009_, _07005_);
  or (_07011_, _07010_, _02168_);
  and (_07012_, _02044_, _01644_);
  not (_07013_, _07012_);
  not (_07014_, _02168_);
  or (_07015_, _04779_, _07014_);
  and (_07016_, _07015_, _07013_);
  and (_07017_, _07016_, _07011_);
  and (_07018_, _01790_, \oc8051_golden_model_1.ACC [7]);
  nor (_07019_, _01790_, \oc8051_golden_model_1.ACC [7]);
  nor (_07020_, _07019_, _07018_);
  and (_07021_, _07012_, _07020_);
  or (_07022_, _07021_, _02079_);
  or (_07023_, _07022_, _07017_);
  and (_07024_, _07023_, _06471_);
  or (_07025_, _07024_, _02167_);
  and (_07026_, _01631_, _01533_);
  not (_07027_, _07026_);
  or (_07028_, _06464_, _02912_);
  and (_07029_, _07028_, _07027_);
  and (_07030_, _07029_, _07025_);
  and (_07031_, _01882_, _01631_);
  and (_07032_, _06407_, _07026_);
  or (_07033_, _07032_, _07031_);
  or (_07034_, _07033_, _07030_);
  not (_07035_, _02178_);
  not (_07036_, _07031_);
  or (_07037_, _07036_, _07007_);
  and (_07038_, _07037_, _07035_);
  and (_07039_, _07038_, _07034_);
  and (_07040_, _02044_, _01631_);
  nor (_07041_, _07040_, _02178_);
  not (_07042_, _07041_);
  or (_07043_, _07040_, _04777_);
  and (_07044_, _07043_, _07042_);
  or (_07045_, _07044_, _07039_);
  not (_07046_, _07040_);
  or (_07047_, _07046_, _07018_);
  and (_07048_, _07047_, _02176_);
  and (_07049_, _07048_, _07045_);
  or (_07050_, _07049_, _06468_);
  nor (_07051_, _06452_, _02595_);
  not (_07052_, _07051_);
  and (_07053_, _07052_, _07050_);
  and (_07054_, _06454_, _01647_);
  or (_07055_, _07054_, _02594_);
  nor (_07056_, _07052_, _06406_);
  or (_07057_, _07056_, _07055_);
  or (_07058_, _07057_, _07053_);
  and (_07059_, _01972_, _01647_);
  not (_07060_, _07059_);
  nand (_07061_, _07055_, _06406_);
  and (_07062_, _07061_, _07060_);
  and (_07063_, _07062_, _07058_);
  nor (_07064_, _06406_, _07060_);
  or (_07065_, _07064_, _06462_);
  or (_07066_, _07065_, _07063_);
  and (_07067_, _07066_, _06463_);
  or (_07068_, _07067_, _02171_);
  and (_07069_, _02044_, _01647_);
  not (_07070_, _07069_);
  nand (_07071_, _04778_, _02171_);
  and (_07072_, _07071_, _07070_);
  and (_07073_, _07072_, _07068_);
  nor (_07074_, _07070_, _07019_);
  or (_07075_, _07074_, _07073_);
  and (_07076_, _07075_, _04788_);
  nor (_07077_, _04770_, _06472_);
  nor (_07078_, _07077_, _06464_);
  nor (_07079_, _07078_, _04788_);
  nor (_07080_, _06452_, _02600_);
  nor (_07081_, _07080_, _02699_);
  and (_07082_, _02049_, _01635_);
  not (_07083_, _07082_);
  and (_07084_, _07083_, _07081_);
  not (_07085_, _07084_);
  or (_07086_, _07085_, _07079_);
  or (_07087_, _07086_, _07076_);
  and (_07088_, _06713_, \oc8051_golden_model_1.ACC [6]);
  and (_07089_, _06717_, \oc8051_golden_model_1.ACC [5]);
  and (_07090_, _06723_, \oc8051_golden_model_1.ACC [4]);
  and (_07091_, _06736_, \oc8051_golden_model_1.ACC [3]);
  and (_07092_, _06741_, \oc8051_golden_model_1.ACC [2]);
  and (_07093_, _06748_, \oc8051_golden_model_1.ACC [1]);
  nor (_07094_, _06750_, _06749_);
  and (_07095_, _06752_, \oc8051_golden_model_1.ACC [0]);
  not (_07096_, _07095_);
  nor (_07097_, _07096_, _07094_);
  nor (_07098_, _07097_, _07093_);
  nor (_07099_, _07098_, _06744_);
  nor (_07100_, _07099_, _07092_);
  nor (_07101_, _07100_, _06739_);
  or (_07102_, _07101_, _07091_);
  and (_07103_, _07102_, _06730_);
  nor (_07104_, _07103_, _07090_);
  nor (_07105_, _07104_, _06727_);
  or (_07106_, _07105_, _07089_);
  and (_07107_, _07106_, _06764_);
  nor (_07108_, _07107_, _07088_);
  nor (_07109_, _07108_, _06710_);
  and (_07110_, _07108_, _06710_);
  nor (_07111_, _07110_, _07109_);
  or (_07112_, _07111_, _07084_);
  and (_07113_, _07112_, _07087_);
  and (_07114_, _01882_, _01635_);
  or (_07115_, _07114_, _07113_);
  not (_07116_, _07114_);
  and (_07117_, _06552_, \oc8051_golden_model_1.ACC [6]);
  and (_07118_, _06557_, \oc8051_golden_model_1.ACC [5]);
  and (_07119_, _06563_, \oc8051_golden_model_1.ACC [4]);
  and (_07120_, _06575_, \oc8051_golden_model_1.ACC [3]);
  and (_07121_, _06580_, \oc8051_golden_model_1.ACC [2]);
  and (_07122_, _06587_, \oc8051_golden_model_1.ACC [1]);
  nor (_07123_, _06589_, _06588_);
  and (_07124_, _06591_, \oc8051_golden_model_1.ACC [0]);
  not (_07125_, _07124_);
  nor (_07126_, _07125_, _07123_);
  nor (_07127_, _07126_, _07122_);
  nor (_07128_, _07127_, _06583_);
  nor (_07129_, _07128_, _07121_);
  nor (_07130_, _07129_, _06578_);
  or (_07131_, _07130_, _07120_);
  and (_07132_, _07131_, _06570_);
  nor (_07133_, _07132_, _07119_);
  nor (_07134_, _07133_, _06567_);
  or (_07135_, _07134_, _07118_);
  and (_07136_, _07135_, _06603_);
  nor (_07137_, _07136_, _07117_);
  nor (_07138_, _07137_, _06548_);
  and (_07139_, _07137_, _06548_);
  nor (_07140_, _07139_, _07138_);
  or (_07141_, _07140_, _07116_);
  and (_07142_, _07141_, _02165_);
  and (_07143_, _07142_, _07115_);
  and (_07144_, _02044_, _01635_);
  nor (_07145_, _07144_, _02164_);
  not (_07146_, _07145_);
  and (_07147_, _06896_, \oc8051_golden_model_1.ACC [6]);
  and (_07148_, _06902_, \oc8051_golden_model_1.ACC [5]);
  and (_07149_, _06908_, \oc8051_golden_model_1.ACC [4]);
  and (_07150_, _06914_, \oc8051_golden_model_1.ACC [3]);
  and (_07151_, _06918_, \oc8051_golden_model_1.ACC [2]);
  and (_07152_, _06927_, \oc8051_golden_model_1.ACC [1]);
  nor (_07153_, _06928_, _06929_);
  and (_07154_, _06931_, \oc8051_golden_model_1.ACC [0]);
  not (_07155_, _07154_);
  nor (_07156_, _07155_, _07153_);
  nor (_07157_, _07156_, _07152_);
  nor (_07158_, _07157_, _06924_);
  nor (_07159_, _07158_, _07151_);
  nor (_07160_, _07159_, _06922_);
  or (_07161_, _07160_, _07150_);
  and (_07162_, _07161_, _06911_);
  nor (_07164_, _07162_, _07149_);
  nor (_07165_, _07164_, _06905_);
  or (_07166_, _07165_, _07148_);
  and (_07167_, _07166_, _06944_);
  nor (_07168_, _07167_, _07147_);
  nor (_07169_, _07168_, _06893_);
  and (_07170_, _07168_, _06893_);
  nor (_07171_, _07170_, _07169_);
  or (_07172_, _07171_, _07144_);
  and (_07173_, _07172_, _07146_);
  or (_07174_, _07173_, _07143_);
  and (_07175_, _01635_, _01543_);
  not (_07176_, _07175_);
  not (_07177_, _07144_);
  and (_07178_, _06489_, \oc8051_golden_model_1.ACC [6]);
  nor (_07179_, _06490_, _06491_);
  and (_07180_, _06494_, \oc8051_golden_model_1.ACC [5]);
  and (_07181_, _06498_, \oc8051_golden_model_1.ACC [4]);
  and (_07182_, _06508_, \oc8051_golden_model_1.ACC [3]);
  and (_07183_, _06513_, \oc8051_golden_model_1.ACC [2]);
  and (_07184_, _06521_, \oc8051_golden_model_1.ACC [1]);
  nor (_07185_, _06523_, _06522_);
  nor (_07186_, _06526_, _01710_);
  not (_07187_, _07186_);
  nor (_07188_, _07187_, _07185_);
  nor (_07189_, _07188_, _07184_);
  nor (_07190_, _07189_, _06516_);
  nor (_07191_, _07190_, _07183_);
  nor (_07192_, _07191_, _06511_);
  or (_07193_, _07192_, _07182_);
  and (_07194_, _07193_, _06505_);
  nor (_07195_, _07194_, _07181_);
  nor (_07196_, _07195_, _06502_);
  nor (_07197_, _07196_, _07180_);
  nor (_07198_, _07197_, _07179_);
  nor (_07199_, _07198_, _07178_);
  nor (_07200_, _07199_, _06486_);
  and (_07201_, _07199_, _06486_);
  nor (_07202_, _07201_, _07200_);
  or (_07203_, _07202_, _07177_);
  and (_07204_, _07203_, _07176_);
  and (_07205_, _07204_, _07174_);
  nand (_07206_, _07175_, \oc8051_golden_model_1.ACC [6]);
  nand (_07207_, _07206_, _06458_);
  or (_07208_, _07207_, _07205_);
  and (_07209_, _07208_, _06460_);
  and (_07210_, _01882_, _01652_);
  or (_07211_, _07210_, _07209_);
  not (_07212_, _07210_);
  and (_07213_, _04861_, \oc8051_golden_model_1.ACC [6]);
  nor (_07214_, _04861_, \oc8051_golden_model_1.ACC [6]);
  nor (_07215_, _07213_, _07214_);
  and (_07216_, _05090_, \oc8051_golden_model_1.ACC [5]);
  nor (_07217_, _05090_, \oc8051_golden_model_1.ACC [5]);
  nor (_07218_, _07217_, _07216_);
  not (_07219_, _07218_);
  and (_07220_, _05135_, \oc8051_golden_model_1.ACC [4]);
  nor (_07221_, _05135_, \oc8051_golden_model_1.ACC [4]);
  nor (_07222_, _07220_, _07221_);
  nor (_07223_, _04998_, \oc8051_golden_model_1.ACC [3]);
  not (_07224_, _07223_);
  and (_07225_, _04998_, \oc8051_golden_model_1.ACC [3]);
  not (_07226_, _07225_);
  and (_07227_, _05043_, \oc8051_golden_model_1.ACC [2]);
  nor (_07228_, _05043_, \oc8051_golden_model_1.ACC [2]);
  nor (_07229_, _07227_, _07228_);
  not (_07230_, _07229_);
  and (_07231_, _04907_, \oc8051_golden_model_1.ACC [1]);
  nor (_07232_, _04907_, \oc8051_golden_model_1.ACC [1]);
  nor (_07233_, _07231_, _07232_);
  and (_07234_, _04952_, \oc8051_golden_model_1.ACC [0]);
  and (_07235_, _07234_, _07233_);
  nor (_07236_, _07235_, _07231_);
  nor (_07237_, _07236_, _07230_);
  nor (_07238_, _07237_, _07227_);
  nand (_07239_, _07238_, _07226_);
  and (_07240_, _07239_, _07224_);
  and (_07241_, _07240_, _07222_);
  nor (_07242_, _07241_, _07220_);
  nor (_07243_, _07242_, _07219_);
  or (_07244_, _07243_, _07216_);
  and (_07245_, _07244_, _07215_);
  nor (_07246_, _07245_, _07213_);
  nor (_07247_, _07246_, _07008_);
  and (_07248_, _07246_, _07008_);
  or (_07249_, _07248_, _07247_);
  or (_07250_, _07249_, _07212_);
  and (_07251_, _07250_, _01891_);
  and (_07252_, _07251_, _07211_);
  and (_07253_, _02044_, _01652_);
  nor (_07254_, _07253_, _01890_);
  not (_07255_, _07254_);
  not (_07256_, _07253_);
  and (_07257_, _04528_, _04776_);
  nor (_07258_, _04528_, _04776_);
  nor (_07259_, _07258_, _07257_);
  nor (_07260_, _06791_, _06026_);
  and (_07261_, _06791_, \oc8051_golden_model_1.ACC [6]);
  nor (_07262_, _06791_, \oc8051_golden_model_1.ACC [6]);
  nor (_07263_, _07262_, _07261_);
  not (_07264_, _07263_);
  nor (_07265_, _06867_, _06079_);
  nor (_07266_, _06867_, \oc8051_golden_model_1.ACC [5]);
  and (_07267_, _06867_, \oc8051_golden_model_1.ACC [5]);
  nor (_07268_, _07267_, _07266_);
  nor (_07269_, _06884_, _06085_);
  and (_07270_, _06884_, \oc8051_golden_model_1.ACC [4]);
  nor (_07271_, _06884_, \oc8051_golden_model_1.ACC [4]);
  nor (_07272_, _07271_, _07270_);
  not (_07273_, _07272_);
  nand (_07274_, _06804_, _01689_);
  or (_07275_, _06804_, _01689_);
  nor (_07276_, _06816_, _06184_);
  and (_07277_, _06816_, \oc8051_golden_model_1.ACC [2]);
  nor (_07278_, _06816_, \oc8051_golden_model_1.ACC [2]);
  nor (_07279_, _07278_, _07277_);
  nor (_07280_, _06838_, _01613_);
  nor (_07281_, _06838_, \oc8051_golden_model_1.ACC [1]);
  and (_07282_, _06838_, \oc8051_golden_model_1.ACC [1]);
  nor (_07283_, _07282_, _07281_);
  nor (_07284_, _06850_, _01710_);
  not (_07285_, _07284_);
  nor (_07286_, _07285_, _07283_);
  nor (_07287_, _07286_, _07280_);
  nor (_07288_, _07287_, _07279_);
  nor (_07289_, _07288_, _07276_);
  nand (_07290_, _07289_, _07275_);
  and (_07291_, _07290_, _07274_);
  and (_07292_, _07291_, _07273_);
  nor (_07293_, _07292_, _07269_);
  nor (_07294_, _07293_, _07268_);
  or (_07295_, _07294_, _07265_);
  and (_07296_, _07295_, _07264_);
  nor (_07297_, _07296_, _07260_);
  nor (_07298_, _07297_, _07259_);
  and (_07299_, _07297_, _07259_);
  nor (_07300_, _07299_, _07298_);
  nand (_07301_, _07300_, _07256_);
  and (_07302_, _07301_, _07255_);
  or (_07303_, _07302_, _07252_);
  and (_07304_, _01652_, _01543_);
  not (_07305_, _07304_);
  nor (_07306_, _01922_, _06026_);
  and (_07307_, _01922_, _06026_);
  nor (_07308_, _07307_, _07306_);
  nor (_07309_, _02252_, _06079_);
  and (_07310_, _02252_, _06079_);
  nor (_07311_, _01855_, _06085_);
  and (_07312_, _01855_, _06085_);
  nor (_07313_, _07312_, _07311_);
  nor (_07314_, _01954_, _01689_);
  and (_07315_, _01954_, _01689_);
  nor (_07316_, _02294_, _06184_);
  and (_07317_, _02294_, _06184_);
  nor (_07318_, _07317_, _07316_);
  not (_07319_, _07318_);
  nor (_07320_, _01822_, _01613_);
  and (_07321_, _01822_, _01613_);
  nor (_07322_, _07321_, _07320_);
  nor (_07323_, _02441_, _01710_);
  and (_07324_, _07323_, _07322_);
  nor (_07325_, _07324_, _07320_);
  nor (_07326_, _07325_, _07319_);
  nor (_07327_, _07326_, _07316_);
  nor (_07328_, _07327_, _07315_);
  or (_07329_, _07328_, _07314_);
  and (_07330_, _07329_, _07313_);
  nor (_07331_, _07330_, _07311_);
  nor (_07332_, _07331_, _07310_);
  or (_07333_, _07332_, _07309_);
  and (_07334_, _07333_, _07308_);
  nor (_07335_, _07334_, _07306_);
  nor (_07336_, _07335_, _07020_);
  and (_07337_, _07335_, _07020_);
  or (_07338_, _07337_, _07336_);
  or (_07339_, _07338_, _07256_);
  and (_07340_, _07339_, _07305_);
  and (_07341_, _07340_, _07303_);
  and (_07342_, _07304_, \oc8051_golden_model_1.ACC [6]);
  or (_07343_, _07342_, _02201_);
  or (_07344_, _07343_, _07341_);
  and (_07345_, _02044_, _01641_);
  not (_07346_, _07345_);
  nand (_07347_, _06638_, _02201_);
  and (_07348_, _07347_, _07346_);
  and (_07349_, _07348_, _07344_);
  and (_07350_, _01641_, _01543_);
  nor (_07351_, \oc8051_golden_model_1.ACC [0], \oc8051_golden_model_1.ACC [1]);
  and (_07352_, _07351_, _06125_);
  and (_07353_, _07352_, _06043_);
  and (_07354_, _07353_, _06026_);
  nor (_07355_, _07354_, _04776_);
  and (_07356_, _07354_, _04776_);
  nor (_07357_, _07356_, _07355_);
  nor (_07358_, _07357_, _07346_);
  or (_07359_, _07358_, _07350_);
  or (_07360_, _07359_, _07349_);
  nand (_07361_, _07350_, _06518_);
  and (_07362_, _07361_, _01887_);
  and (_07363_, _07362_, _07360_);
  nor (_07364_, _06687_, _01887_);
  or (_07365_, _07364_, _01537_);
  or (_07366_, _07365_, _07363_);
  and (_07367_, _02044_, _01403_);
  not (_07368_, _07367_);
  and (_07369_, _04264_, _03680_);
  nor (_07370_, _07369_, _06464_);
  nand (_07371_, _07370_, _01537_);
  and (_07372_, _07371_, _07368_);
  and (_07373_, _07372_, _07366_);
  and (_07374_, _01543_, _01403_);
  and (_07375_, \oc8051_golden_model_1.ACC [0], \oc8051_golden_model_1.ACC [1]);
  nand (_07376_, _07375_, _06126_);
  nor (_07377_, _07376_, _06085_);
  and (_07378_, _07377_, \oc8051_golden_model_1.ACC [5]);
  and (_07379_, _07378_, \oc8051_golden_model_1.ACC [6]);
  nor (_07380_, _07379_, \oc8051_golden_model_1.ACC [7]);
  and (_07381_, _07379_, \oc8051_golden_model_1.ACC [7]);
  nor (_07382_, _07381_, _07380_);
  and (_07383_, _07382_, _07367_);
  or (_07384_, _07383_, _07374_);
  or (_07385_, _07384_, _07373_);
  nand (_07386_, _07374_, _01710_);
  and (_07387_, _07386_, _38087_);
  and (_07388_, _07387_, _07385_);
  or (_07389_, _07388_, _06405_);
  and (_37139_, _07389_, _37580_);
  or (_07390_, _38087_, \oc8051_golden_model_1.DPL [7]);
  and (_07391_, _07390_, _37580_);
  not (_07392_, \oc8051_golden_model_1.DPL [7]);
  nor (_07393_, _03856_, _07392_);
  and (_07394_, _04779_, _03856_);
  or (_07395_, _07394_, _07393_);
  and (_07396_, _07395_, _02167_);
  not (_07397_, _03856_);
  nor (_07398_, _07397_, _03616_);
  or (_07399_, _07398_, _07393_);
  or (_07400_, _07399_, _05249_);
  not (_07401_, _02080_);
  and (_07402_, _04496_, _03856_);
  or (_07403_, _07402_, _07393_);
  or (_07404_, _07403_, _02814_);
  and (_07405_, _03748_, \oc8051_golden_model_1.ACC [7]);
  or (_07406_, _07405_, _07393_);
  and (_07407_, _07406_, _02817_);
  nor (_07408_, _02817_, _07392_);
  or (_07409_, _07408_, _02001_);
  or (_07410_, _07409_, _07407_);
  and (_07411_, _07410_, _02840_);
  and (_07412_, _07411_, _07404_);
  and (_07413_, _07399_, _01999_);
  or (_07414_, _07413_, _02006_);
  or (_07415_, _07414_, _07412_);
  and (_07416_, _01965_, _01543_);
  not (_07417_, _07416_);
  or (_07418_, _07406_, _02021_);
  and (_07419_, _07418_, _07417_);
  and (_07420_, _07419_, _07415_);
  and (_07421_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.DPL [0]);
  and (_07422_, _07421_, \oc8051_golden_model_1.DPL [2]);
  and (_07423_, _07422_, \oc8051_golden_model_1.DPL [3]);
  and (_07424_, _07423_, \oc8051_golden_model_1.DPL [4]);
  and (_07425_, _07424_, \oc8051_golden_model_1.DPL [5]);
  and (_07426_, _07425_, \oc8051_golden_model_1.DPL [6]);
  nor (_07427_, _07426_, \oc8051_golden_model_1.DPL [7]);
  and (_07428_, _07426_, \oc8051_golden_model_1.DPL [7]);
  nor (_07429_, _07428_, _07427_);
  and (_07430_, _07429_, _07416_);
  or (_07431_, _07430_, _07420_);
  and (_07432_, _07431_, _07401_);
  nor (_07433_, _04307_, _07401_);
  or (_07434_, _07433_, _05994_);
  or (_07435_, _07434_, _07432_);
  and (_07436_, _07435_, _07400_);
  or (_07437_, _07436_, _02528_);
  or (_07438_, _07393_, _02888_);
  and (_07439_, _04483_, _03748_);
  or (_07440_, _07439_, _07438_);
  and (_07441_, _07440_, _02043_);
  and (_07442_, _07441_, _07437_);
  not (_07443_, _03748_);
  nor (_07444_, _04753_, _07443_);
  or (_07445_, _07444_, _07393_);
  and (_07446_, _07445_, _01602_);
  or (_07447_, _07446_, _01869_);
  or (_07448_, _07447_, _07442_);
  and (_07449_, _04560_, _03748_);
  or (_07450_, _07449_, _07393_);
  or (_07451_, _07450_, _01870_);
  and (_07452_, _07451_, _07448_);
  or (_07453_, _07452_, _02079_);
  and (_07454_, _04771_, _03856_);
  or (_07455_, _07393_, _02166_);
  or (_07456_, _07455_, _07454_);
  and (_07457_, _07456_, _02912_);
  and (_07458_, _07457_, _07453_);
  or (_07459_, _07458_, _07396_);
  and (_07460_, _07459_, _02176_);
  or (_07461_, _07393_, _03755_);
  and (_07462_, _07450_, _02072_);
  and (_07463_, _07462_, _07461_);
  or (_07464_, _07463_, _07460_);
  and (_07465_, _07464_, _02907_);
  and (_07466_, _07406_, _02177_);
  and (_07467_, _07466_, _07461_);
  or (_07468_, _07467_, _02071_);
  or (_07469_, _07468_, _07465_);
  nor (_07470_, _04770_, _07397_);
  or (_07471_, _07393_, _04788_);
  or (_07472_, _07471_, _07470_);
  and (_07473_, _07472_, _04793_);
  and (_07474_, _07473_, _07469_);
  nor (_07475_, _04778_, _07397_);
  or (_07476_, _07475_, _07393_);
  and (_07477_, _07476_, _02173_);
  or (_07478_, _07477_, _02201_);
  or (_07479_, _07478_, _07474_);
  or (_07480_, _07403_, _02303_);
  and (_07481_, _07480_, _01538_);
  and (_07482_, _07481_, _07479_);
  and (_07483_, _04264_, _03856_);
  or (_07484_, _07483_, _07393_);
  and (_07485_, _07484_, _01537_);
  or (_07486_, _07485_, _38088_);
  or (_07487_, _07486_, _07482_);
  and (_37140_, _07487_, _07391_);
  or (_07488_, _38087_, \oc8051_golden_model_1.DPH [7]);
  and (_07489_, _07488_, _37580_);
  not (_07490_, \oc8051_golden_model_1.DPH [7]);
  nor (_07491_, _03850_, _07490_);
  and (_07492_, _04779_, _03850_);
  or (_07493_, _07492_, _07491_);
  and (_07494_, _07493_, _02167_);
  not (_07495_, _03850_);
  nor (_07496_, _07495_, _03616_);
  or (_07497_, _07496_, _07491_);
  or (_07498_, _07497_, _05249_);
  and (_07499_, _04496_, _03850_);
  or (_07500_, _07499_, _07491_);
  or (_07501_, _07500_, _02814_);
  and (_07502_, _03741_, \oc8051_golden_model_1.ACC [7]);
  or (_07503_, _07502_, _07491_);
  and (_07504_, _07503_, _02817_);
  nor (_07505_, _02817_, _07490_);
  or (_07506_, _07505_, _02001_);
  or (_07507_, _07506_, _07504_);
  and (_07508_, _07507_, _02840_);
  and (_07509_, _07508_, _07501_);
  and (_07510_, _07497_, _01999_);
  or (_07511_, _07510_, _02006_);
  or (_07512_, _07511_, _07509_);
  or (_07513_, _07503_, _02021_);
  and (_07514_, _07513_, _07417_);
  and (_07515_, _07514_, _07512_);
  not (_07516_, \oc8051_golden_model_1.DPH [2]);
  and (_07517_, _07428_, \oc8051_golden_model_1.DPH [0]);
  nand (_07518_, _07517_, \oc8051_golden_model_1.DPH [1]);
  nor (_07519_, _07518_, _07516_);
  and (_07520_, _07519_, \oc8051_golden_model_1.DPH [3]);
  and (_07521_, _07520_, \oc8051_golden_model_1.DPH [4]);
  and (_07522_, _07521_, \oc8051_golden_model_1.DPH [5]);
  and (_07523_, _07522_, \oc8051_golden_model_1.DPH [6]);
  and (_07524_, _07523_, _07490_);
  nor (_07525_, _07523_, _07490_);
  or (_07526_, _07525_, _07524_);
  and (_07527_, _07526_, _07416_);
  or (_07528_, _07527_, _07515_);
  and (_07529_, _07528_, _07401_);
  and (_07530_, _02080_, _01790_);
  or (_07531_, _07530_, _05994_);
  or (_07532_, _07531_, _07529_);
  and (_07533_, _07532_, _07498_);
  or (_07534_, _07533_, _02528_);
  or (_07535_, _07491_, _02888_);
  and (_07536_, _04483_, _03741_);
  or (_07537_, _07536_, _07535_);
  and (_07538_, _07537_, _02043_);
  and (_07539_, _07538_, _07534_);
  not (_07540_, _03741_);
  nor (_07541_, _04753_, _07540_);
  or (_07542_, _07541_, _07491_);
  and (_07543_, _07542_, _01602_);
  or (_07544_, _07543_, _01869_);
  or (_07545_, _07544_, _07539_);
  and (_07546_, _04560_, _03741_);
  or (_07547_, _07546_, _07491_);
  or (_07548_, _07547_, _01870_);
  and (_07549_, _07548_, _07545_);
  or (_07550_, _07549_, _02079_);
  and (_07551_, _04771_, _03850_);
  or (_07552_, _07491_, _02166_);
  or (_07553_, _07552_, _07551_);
  and (_07554_, _07553_, _02912_);
  and (_07555_, _07554_, _07550_);
  or (_07556_, _07555_, _07494_);
  and (_07557_, _07556_, _02176_);
  or (_07558_, _07491_, _03755_);
  and (_07559_, _07547_, _02072_);
  and (_07560_, _07559_, _07558_);
  or (_07561_, _07560_, _07557_);
  and (_07562_, _07561_, _02907_);
  and (_07563_, _07503_, _02177_);
  and (_07564_, _07563_, _07558_);
  or (_07565_, _07564_, _02071_);
  or (_07566_, _07565_, _07562_);
  nor (_07567_, _04770_, _07495_);
  or (_07568_, _07491_, _04788_);
  or (_07569_, _07568_, _07567_);
  and (_07570_, _07569_, _04793_);
  and (_07571_, _07570_, _07566_);
  nor (_07572_, _04778_, _07495_);
  or (_07573_, _07572_, _07491_);
  and (_07574_, _07573_, _02173_);
  or (_07575_, _07574_, _02201_);
  or (_07576_, _07575_, _07571_);
  or (_07577_, _07500_, _02303_);
  and (_07578_, _07577_, _01538_);
  and (_07579_, _07578_, _07576_);
  and (_07580_, _04264_, _03850_);
  or (_07581_, _07580_, _07491_);
  and (_07582_, _07581_, _01537_);
  or (_07583_, _07582_, _38088_);
  or (_07584_, _07583_, _07579_);
  and (_37141_, _07584_, _07489_);
  and (_07585_, _38088_, \oc8051_golden_model_1.IE [7]);
  not (_07586_, _03633_);
  and (_07587_, _07586_, \oc8051_golden_model_1.IE [7]);
  and (_07588_, _04779_, _03633_);
  or (_07589_, _07588_, _07587_);
  and (_07590_, _07589_, _02167_);
  nor (_07591_, _07586_, _03616_);
  or (_07592_, _07591_, _07587_);
  or (_07593_, _07592_, _05249_);
  not (_07594_, _04333_);
  and (_07595_, _07594_, \oc8051_golden_model_1.IE [7]);
  and (_07596_, _04364_, _04333_);
  or (_07597_, _07596_, _07595_);
  and (_07598_, _07597_, _01997_);
  and (_07599_, _04496_, _03633_);
  or (_07600_, _07599_, _07587_);
  or (_07601_, _07600_, _02814_);
  and (_07602_, _03633_, \oc8051_golden_model_1.ACC [7]);
  or (_07603_, _07602_, _07587_);
  and (_07604_, _07603_, _02817_);
  and (_07605_, _02818_, \oc8051_golden_model_1.IE [7]);
  or (_07606_, _07605_, _02001_);
  or (_07607_, _07606_, _07604_);
  and (_07608_, _07607_, _02024_);
  and (_07609_, _07608_, _07601_);
  and (_07610_, _04368_, _04333_);
  or (_07611_, _07610_, _07595_);
  and (_07612_, _07611_, _02007_);
  or (_07613_, _07612_, _01999_);
  or (_07614_, _07613_, _07609_);
  or (_07615_, _07592_, _02840_);
  and (_07616_, _07615_, _07614_);
  or (_07617_, _07616_, _02006_);
  or (_07618_, _07603_, _02021_);
  and (_07619_, _07618_, _02025_);
  and (_07620_, _07619_, _07617_);
  or (_07621_, _07620_, _07598_);
  and (_07622_, _07621_, _02861_);
  and (_07623_, _04534_, _04333_);
  or (_07624_, _07623_, _07595_);
  and (_07625_, _07624_, _01991_);
  or (_07626_, _07625_, _07622_);
  and (_07627_, _07626_, _02408_);
  nor (_07628_, _04351_, _07594_);
  or (_07629_, _07628_, _07595_);
  and (_07630_, _07629_, _01875_);
  or (_07631_, _07630_, _05994_);
  or (_07632_, _07631_, _07627_);
  and (_07633_, _07632_, _07593_);
  or (_07634_, _07633_, _02528_);
  and (_07635_, _04483_, _03633_);
  or (_07636_, _07587_, _02888_);
  or (_07637_, _07636_, _07635_);
  and (_07638_, _07637_, _02043_);
  and (_07639_, _07638_, _07634_);
  nor (_07640_, _04753_, _07586_);
  or (_07641_, _07640_, _07587_);
  and (_07642_, _07641_, _01602_);
  or (_07643_, _07642_, _01869_);
  or (_07644_, _07643_, _07639_);
  and (_07645_, _04560_, _03633_);
  or (_07646_, _07645_, _07587_);
  or (_07647_, _07646_, _01870_);
  and (_07648_, _07647_, _07644_);
  or (_07649_, _07648_, _02079_);
  and (_07650_, _04771_, _03633_);
  or (_07651_, _07587_, _02166_);
  or (_07652_, _07651_, _07650_);
  and (_07653_, _07652_, _02912_);
  and (_07654_, _07653_, _07649_);
  or (_07655_, _07654_, _07590_);
  and (_07656_, _07655_, _02176_);
  or (_07657_, _07587_, _03755_);
  and (_07658_, _07646_, _02072_);
  and (_07659_, _07658_, _07657_);
  or (_07660_, _07659_, _07656_);
  and (_07661_, _07660_, _02907_);
  and (_07662_, _07603_, _02177_);
  and (_07663_, _07662_, _07657_);
  or (_07664_, _07663_, _02071_);
  or (_07665_, _07664_, _07661_);
  nor (_07666_, _04770_, _07586_);
  or (_07667_, _07587_, _04788_);
  or (_07668_, _07667_, _07666_);
  and (_07669_, _07668_, _04793_);
  and (_07670_, _07669_, _07665_);
  nor (_07671_, _04778_, _07586_);
  or (_07672_, _07671_, _07587_);
  and (_07673_, _07672_, _02173_);
  or (_07674_, _07673_, _02201_);
  or (_07675_, _07674_, _07670_);
  or (_07676_, _07600_, _02303_);
  and (_07677_, _07676_, _01887_);
  and (_07678_, _07677_, _07675_);
  and (_07679_, _07597_, _01860_);
  or (_07680_, _07679_, _01537_);
  or (_07681_, _07680_, _07678_);
  and (_07682_, _04264_, _03633_);
  or (_07683_, _07587_, _01538_);
  or (_07684_, _07683_, _07682_);
  and (_07685_, _07684_, _38087_);
  and (_07686_, _07685_, _07681_);
  or (_07687_, _07686_, _07585_);
  and (_37142_, _07687_, _37580_);
  and (_07688_, _38088_, \oc8051_golden_model_1.IP [7]);
  not (_07689_, _03670_);
  and (_07690_, _07689_, \oc8051_golden_model_1.IP [7]);
  and (_07691_, _04779_, _03670_);
  or (_07692_, _07691_, _07690_);
  and (_07693_, _07692_, _02167_);
  nor (_07694_, _07689_, _03616_);
  or (_07695_, _07694_, _07690_);
  or (_07696_, _07695_, _05249_);
  not (_07697_, _04324_);
  and (_07698_, _07697_, \oc8051_golden_model_1.IP [7]);
  and (_07699_, _04364_, _04324_);
  or (_07700_, _07699_, _07698_);
  and (_07701_, _07700_, _01997_);
  and (_07702_, _04496_, _03670_);
  or (_07703_, _07702_, _07690_);
  or (_07704_, _07703_, _02814_);
  and (_07705_, _03670_, \oc8051_golden_model_1.ACC [7]);
  or (_07706_, _07705_, _07690_);
  and (_07707_, _07706_, _02817_);
  and (_07708_, _02818_, \oc8051_golden_model_1.IP [7]);
  or (_07709_, _07708_, _02001_);
  or (_07710_, _07709_, _07707_);
  and (_07711_, _07710_, _02024_);
  and (_07712_, _07711_, _07704_);
  and (_07713_, _04368_, _04324_);
  or (_07714_, _07713_, _07698_);
  and (_07715_, _07714_, _02007_);
  or (_07716_, _07715_, _01999_);
  or (_07717_, _07716_, _07712_);
  or (_07718_, _07695_, _02840_);
  and (_07719_, _07718_, _07717_);
  or (_07720_, _07719_, _02006_);
  or (_07721_, _07706_, _02021_);
  and (_07722_, _07721_, _02025_);
  and (_07723_, _07722_, _07720_);
  or (_07724_, _07723_, _07701_);
  and (_07725_, _07724_, _02861_);
  and (_07726_, _04534_, _04324_);
  or (_07727_, _07726_, _07698_);
  and (_07728_, _07727_, _01991_);
  or (_07729_, _07728_, _07725_);
  and (_07730_, _07729_, _02408_);
  nor (_07731_, _04351_, _07697_);
  or (_07732_, _07731_, _07698_);
  and (_07733_, _07732_, _01875_);
  or (_07734_, _07733_, _05994_);
  or (_07735_, _07734_, _07730_);
  and (_07736_, _07735_, _07696_);
  or (_07737_, _07736_, _02528_);
  and (_07738_, _04483_, _03670_);
  or (_07739_, _07690_, _02888_);
  or (_07740_, _07739_, _07738_);
  and (_07741_, _07740_, _02043_);
  and (_07742_, _07741_, _07737_);
  nor (_07743_, _04753_, _07689_);
  or (_07744_, _07743_, _07690_);
  and (_07745_, _07744_, _01602_);
  or (_07746_, _07745_, _01869_);
  or (_07747_, _07746_, _07742_);
  and (_07748_, _04560_, _03670_);
  or (_07749_, _07748_, _07690_);
  or (_07750_, _07749_, _01870_);
  and (_07751_, _07750_, _07747_);
  or (_07752_, _07751_, _02079_);
  and (_07753_, _04771_, _03670_);
  or (_07754_, _07690_, _02166_);
  or (_07755_, _07754_, _07753_);
  and (_07756_, _07755_, _02912_);
  and (_07757_, _07756_, _07752_);
  or (_07758_, _07757_, _07693_);
  and (_07759_, _07758_, _02176_);
  or (_07760_, _07690_, _03755_);
  and (_07761_, _07749_, _02072_);
  and (_07762_, _07761_, _07760_);
  or (_07763_, _07762_, _07759_);
  and (_07764_, _07763_, _02907_);
  and (_07765_, _07706_, _02177_);
  and (_07766_, _07765_, _07760_);
  or (_07767_, _07766_, _02071_);
  or (_07768_, _07767_, _07764_);
  nor (_07769_, _04770_, _07689_);
  or (_07770_, _07690_, _04788_);
  or (_07771_, _07770_, _07769_);
  and (_07772_, _07771_, _04793_);
  and (_07773_, _07772_, _07768_);
  nor (_07774_, _04778_, _07689_);
  or (_07775_, _07774_, _07690_);
  and (_07776_, _07775_, _02173_);
  or (_07777_, _07776_, _02201_);
  or (_07778_, _07777_, _07773_);
  or (_07779_, _07703_, _02303_);
  and (_07780_, _07779_, _01887_);
  and (_07781_, _07780_, _07778_);
  and (_07782_, _07700_, _01860_);
  or (_07783_, _07782_, _01537_);
  or (_07784_, _07783_, _07781_);
  and (_07785_, _04264_, _03670_);
  or (_07786_, _07690_, _01538_);
  or (_07787_, _07786_, _07785_);
  and (_07788_, _07787_, _38087_);
  and (_07789_, _07788_, _07784_);
  or (_07790_, _07789_, _07688_);
  and (_37143_, _07790_, _37580_);
  not (_07791_, _03737_);
  and (_07792_, _07791_, \oc8051_golden_model_1.P0 [7]);
  and (_07793_, _04779_, _03832_);
  or (_07794_, _07793_, _07792_);
  and (_07795_, _07794_, _02167_);
  not (_07796_, _03832_);
  nor (_07797_, _07796_, _03616_);
  or (_07798_, _07797_, _07792_);
  or (_07799_, _07798_, _05249_);
  not (_07800_, _03656_);
  and (_07801_, _07800_, \oc8051_golden_model_1.P0 [7]);
  and (_07802_, _04364_, _03656_);
  or (_07803_, _07802_, _07801_);
  and (_07804_, _07803_, _01997_);
  and (_07805_, _04496_, _03832_);
  or (_07806_, _07805_, _07792_);
  or (_07807_, _07806_, _02814_);
  and (_07808_, _03737_, \oc8051_golden_model_1.ACC [7]);
  or (_07809_, _07808_, _07792_);
  and (_07810_, _07809_, _02817_);
  and (_07811_, _02818_, \oc8051_golden_model_1.P0 [7]);
  or (_07812_, _07811_, _02001_);
  or (_07813_, _07812_, _07810_);
  and (_07814_, _07813_, _02024_);
  and (_07815_, _07814_, _07807_);
  and (_07816_, _04368_, _03656_);
  or (_07817_, _07816_, _07801_);
  and (_07818_, _07817_, _02007_);
  or (_07819_, _07818_, _01999_);
  or (_07820_, _07819_, _07815_);
  or (_07821_, _07798_, _02840_);
  and (_07822_, _07821_, _07820_);
  or (_07823_, _07822_, _02006_);
  or (_07824_, _07809_, _02021_);
  and (_07825_, _07824_, _02025_);
  and (_07826_, _07825_, _07823_);
  or (_07827_, _07826_, _07804_);
  and (_07828_, _07827_, _02861_);
  or (_07829_, _07801_, _04533_);
  and (_07830_, _07829_, _01991_);
  and (_07831_, _07830_, _07817_);
  or (_07832_, _07831_, _07828_);
  and (_07833_, _07832_, _02408_);
  or (_07834_, _04364_, _04350_);
  and (_07835_, _07834_, _03656_);
  or (_07836_, _07835_, _07801_);
  and (_07837_, _07836_, _01875_);
  or (_07838_, _07837_, _05994_);
  or (_07839_, _07838_, _07833_);
  and (_07840_, _07839_, _07799_);
  or (_07841_, _07840_, _02528_);
  or (_07842_, _07792_, _02888_);
  and (_07843_, _04483_, _03737_);
  or (_07844_, _07843_, _07842_);
  and (_07845_, _07844_, _02043_);
  and (_07846_, _07845_, _07841_);
  and (_07847_, _04675_, \oc8051_golden_model_1.P2 [7]);
  and (_07848_, _04703_, \oc8051_golden_model_1.P0 [7]);
  or (_07849_, _07848_, _04682_);
  or (_07850_, _07849_, _07847_);
  and (_07851_, _04706_, \oc8051_golden_model_1.P1 [7]);
  and (_07852_, _04710_, \oc8051_golden_model_1.P3 [7]);
  or (_07853_, _07852_, _07851_);
  nor (_07854_, _07853_, _04687_);
  nand (_07855_, _07854_, _04702_);
  nor (_07856_, _07855_, _07850_);
  and (_07857_, _07856_, _04669_);
  nand (_07858_, _07857_, _04750_);
  or (_07859_, _07858_, _04561_);
  and (_07860_, _07859_, _03832_);
  or (_07861_, _07860_, _07792_);
  and (_07862_, _07861_, _01602_);
  or (_07863_, _07862_, _01869_);
  or (_07864_, _07863_, _07846_);
  and (_07865_, _04560_, _03737_);
  or (_07866_, _07865_, _07792_);
  or (_07867_, _07866_, _01870_);
  and (_07868_, _07867_, _07864_);
  or (_07869_, _07868_, _02079_);
  and (_07870_, _04771_, _03832_);
  or (_07871_, _07792_, _02166_);
  or (_07872_, _07871_, _07870_);
  and (_07873_, _07872_, _02912_);
  and (_07874_, _07873_, _07869_);
  or (_07875_, _07874_, _07795_);
  and (_07876_, _07875_, _02176_);
  or (_07877_, _07792_, _03755_);
  and (_07878_, _07866_, _02072_);
  and (_07879_, _07878_, _07877_);
  or (_07880_, _07879_, _07876_);
  and (_07881_, _07880_, _02907_);
  and (_07882_, _07809_, _02177_);
  and (_07883_, _07882_, _07877_);
  or (_07884_, _07883_, _02071_);
  or (_07885_, _07884_, _07881_);
  nor (_07886_, _04770_, _07796_);
  or (_07887_, _07792_, _04788_);
  or (_07888_, _07887_, _07886_);
  and (_07889_, _07888_, _04793_);
  and (_07890_, _07889_, _07885_);
  nor (_07891_, _04778_, _07796_);
  or (_07892_, _07891_, _07792_);
  and (_07893_, _07892_, _02173_);
  or (_07894_, _07893_, _02201_);
  or (_07895_, _07894_, _07890_);
  or (_07896_, _07806_, _02303_);
  and (_07897_, _07896_, _01887_);
  and (_07898_, _07897_, _07895_);
  and (_07899_, _07803_, _01860_);
  or (_07900_, _07899_, _01537_);
  or (_07901_, _07900_, _07898_);
  and (_07902_, _04264_, _03832_);
  or (_07903_, _07792_, _01538_);
  or (_07904_, _07903_, _07902_);
  and (_07905_, _07904_, _38087_);
  and (_07906_, _07905_, _07901_);
  nor (_07907_, \oc8051_golden_model_1.P0 [7], rst);
  nor (_07908_, _07907_, _03183_);
  or (_37145_, _07908_, _07906_);
  not (_07909_, _03698_);
  and (_07910_, _07909_, \oc8051_golden_model_1.P1 [7]);
  and (_07911_, _04779_, _03698_);
  or (_07912_, _07911_, _07910_);
  and (_07913_, _07912_, _02167_);
  nor (_07914_, _07909_, _03616_);
  or (_07915_, _07914_, _07910_);
  or (_07916_, _07915_, _05249_);
  not (_07917_, _04336_);
  and (_07918_, _07917_, \oc8051_golden_model_1.P1 [7]);
  and (_07919_, _04364_, _04336_);
  or (_07920_, _07919_, _07918_);
  and (_07921_, _07920_, _01997_);
  and (_07922_, _04496_, _03698_);
  or (_07923_, _07922_, _07910_);
  or (_07924_, _07923_, _02814_);
  and (_07925_, _03698_, \oc8051_golden_model_1.ACC [7]);
  or (_07926_, _07925_, _07910_);
  and (_07927_, _07926_, _02817_);
  and (_07928_, _02818_, \oc8051_golden_model_1.P1 [7]);
  or (_07929_, _07928_, _02001_);
  or (_07930_, _07929_, _07927_);
  and (_07931_, _07930_, _02024_);
  and (_07932_, _07931_, _07924_);
  and (_07933_, _04368_, _04336_);
  or (_07934_, _07933_, _07918_);
  and (_07935_, _07934_, _02007_);
  or (_07936_, _07935_, _01999_);
  or (_07937_, _07936_, _07932_);
  or (_07938_, _07915_, _02840_);
  and (_07939_, _07938_, _07937_);
  or (_07940_, _07939_, _02006_);
  or (_07941_, _07926_, _02021_);
  and (_07942_, _07941_, _02025_);
  and (_07943_, _07942_, _07940_);
  or (_07944_, _07943_, _07921_);
  and (_07945_, _07944_, _02861_);
  and (_07946_, _04534_, _04336_);
  or (_07947_, _07946_, _07918_);
  and (_07948_, _07947_, _01991_);
  or (_07949_, _07948_, _07945_);
  and (_07950_, _07949_, _02408_);
  and (_07951_, _07834_, _04336_);
  or (_07952_, _07951_, _07918_);
  and (_07953_, _07952_, _01875_);
  or (_07954_, _07953_, _05994_);
  or (_07955_, _07954_, _07950_);
  and (_07956_, _07955_, _07916_);
  or (_07957_, _07956_, _02528_);
  and (_07958_, _04483_, _03698_);
  or (_07959_, _07910_, _02888_);
  or (_07960_, _07959_, _07958_);
  and (_07961_, _07960_, _02043_);
  and (_07962_, _07961_, _07957_);
  and (_07963_, _07859_, _03698_);
  or (_07964_, _07963_, _07910_);
  and (_07965_, _07964_, _01602_);
  or (_07966_, _07965_, _01869_);
  or (_07967_, _07966_, _07962_);
  and (_07968_, _04560_, _03698_);
  or (_07969_, _07968_, _07910_);
  or (_07970_, _07969_, _01870_);
  and (_07971_, _07970_, _07967_);
  or (_07972_, _07971_, _02079_);
  and (_07973_, _04771_, _03698_);
  or (_07974_, _07910_, _02166_);
  or (_07975_, _07974_, _07973_);
  and (_07976_, _07975_, _02912_);
  and (_07977_, _07976_, _07972_);
  or (_07978_, _07977_, _07913_);
  and (_07979_, _07978_, _02176_);
  or (_07980_, _07910_, _03755_);
  and (_07981_, _07969_, _02072_);
  and (_07982_, _07981_, _07980_);
  or (_07983_, _07982_, _07979_);
  and (_07984_, _07983_, _02907_);
  and (_07985_, _07926_, _02177_);
  and (_07986_, _07985_, _07980_);
  or (_07987_, _07986_, _02071_);
  or (_07988_, _07987_, _07984_);
  nor (_07989_, _04770_, _07909_);
  or (_07990_, _07910_, _04788_);
  or (_07991_, _07990_, _07989_);
  and (_07992_, _07991_, _04793_);
  and (_07993_, _07992_, _07988_);
  nor (_07994_, _04778_, _07909_);
  or (_07995_, _07994_, _07910_);
  and (_07996_, _07995_, _02173_);
  or (_07997_, _07996_, _02201_);
  or (_07998_, _07997_, _07993_);
  or (_07999_, _07923_, _02303_);
  and (_08000_, _07999_, _01887_);
  and (_08001_, _08000_, _07998_);
  and (_08002_, _07920_, _01860_);
  or (_08003_, _08002_, _01537_);
  or (_08004_, _08003_, _08001_);
  and (_08005_, _04264_, _03698_);
  or (_08006_, _07910_, _01538_);
  or (_08007_, _08006_, _08005_);
  and (_08008_, _08007_, _38087_);
  and (_08009_, _08008_, _08004_);
  nor (_08010_, \oc8051_golden_model_1.P1 [7], rst);
  nor (_08011_, _08010_, _03183_);
  or (_37146_, _08011_, _08009_);
  not (_08012_, _03665_);
  and (_08013_, _08012_, \oc8051_golden_model_1.P2 [7]);
  and (_08014_, _04779_, _03665_);
  or (_08015_, _08014_, _08013_);
  and (_08016_, _08015_, _02167_);
  nor (_08017_, _08012_, _03616_);
  or (_08018_, _08017_, _08013_);
  or (_08019_, _08018_, _05249_);
  not (_08020_, _04342_);
  and (_08021_, _08020_, \oc8051_golden_model_1.P2 [7]);
  and (_08022_, _04364_, _04342_);
  or (_08023_, _08022_, _08021_);
  and (_08024_, _08023_, _01997_);
  and (_08025_, _04496_, _03665_);
  or (_08026_, _08025_, _08013_);
  or (_08027_, _08026_, _02814_);
  and (_08028_, _03665_, \oc8051_golden_model_1.ACC [7]);
  or (_08029_, _08028_, _08013_);
  and (_08030_, _08029_, _02817_);
  and (_08031_, _02818_, \oc8051_golden_model_1.P2 [7]);
  or (_08032_, _08031_, _02001_);
  or (_08033_, _08032_, _08030_);
  and (_08034_, _08033_, _02024_);
  and (_08035_, _08034_, _08027_);
  and (_08036_, _04368_, _04342_);
  or (_08037_, _08036_, _08021_);
  and (_08038_, _08037_, _02007_);
  or (_08039_, _08038_, _01999_);
  or (_08040_, _08039_, _08035_);
  or (_08041_, _08018_, _02840_);
  and (_08042_, _08041_, _08040_);
  or (_08043_, _08042_, _02006_);
  or (_08044_, _08029_, _02021_);
  and (_08045_, _08044_, _02025_);
  and (_08046_, _08045_, _08043_);
  or (_08047_, _08046_, _08024_);
  and (_08048_, _08047_, _02861_);
  or (_08049_, _08021_, _04533_);
  and (_08050_, _08049_, _01991_);
  and (_08051_, _08050_, _08037_);
  or (_08052_, _08051_, _08048_);
  and (_08053_, _08052_, _02408_);
  and (_08054_, _07834_, _04342_);
  or (_08055_, _08054_, _08021_);
  and (_08056_, _08055_, _01875_);
  or (_08057_, _08056_, _05994_);
  or (_08058_, _08057_, _08053_);
  and (_08059_, _08058_, _08019_);
  or (_08060_, _08059_, _02528_);
  and (_08061_, _04483_, _03665_);
  or (_08062_, _08013_, _02888_);
  or (_08063_, _08062_, _08061_);
  and (_08064_, _08063_, _02043_);
  and (_08065_, _08064_, _08060_);
  and (_08066_, _07859_, _03665_);
  or (_08067_, _08066_, _08013_);
  and (_08068_, _08067_, _01602_);
  or (_08069_, _08068_, _01869_);
  or (_08070_, _08069_, _08065_);
  and (_08071_, _04560_, _03665_);
  or (_08072_, _08071_, _08013_);
  or (_08073_, _08072_, _01870_);
  and (_08074_, _08073_, _08070_);
  or (_08075_, _08074_, _02079_);
  and (_08076_, _04771_, _03665_);
  or (_08077_, _08013_, _02166_);
  or (_08078_, _08077_, _08076_);
  and (_08079_, _08078_, _02912_);
  and (_08080_, _08079_, _08075_);
  or (_08081_, _08080_, _08016_);
  and (_08082_, _08081_, _02176_);
  or (_08083_, _08013_, _03755_);
  and (_08084_, _08072_, _02072_);
  and (_08085_, _08084_, _08083_);
  or (_08086_, _08085_, _08082_);
  and (_08087_, _08086_, _02907_);
  and (_08088_, _08029_, _02177_);
  and (_08089_, _08088_, _08083_);
  or (_08090_, _08089_, _02071_);
  or (_08091_, _08090_, _08087_);
  nor (_08092_, _04770_, _08012_);
  or (_08093_, _08013_, _04788_);
  or (_08094_, _08093_, _08092_);
  and (_08095_, _08094_, _04793_);
  and (_08096_, _08095_, _08091_);
  nor (_08097_, _04778_, _08012_);
  or (_08098_, _08097_, _08013_);
  and (_08099_, _08098_, _02173_);
  or (_08100_, _08099_, _02201_);
  or (_08101_, _08100_, _08096_);
  or (_08102_, _08026_, _02303_);
  and (_08103_, _08102_, _01887_);
  and (_08104_, _08103_, _08101_);
  and (_08105_, _08023_, _01860_);
  or (_08106_, _08105_, _01537_);
  or (_08107_, _08106_, _08104_);
  and (_08108_, _04264_, _03665_);
  or (_08109_, _08013_, _01538_);
  or (_08110_, _08109_, _08108_);
  and (_08111_, _08110_, _38087_);
  and (_08112_, _08111_, _08107_);
  nor (_08113_, \oc8051_golden_model_1.P2 [7], rst);
  nor (_08114_, _08113_, _03183_);
  or (_37147_, _08114_, _08112_);
  not (_08115_, _03646_);
  and (_08116_, _08115_, \oc8051_golden_model_1.P3 [7]);
  and (_08117_, _04779_, _03646_);
  or (_08118_, _08117_, _08116_);
  and (_08119_, _08118_, _02167_);
  nor (_08120_, _08115_, _03616_);
  or (_08121_, _08120_, _08116_);
  or (_08122_, _08121_, _05249_);
  not (_08123_, _04338_);
  and (_08124_, _08123_, \oc8051_golden_model_1.P3 [7]);
  and (_08125_, _04364_, _04338_);
  or (_08126_, _08125_, _08124_);
  and (_08127_, _08126_, _01997_);
  and (_08128_, _04496_, _03646_);
  or (_08129_, _08128_, _08116_);
  or (_08130_, _08129_, _02814_);
  and (_08131_, _03646_, \oc8051_golden_model_1.ACC [7]);
  or (_08132_, _08131_, _08116_);
  and (_08133_, _08132_, _02817_);
  and (_08134_, _02818_, \oc8051_golden_model_1.P3 [7]);
  or (_08135_, _08134_, _02001_);
  or (_08136_, _08135_, _08133_);
  and (_08137_, _08136_, _02024_);
  and (_08138_, _08137_, _08130_);
  and (_08139_, _04368_, _04338_);
  or (_08140_, _08139_, _08124_);
  and (_08141_, _08140_, _02007_);
  or (_08142_, _08141_, _01999_);
  or (_08143_, _08142_, _08138_);
  or (_08144_, _08121_, _02840_);
  and (_08145_, _08144_, _08143_);
  or (_08146_, _08145_, _02006_);
  or (_08147_, _08132_, _02021_);
  and (_08148_, _08147_, _02025_);
  and (_08149_, _08148_, _08146_);
  or (_08150_, _08149_, _08127_);
  and (_08151_, _08150_, _02861_);
  or (_08152_, _08124_, _04533_);
  and (_08153_, _08152_, _01991_);
  and (_08154_, _08153_, _08140_);
  or (_08155_, _08154_, _08151_);
  and (_08156_, _08155_, _02408_);
  and (_08157_, _07834_, _04338_);
  or (_08158_, _08157_, _08124_);
  and (_08159_, _08158_, _01875_);
  or (_08160_, _08159_, _05994_);
  or (_08161_, _08160_, _08156_);
  and (_08162_, _08161_, _08122_);
  or (_08163_, _08162_, _02528_);
  and (_08164_, _04483_, _03646_);
  or (_08165_, _08116_, _02888_);
  or (_08166_, _08165_, _08164_);
  and (_08167_, _08166_, _02043_);
  and (_08168_, _08167_, _08163_);
  and (_08169_, _07859_, _03646_);
  or (_08170_, _08169_, _08116_);
  and (_08171_, _08170_, _01602_);
  or (_08172_, _08171_, _01869_);
  or (_08173_, _08172_, _08168_);
  and (_08174_, _04560_, _03646_);
  or (_08175_, _08174_, _08116_);
  or (_08176_, _08175_, _01870_);
  and (_08177_, _08176_, _08173_);
  or (_08178_, _08177_, _02079_);
  and (_08179_, _04771_, _03646_);
  or (_08180_, _08116_, _02166_);
  or (_08181_, _08180_, _08179_);
  and (_08182_, _08181_, _02912_);
  and (_08183_, _08182_, _08178_);
  or (_08184_, _08183_, _08119_);
  and (_08185_, _08184_, _02176_);
  or (_08186_, _08116_, _03755_);
  and (_08187_, _08175_, _02072_);
  and (_08188_, _08187_, _08186_);
  or (_08189_, _08188_, _08185_);
  and (_08190_, _08189_, _02907_);
  and (_08191_, _08132_, _02177_);
  and (_08192_, _08191_, _08186_);
  or (_08193_, _08192_, _02071_);
  or (_08194_, _08193_, _08190_);
  nor (_08195_, _04770_, _08115_);
  or (_08196_, _08116_, _04788_);
  or (_08197_, _08196_, _08195_);
  and (_08198_, _08197_, _04793_);
  and (_08199_, _08198_, _08194_);
  nor (_08200_, _04778_, _08115_);
  or (_08201_, _08200_, _08116_);
  and (_08202_, _08201_, _02173_);
  or (_08203_, _08202_, _02201_);
  or (_08204_, _08203_, _08199_);
  or (_08205_, _08129_, _02303_);
  and (_08206_, _08205_, _01887_);
  and (_08207_, _08206_, _08204_);
  and (_08209_, _08126_, _01860_);
  or (_08210_, _08209_, _01537_);
  or (_08211_, _08210_, _08207_);
  and (_08212_, _04264_, _03646_);
  or (_08213_, _08116_, _01538_);
  or (_08214_, _08213_, _08212_);
  and (_08215_, _08214_, _38087_);
  and (_08216_, _08215_, _08211_);
  nor (_08217_, \oc8051_golden_model_1.P3 [7], rst);
  nor (_08218_, _08217_, _03183_);
  or (_37148_, _08218_, _08216_);
  nor (_08219_, _38087_, _06518_);
  nor (_08220_, _04321_, _06518_);
  and (_08221_, _04364_, _04321_);
  or (_08222_, _08221_, _08220_);
  or (_08223_, _08222_, _01887_);
  not (_08224_, _07018_);
  or (_08225_, _07335_, _07019_);
  and (_08226_, _08225_, _07253_);
  nand (_08227_, _08226_, _08224_);
  nor (_08228_, _03676_, _06518_);
  and (_08229_, _04779_, _03676_);
  or (_08230_, _08229_, _08228_);
  and (_08231_, _08230_, _02167_);
  not (_08232_, _03676_);
  nor (_08233_, _04753_, _08232_);
  or (_08234_, _08233_, _08228_);
  and (_08235_, _08234_, _01602_);
  nor (_08236_, _08232_, _03616_);
  or (_08237_, _08236_, _08228_);
  or (_08238_, _08237_, _05249_);
  and (_08239_, _06553_, _06548_);
  nor (_08240_, _08239_, _06546_);
  nand (_08241_, _06602_, _06548_);
  or (_08242_, _08241_, _06600_);
  and (_08243_, _08242_, _08240_);
  and (_08244_, _06542_, _04483_);
  not (_08245_, _06609_);
  or (_08246_, _08245_, _08244_);
  or (_08247_, _08246_, _08243_);
  not (_08248_, _01966_);
  not (_08249_, _01967_);
  not (_08250_, _03855_);
  and (_08251_, _04331_, \oc8051_golden_model_1.SCON [2]);
  not (_08252_, _08251_);
  and (_08253_, _04333_, \oc8051_golden_model_1.IE [2]);
  and (_08254_, _04326_, \oc8051_golden_model_1.ACC [2]);
  nor (_08255_, _08254_, _08253_);
  and (_08256_, _08255_, _08252_);
  and (_08257_, _04321_, \oc8051_golden_model_1.PSW [2]);
  and (_08258_, _04318_, \oc8051_golden_model_1.B [2]);
  nor (_08259_, _08258_, _08257_);
  and (_08260_, _04315_, \oc8051_golden_model_1.TCON [2]);
  and (_08261_, _04324_, \oc8051_golden_model_1.IP [2]);
  nor (_08262_, _08261_, _08260_);
  and (_08263_, _08262_, _08259_);
  and (_08264_, _08263_, _08256_);
  and (_08265_, _03656_, \oc8051_golden_model_1.P0INREG [2]);
  and (_08266_, _04342_, \oc8051_golden_model_1.P2INREG [2]);
  nor (_08267_, _08266_, _08265_);
  and (_08268_, _04336_, \oc8051_golden_model_1.P1INREG [2]);
  and (_08269_, _04338_, \oc8051_golden_model_1.P3INREG [2]);
  nor (_08270_, _08269_, _08268_);
  and (_08271_, _08270_, _08267_);
  and (_08272_, _08271_, _08264_);
  and (_08273_, _08272_, _04108_);
  nor (_08274_, _08273_, _08250_);
  not (_08275_, _03619_);
  and (_08276_, _04315_, \oc8051_golden_model_1.TCON [1]);
  and (_08277_, _04318_, \oc8051_golden_model_1.B [1]);
  nor (_08278_, _08277_, _08276_);
  and (_08279_, _04321_, \oc8051_golden_model_1.PSW [1]);
  not (_08280_, _08279_);
  and (_08281_, _04324_, \oc8051_golden_model_1.IP [1]);
  and (_08282_, _04326_, \oc8051_golden_model_1.ACC [1]);
  nor (_08283_, _08282_, _08281_);
  and (_08284_, _08283_, _08280_);
  and (_08285_, _08284_, _08278_);
  and (_08286_, _04331_, \oc8051_golden_model_1.SCON [1]);
  and (_08287_, _04333_, \oc8051_golden_model_1.IE [1]);
  nor (_08288_, _08287_, _08286_);
  and (_08289_, _03656_, \oc8051_golden_model_1.P0INREG [1]);
  and (_08290_, _04342_, \oc8051_golden_model_1.P2INREG [1]);
  nor (_08291_, _08290_, _08289_);
  and (_08292_, _04336_, \oc8051_golden_model_1.P1INREG [1]);
  and (_08293_, _04338_, \oc8051_golden_model_1.P3INREG [1]);
  nor (_08294_, _08293_, _08292_);
  and (_08295_, _08294_, _08291_);
  and (_08296_, _08295_, _08288_);
  and (_08297_, _08296_, _08285_);
  and (_08298_, _08297_, _04015_);
  nor (_08299_, _08298_, _08275_);
  nor (_08300_, _08299_, _08274_);
  and (_08301_, _03627_, _03391_);
  not (_08302_, _08301_);
  and (_08303_, _04331_, \oc8051_golden_model_1.SCON [4]);
  not (_08304_, _08303_);
  and (_08306_, _04315_, \oc8051_golden_model_1.TCON [4]);
  and (_08307_, _04333_, \oc8051_golden_model_1.IE [4]);
  nor (_08309_, _08307_, _08306_);
  and (_08310_, _08309_, _08304_);
  and (_08312_, _04321_, \oc8051_golden_model_1.PSW [4]);
  and (_08313_, _04318_, \oc8051_golden_model_1.B [4]);
  nor (_08315_, _08313_, _08312_);
  and (_08316_, _04324_, \oc8051_golden_model_1.IP [4]);
  and (_08317_, _04326_, \oc8051_golden_model_1.ACC [4]);
  nor (_08318_, _08317_, _08316_);
  and (_08319_, _08318_, _08315_);
  and (_08320_, _03656_, \oc8051_golden_model_1.P0INREG [4]);
  and (_08321_, _04342_, \oc8051_golden_model_1.P2INREG [4]);
  nor (_08322_, _08321_, _08320_);
  and (_08323_, _04336_, \oc8051_golden_model_1.P1INREG [4]);
  and (_08324_, _04338_, \oc8051_golden_model_1.P3INREG [4]);
  nor (_08325_, _08324_, _08323_);
  and (_08326_, _08325_, _08322_);
  and (_08327_, _08326_, _08319_);
  and (_08328_, _08327_, _08310_);
  and (_08329_, _08328_, _04212_);
  nor (_08330_, _08329_, _08302_);
  nor (_08331_, _04348_, _04367_);
  nor (_08332_, _08331_, _08330_);
  and (_08333_, _08332_, _08300_);
  not (_08334_, _03628_);
  and (_08335_, _04315_, \oc8051_golden_model_1.TCON [0]);
  and (_08336_, _04318_, \oc8051_golden_model_1.B [0]);
  nor (_08337_, _08336_, _08335_);
  and (_08338_, _04321_, \oc8051_golden_model_1.PSW [0]);
  not (_08339_, _08338_);
  and (_08340_, _04324_, \oc8051_golden_model_1.IP [0]);
  and (_08341_, _04326_, \oc8051_golden_model_1.ACC [0]);
  nor (_08342_, _08341_, _08340_);
  and (_08343_, _08342_, _08339_);
  and (_08344_, _08343_, _08337_);
  and (_08345_, _04331_, \oc8051_golden_model_1.SCON [0]);
  and (_08346_, _04333_, \oc8051_golden_model_1.IE [0]);
  nor (_08347_, _08346_, _08345_);
  and (_08348_, _03656_, \oc8051_golden_model_1.P0INREG [0]);
  and (_08349_, _04342_, \oc8051_golden_model_1.P2INREG [0]);
  nor (_08350_, _08349_, _08348_);
  and (_08351_, _04336_, \oc8051_golden_model_1.P1INREG [0]);
  and (_08352_, _04338_, \oc8051_golden_model_1.P3INREG [0]);
  nor (_08353_, _08352_, _08351_);
  and (_08354_, _08353_, _08350_);
  and (_08355_, _08354_, _08347_);
  and (_08356_, _08355_, _08344_);
  and (_08357_, _08356_, _04059_);
  nor (_08358_, _08357_, _08334_);
  and (_08359_, _03728_, _03391_);
  not (_08360_, _08359_);
  and (_08361_, _04315_, \oc8051_golden_model_1.TCON [6]);
  and (_08362_, _04326_, \oc8051_golden_model_1.ACC [6]);
  nor (_08363_, _08362_, _08361_);
  and (_08364_, _04324_, \oc8051_golden_model_1.IP [6]);
  not (_08365_, _08364_);
  and (_08366_, _04321_, \oc8051_golden_model_1.PSW [6]);
  and (_08367_, _04318_, \oc8051_golden_model_1.B [6]);
  nor (_08368_, _08367_, _08366_);
  and (_08369_, _08368_, _08365_);
  and (_08370_, _08369_, _08363_);
  and (_08371_, _04331_, \oc8051_golden_model_1.SCON [6]);
  and (_08372_, _04333_, \oc8051_golden_model_1.IE [6]);
  nor (_08373_, _08372_, _08371_);
  and (_08374_, _03656_, \oc8051_golden_model_1.P0INREG [6]);
  and (_08375_, _04342_, \oc8051_golden_model_1.P2INREG [6]);
  nor (_08376_, _08375_, _08374_);
  and (_08377_, _04336_, \oc8051_golden_model_1.P1INREG [6]);
  and (_08378_, _04338_, \oc8051_golden_model_1.P3INREG [6]);
  nor (_08379_, _08378_, _08377_);
  and (_08380_, _08379_, _08376_);
  and (_08381_, _08380_, _08373_);
  and (_08382_, _08381_, _08370_);
  and (_08383_, _08382_, _03809_);
  nor (_08384_, _08383_, _08360_);
  nor (_08385_, _08384_, _08358_);
  not (_08386_, _03849_);
  and (_08387_, _04315_, \oc8051_golden_model_1.TCON [3]);
  and (_08388_, _04318_, \oc8051_golden_model_1.B [3]);
  nor (_08389_, _08388_, _08387_);
  and (_08390_, _04321_, \oc8051_golden_model_1.PSW [3]);
  not (_08391_, _08390_);
  and (_08392_, _04324_, \oc8051_golden_model_1.IP [3]);
  and (_08393_, _04326_, \oc8051_golden_model_1.ACC [3]);
  nor (_08394_, _08393_, _08392_);
  and (_08395_, _08394_, _08391_);
  and (_08396_, _08395_, _08389_);
  and (_08397_, _04331_, \oc8051_golden_model_1.SCON [3]);
  and (_08398_, _04333_, \oc8051_golden_model_1.IE [3]);
  nor (_08399_, _08398_, _08397_);
  and (_08400_, _03656_, \oc8051_golden_model_1.P0INREG [3]);
  and (_08401_, _04342_, \oc8051_golden_model_1.P2INREG [3]);
  nor (_08402_, _08401_, _08400_);
  and (_08403_, _04336_, \oc8051_golden_model_1.P1INREG [3]);
  and (_08404_, _04338_, \oc8051_golden_model_1.P3INREG [3]);
  nor (_08405_, _08404_, _08403_);
  and (_08406_, _08405_, _08402_);
  and (_08407_, _08406_, _08399_);
  and (_08408_, _08407_, _08396_);
  and (_08409_, _08408_, _03966_);
  nor (_08410_, _08409_, _08386_);
  and (_08411_, _03618_, _03391_);
  not (_08412_, _08411_);
  and (_08413_, _04315_, \oc8051_golden_model_1.TCON [5]);
  and (_08414_, _04326_, \oc8051_golden_model_1.ACC [5]);
  nor (_08415_, _08414_, _08413_);
  and (_08416_, _04321_, \oc8051_golden_model_1.PSW [5]);
  not (_08417_, _08416_);
  and (_08418_, _04324_, \oc8051_golden_model_1.IP [5]);
  and (_08419_, _04318_, \oc8051_golden_model_1.B [5]);
  nor (_08420_, _08419_, _08418_);
  and (_08421_, _08420_, _08417_);
  and (_08422_, _08421_, _08415_);
  and (_08423_, _04331_, \oc8051_golden_model_1.SCON [5]);
  and (_08424_, _04333_, \oc8051_golden_model_1.IE [5]);
  nor (_08425_, _08424_, _08423_);
  and (_08426_, _03656_, \oc8051_golden_model_1.P0INREG [5]);
  and (_08427_, _04342_, \oc8051_golden_model_1.P2INREG [5]);
  nor (_08428_, _08427_, _08426_);
  and (_08429_, _04336_, \oc8051_golden_model_1.P1INREG [5]);
  and (_08430_, _04338_, \oc8051_golden_model_1.P3INREG [5]);
  nor (_08431_, _08430_, _08429_);
  and (_08432_, _08431_, _08428_);
  and (_08433_, _08432_, _08425_);
  and (_08434_, _08433_, _08422_);
  and (_08435_, _08434_, _03917_);
  nor (_08436_, _08435_, _08412_);
  nor (_08437_, _08436_, _08410_);
  and (_08438_, _08437_, _08385_);
  and (_08439_, _08438_, _08333_);
  nor (_08440_, _08439_, _08249_);
  nor (_08441_, _02045_, _01995_);
  or (_08442_, _04998_, _01954_);
  or (_08443_, _05043_, _02294_);
  not (_08444_, _08443_);
  nand (_08445_, _04998_, _01954_);
  nand (_08446_, _08445_, _08444_);
  nand (_08447_, _08446_, _08442_);
  nor (_08448_, _04907_, _01822_);
  nand (_08449_, _04952_, _02441_);
  nor (_08450_, _04907_, _01823_);
  and (_08451_, _04907_, _01823_);
  or (_08452_, _08451_, _08450_);
  and (_08453_, _08452_, _08449_);
  or (_08454_, _08453_, _08448_);
  and (_08455_, _08445_, _08442_);
  nand (_08456_, _05043_, _02294_);
  and (_08457_, _08456_, _08455_);
  and (_08458_, _08457_, _08443_);
  and (_08459_, _08458_, _08454_);
  or (_08460_, _08459_, _08447_);
  or (_08461_, _05135_, _01855_);
  or (_08462_, _05090_, _02252_);
  nand (_08463_, _05090_, _02252_);
  and (_08464_, _08463_, _08462_);
  and (_08465_, _08464_, _08461_);
  nand (_08466_, _05135_, _01855_);
  nand (_08468_, _04861_, _01922_);
  or (_08470_, _04861_, _01922_);
  or (_08472_, _04483_, _03673_);
  and (_08474_, _08472_, _04544_);
  and (_08476_, _08474_, _08470_);
  and (_08478_, _08476_, _08468_);
  and (_08480_, _08478_, _08466_);
  and (_08482_, _08480_, _08465_);
  and (_08484_, _08482_, _08460_);
  nand (_08485_, _08461_, _08462_);
  and (_08486_, _08478_, _08485_);
  and (_08487_, _08486_, _08463_);
  not (_08488_, _08470_);
  nand (_08489_, _08474_, _08488_);
  nand (_08490_, _08489_, _08472_);
  or (_08491_, _08490_, _08487_);
  or (_08492_, _08491_, _08484_);
  and (_08493_, _01882_, _01990_);
  not (_08494_, _08493_);
  or (_08495_, _04952_, _02441_);
  and (_08496_, _08458_, _08453_);
  and (_08497_, _08496_, _08495_);
  and (_08498_, _08497_, _08482_);
  nor (_08499_, _08498_, _08494_);
  and (_08500_, _08499_, _08492_);
  and (_08501_, _04496_, _03676_);
  or (_08502_, _08501_, _08228_);
  or (_08503_, _08502_, _02814_);
  and (_08504_, _03676_, \oc8051_golden_model_1.ACC [7]);
  or (_08505_, _08504_, _08228_);
  and (_08506_, _08505_, _02817_);
  nor (_08507_, _02817_, _06518_);
  or (_08508_, _08507_, _02001_);
  or (_08509_, _08508_, _08506_);
  and (_08510_, _08509_, _06642_);
  and (_08511_, _08510_, _08503_);
  nor (_08512_, _06647_, \oc8051_golden_model_1.PSW [7]);
  not (_08513_, _08512_);
  nor (_08514_, _08513_, _06657_);
  nor (_08515_, _08514_, _06642_);
  and (_08516_, _01881_, _01543_);
  not (_08517_, _08516_);
  nand (_08518_, _08517_, _02008_);
  or (_08519_, _08518_, _08515_);
  or (_08520_, _08519_, _08511_);
  and (_08521_, _04368_, _04321_);
  or (_08522_, _08521_, _08220_);
  or (_08523_, _08522_, _02024_);
  or (_08524_, _08237_, _02840_);
  and (_08525_, _08524_, _08523_);
  and (_08526_, _08525_, _08520_);
  or (_08527_, _08526_, _02006_);
  or (_08528_, _08505_, _02021_);
  and (_08529_, _01877_, _01543_);
  nor (_08530_, _08529_, _01997_);
  and (_08531_, _08530_, _08528_);
  and (_08532_, _08531_, _08527_);
  and (_08533_, _08222_, _01997_);
  not (_08534_, _02050_);
  and (_08535_, _01983_, _01990_);
  not (_08536_, _08535_);
  and (_08537_, _08536_, _02068_);
  and (_08538_, _08537_, _08534_);
  not (_08539_, _08538_);
  or (_08540_, _08539_, _08533_);
  or (_08541_, _08540_, _08532_);
  or (_08542_, _03916_, _03630_);
  and (_08543_, _03616_, _01790_);
  not (_08544_, _08543_);
  and (_08545_, _08544_, _03617_);
  nor (_08546_, _03808_, _03379_);
  and (_08547_, _03808_, _03379_);
  nor (_08548_, _08547_, _08546_);
  and (_08549_, _08548_, _08545_);
  and (_08550_, _03916_, _03630_);
  and (_08551_, _04211_, _03622_);
  nor (_08552_, _04211_, _03622_);
  or (_08553_, _08552_, _08551_);
  nor (_08554_, _08553_, _08550_);
  and (_08555_, _08554_, _08549_);
  and (_08556_, _08555_, _08542_);
  or (_08557_, _03028_, _02441_);
  and (_08558_, _03268_, _01955_);
  and (_08559_, _03455_, _03391_);
  nor (_08560_, _08559_, _08558_);
  or (_08561_, _03268_, _01955_);
  or (_08562_, _03455_, _03391_);
  and (_08563_, _08562_, _08561_);
  and (_08564_, _08563_, _08560_);
  or (_08565_, _02811_, _01823_);
  or (_08566_, _03042_, _02584_);
  nand (_08567_, _02811_, _01823_);
  and (_08568_, _08567_, _08566_);
  and (_08569_, _08568_, _08565_);
  and (_08570_, _08569_, _08564_);
  and (_08571_, _08570_, _08557_);
  and (_08572_, _08571_, _08556_);
  not (_08573_, _08572_);
  nand (_08574_, _08565_, _08566_);
  nand (_08575_, _08567_, _08574_);
  and (_08576_, _08575_, _08564_);
  and (_08577_, _08561_, _08559_);
  or (_08578_, _08577_, _08558_);
  or (_08579_, _08578_, _08576_);
  and (_08580_, _08579_, _08556_);
  or (_08581_, _08550_, _08551_);
  and (_08582_, _08581_, _08549_);
  and (_08583_, _08582_, _08542_);
  and (_08584_, _08547_, _03617_);
  or (_08585_, _08584_, _08543_);
  or (_08586_, _08585_, _08583_);
  or (_08587_, _08586_, _08580_);
  and (_08588_, _08587_, _08573_);
  or (_08589_, _08588_, _08538_);
  and (_08590_, _08589_, _08494_);
  and (_08591_, _08590_, _08541_);
  or (_08592_, _08591_, _08500_);
  and (_08593_, _08592_, _08441_);
  nor (_08594_, _06804_, \oc8051_golden_model_1.ACC [3]);
  and (_08595_, _06804_, \oc8051_golden_model_1.ACC [3]);
  nor (_08596_, _08595_, _08594_);
  and (_08597_, _08596_, _07279_);
  not (_08598_, _07283_);
  and (_08599_, _06850_, \oc8051_golden_model_1.ACC [0]);
  nor (_08600_, _08599_, _08598_);
  or (_08601_, _08600_, _07281_);
  and (_08602_, _08601_, _08597_);
  not (_08603_, _08595_);
  and (_08604_, _07278_, _08603_);
  or (_08605_, _08604_, _08594_);
  or (_08606_, _08605_, _08602_);
  and (_08607_, _07268_, _07272_);
  not (_08608_, _07259_);
  and (_08609_, _07263_, _08608_);
  and (_08610_, _08609_, _08607_);
  and (_08611_, _08610_, _08606_);
  not (_08612_, _07267_);
  or (_08613_, _07271_, _07266_);
  and (_08614_, _08613_, _08612_);
  and (_08615_, _08609_, _08614_);
  nor (_08616_, _04528_, \oc8051_golden_model_1.ACC [7]);
  and (_08617_, _07262_, _08608_);
  or (_08618_, _08617_, _08616_);
  or (_08619_, _08618_, _08615_);
  or (_08620_, _08619_, _08611_);
  nor (_08621_, _06850_, \oc8051_golden_model_1.ACC [0]);
  nor (_08622_, _08599_, _08621_);
  and (_08623_, _08622_, _07283_);
  and (_08624_, _08623_, _08597_);
  and (_08625_, _08610_, _08624_);
  nor (_08626_, _08625_, _02444_);
  and (_08627_, _08626_, _08620_);
  and (_08628_, _01990_, _01543_);
  nor (_08629_, _07314_, _07315_);
  nor (_08630_, _08629_, _07318_);
  nor (_08631_, _01822_, \oc8051_golden_model_1.ACC [1]);
  and (_08632_, _01822_, \oc8051_golden_model_1.ACC [1]);
  and (_08633_, _02441_, \oc8051_golden_model_1.ACC [0]);
  nor (_08634_, _08633_, _08632_);
  or (_08635_, _08634_, _08631_);
  and (_08636_, _08635_, _08630_);
  nand (_08637_, _01954_, \oc8051_golden_model_1.ACC [3]);
  nor (_08638_, _01954_, \oc8051_golden_model_1.ACC [3]);
  nor (_08639_, _02294_, \oc8051_golden_model_1.ACC [2]);
  or (_08640_, _08639_, _08638_);
  and (_08641_, _08640_, _08637_);
  or (_08642_, _08641_, _08636_);
  nor (_08643_, _07310_, _07309_);
  nor (_08644_, _08643_, _07313_);
  nor (_08645_, _07308_, _07020_);
  and (_08646_, _08645_, _08644_);
  and (_08647_, _08646_, _08642_);
  nand (_08648_, _02252_, \oc8051_golden_model_1.ACC [5]);
  nor (_08649_, _02252_, \oc8051_golden_model_1.ACC [5]);
  nor (_08650_, _01855_, \oc8051_golden_model_1.ACC [4]);
  or (_08651_, _08650_, _08649_);
  and (_08652_, _08651_, _08648_);
  and (_08653_, _08645_, _08652_);
  and (_08654_, _01790_, _04776_);
  or (_08655_, _01922_, \oc8051_golden_model_1.ACC [6]);
  nor (_08656_, _08655_, _07020_);
  or (_08657_, _08656_, _08654_);
  or (_08658_, _08657_, _08653_);
  or (_08659_, _08658_, _08647_);
  and (_08660_, _02441_, _01710_);
  nor (_08661_, _08660_, _07323_);
  nor (_08662_, _08661_, _07322_);
  and (_08663_, _08662_, _08630_);
  and (_08664_, _08663_, _08646_);
  nor (_08665_, _08664_, _02046_);
  and (_08666_, _08665_, _08659_);
  or (_08667_, _08666_, _08628_);
  or (_08668_, _08667_, _08627_);
  or (_08669_, _08668_, _08593_);
  nand (_08670_, _08628_, \oc8051_golden_model_1.PSW [7]);
  and (_08671_, _08670_, _02861_);
  and (_08672_, _08671_, _08669_);
  or (_08673_, _08220_, _04533_);
  and (_08674_, _08673_, _01991_);
  and (_08675_, _08674_, _08522_);
  or (_08676_, _08675_, _01992_);
  or (_08677_, _08676_, _08672_);
  nor (_08678_, _05279_, _01967_);
  and (_08679_, _03656_, \oc8051_golden_model_1.P0 [2]);
  and (_08680_, _04338_, \oc8051_golden_model_1.P3 [2]);
  nor (_08681_, _08680_, _08679_);
  and (_08682_, _04336_, \oc8051_golden_model_1.P1 [2]);
  and (_08683_, _04342_, \oc8051_golden_model_1.P2 [2]);
  nor (_08684_, _08683_, _08682_);
  and (_08685_, _08684_, _08681_);
  and (_08686_, _08685_, _08264_);
  and (_08687_, _08686_, _04108_);
  nor (_08688_, _08687_, _08250_);
  and (_08689_, _04342_, \oc8051_golden_model_1.P2 [1]);
  and (_08690_, _04338_, \oc8051_golden_model_1.P3 [1]);
  nor (_08691_, _08690_, _08689_);
  and (_08692_, _03656_, \oc8051_golden_model_1.P0 [1]);
  and (_08693_, _04336_, \oc8051_golden_model_1.P1 [1]);
  nor (_08694_, _08693_, _08692_);
  and (_08695_, _08694_, _08691_);
  and (_08696_, _08695_, _08288_);
  and (_08697_, _08696_, _08285_);
  and (_08698_, _08697_, _04015_);
  nor (_08699_, _08698_, _08275_);
  nor (_08700_, _08699_, _08688_);
  and (_08701_, _04342_, \oc8051_golden_model_1.P2 [4]);
  and (_08702_, _04338_, \oc8051_golden_model_1.P3 [4]);
  nor (_08703_, _08702_, _08701_);
  and (_08704_, _03656_, \oc8051_golden_model_1.P0 [4]);
  and (_08705_, _04336_, \oc8051_golden_model_1.P1 [4]);
  nor (_08706_, _08705_, _08704_);
  and (_08707_, _08706_, _08703_);
  and (_08708_, _08707_, _08319_);
  and (_08709_, _08708_, _08310_);
  and (_08710_, _08709_, _04212_);
  nor (_08711_, _08302_, _08710_);
  nor (_08712_, _08711_, _04532_);
  and (_08713_, _08712_, _08700_);
  and (_08714_, _04342_, \oc8051_golden_model_1.P2 [0]);
  and (_08715_, _04338_, \oc8051_golden_model_1.P3 [0]);
  nor (_08716_, _08715_, _08714_);
  and (_08717_, _03656_, \oc8051_golden_model_1.P0 [0]);
  and (_08718_, _04336_, \oc8051_golden_model_1.P1 [0]);
  nor (_08719_, _08718_, _08717_);
  and (_08720_, _08719_, _08716_);
  and (_08721_, _08720_, _08347_);
  and (_08722_, _08721_, _08344_);
  and (_08723_, _08722_, _04059_);
  nor (_08724_, _08723_, _08334_);
  and (_08725_, _04342_, \oc8051_golden_model_1.P2 [6]);
  and (_08726_, _04338_, \oc8051_golden_model_1.P3 [6]);
  nor (_08727_, _08726_, _08725_);
  and (_08728_, _03656_, \oc8051_golden_model_1.P0 [6]);
  and (_08729_, _04336_, \oc8051_golden_model_1.P1 [6]);
  nor (_08730_, _08729_, _08728_);
  and (_08731_, _08730_, _08727_);
  and (_08732_, _08731_, _08373_);
  and (_08733_, _08732_, _08370_);
  and (_08734_, _08733_, _03809_);
  nor (_08735_, _08360_, _08734_);
  nor (_08736_, _08735_, _08724_);
  and (_08737_, _04342_, \oc8051_golden_model_1.P2 [3]);
  and (_08738_, _04338_, \oc8051_golden_model_1.P3 [3]);
  nor (_08739_, _08738_, _08737_);
  and (_08740_, _03656_, \oc8051_golden_model_1.P0 [3]);
  and (_08741_, _04336_, \oc8051_golden_model_1.P1 [3]);
  nor (_08742_, _08741_, _08740_);
  and (_08743_, _08742_, _08739_);
  and (_08744_, _08743_, _08399_);
  and (_08745_, _08744_, _08396_);
  and (_08746_, _08745_, _03966_);
  nor (_08747_, _08746_, _08386_);
  and (_08748_, _04342_, \oc8051_golden_model_1.P2 [5]);
  and (_08749_, _04338_, \oc8051_golden_model_1.P3 [5]);
  nor (_08750_, _08749_, _08748_);
  and (_08751_, _03656_, \oc8051_golden_model_1.P0 [5]);
  and (_08752_, _04336_, \oc8051_golden_model_1.P1 [5]);
  nor (_08753_, _08752_, _08751_);
  and (_08754_, _08753_, _08750_);
  and (_08755_, _08754_, _08425_);
  and (_08756_, _08755_, _08422_);
  and (_08757_, _08756_, _03917_);
  nor (_08758_, _08412_, _08757_);
  nor (_08759_, _08758_, _08747_);
  and (_08760_, _08759_, _08736_);
  and (_08761_, _08760_, _08713_);
  nand (_08762_, _08761_, \oc8051_golden_model_1.PSW [7]);
  nand (_08763_, _08762_, _01992_);
  and (_08764_, _08763_, _08678_);
  and (_08765_, _08764_, _08677_);
  or (_08766_, _08765_, _08440_);
  and (_08767_, _08766_, _08248_);
  and (_08768_, _01977_, _01548_);
  not (_08769_, _08768_);
  or (_08770_, _03122_, _02372_);
  and (_08771_, _08770_, _08769_);
  not (_08772_, _08771_);
  or (_08773_, _08761_, \oc8051_golden_model_1.PSW [7]);
  and (_08774_, _08773_, _01966_);
  or (_08775_, _08774_, _08772_);
  or (_08776_, _08775_, _08767_);
  and (_08777_, _01972_, _01548_);
  not (_08778_, _08777_);
  nor (_08779_, _03808_, _03616_);
  and (_08780_, _06703_, _08779_);
  and (_08781_, _06714_, _06710_);
  nor (_08782_, _08781_, _06708_);
  nand (_08783_, _06763_, _06710_);
  or (_08784_, _08783_, _06761_);
  and (_08785_, _08784_, _08782_);
  or (_08786_, _08785_, _08780_);
  and (_08787_, _08786_, _08778_);
  or (_08788_, _08787_, _06700_);
  and (_08789_, _08788_, _08776_);
  and (_08790_, _08786_, _08777_);
  or (_08791_, _08790_, _06609_);
  or (_08792_, _08791_, _08789_);
  and (_08793_, _08792_, _08247_);
  or (_08794_, _08793_, _01963_);
  and (_08795_, _06897_, _06893_);
  nor (_08796_, _08795_, _06891_);
  nand (_08797_, _06943_, _06893_);
  or (_08798_, _08797_, _06941_);
  and (_08799_, _08798_, _08796_);
  not (_08800_, _04528_);
  and (_08801_, _06887_, _08800_);
  or (_08802_, _08801_, _02036_);
  or (_08803_, _08802_, _08799_);
  and (_08804_, _08803_, _06777_);
  and (_08805_, _08804_, _08794_);
  and (_08806_, _06478_, _03682_);
  and (_08807_, _06490_, _06486_);
  nor (_08808_, _08807_, _06484_);
  nand (_08809_, _07179_, _06486_);
  or (_08810_, _08809_, _06535_);
  and (_08811_, _08810_, _08808_);
  or (_08812_, _08811_, _08806_);
  and (_08813_, _08812_, _06476_);
  or (_08814_, _08813_, _05994_);
  or (_08815_, _08814_, _08805_);
  and (_08816_, _08815_, _08238_);
  or (_08817_, _08816_, _02528_);
  and (_08818_, _04483_, _03676_);
  or (_08819_, _08228_, _02888_);
  or (_08820_, _08819_, _08818_);
  and (_08821_, _08820_, _02043_);
  and (_08822_, _08821_, _08817_);
  or (_08823_, _08822_, _08235_);
  nor (_08824_, _06008_, _01959_);
  and (_08825_, _08824_, _08823_);
  nor (_08826_, _08761_, _06518_);
  and (_08827_, _08826_, _01959_);
  or (_08828_, _08827_, _01869_);
  or (_08829_, _08828_, _08825_);
  and (_08830_, _04560_, _03676_);
  or (_08831_, _08830_, _08228_);
  or (_08832_, _08831_, _01870_);
  and (_08833_, _08832_, _08829_);
  or (_08834_, _08833_, _01958_);
  nand (_08835_, _08761_, _06518_);
  or (_08836_, _08835_, _02576_);
  and (_08837_, _08836_, _08834_);
  or (_08838_, _08837_, _02079_);
  and (_08839_, _04771_, _03676_);
  or (_08840_, _08228_, _02166_);
  or (_08841_, _08840_, _08839_);
  and (_08842_, _08841_, _02912_);
  and (_08843_, _08842_, _08838_);
  or (_08844_, _08843_, _08231_);
  and (_08845_, _08844_, _02176_);
  or (_08846_, _08228_, _03755_);
  and (_08847_, _08831_, _02072_);
  and (_08848_, _08847_, _08846_);
  or (_08849_, _08848_, _08845_);
  and (_08850_, _08849_, _02907_);
  and (_08851_, _08505_, _02177_);
  and (_08852_, _08851_, _08846_);
  or (_08853_, _08852_, _02071_);
  or (_08854_, _08853_, _08850_);
  nor (_08855_, _04770_, _08232_);
  or (_08856_, _08228_, _04788_);
  or (_08857_, _08856_, _08855_);
  and (_08858_, _08857_, _04793_);
  and (_08859_, _08858_, _08854_);
  nor (_08860_, _04778_, _08232_);
  or (_08861_, _08860_, _08228_);
  and (_08862_, _08861_, _02173_);
  or (_08863_, _08862_, _07085_);
  or (_08864_, _08863_, _08859_);
  nor (_08865_, _06707_, _04776_);
  or (_08866_, _08865_, _07109_);
  or (_08867_, _08866_, _08780_);
  or (_08868_, _08867_, _07084_);
  and (_08870_, _08868_, _08864_);
  or (_08871_, _08870_, _07114_);
  and (_08872_, _06545_, \oc8051_golden_model_1.ACC [7]);
  or (_08873_, _08872_, _07138_);
  or (_08874_, _07116_, _08244_);
  or (_08875_, _08874_, _08873_);
  and (_08876_, _08875_, _02165_);
  and (_08877_, _08876_, _08871_);
  nor (_08878_, _06890_, _04776_);
  or (_08879_, _08878_, _07169_);
  or (_08881_, _08879_, _08801_);
  and (_08882_, _08881_, _02164_);
  or (_08883_, _08882_, _07144_);
  or (_08884_, _08883_, _08877_);
  and (_08885_, _06483_, \oc8051_golden_model_1.ACC [7]);
  or (_08886_, _08885_, _07200_);
  or (_08887_, _07177_, _08806_);
  or (_08888_, _08887_, _08886_);
  and (_08889_, _08888_, _07176_);
  and (_08890_, _08889_, _08884_);
  nand (_08892_, _07175_, \oc8051_golden_model_1.ACC [7]);
  nand (_08893_, _08892_, _06458_);
  or (_08894_, _08893_, _08890_);
  and (_08895_, _06445_, _06408_);
  not (_08896_, _06406_);
  or (_08897_, _06410_, _06407_);
  and (_08898_, _08897_, _08896_);
  or (_08899_, _08898_, _06458_);
  or (_08900_, _08899_, _08895_);
  and (_08901_, _08900_, _08894_);
  or (_08903_, _08901_, _07210_);
  and (_08904_, _07245_, _07008_);
  not (_08905_, _06461_);
  or (_08906_, _07213_, _07007_);
  and (_08907_, _08906_, _08905_);
  or (_08908_, _08907_, _07212_);
  or (_08909_, _08908_, _08904_);
  and (_08910_, _08909_, _01891_);
  and (_08911_, _08910_, _08903_);
  not (_08912_, _07257_);
  not (_08914_, _07258_);
  nand (_08915_, _07297_, _08914_);
  and (_08916_, _08915_, _01890_);
  and (_08917_, _08916_, _08912_);
  or (_08918_, _08917_, _07253_);
  or (_08919_, _08918_, _08911_);
  and (_08920_, _08919_, _08227_);
  or (_08921_, _08920_, _02201_);
  not (_08922_, _07350_);
  or (_08923_, _08502_, _02303_);
  and (_08925_, _08923_, _08922_);
  and (_08926_, _08925_, _08921_);
  and (_08927_, _07350_, \oc8051_golden_model_1.ACC [0]);
  or (_08928_, _08927_, _01860_);
  or (_08929_, _08928_, _08926_);
  and (_08930_, _08929_, _08223_);
  or (_08931_, _08930_, _01537_);
  and (_08932_, _04264_, _03676_);
  or (_08933_, _08228_, _01538_);
  or (_08934_, _08933_, _08932_);
  and (_08936_, _08934_, _38087_);
  and (_08937_, _08936_, _08931_);
  or (_08938_, _08937_, _08219_);
  and (_37149_, _08938_, _37580_);
  or (_08939_, _38087_, \oc8051_golden_model_1.PCON [7]);
  and (_08940_, _08939_, _37580_);
  not (_08941_, _03662_);
  and (_08942_, _08941_, \oc8051_golden_model_1.PCON [7]);
  and (_08943_, _04779_, _03662_);
  or (_08944_, _08943_, _08942_);
  and (_08945_, _08944_, _02167_);
  nor (_08946_, _08941_, _03616_);
  or (_08947_, _08946_, _08942_);
  or (_08948_, _08947_, _05249_);
  and (_08949_, _04496_, _03662_);
  or (_08950_, _08949_, _08942_);
  or (_08951_, _08950_, _02814_);
  and (_08952_, _03662_, \oc8051_golden_model_1.ACC [7]);
  or (_08953_, _08952_, _08942_);
  and (_08954_, _08953_, _02817_);
  and (_08955_, _02818_, \oc8051_golden_model_1.PCON [7]);
  or (_08956_, _08955_, _02001_);
  or (_08957_, _08956_, _08954_);
  and (_08958_, _08957_, _02840_);
  and (_08959_, _08958_, _08951_);
  and (_08960_, _08947_, _01999_);
  or (_08961_, _08960_, _08959_);
  and (_08962_, _08961_, _02021_);
  and (_08963_, _08953_, _02006_);
  or (_08964_, _08963_, _05994_);
  or (_08965_, _08964_, _08962_);
  and (_08966_, _08965_, _08948_);
  or (_08967_, _08966_, _02528_);
  and (_08968_, _04483_, _03662_);
  or (_08969_, _08942_, _02888_);
  or (_08970_, _08969_, _08968_);
  and (_08971_, _08970_, _02043_);
  and (_08972_, _08971_, _08967_);
  nor (_08973_, _04753_, _08941_);
  or (_08974_, _08973_, _08942_);
  and (_08975_, _08974_, _01602_);
  or (_08976_, _08975_, _01869_);
  or (_08977_, _08976_, _08972_);
  and (_08978_, _04560_, _03662_);
  or (_08979_, _08978_, _08942_);
  or (_08980_, _08979_, _01870_);
  and (_08981_, _08980_, _08977_);
  or (_08982_, _08981_, _02079_);
  and (_08983_, _04771_, _03662_);
  or (_08984_, _08942_, _02166_);
  or (_08985_, _08984_, _08983_);
  and (_08986_, _08985_, _02912_);
  and (_08987_, _08986_, _08982_);
  or (_08988_, _08987_, _08945_);
  and (_08989_, _08988_, _02176_);
  or (_08990_, _08942_, _03755_);
  and (_08991_, _08979_, _02072_);
  and (_08992_, _08991_, _08990_);
  or (_08993_, _08992_, _08989_);
  and (_08994_, _08993_, _02907_);
  and (_08995_, _08953_, _02177_);
  and (_08996_, _08995_, _08990_);
  or (_08997_, _08996_, _02071_);
  or (_08998_, _08997_, _08994_);
  nor (_08999_, _04770_, _08941_);
  or (_09000_, _08942_, _04788_);
  or (_09001_, _09000_, _08999_);
  and (_09002_, _09001_, _04793_);
  and (_09003_, _09002_, _08998_);
  nor (_09004_, _04778_, _08941_);
  or (_09005_, _09004_, _08942_);
  and (_09006_, _09005_, _02173_);
  or (_09007_, _09006_, _02201_);
  or (_09008_, _09007_, _09003_);
  or (_09009_, _08950_, _02303_);
  and (_09010_, _09009_, _01538_);
  and (_09011_, _09010_, _09008_);
  and (_09012_, _04264_, _03662_);
  or (_09013_, _09012_, _08942_);
  and (_09014_, _09013_, _01537_);
  or (_09015_, _09014_, _38088_);
  or (_09016_, _09015_, _09011_);
  and (_37150_, _09016_, _08940_);
  or (_09017_, _38087_, \oc8051_golden_model_1.SBUF [7]);
  and (_09018_, _09017_, _37580_);
  not (_09019_, _03625_);
  and (_09020_, _09019_, \oc8051_golden_model_1.SBUF [7]);
  and (_09021_, _04779_, _03625_);
  or (_09022_, _09021_, _09020_);
  and (_09023_, _09022_, _02167_);
  and (_09024_, _04496_, _03625_);
  or (_09025_, _09024_, _09020_);
  or (_09026_, _09025_, _02814_);
  and (_09027_, _03625_, \oc8051_golden_model_1.ACC [7]);
  or (_09028_, _09027_, _09020_);
  and (_09029_, _09028_, _02817_);
  and (_09030_, _02818_, \oc8051_golden_model_1.SBUF [7]);
  or (_09031_, _09030_, _02001_);
  or (_09032_, _09031_, _09029_);
  and (_09033_, _09032_, _02840_);
  and (_09034_, _09033_, _09026_);
  nor (_09035_, _09019_, _03616_);
  or (_09036_, _09035_, _09020_);
  and (_09037_, _09036_, _01999_);
  or (_09038_, _09037_, _09034_);
  and (_09039_, _09038_, _02021_);
  and (_09040_, _09028_, _02006_);
  or (_09041_, _09040_, _05994_);
  or (_09042_, _09041_, _09039_);
  or (_09043_, _09036_, _05249_);
  and (_09044_, _09043_, _09042_);
  or (_09045_, _09044_, _02528_);
  and (_09046_, _04483_, _03625_);
  or (_09047_, _09020_, _02888_);
  or (_09048_, _09047_, _09046_);
  and (_09049_, _09048_, _02043_);
  and (_09050_, _09049_, _09045_);
  nor (_09051_, _04753_, _09019_);
  or (_09052_, _09051_, _09020_);
  and (_09053_, _09052_, _01602_);
  or (_09054_, _09053_, _01869_);
  or (_09055_, _09054_, _09050_);
  and (_09056_, _04560_, _03625_);
  or (_09057_, _09056_, _09020_);
  or (_09058_, _09057_, _01870_);
  and (_09059_, _09058_, _09055_);
  or (_09060_, _09059_, _02079_);
  and (_09061_, _04771_, _03625_);
  or (_09062_, _09020_, _02166_);
  or (_09063_, _09062_, _09061_);
  and (_09064_, _09063_, _02912_);
  and (_09065_, _09064_, _09060_);
  or (_09066_, _09065_, _09023_);
  and (_09067_, _09066_, _02176_);
  or (_09068_, _09020_, _03755_);
  and (_09069_, _09057_, _02072_);
  and (_09070_, _09069_, _09068_);
  or (_09071_, _09070_, _09067_);
  and (_09072_, _09071_, _02907_);
  and (_09073_, _09028_, _02177_);
  and (_09074_, _09073_, _09068_);
  or (_09075_, _09074_, _02071_);
  or (_09076_, _09075_, _09072_);
  nor (_09077_, _04770_, _09019_);
  or (_09078_, _09020_, _04788_);
  or (_09079_, _09078_, _09077_);
  and (_09080_, _09079_, _04793_);
  and (_09081_, _09080_, _09076_);
  nor (_09082_, _04778_, _09019_);
  or (_09083_, _09082_, _09020_);
  and (_09084_, _09083_, _02173_);
  or (_09085_, _09084_, _02201_);
  or (_09086_, _09085_, _09081_);
  or (_09087_, _09025_, _02303_);
  and (_09088_, _09087_, _01538_);
  and (_09089_, _09088_, _09086_);
  and (_09090_, _04264_, _03625_);
  or (_09091_, _09090_, _09020_);
  and (_09092_, _09091_, _01537_);
  or (_09093_, _09092_, _38088_);
  or (_09094_, _09093_, _09089_);
  and (_37151_, _09094_, _09018_);
  and (_09095_, _38088_, \oc8051_golden_model_1.SCON [7]);
  not (_09096_, _03716_);
  and (_09097_, _09096_, \oc8051_golden_model_1.SCON [7]);
  and (_09098_, _04779_, _03716_);
  or (_09099_, _09098_, _09097_);
  and (_09100_, _09099_, _02167_);
  nor (_09101_, _09096_, _03616_);
  or (_09102_, _09101_, _09097_);
  or (_09103_, _09102_, _05249_);
  not (_09104_, _04331_);
  and (_09105_, _09104_, \oc8051_golden_model_1.SCON [7]);
  and (_09106_, _04364_, _04331_);
  or (_09107_, _09106_, _09105_);
  and (_09108_, _09107_, _01997_);
  and (_09109_, _04496_, _03716_);
  or (_09110_, _09109_, _09097_);
  or (_09111_, _09110_, _02814_);
  and (_09112_, _03716_, \oc8051_golden_model_1.ACC [7]);
  or (_09113_, _09112_, _09097_);
  and (_09114_, _09113_, _02817_);
  and (_09115_, _02818_, \oc8051_golden_model_1.SCON [7]);
  or (_09116_, _09115_, _02001_);
  or (_09117_, _09116_, _09114_);
  and (_09118_, _09117_, _02024_);
  and (_09119_, _09118_, _09111_);
  and (_09120_, _04368_, _04331_);
  or (_09121_, _09120_, _09105_);
  and (_09122_, _09121_, _02007_);
  or (_09123_, _09122_, _01999_);
  or (_09124_, _09123_, _09119_);
  or (_09125_, _09102_, _02840_);
  and (_09126_, _09125_, _09124_);
  or (_09127_, _09126_, _02006_);
  or (_09128_, _09113_, _02021_);
  and (_09129_, _09128_, _02025_);
  and (_09130_, _09129_, _09127_);
  or (_09131_, _09130_, _09108_);
  and (_09132_, _09131_, _02861_);
  or (_09133_, _09105_, _04533_);
  and (_09134_, _09133_, _01991_);
  and (_09135_, _09134_, _09121_);
  or (_09136_, _09135_, _09132_);
  and (_09137_, _09136_, _02408_);
  nor (_09138_, _04351_, _09104_);
  or (_09139_, _09138_, _09105_);
  and (_09140_, _09139_, _01875_);
  or (_09141_, _09140_, _05994_);
  or (_09142_, _09141_, _09137_);
  and (_09143_, _09142_, _09103_);
  or (_09144_, _09143_, _02528_);
  and (_09145_, _04483_, _03716_);
  or (_09146_, _09097_, _02888_);
  or (_09147_, _09146_, _09145_);
  and (_09148_, _09147_, _02043_);
  and (_09149_, _09148_, _09144_);
  nor (_09150_, _04753_, _09096_);
  or (_09151_, _09150_, _09097_);
  and (_09152_, _09151_, _01602_);
  or (_09153_, _09152_, _01869_);
  or (_09154_, _09153_, _09149_);
  and (_09155_, _04560_, _03716_);
  or (_09156_, _09155_, _09097_);
  or (_09157_, _09156_, _01870_);
  and (_09158_, _09157_, _09154_);
  or (_09159_, _09158_, _02079_);
  and (_09160_, _04771_, _03716_);
  or (_09161_, _09097_, _02166_);
  or (_09162_, _09161_, _09160_);
  and (_09163_, _09162_, _02912_);
  and (_09164_, _09163_, _09159_);
  or (_09165_, _09164_, _09100_);
  and (_09166_, _09165_, _02176_);
  or (_09167_, _09097_, _03755_);
  and (_09168_, _09156_, _02072_);
  and (_09169_, _09168_, _09167_);
  or (_09170_, _09169_, _09166_);
  and (_09171_, _09170_, _02907_);
  and (_09172_, _09113_, _02177_);
  and (_09173_, _09172_, _09167_);
  or (_09174_, _09173_, _02071_);
  or (_09175_, _09174_, _09171_);
  nor (_09176_, _04770_, _09096_);
  or (_09177_, _09097_, _04788_);
  or (_09178_, _09177_, _09176_);
  and (_09179_, _09178_, _04793_);
  and (_09180_, _09179_, _09175_);
  nor (_09181_, _04778_, _09096_);
  or (_09182_, _09181_, _09097_);
  and (_09183_, _09182_, _02173_);
  or (_09184_, _09183_, _02201_);
  or (_09185_, _09184_, _09180_);
  or (_09186_, _09110_, _02303_);
  and (_09187_, _09186_, _01887_);
  and (_09188_, _09187_, _09185_);
  and (_09189_, _09107_, _01860_);
  or (_09190_, _09189_, _01537_);
  or (_09191_, _09190_, _09188_);
  and (_09192_, _04264_, _03716_);
  or (_09193_, _09097_, _01538_);
  or (_09194_, _09193_, _09192_);
  and (_09195_, _09194_, _38087_);
  and (_09196_, _09195_, _09191_);
  or (_09197_, _09196_, _09095_);
  and (_37152_, _09197_, _37580_);
  not (_09198_, \oc8051_golden_model_1.SP [7]);
  nor (_09199_, _38087_, _09198_);
  and (_09200_, _03549_, \oc8051_golden_model_1.SP [4]);
  and (_09201_, _09200_, \oc8051_golden_model_1.SP [5]);
  and (_09202_, _09201_, \oc8051_golden_model_1.SP [6]);
  or (_09203_, _09202_, \oc8051_golden_model_1.SP [7]);
  nand (_09204_, _09202_, \oc8051_golden_model_1.SP [7]);
  and (_09205_, _09204_, _09203_);
  or (_09206_, _09205_, _02942_);
  nor (_09207_, _03745_, _09198_);
  and (_09208_, _04779_, _03853_);
  or (_09209_, _09208_, _09207_);
  and (_09210_, _09209_, _02167_);
  and (_09211_, _05249_, _02888_);
  not (_09212_, _09211_);
  not (_09213_, _03853_);
  nor (_09214_, _09213_, _03616_);
  or (_09215_, _09207_, _02528_);
  or (_09216_, _09215_, _09214_);
  and (_09217_, _09216_, _09212_);
  and (_09218_, _04496_, _03853_);
  or (_09219_, _09218_, _09207_);
  or (_09220_, _09219_, _02814_);
  and (_09221_, _03745_, \oc8051_golden_model_1.ACC [7]);
  or (_09222_, _09221_, _09207_);
  and (_09223_, _09222_, _02817_);
  nor (_09224_, _02817_, _02823_);
  and (_09225_, _09224_, \oc8051_golden_model_1.SP [7]);
  and (_09226_, _09205_, _02823_);
  or (_09227_, _09226_, _02001_);
  or (_09228_, _09227_, _09225_);
  or (_09229_, _09228_, _09223_);
  and (_09230_, _09229_, _01558_);
  and (_09231_, _09230_, _09220_);
  and (_09232_, _09205_, _03279_);
  or (_09233_, _09232_, _01999_);
  or (_09234_, _09233_, _09231_);
  not (_09235_, \oc8051_golden_model_1.SP [6]);
  not (_09236_, \oc8051_golden_model_1.SP [5]);
  not (_09237_, \oc8051_golden_model_1.SP [4]);
  and (_09238_, _04399_, _09237_);
  and (_09239_, _09238_, _09236_);
  and (_09240_, _09239_, _09235_);
  and (_09241_, _09240_, _01864_);
  nor (_09242_, _09241_, _09198_);
  and (_09243_, _09241_, _09198_);
  nor (_09244_, _09243_, _09242_);
  nand (_09245_, _09244_, _01999_);
  and (_09246_, _09245_, _09234_);
  or (_09247_, _09246_, _02006_);
  or (_09248_, _09222_, _02021_);
  and (_09249_, _09248_, _01880_);
  and (_09250_, _09249_, _09247_);
  and (_09251_, _09202_, \oc8051_golden_model_1.SP [0]);
  or (_09252_, _09251_, \oc8051_golden_model_1.SP [7]);
  nand (_09253_, _09251_, \oc8051_golden_model_1.SP [7]);
  and (_09254_, _09253_, _09252_);
  and (_09255_, _09254_, _01878_);
  or (_09256_, _09255_, _03132_);
  or (_09257_, _09256_, _09250_);
  or (_09258_, _09205_, _03133_);
  and (_09259_, _09258_, _05249_);
  and (_09260_, _09259_, _09257_);
  or (_09261_, _09260_, _09217_);
  or (_09262_, _09207_, _02888_);
  and (_09263_, _04483_, _03745_);
  or (_09264_, _09263_, _09262_);
  and (_09265_, _09264_, _02043_);
  and (_09266_, _09265_, _09261_);
  nor (_09267_, _04753_, _09213_);
  or (_09268_, _09267_, _09207_);
  and (_09269_, _09268_, _01602_);
  or (_09270_, _09269_, _01869_);
  or (_09271_, _09270_, _09266_);
  and (_09272_, _04560_, _03745_);
  or (_09273_, _09272_, _09207_);
  or (_09274_, _09273_, _01870_);
  and (_09275_, _09274_, _09271_);
  or (_09276_, _09275_, _01638_);
  not (_09277_, _01638_);
  or (_09278_, _09205_, _09277_);
  and (_09279_, _09278_, _09276_);
  or (_09280_, _09279_, _02079_);
  and (_09281_, _04771_, _03853_);
  or (_09282_, _09207_, _02166_);
  or (_09283_, _09282_, _09281_);
  and (_09284_, _09283_, _02912_);
  and (_09285_, _09284_, _09280_);
  or (_09286_, _09285_, _09210_);
  and (_09287_, _09286_, _02176_);
  or (_09288_, _09207_, _03755_);
  and (_09289_, _09273_, _02072_);
  and (_09290_, _09289_, _09288_);
  or (_09291_, _09290_, _09287_);
  nor (_09292_, _02177_, _01632_);
  and (_09293_, _09292_, _09291_);
  and (_09294_, _09222_, _02177_);
  and (_09295_, _09294_, _09288_);
  and (_09296_, _09205_, _01632_);
  or (_09297_, _09296_, _02071_);
  or (_09298_, _09297_, _09295_);
  or (_09299_, _09298_, _09293_);
  nor (_09300_, _04770_, _09213_);
  or (_09301_, _09207_, _04788_);
  or (_09302_, _09301_, _09300_);
  and (_09303_, _09302_, _09299_);
  or (_09304_, _09303_, _02173_);
  not (_09305_, _02185_);
  nor (_09306_, _04778_, _09213_);
  or (_09307_, _09207_, _04793_);
  or (_09308_, _09307_, _09306_);
  and (_09309_, _09308_, _09305_);
  and (_09310_, _09309_, _09304_);
  or (_09311_, _09240_, \oc8051_golden_model_1.SP [7]);
  nand (_09312_, _09240_, \oc8051_golden_model_1.SP [7]);
  and (_09313_, _09312_, _09311_);
  and (_09314_, _09313_, _02185_);
  or (_09315_, _09314_, _01636_);
  or (_09316_, _09315_, _09310_);
  or (_09317_, _09205_, _04799_);
  and (_09318_, _09317_, _09316_);
  or (_09319_, _09318_, _01888_);
  or (_09320_, _09313_, _01889_);
  and (_09321_, _09320_, _02303_);
  and (_09322_, _09321_, _09319_);
  and (_09323_, _09219_, _02201_);
  or (_09324_, _09323_, _03370_);
  or (_09325_, _09324_, _09322_);
  and (_09326_, _09325_, _09206_);
  or (_09327_, _09326_, _01537_);
  and (_09328_, _04264_, _03853_);
  or (_09329_, _09207_, _01538_);
  or (_09330_, _09329_, _09328_);
  and (_09331_, _09330_, _38087_);
  and (_09332_, _09331_, _09327_);
  or (_09333_, _09332_, _09199_);
  and (_37153_, _09333_, _37580_);
  and (_09334_, _38088_, \oc8051_golden_model_1.TCON [7]);
  not (_09335_, _03693_);
  and (_09336_, _09335_, \oc8051_golden_model_1.TCON [7]);
  and (_09337_, _04779_, _03693_);
  or (_09338_, _09337_, _09336_);
  and (_09339_, _09338_, _02167_);
  nor (_09340_, _09335_, _03616_);
  or (_09341_, _09340_, _09336_);
  or (_09342_, _09341_, _05249_);
  not (_09343_, _04315_);
  and (_09344_, _09343_, \oc8051_golden_model_1.TCON [7]);
  and (_09345_, _04364_, _04315_);
  or (_09346_, _09345_, _09344_);
  and (_09347_, _09346_, _01997_);
  and (_09348_, _04496_, _03693_);
  or (_09349_, _09348_, _09336_);
  or (_09350_, _09349_, _02814_);
  and (_09351_, _03693_, \oc8051_golden_model_1.ACC [7]);
  or (_09352_, _09351_, _09336_);
  and (_09353_, _09352_, _02817_);
  and (_09354_, _02818_, \oc8051_golden_model_1.TCON [7]);
  or (_09355_, _09354_, _02001_);
  or (_09356_, _09355_, _09353_);
  and (_09357_, _09356_, _02024_);
  and (_09358_, _09357_, _09350_);
  and (_09359_, _04368_, _04315_);
  or (_09360_, _09359_, _09344_);
  and (_09361_, _09360_, _02007_);
  or (_09362_, _09361_, _01999_);
  or (_09363_, _09362_, _09358_);
  or (_09364_, _09341_, _02840_);
  and (_09365_, _09364_, _09363_);
  or (_09366_, _09365_, _02006_);
  or (_09367_, _09352_, _02021_);
  and (_09368_, _09367_, _02025_);
  and (_09369_, _09368_, _09366_);
  or (_09370_, _09369_, _09347_);
  and (_09371_, _09370_, _02861_);
  or (_09372_, _09344_, _04533_);
  and (_09373_, _09372_, _01991_);
  and (_09374_, _09373_, _09360_);
  or (_09375_, _09374_, _09371_);
  and (_09376_, _09375_, _02408_);
  nor (_09377_, _04351_, _09343_);
  or (_09378_, _09377_, _09344_);
  and (_09379_, _09378_, _01875_);
  or (_09380_, _09379_, _05994_);
  or (_09381_, _09380_, _09376_);
  and (_09382_, _09381_, _09342_);
  or (_09383_, _09382_, _02528_);
  and (_09384_, _04483_, _03693_);
  or (_09385_, _09336_, _02888_);
  or (_09386_, _09385_, _09384_);
  and (_09387_, _09386_, _02043_);
  and (_09388_, _09387_, _09383_);
  nor (_09389_, _04753_, _09335_);
  or (_09390_, _09389_, _09336_);
  and (_09391_, _09390_, _01602_);
  or (_09392_, _09391_, _01869_);
  or (_09393_, _09392_, _09388_);
  and (_09394_, _04560_, _03693_);
  or (_09395_, _09394_, _09336_);
  or (_09396_, _09395_, _01870_);
  and (_09397_, _09396_, _09393_);
  or (_09398_, _09397_, _02079_);
  and (_09399_, _04771_, _03693_);
  or (_09400_, _09336_, _02166_);
  or (_09401_, _09400_, _09399_);
  and (_09402_, _09401_, _02912_);
  and (_09403_, _09402_, _09398_);
  or (_09404_, _09403_, _09339_);
  and (_09405_, _09404_, _02176_);
  or (_09406_, _09336_, _03755_);
  and (_09407_, _09395_, _02072_);
  and (_09408_, _09407_, _09406_);
  or (_09409_, _09408_, _09405_);
  and (_09410_, _09409_, _02907_);
  and (_09411_, _09352_, _02177_);
  and (_09412_, _09411_, _09406_);
  or (_09413_, _09412_, _02071_);
  or (_09414_, _09413_, _09410_);
  nor (_09415_, _04770_, _09335_);
  or (_09416_, _09336_, _04788_);
  or (_09417_, _09416_, _09415_);
  and (_09418_, _09417_, _04793_);
  and (_09419_, _09418_, _09414_);
  nor (_09420_, _04778_, _09335_);
  or (_09421_, _09420_, _09336_);
  and (_09422_, _09421_, _02173_);
  or (_09423_, _09422_, _02201_);
  or (_09424_, _09423_, _09419_);
  or (_09425_, _09349_, _02303_);
  and (_09426_, _09425_, _01887_);
  and (_09427_, _09426_, _09424_);
  and (_09428_, _09346_, _01860_);
  or (_09429_, _09428_, _01537_);
  or (_09430_, _09429_, _09427_);
  and (_09431_, _04264_, _03693_);
  or (_09432_, _09336_, _01538_);
  or (_09433_, _09432_, _09431_);
  and (_09434_, _09433_, _38087_);
  and (_09435_, _09434_, _09430_);
  or (_09436_, _09435_, _09334_);
  and (_37154_, _09436_, _37580_);
  or (_09437_, _38087_, \oc8051_golden_model_1.TH0 [7]);
  and (_09438_, _09437_, _37580_);
  not (_09439_, _03691_);
  and (_09440_, _09439_, \oc8051_golden_model_1.TH0 [7]);
  and (_09441_, _04779_, _03691_);
  or (_09442_, _09441_, _09440_);
  and (_09443_, _09442_, _02167_);
  and (_09444_, _04496_, _03691_);
  or (_09445_, _09444_, _09440_);
  or (_09446_, _09445_, _02814_);
  and (_09447_, _03691_, \oc8051_golden_model_1.ACC [7]);
  or (_09448_, _09447_, _09440_);
  and (_09449_, _09448_, _02817_);
  and (_09450_, _02818_, \oc8051_golden_model_1.TH0 [7]);
  or (_09451_, _09450_, _02001_);
  or (_09452_, _09451_, _09449_);
  and (_09453_, _09452_, _02840_);
  and (_09454_, _09453_, _09446_);
  nor (_09455_, _09439_, _03616_);
  or (_09456_, _09455_, _09440_);
  and (_09457_, _09456_, _01999_);
  or (_09458_, _09457_, _09454_);
  and (_09459_, _09458_, _02021_);
  and (_09460_, _09448_, _02006_);
  or (_09461_, _09460_, _05994_);
  or (_09462_, _09461_, _09459_);
  or (_09463_, _09456_, _05249_);
  and (_09464_, _09463_, _09462_);
  or (_09465_, _09464_, _02528_);
  and (_09466_, _04483_, _03691_);
  or (_09467_, _09440_, _02888_);
  or (_09468_, _09467_, _09466_);
  and (_09469_, _09468_, _02043_);
  and (_09470_, _09469_, _09465_);
  nor (_09471_, _04753_, _09439_);
  or (_09472_, _09471_, _09440_);
  and (_09473_, _09472_, _01602_);
  or (_09474_, _09473_, _01869_);
  or (_09475_, _09474_, _09470_);
  and (_09476_, _04560_, _03691_);
  or (_09477_, _09476_, _09440_);
  or (_09478_, _09477_, _01870_);
  and (_09479_, _09478_, _09475_);
  or (_09480_, _09479_, _02079_);
  and (_09481_, _04771_, _03691_);
  or (_09482_, _09440_, _02166_);
  or (_09483_, _09482_, _09481_);
  and (_09484_, _09483_, _02912_);
  and (_09485_, _09484_, _09480_);
  or (_09486_, _09485_, _09443_);
  and (_09487_, _09486_, _02176_);
  or (_09488_, _09440_, _03755_);
  and (_09489_, _09477_, _02072_);
  and (_09490_, _09489_, _09488_);
  or (_09491_, _09490_, _09487_);
  and (_09492_, _09491_, _02907_);
  and (_09493_, _09448_, _02177_);
  and (_09494_, _09493_, _09488_);
  or (_09495_, _09494_, _02071_);
  or (_09496_, _09495_, _09492_);
  nor (_09497_, _04770_, _09439_);
  or (_09498_, _09440_, _04788_);
  or (_09499_, _09498_, _09497_);
  and (_09500_, _09499_, _04793_);
  and (_09501_, _09500_, _09496_);
  nor (_09502_, _04778_, _09439_);
  or (_09503_, _09502_, _09440_);
  and (_09504_, _09503_, _02173_);
  or (_09505_, _09504_, _02201_);
  or (_09506_, _09505_, _09501_);
  or (_09507_, _09445_, _02303_);
  and (_09508_, _09507_, _01538_);
  and (_09509_, _09508_, _09506_);
  and (_09510_, _04264_, _03691_);
  or (_09511_, _09510_, _09440_);
  and (_09512_, _09511_, _01537_);
  or (_09513_, _09512_, _38088_);
  or (_09514_, _09513_, _09509_);
  and (_37156_, _09514_, _09438_);
  or (_09515_, _38087_, \oc8051_golden_model_1.TH1 [7]);
  and (_09516_, _09515_, _37580_);
  not (_09517_, _03722_);
  and (_09518_, _09517_, \oc8051_golden_model_1.TH1 [7]);
  and (_09519_, _04779_, _03722_);
  or (_09520_, _09519_, _09518_);
  and (_09521_, _09520_, _02167_);
  nor (_09522_, _09517_, _03616_);
  or (_09523_, _09522_, _09518_);
  or (_09524_, _09523_, _05249_);
  and (_09525_, _04496_, _03722_);
  or (_09526_, _09525_, _09518_);
  or (_09527_, _09526_, _02814_);
  and (_09528_, _03722_, \oc8051_golden_model_1.ACC [7]);
  or (_09529_, _09528_, _09518_);
  and (_09530_, _09529_, _02817_);
  and (_09531_, _02818_, \oc8051_golden_model_1.TH1 [7]);
  or (_09532_, _09531_, _02001_);
  or (_09533_, _09532_, _09530_);
  and (_09534_, _09533_, _02840_);
  and (_09535_, _09534_, _09527_);
  and (_09536_, _09523_, _01999_);
  or (_09537_, _09536_, _09535_);
  and (_09538_, _09537_, _02021_);
  and (_09539_, _09529_, _02006_);
  or (_09540_, _09539_, _05994_);
  or (_09541_, _09540_, _09538_);
  and (_09542_, _09541_, _09524_);
  or (_09543_, _09542_, _02528_);
  and (_09544_, _04483_, _03722_);
  or (_09545_, _09518_, _02888_);
  or (_09546_, _09545_, _09544_);
  and (_09547_, _09546_, _02043_);
  and (_09548_, _09547_, _09543_);
  nor (_09549_, _04753_, _09517_);
  or (_09550_, _09549_, _09518_);
  and (_09551_, _09550_, _01602_);
  or (_09552_, _09551_, _01869_);
  or (_09553_, _09552_, _09548_);
  and (_09554_, _04560_, _03722_);
  or (_09555_, _09554_, _09518_);
  or (_09556_, _09555_, _01870_);
  and (_09557_, _09556_, _09553_);
  or (_09558_, _09557_, _02079_);
  and (_09559_, _04771_, _03722_);
  or (_09560_, _09518_, _02166_);
  or (_09561_, _09560_, _09559_);
  and (_09562_, _09561_, _02912_);
  and (_09563_, _09562_, _09558_);
  or (_09564_, _09563_, _09521_);
  and (_09565_, _09564_, _02176_);
  or (_09566_, _09518_, _03755_);
  and (_09567_, _09555_, _02072_);
  and (_09568_, _09567_, _09566_);
  or (_09569_, _09568_, _09565_);
  and (_09570_, _09569_, _02907_);
  and (_09571_, _09529_, _02177_);
  and (_09572_, _09571_, _09566_);
  or (_09573_, _09572_, _02071_);
  or (_09574_, _09573_, _09570_);
  nor (_09575_, _04770_, _09517_);
  or (_09576_, _09518_, _04788_);
  or (_09577_, _09576_, _09575_);
  and (_09578_, _09577_, _04793_);
  and (_09579_, _09578_, _09574_);
  nor (_09580_, _04778_, _09517_);
  or (_09581_, _09580_, _09518_);
  and (_09582_, _09581_, _02173_);
  or (_09583_, _09582_, _02201_);
  or (_09584_, _09583_, _09579_);
  or (_09585_, _09526_, _02303_);
  and (_09586_, _09585_, _01538_);
  and (_09587_, _09586_, _09584_);
  and (_09588_, _04264_, _03722_);
  or (_09589_, _09588_, _09518_);
  and (_09590_, _09589_, _01537_);
  or (_09591_, _09590_, _38088_);
  or (_09592_, _09591_, _09587_);
  and (_37157_, _09592_, _09516_);
  or (_09593_, _38087_, \oc8051_golden_model_1.TL0 [7]);
  and (_09594_, _09593_, _37580_);
  not (_09595_, _03730_);
  and (_09596_, _09595_, \oc8051_golden_model_1.TL0 [7]);
  and (_09597_, _04779_, _03730_);
  or (_09598_, _09597_, _09596_);
  and (_09599_, _09598_, _02167_);
  and (_09600_, _04496_, _03730_);
  or (_09601_, _09600_, _09596_);
  or (_09602_, _09601_, _02814_);
  and (_09603_, _03730_, \oc8051_golden_model_1.ACC [7]);
  or (_09604_, _09603_, _09596_);
  and (_09605_, _09604_, _02817_);
  and (_09606_, _02818_, \oc8051_golden_model_1.TL0 [7]);
  or (_09607_, _09606_, _02001_);
  or (_09608_, _09607_, _09605_);
  and (_09609_, _09608_, _02840_);
  and (_09610_, _09609_, _09602_);
  nor (_09611_, _09595_, _03616_);
  or (_09612_, _09611_, _09596_);
  and (_09613_, _09612_, _01999_);
  or (_09614_, _09613_, _09610_);
  and (_09615_, _09614_, _02021_);
  and (_09616_, _09604_, _02006_);
  or (_09617_, _09616_, _05994_);
  or (_09618_, _09617_, _09615_);
  or (_09619_, _09612_, _05249_);
  and (_09620_, _09619_, _09618_);
  or (_09621_, _09620_, _02528_);
  and (_09622_, _04483_, _03730_);
  or (_09623_, _09596_, _02888_);
  or (_09624_, _09623_, _09622_);
  and (_09625_, _09624_, _02043_);
  and (_09626_, _09625_, _09621_);
  nor (_09627_, _04753_, _09595_);
  or (_09628_, _09627_, _09596_);
  and (_09629_, _09628_, _01602_);
  or (_09630_, _09629_, _01869_);
  or (_09631_, _09630_, _09626_);
  and (_09632_, _04560_, _03730_);
  or (_09633_, _09632_, _09596_);
  or (_09634_, _09633_, _01870_);
  and (_09635_, _09634_, _09631_);
  or (_09636_, _09635_, _02079_);
  and (_09637_, _04771_, _03730_);
  or (_09638_, _09596_, _02166_);
  or (_09639_, _09638_, _09637_);
  and (_09640_, _09639_, _02912_);
  and (_09641_, _09640_, _09636_);
  or (_09642_, _09641_, _09599_);
  and (_09643_, _09642_, _02176_);
  or (_09644_, _09596_, _03755_);
  and (_09645_, _09633_, _02072_);
  and (_09646_, _09645_, _09644_);
  or (_09647_, _09646_, _09643_);
  and (_09648_, _09647_, _02907_);
  and (_09649_, _09604_, _02177_);
  and (_09650_, _09649_, _09644_);
  or (_09651_, _09650_, _02071_);
  or (_09652_, _09651_, _09648_);
  nor (_09653_, _04770_, _09595_);
  or (_09654_, _09596_, _04788_);
  or (_09655_, _09654_, _09653_);
  and (_09656_, _09655_, _04793_);
  and (_09657_, _09656_, _09652_);
  nor (_09658_, _04778_, _09595_);
  or (_09659_, _09658_, _09596_);
  and (_09660_, _09659_, _02173_);
  or (_09661_, _09660_, _02201_);
  or (_09662_, _09661_, _09657_);
  or (_09663_, _09601_, _02303_);
  and (_09664_, _09663_, _01538_);
  and (_09665_, _09664_, _09662_);
  and (_09666_, _04264_, _03730_);
  or (_09667_, _09666_, _09596_);
  and (_09668_, _09667_, _01537_);
  or (_09669_, _09668_, _38088_);
  or (_09670_, _09669_, _09665_);
  and (_37158_, _09670_, _09594_);
  or (_09671_, _38087_, \oc8051_golden_model_1.TL1 [7]);
  and (_09672_, _09671_, _37580_);
  not (_09673_, _03708_);
  and (_09674_, _09673_, \oc8051_golden_model_1.TL1 [7]);
  and (_09675_, _04779_, _03845_);
  or (_09676_, _09675_, _09674_);
  and (_09677_, _09676_, _02167_);
  not (_09678_, _03845_);
  nor (_09679_, _09678_, _03616_);
  or (_09680_, _09679_, _09674_);
  or (_09681_, _09680_, _05249_);
  and (_09682_, _04496_, _03845_);
  or (_09683_, _09682_, _09674_);
  or (_09684_, _09683_, _02814_);
  and (_09685_, _03708_, \oc8051_golden_model_1.ACC [7]);
  or (_09686_, _09685_, _09674_);
  and (_09687_, _09686_, _02817_);
  and (_09688_, _02818_, \oc8051_golden_model_1.TL1 [7]);
  or (_09689_, _09688_, _02001_);
  or (_09690_, _09689_, _09687_);
  and (_09691_, _09690_, _02840_);
  and (_09692_, _09691_, _09684_);
  and (_09693_, _09680_, _01999_);
  or (_09694_, _09693_, _09692_);
  and (_09695_, _09694_, _02021_);
  and (_09696_, _09686_, _02006_);
  or (_09697_, _09696_, _05994_);
  or (_09698_, _09697_, _09695_);
  and (_09699_, _09698_, _09681_);
  or (_09700_, _09699_, _02528_);
  or (_09701_, _09674_, _02888_);
  and (_09702_, _04483_, _03708_);
  or (_09703_, _09702_, _09701_);
  and (_09704_, _09703_, _02043_);
  and (_09705_, _09704_, _09700_);
  nor (_09706_, _04753_, _09673_);
  or (_09707_, _09706_, _09674_);
  and (_09708_, _09707_, _01602_);
  or (_09709_, _09708_, _01869_);
  or (_09710_, _09709_, _09705_);
  and (_09711_, _04560_, _03708_);
  or (_09712_, _09711_, _09674_);
  or (_09713_, _09712_, _01870_);
  and (_09714_, _09713_, _09710_);
  or (_09715_, _09714_, _02079_);
  and (_09716_, _04771_, _03845_);
  or (_09717_, _09674_, _02166_);
  or (_09718_, _09717_, _09716_);
  and (_09719_, _09718_, _02912_);
  and (_09720_, _09719_, _09715_);
  or (_09721_, _09720_, _09677_);
  and (_09722_, _09721_, _02176_);
  or (_09723_, _09674_, _03755_);
  and (_09724_, _09712_, _02072_);
  and (_09725_, _09724_, _09723_);
  or (_09726_, _09725_, _09722_);
  and (_09727_, _09726_, _02907_);
  and (_09728_, _09686_, _02177_);
  and (_09729_, _09728_, _09723_);
  or (_09730_, _09729_, _02071_);
  or (_09731_, _09730_, _09727_);
  nor (_09732_, _04770_, _09678_);
  or (_09733_, _09674_, _04788_);
  or (_09734_, _09733_, _09732_);
  and (_09735_, _09734_, _04793_);
  and (_09736_, _09735_, _09731_);
  nor (_09737_, _04778_, _09678_);
  or (_09738_, _09737_, _09674_);
  and (_09739_, _09738_, _02173_);
  or (_09740_, _09739_, _02201_);
  or (_09741_, _09740_, _09736_);
  or (_09742_, _09683_, _02303_);
  and (_09743_, _09742_, _01538_);
  and (_09744_, _09743_, _09741_);
  and (_09745_, _04264_, _03845_);
  or (_09746_, _09745_, _09674_);
  and (_09747_, _09746_, _01537_);
  or (_09748_, _09747_, _38088_);
  or (_09749_, _09748_, _09744_);
  and (_37159_, _09749_, _09672_);
  or (_09750_, _38087_, \oc8051_golden_model_1.TMOD [7]);
  and (_09751_, _09750_, _37580_);
  not (_09752_, _03726_);
  and (_09753_, _09752_, \oc8051_golden_model_1.TMOD [7]);
  and (_09754_, _04779_, _03726_);
  or (_09755_, _09754_, _09753_);
  and (_09756_, _09755_, _02167_);
  nor (_09757_, _09752_, _03616_);
  or (_09758_, _09757_, _09753_);
  or (_09759_, _09758_, _05249_);
  and (_09760_, _04496_, _03726_);
  or (_09761_, _09760_, _09753_);
  or (_09762_, _09761_, _02814_);
  and (_09763_, _03726_, \oc8051_golden_model_1.ACC [7]);
  or (_09764_, _09763_, _09753_);
  and (_09765_, _09764_, _02817_);
  and (_09766_, _02818_, \oc8051_golden_model_1.TMOD [7]);
  or (_09767_, _09766_, _02001_);
  or (_09768_, _09767_, _09765_);
  and (_09769_, _09768_, _02840_);
  and (_09770_, _09769_, _09762_);
  and (_09771_, _09758_, _01999_);
  or (_09772_, _09771_, _09770_);
  and (_09773_, _09772_, _02021_);
  and (_09774_, _09764_, _02006_);
  or (_09775_, _09774_, _05994_);
  or (_09776_, _09775_, _09773_);
  and (_09777_, _09776_, _09759_);
  or (_09778_, _09777_, _02528_);
  and (_09779_, _04483_, _03726_);
  or (_09780_, _09753_, _02888_);
  or (_09781_, _09780_, _09779_);
  and (_09782_, _09781_, _02043_);
  and (_09783_, _09782_, _09778_);
  nor (_09784_, _04753_, _09752_);
  or (_09785_, _09784_, _09753_);
  and (_09786_, _09785_, _01602_);
  or (_09787_, _09786_, _01869_);
  or (_09788_, _09787_, _09783_);
  and (_09789_, _04560_, _03726_);
  or (_09790_, _09789_, _09753_);
  or (_09791_, _09790_, _01870_);
  and (_09792_, _09791_, _09788_);
  or (_09793_, _09792_, _02079_);
  and (_09794_, _04771_, _03726_);
  or (_09795_, _09753_, _02166_);
  or (_09796_, _09795_, _09794_);
  and (_09797_, _09796_, _02912_);
  and (_09798_, _09797_, _09793_);
  or (_09799_, _09798_, _09756_);
  and (_09800_, _09799_, _02176_);
  or (_09801_, _09753_, _03755_);
  and (_09802_, _09790_, _02072_);
  and (_09803_, _09802_, _09801_);
  or (_09804_, _09803_, _09800_);
  and (_09805_, _09804_, _02907_);
  and (_09806_, _09764_, _02177_);
  and (_09807_, _09806_, _09801_);
  or (_09808_, _09807_, _02071_);
  or (_09809_, _09808_, _09805_);
  nor (_09810_, _04770_, _09752_);
  or (_09811_, _09753_, _04788_);
  or (_09812_, _09811_, _09810_);
  and (_09813_, _09812_, _04793_);
  and (_09814_, _09813_, _09809_);
  nor (_09815_, _04778_, _09752_);
  or (_09816_, _09815_, _09753_);
  and (_09817_, _09816_, _02173_);
  or (_09818_, _09817_, _02201_);
  or (_09819_, _09818_, _09814_);
  or (_09820_, _09761_, _02303_);
  and (_09821_, _09820_, _01538_);
  and (_09822_, _09821_, _09819_);
  and (_09823_, _04264_, _03726_);
  or (_09824_, _09823_, _09753_);
  and (_09825_, _09824_, _01537_);
  or (_09826_, _09825_, _38088_);
  or (_09827_, _09826_, _09822_);
  and (_37160_, _09827_, _09751_);
  and (_09828_, _38088_, \oc8051_golden_model_1.PC [15]);
  and (_09829_, _01859_, _01403_);
  not (_09830_, _01267_);
  and (_09831_, _04268_, _09830_);
  and (_09832_, _09831_, \oc8051_golden_model_1.PC [6]);
  and (_09833_, _09832_, \oc8051_golden_model_1.PC [7]);
  and (_09834_, _09833_, \oc8051_golden_model_1.PC [8]);
  and (_09835_, _09834_, \oc8051_golden_model_1.PC [9]);
  and (_09836_, _09835_, \oc8051_golden_model_1.PC [10]);
  and (_09837_, _09836_, \oc8051_golden_model_1.PC [11]);
  and (_09838_, _09837_, \oc8051_golden_model_1.PC [12]);
  and (_09839_, _09838_, \oc8051_golden_model_1.PC [13]);
  and (_09840_, _09839_, \oc8051_golden_model_1.PC [14]);
  or (_09841_, _09840_, \oc8051_golden_model_1.PC [15]);
  nand (_09842_, _09840_, \oc8051_golden_model_1.PC [15]);
  and (_09843_, _09842_, _09841_);
  and (_09844_, _07212_, _06458_);
  or (_09845_, _09844_, _09843_);
  and (_09846_, _07116_, _07084_);
  or (_09847_, _09846_, _09843_);
  and (_09848_, _01859_, _01647_);
  not (_09849_, _09848_);
  nor (_09850_, _02173_, _01648_);
  or (_09851_, _09850_, _05212_);
  and (_09852_, _09851_, _09849_);
  nor (_09853_, _07069_, _02171_);
  not (_09854_, _09853_);
  not (_09855_, _06462_);
  nand (_09856_, _02049_, _01647_);
  and (_09857_, _09856_, _09855_);
  and (_09858_, _01977_, _01647_);
  not (_09859_, _09858_);
  and (_09860_, _09859_, _02730_);
  and (_09861_, _09860_, _09857_);
  or (_09862_, _09861_, _09843_);
  or (_09863_, _07031_, _07026_);
  not (_09864_, _09863_);
  or (_09865_, _09864_, _09843_);
  and (_09866_, _05228_, _01602_);
  not (_09867_, _08628_);
  and (_09868_, _05212_, _02006_);
  and (_09869_, _02008_, _01558_);
  or (_09870_, _09869_, _05212_);
  nor (_09871_, _08516_, _06636_);
  and (_09872_, _03862_, _03754_);
  and (_09873_, _09872_, _04487_);
  and (_09874_, _04106_, _04057_);
  and (_09875_, _04490_, _09874_);
  nand (_09876_, _09875_, _09873_);
  or (_09877_, _09876_, _05228_);
  nor (_09878_, _05217_, \oc8051_golden_model_1.PC [14]);
  nor (_09879_, _09878_, _05218_);
  nand (_09880_, _09879_, _04560_);
  or (_09881_, _09879_, _04560_);
  and (_09882_, _09881_, _09880_);
  not (_09883_, \oc8051_golden_model_1.PC [13]);
  and (_09884_, \oc8051_golden_model_1.PC [11], \oc8051_golden_model_1.PC [10]);
  and (_09885_, _09884_, _05196_);
  and (_09886_, _09885_, _04271_);
  and (_09887_, _09886_, \oc8051_golden_model_1.PC [12]);
  nor (_09888_, _09887_, _09883_);
  and (_09889_, _09887_, _09883_);
  or (_09890_, _09889_, _09888_);
  not (_09891_, _09890_);
  nor (_09892_, _09891_, _04307_);
  and (_09893_, _09891_, _04307_);
  nor (_09894_, _05215_, \oc8051_golden_model_1.PC [12]);
  nor (_09895_, _09894_, _05216_);
  nand (_09896_, _09895_, _04560_);
  not (_09897_, \oc8051_golden_model_1.PC [11]);
  nor (_09898_, _05214_, _09897_);
  and (_09899_, _05214_, _09897_);
  or (_09900_, _09899_, _09898_);
  not (_09901_, _09900_);
  nor (_09902_, _09901_, _04307_);
  and (_09903_, _09901_, _04307_);
  nor (_09904_, _09903_, _09902_);
  nor (_09905_, _05221_, \oc8051_golden_model_1.PC [10]);
  nor (_09906_, _09905_, _05214_);
  and (_09907_, _09906_, _04560_);
  nor (_09908_, _09906_, _04560_);
  nor (_09909_, _09908_, _09907_);
  and (_09910_, _09909_, _09904_);
  nor (_09911_, _05220_, \oc8051_golden_model_1.PC [9]);
  nor (_09912_, _09911_, _05221_);
  not (_09913_, _09912_);
  nor (_09914_, _09913_, _04307_);
  and (_09915_, _09913_, _04307_);
  nor (_09916_, _09915_, _09914_);
  not (_09917_, _09916_);
  nor (_09918_, _04307_, _04275_);
  and (_09919_, _04307_, _04275_);
  not (_09920_, _04594_);
  and (_09921_, _04267_, _04268_);
  nor (_09922_, _09921_, \oc8051_golden_model_1.PC [6]);
  nor (_09923_, _09922_, _04272_);
  nand (_09924_, _09923_, _09920_);
  or (_09925_, _09923_, _09920_);
  and (_09926_, _09925_, _09924_);
  and (_09927_, _04267_, \oc8051_golden_model_1.PC [4]);
  nor (_09928_, _09927_, \oc8051_golden_model_1.PC [5]);
  nor (_09929_, _09928_, _09921_);
  not (_09930_, _09929_);
  nor (_09931_, _09930_, _04626_);
  and (_09932_, _09930_, _04626_);
  nor (_09933_, _04267_, \oc8051_golden_model_1.PC [4]);
  nor (_09934_, _09933_, _09927_);
  nand (_09935_, _09934_, _04694_);
  nor (_09936_, _04266_, \oc8051_golden_model_1.PC [3]);
  nor (_09937_, _09936_, _04267_);
  not (_09938_, _09937_);
  nor (_09939_, _09938_, _02159_);
  and (_09940_, _09938_, _02159_);
  nor (_09941_, _01284_, \oc8051_golden_model_1.PC [2]);
  nor (_09942_, _09941_, _04266_);
  not (_09943_, _09942_);
  nor (_09944_, _09943_, _02338_);
  nor (_09945_, _02687_, _01723_);
  nor (_09946_, _02568_, \oc8051_golden_model_1.PC [0]);
  and (_09947_, _02687_, _01723_);
  nor (_09948_, _09947_, _09945_);
  and (_09949_, _09948_, _09946_);
  nor (_09950_, _09949_, _09945_);
  not (_09951_, _09950_);
  and (_09952_, _09943_, _02338_);
  nor (_09953_, _09952_, _09944_);
  and (_09954_, _09953_, _09951_);
  nor (_09955_, _09954_, _09944_);
  nor (_09956_, _09955_, _09940_);
  or (_09957_, _09956_, _09939_);
  or (_09958_, _09934_, _04694_);
  and (_09959_, _09958_, _09935_);
  nand (_09960_, _09959_, _09957_);
  and (_09961_, _09960_, _09935_);
  nor (_09962_, _09961_, _09932_);
  or (_09963_, _09962_, _09931_);
  nand (_09964_, _09963_, _09926_);
  and (_09965_, _09964_, _09924_);
  nor (_09966_, _09965_, _09919_);
  or (_09967_, _09966_, _09918_);
  nor (_09968_, _04271_, \oc8051_golden_model_1.PC [8]);
  nor (_09969_, _09968_, _05220_);
  and (_09970_, _09969_, _04560_);
  nor (_09971_, _09969_, _04560_);
  nor (_09972_, _09971_, _09970_);
  nand (_09973_, _09972_, _09967_);
  nor (_09974_, _09973_, _09917_);
  and (_09975_, _09974_, _09910_);
  or (_09976_, _09970_, _09914_);
  and (_09977_, _09976_, _09910_);
  or (_09978_, _09907_, _09902_);
  or (_09979_, _09978_, _09977_);
  or (_09980_, _09979_, _09975_);
  or (_09981_, _09895_, _04560_);
  and (_09982_, _09981_, _09896_);
  nand (_09983_, _09982_, _09980_);
  and (_09984_, _09983_, _09896_);
  nor (_09985_, _09984_, _09893_);
  or (_09986_, _09985_, _09892_);
  nand (_09987_, _09986_, _09882_);
  and (_09988_, _09987_, _09880_);
  not (_09989_, _05228_);
  and (_09990_, _09989_, _04307_);
  nor (_09991_, _09989_, _04307_);
  nor (_09992_, _09991_, _09990_);
  and (_09993_, _09992_, _09988_);
  nor (_09994_, _09992_, _09988_);
  or (_09995_, _09994_, _09993_);
  and (_09996_, _09875_, _09873_);
  or (_09997_, _09996_, _09995_);
  and (_09998_, _09997_, _02001_);
  and (_09999_, _09998_, _09877_);
  nor (_10000_, _05201_, \oc8051_golden_model_1.PC [14]);
  nor (_10001_, _10000_, _05202_);
  nand (_10002_, _10001_, _01790_);
  or (_10003_, _10001_, _01790_);
  and (_10004_, _10003_, _10002_);
  and (_10005_, _09885_, _04385_);
  and (_10006_, _10005_, \oc8051_golden_model_1.PC [12]);
  nor (_10007_, _10006_, _09883_);
  and (_10008_, _10006_, _09883_);
  or (_10009_, _10008_, _10007_);
  and (_10010_, _10009_, _01790_);
  nor (_10011_, _10009_, _01790_);
  nor (_10012_, _05199_, \oc8051_golden_model_1.PC [12]);
  nor (_10013_, _10012_, _05200_);
  nand (_10014_, _10013_, _01790_);
  nor (_10015_, _05198_, _09897_);
  and (_10016_, _05198_, _09897_);
  or (_10017_, _10016_, _10015_);
  and (_10018_, _10017_, _01790_);
  nor (_10019_, _10017_, _01790_);
  nor (_10020_, _05205_, \oc8051_golden_model_1.PC [10]);
  nor (_10021_, _10020_, _05198_);
  nand (_10022_, _10021_, _01790_);
  or (_10023_, _10021_, _01790_);
  and (_10024_, _10023_, _10022_);
  nor (_10025_, _05204_, \oc8051_golden_model_1.PC [9]);
  nor (_10026_, _10025_, _05205_);
  and (_10027_, _10026_, _01790_);
  nor (_10028_, _10026_, _01790_);
  nor (_10029_, _04385_, \oc8051_golden_model_1.PC [8]);
  nor (_10030_, _10029_, _05204_);
  nand (_10031_, _10030_, _01790_);
  and (_10032_, _04387_, _01790_);
  nor (_10033_, _04387_, _01790_);
  and (_10034_, _04268_, _01680_);
  nor (_10035_, _10034_, \oc8051_golden_model_1.PC [6]);
  nor (_10036_, _10035_, _04384_);
  not (_10037_, _10036_);
  or (_10038_, _10037_, _01922_);
  nand (_10039_, _10037_, _01922_);
  and (_10040_, _10039_, _10038_);
  and (_10041_, _01680_, \oc8051_golden_model_1.PC [4]);
  nor (_10042_, _10041_, \oc8051_golden_model_1.PC [5]);
  nor (_10043_, _10042_, _10034_);
  not (_10044_, _10043_);
  nor (_10045_, _10044_, _02252_);
  and (_10046_, _10044_, _02252_);
  nor (_10047_, _01680_, \oc8051_golden_model_1.PC [4]);
  nor (_10048_, _10047_, _10041_);
  not (_10049_, _10048_);
  or (_10050_, _10049_, _01855_);
  nor (_10051_, _01954_, _01683_);
  and (_10052_, _01954_, _01683_);
  nor (_10053_, _02294_, _01554_);
  nor (_10054_, _01822_, \oc8051_golden_model_1.PC [1]);
  nor (_10055_, _02441_, _01280_);
  and (_10056_, _01822_, \oc8051_golden_model_1.PC [1]);
  nor (_10057_, _10056_, _10054_);
  and (_10058_, _10057_, _10055_);
  nor (_10059_, _10058_, _10054_);
  not (_10060_, _10059_);
  and (_10061_, _02294_, _01554_);
  nor (_10062_, _10061_, _10053_);
  and (_10063_, _10062_, _10060_);
  nor (_10064_, _10063_, _10053_);
  nor (_10065_, _10064_, _10052_);
  or (_10066_, _10065_, _10051_);
  nand (_10067_, _10049_, _01855_);
  and (_10068_, _10067_, _10050_);
  nand (_10069_, _10068_, _10066_);
  and (_10070_, _10069_, _10050_);
  nor (_10071_, _10070_, _10046_);
  or (_10072_, _10071_, _10045_);
  nand (_10073_, _10072_, _10040_);
  and (_10074_, _10073_, _10038_);
  nor (_10075_, _10074_, _10033_);
  or (_10076_, _10075_, _10032_);
  or (_10077_, _10030_, _01790_);
  and (_10078_, _10077_, _10031_);
  nand (_10079_, _10078_, _10076_);
  and (_10080_, _10079_, _10031_);
  nor (_10081_, _10080_, _10028_);
  or (_10082_, _10081_, _10027_);
  nand (_10083_, _10082_, _10024_);
  and (_10084_, _10083_, _10022_);
  nor (_10085_, _10084_, _10019_);
  or (_10086_, _10085_, _10018_);
  or (_10087_, _10013_, _01790_);
  and (_10088_, _10087_, _10014_);
  nand (_10089_, _10088_, _10086_);
  and (_10090_, _10089_, _10014_);
  nor (_10091_, _10090_, _10011_);
  or (_10092_, _10091_, _10010_);
  nand (_10093_, _10092_, _10004_);
  and (_10094_, _10093_, _10002_);
  nor (_10095_, _05212_, _01790_);
  and (_10096_, _05212_, _01790_);
  nor (_10097_, _10096_, _10095_);
  and (_10098_, _10097_, _10094_);
  nor (_10099_, _10097_, _10094_);
  or (_10100_, _10099_, _10098_);
  and (_10101_, _04373_, _04371_);
  and (_10102_, _03028_, _02811_);
  and (_10103_, _03808_, _03616_);
  and (_10104_, _10103_, _10102_);
  nand (_10105_, _10104_, _10101_);
  and (_10106_, _10105_, _10100_);
  and (_10107_, _10104_, _10101_);
  and (_10108_, _10107_, _05212_);
  or (_10109_, _10108_, _04381_);
  or (_10110_, _10109_, _10106_);
  nor (_10111_, _01882_, _01533_);
  nor (_10112_, _10111_, _01561_);
  not (_10113_, _10112_);
  or (_10114_, _10113_, _09843_);
  or (_10115_, _10112_, \oc8051_golden_model_1.PC [15]);
  and (_10116_, _10115_, _02818_);
  and (_10117_, _10116_, _10114_);
  and (_10118_, _05212_, _02817_);
  or (_10119_, _10118_, _06625_);
  or (_10120_, _10119_, _10117_);
  not (_10121_, _06625_);
  or (_10122_, _09843_, _10121_);
  and (_10123_, _10122_, _01562_);
  and (_10124_, _10123_, _10120_);
  or (_10125_, _06629_, _02823_);
  or (_10126_, _06629_, _05212_);
  and (_10127_, _10126_, _10125_);
  or (_10128_, _10127_, _10124_);
  not (_10129_, _06629_);
  or (_10130_, _09843_, _10129_);
  and (_10131_, _10130_, _06618_);
  and (_10132_, _10131_, _10128_);
  and (_10133_, _05212_, _02003_);
  or (_10134_, _10133_, _06616_);
  or (_10135_, _10134_, _10132_);
  not (_10136_, _06616_);
  or (_10137_, _09843_, _10136_);
  and (_10138_, _10137_, _01568_);
  and (_10139_, _10138_, _10135_);
  not (_10140_, _01568_);
  and (_10141_, _05212_, _10140_);
  or (_10142_, _10141_, _04380_);
  or (_10143_, _10142_, _10139_);
  nor (_10144_, _02001_, _01883_);
  and (_10145_, _10144_, _10143_);
  and (_10146_, _10145_, _10110_);
  or (_10147_, _10146_, _09999_);
  and (_10148_, _10147_, _09871_);
  not (_10149_, _09869_);
  and (_10150_, _09871_, _04394_);
  not (_10151_, _10150_);
  and (_10152_, _10151_, _09843_);
  or (_10153_, _10152_, _10149_);
  or (_10154_, _10153_, _10148_);
  and (_10155_, _10154_, _09870_);
  and (_10156_, _06613_, _06675_);
  not (_10157_, _10156_);
  or (_10158_, _10157_, _10155_);
  or (_10159_, _10156_, _09843_);
  and (_10160_, _10159_, _02021_);
  and (_10161_, _10160_, _10158_);
  or (_10162_, _10161_, _09868_);
  nor (_10163_, _08529_, _06679_);
  and (_10164_, _10163_, _10162_);
  not (_10165_, _10163_);
  nand (_10166_, _10165_, _09843_);
  not (_10167_, _01574_);
  nor (_10168_, _01878_, _10167_);
  and (_10169_, _10168_, _02025_);
  nand (_10170_, _10169_, _10166_);
  or (_10171_, _10170_, _10164_);
  or (_10172_, _10169_, _05212_);
  and (_10173_, _10172_, _10171_);
  or (_10174_, _10173_, _08539_);
  or (_10175_, _09995_, _08572_);
  nand (_10176_, _08572_, _09989_);
  and (_10177_, _10176_, _10175_);
  or (_10178_, _10177_, _08538_);
  and (_10179_, _10178_, _10174_);
  or (_10180_, _10179_, _08493_);
  nand (_10181_, _08498_, _09989_);
  or (_10182_, _09995_, _08498_);
  and (_10183_, _10182_, _10181_);
  or (_10184_, _10183_, _08494_);
  and (_10185_, _10184_, _10180_);
  and (_10186_, _10185_, _08441_);
  nand (_10187_, _08625_, _09989_);
  or (_10188_, _09995_, _08625_);
  and (_10189_, _10188_, _01995_);
  and (_10190_, _10189_, _10187_);
  or (_10191_, _09995_, _08664_);
  nand (_10192_, _08664_, _09989_);
  and (_10193_, _10192_, _02045_);
  and (_10194_, _10193_, _10191_);
  or (_10195_, _10194_, _10190_);
  or (_10196_, _10195_, _10186_);
  and (_10197_, _10196_, _09867_);
  nand (_10198_, _09843_, _08628_);
  nor (_10199_, _02871_, _03131_);
  and (_10200_, _10199_, _01993_);
  and (_10201_, _10200_, _01989_);
  nand (_10202_, _10201_, _10198_);
  or (_10203_, _10202_, _10197_);
  and (_10204_, _01965_, _01536_);
  not (_10205_, _10204_);
  nor (_10206_, _07416_, _05279_);
  and (_10207_, _10206_, _10205_);
  or (_10208_, _10201_, _05212_);
  and (_10209_, _10208_, _10207_);
  and (_10210_, _10209_, _10203_);
  not (_10211_, _10207_);
  and (_10212_, _10211_, _09843_);
  not (_10213_, _01572_);
  nor (_10214_, _01966_, _10213_);
  and (_10215_, _10214_, _08249_);
  not (_10216_, _10215_);
  or (_10217_, _10216_, _10212_);
  or (_10218_, _10217_, _10210_);
  nor (_10219_, _10111_, _02372_);
  not (_10220_, _10219_);
  or (_10221_, _10215_, _05212_);
  and (_10222_, _10221_, _10220_);
  and (_10223_, _10222_, _10218_);
  and (_10224_, _10219_, _09843_);
  or (_10225_, _10224_, _06776_);
  or (_10226_, _10225_, _10223_);
  or (_10227_, _06775_, _05212_);
  and (_10228_, _10227_, _01550_);
  and (_10229_, _10228_, _10226_);
  and (_10230_, _09843_, _01549_);
  nor (_10231_, _01875_, _01604_);
  not (_10232_, _10231_);
  or (_10233_, _10232_, _10230_);
  or (_10234_, _10233_, _10229_);
  or (_10235_, _10231_, _05212_);
  and (_10236_, _10235_, _07401_);
  and (_10237_, _10236_, _10234_);
  nand (_10238_, _05228_, _02080_);
  nand (_10239_, _10238_, _09211_);
  or (_10240_, _10239_, _10237_);
  or (_10241_, _09211_, _05212_);
  and (_10242_, _10241_, _02043_);
  and (_10243_, _10242_, _10240_);
  or (_10244_, _10243_, _09866_);
  nor (_10245_, _06008_, _01608_);
  and (_10246_, _10245_, _10244_);
  nor (_10247_, _01959_, _01649_);
  not (_10248_, _10247_);
  not (_10249_, _10245_);
  and (_10250_, _10249_, _09843_);
  or (_10251_, _10250_, _10248_);
  or (_10252_, _10251_, _10246_);
  and (_10253_, _01859_, _01601_);
  not (_10254_, _10253_);
  or (_10255_, _10247_, _05212_);
  and (_10256_, _10255_, _10254_);
  and (_10257_, _10256_, _10252_);
  and (_10258_, _10253_, _10100_);
  or (_10259_, _10258_, _04758_);
  or (_10260_, _10259_, _10257_);
  or (_10261_, _05212_, _04757_);
  and (_10262_, _10261_, _01870_);
  and (_10263_, _10262_, _10260_);
  and (_10264_, _05228_, _01869_);
  or (_10265_, _10264_, _06984_);
  or (_10266_, _10265_, _10263_);
  and (_10267_, _01637_, _01543_);
  not (_10268_, _10267_);
  or (_10269_, _06985_, _05212_);
  and (_10270_, _10269_, _10268_);
  and (_10271_, _10270_, _10266_);
  not (_10272_, \oc8051_golden_model_1.DPH [6]);
  and (_10273_, \oc8051_golden_model_1.DPL [7], \oc8051_golden_model_1.ACC [7]);
  nor (_10274_, \oc8051_golden_model_1.DPL [7], \oc8051_golden_model_1.ACC [7]);
  nand (_10275_, \oc8051_golden_model_1.DPL [6], \oc8051_golden_model_1.ACC [6]);
  or (_10276_, \oc8051_golden_model_1.DPL [6], \oc8051_golden_model_1.ACC [6]);
  and (_10277_, _10276_, _10275_);
  and (_10278_, \oc8051_golden_model_1.DPL [5], \oc8051_golden_model_1.ACC [5]);
  nor (_10279_, \oc8051_golden_model_1.DPL [5], \oc8051_golden_model_1.ACC [5]);
  nor (_10280_, _10279_, _10278_);
  and (_10281_, \oc8051_golden_model_1.DPL [4], \oc8051_golden_model_1.ACC [4]);
  nor (_10282_, _01669_, _01665_);
  not (_10283_, _10282_);
  nor (_10284_, \oc8051_golden_model_1.DPL [4], \oc8051_golden_model_1.ACC [4]);
  nor (_10285_, _10284_, _10281_);
  and (_10286_, _10285_, _10283_);
  nor (_10287_, _10286_, _10281_);
  not (_10288_, _10287_);
  and (_10289_, _10288_, _10280_);
  or (_10290_, _10289_, _10278_);
  nand (_10291_, _10290_, _10277_);
  and (_10292_, _10291_, _10275_);
  nor (_10293_, _10292_, _10274_);
  or (_10294_, _10293_, _10273_);
  and (_10295_, _10294_, \oc8051_golden_model_1.DPH [0]);
  and (_10296_, _10295_, \oc8051_golden_model_1.DPH [1]);
  and (_10297_, _10296_, \oc8051_golden_model_1.DPH [2]);
  and (_10298_, _10297_, \oc8051_golden_model_1.DPH [3]);
  and (_10299_, _10298_, \oc8051_golden_model_1.DPH [4]);
  nand (_10300_, _10299_, \oc8051_golden_model_1.DPH [5]);
  nor (_10301_, _10300_, _10272_);
  or (_10302_, _10301_, \oc8051_golden_model_1.DPH [7]);
  nand (_10303_, _10301_, \oc8051_golden_model_1.DPH [7]);
  and (_10304_, _10303_, _10302_);
  and (_10305_, _10304_, _10267_);
  nor (_10306_, _01958_, _01638_);
  not (_10307_, _10306_);
  or (_10308_, _10307_, _10305_);
  or (_10309_, _10308_, _10271_);
  and (_10310_, _01859_, _01637_);
  not (_10311_, _10310_);
  or (_10312_, _10306_, _05212_);
  and (_10313_, _10312_, _10311_);
  and (_10314_, _10313_, _10309_);
  or (_10315_, _10100_, _07356_);
  not (_10316_, _07356_);
  or (_10317_, _10316_, _05212_);
  and (_10318_, _10317_, _10310_);
  and (_10319_, _10318_, _10315_);
  or (_10320_, _10319_, _10314_);
  or (_10321_, _02690_, _01978_);
  and (_10322_, _10321_, _01644_);
  nor (_10323_, _10322_, _06990_);
  nor (_10324_, _05242_, _02371_);
  not (_10325_, _10324_);
  and (_10326_, _10325_, _10323_);
  and (_10327_, _10326_, _07006_);
  and (_10328_, _10327_, _10320_);
  nor (_10329_, _07012_, _02168_);
  not (_10330_, _10329_);
  not (_10331_, _10327_);
  and (_10332_, _10331_, _09843_);
  or (_10333_, _10332_, _10330_);
  or (_10334_, _10333_, _10328_);
  or (_10335_, _10329_, _05212_);
  and (_10336_, _10335_, _02166_);
  and (_10337_, _10336_, _10334_);
  and (_10338_, _05228_, _02079_);
  nor (_10339_, _02167_, _01645_);
  not (_10340_, _10339_);
  or (_10341_, _10340_, _10338_);
  or (_10342_, _10341_, _10337_);
  and (_10343_, _01859_, _01644_);
  not (_10344_, _10343_);
  or (_10345_, _10339_, _05212_);
  and (_10346_, _10345_, _10344_);
  and (_10347_, _10346_, _10342_);
  or (_10348_, _10100_, _10316_);
  or (_10349_, _07356_, _05212_);
  and (_10350_, _10349_, _10343_);
  and (_10351_, _10350_, _10348_);
  or (_10352_, _09863_, _10351_);
  or (_10353_, _10352_, _10347_);
  and (_10354_, _10353_, _09865_);
  or (_10355_, _10354_, _07042_);
  or (_10356_, _07041_, _05212_);
  and (_10357_, _10356_, _02176_);
  and (_10358_, _10357_, _10355_);
  not (_10359_, _09292_);
  and (_10360_, _05228_, _02072_);
  or (_10361_, _10360_, _10359_);
  or (_10362_, _10361_, _10358_);
  and (_10363_, _01859_, _01631_);
  not (_10364_, _10363_);
  or (_10365_, _09292_, _05212_);
  and (_10366_, _10365_, _10364_);
  and (_10367_, _10366_, _10362_);
  not (_10368_, _09861_);
  or (_10369_, _10100_, \oc8051_golden_model_1.PSW [7]);
  or (_10370_, _05212_, _06518_);
  and (_10371_, _10370_, _10363_);
  and (_10372_, _10371_, _10369_);
  or (_10373_, _10372_, _10368_);
  or (_10374_, _10373_, _10367_);
  and (_10375_, _10374_, _09862_);
  or (_10376_, _10375_, _09854_);
  or (_10377_, _09853_, _05212_);
  and (_10378_, _10377_, _04788_);
  and (_10379_, _10378_, _10376_);
  not (_10380_, _09850_);
  and (_10381_, _05228_, _02071_);
  or (_10382_, _10381_, _10380_);
  or (_10383_, _10382_, _10379_);
  and (_10384_, _10383_, _09852_);
  not (_10385_, _09846_);
  or (_10386_, _10100_, _06518_);
  or (_10387_, _05212_, \oc8051_golden_model_1.PSW [7]);
  and (_10388_, _10387_, _09848_);
  and (_10389_, _10388_, _10386_);
  or (_10390_, _10389_, _10385_);
  or (_10391_, _10390_, _10384_);
  and (_10392_, _10391_, _09847_);
  or (_10393_, _10392_, _07146_);
  or (_10394_, _07145_, _05212_);
  and (_10395_, _10394_, _07176_);
  and (_10396_, _10395_, _10393_);
  and (_10397_, _09843_, _07175_);
  or (_10398_, _10397_, _02185_);
  or (_10399_, _10398_, _10396_);
  nand (_10400_, _03616_, _02185_);
  and (_10401_, _10400_, _10399_);
  or (_10402_, _10401_, _01636_);
  not (_10403_, _02083_);
  or (_10404_, _05212_, _04799_);
  and (_10405_, _10404_, _10403_);
  and (_10406_, _10405_, _10402_);
  not (_10407_, _09844_);
  not (_10408_, _08439_);
  or (_10409_, _09995_, _10408_);
  or (_10410_, _08439_, _05228_);
  and (_10411_, _10410_, _02083_);
  and (_10412_, _10411_, _10409_);
  or (_10413_, _10412_, _10407_);
  or (_10414_, _10413_, _10406_);
  and (_10415_, _10414_, _09845_);
  or (_10416_, _10415_, _07255_);
  or (_10417_, _07254_, _05212_);
  and (_10418_, _10417_, _07305_);
  and (_10419_, _10418_, _10416_);
  and (_10420_, _09843_, _07304_);
  or (_10421_, _10420_, _01888_);
  or (_10422_, _10421_, _10419_);
  nand (_10423_, _03616_, _01888_);
  and (_10424_, _10423_, _10422_);
  or (_10425_, _10424_, _01653_);
  not (_10426_, _01653_);
  or (_10427_, _05212_, _10426_);
  and (_10428_, _10427_, _02202_);
  and (_10429_, _10428_, _10425_);
  or (_10430_, _09995_, _08439_);
  nand (_10431_, _08439_, _09989_);
  and (_10432_, _10431_, _10430_);
  and (_10433_, _10432_, _02082_);
  not (_10434_, _01641_);
  nor (_10435_, _10111_, _10434_);
  or (_10436_, _10435_, _10433_);
  or (_10437_, _10436_, _10429_);
  not (_10438_, _10435_);
  or (_10439_, _10438_, _09843_);
  and (_10440_, _10439_, _02303_);
  and (_10441_, _10440_, _10437_);
  nor (_10442_, _07350_, _07345_);
  not (_10443_, _10442_);
  and (_10444_, _05212_, _02201_);
  or (_10445_, _10444_, _10443_);
  or (_10446_, _10445_, _10441_);
  or (_10447_, _09843_, _10442_);
  and (_10448_, _10447_, _05195_);
  and (_10449_, _10448_, _10446_);
  and (_10450_, _02058_, _01790_);
  or (_10451_, _10450_, _01642_);
  or (_10452_, _10451_, _10449_);
  not (_10453_, _01642_);
  or (_10454_, _05212_, _10453_);
  and (_10455_, _10454_, _01887_);
  and (_10456_, _10455_, _10452_);
  and (_10457_, _10432_, _01860_);
  or (_10458_, _05171_, _02952_);
  or (_10459_, _10458_, _10457_);
  or (_10460_, _10459_, _10456_);
  not (_10461_, _10458_);
  or (_10462_, _10461_, _09843_);
  and (_10463_, _10462_, _01538_);
  and (_10464_, _10463_, _10460_);
  nor (_10465_, _07374_, _07367_);
  not (_10466_, _10465_);
  and (_10467_, _05212_, _01537_);
  or (_10468_, _10467_, _10466_);
  or (_10469_, _10468_, _10464_);
  not (_10470_, _02057_);
  or (_10471_, _09843_, _10465_);
  and (_10472_, _10471_, _10470_);
  and (_10473_, _10472_, _10469_);
  and (_10474_, _02057_, _01790_);
  or (_10475_, _10474_, _01651_);
  or (_10476_, _10475_, _10473_);
  not (_10477_, _01651_);
  or (_10478_, _05212_, _10477_);
  and (_10479_, _10478_, _10476_);
  or (_10480_, _10479_, _09829_);
  not (_10481_, _09829_);
  or (_10482_, _09843_, _10481_);
  and (_10483_, _10482_, _38087_);
  and (_10484_, _10483_, _10480_);
  or (_10485_, _10484_, _09828_);
  and (_37162_, _10485_, _37580_);
  and (_10486_, _38088_, \oc8051_golden_model_1.P0INREG [7]);
  or (_10487_, _10486_, _38465_);
  and (_37163_, _10487_, _37580_);
  and (_10488_, _38088_, \oc8051_golden_model_1.P1INREG [7]);
  or (_10489_, _10488_, _38240_);
  and (_37164_, _10489_, _37580_);
  and (_10490_, _38088_, \oc8051_golden_model_1.P2INREG [7]);
  or (_10491_, _10490_, _38199_);
  and (_37165_, _10491_, _37580_);
  and (_10492_, _38088_, \oc8051_golden_model_1.P3INREG [7]);
  or (_10493_, _10492_, _38420_);
  and (_37166_, _10493_, _37580_);
  nand (_10494_, _02058_, \oc8051_golden_model_1.PC [0]);
  and (_10495_, _04106_, _04562_);
  and (_10496_, _10495_, _02910_);
  or (_10497_, _03028_, _02887_);
  nand (_10498_, _06850_, _02503_);
  and (_10499_, _03028_, _02841_);
  or (_10500_, _04381_, _03042_);
  nor (_10501_, _01562_, _01280_);
  and (_10502_, _01562_, \oc8051_golden_model_1.ACC [0]);
  or (_10503_, _10502_, _10501_);
  nor (_10504_, _10503_, _04380_);
  nor (_10505_, _10504_, _02815_);
  and (_10506_, _10505_, _10500_);
  nor (_10507_, _04106_, _02816_);
  or (_10508_, _10507_, _10506_);
  and (_10509_, _10508_, _04366_);
  nand (_10510_, _08723_, _08334_);
  and (_10511_, _10510_, _02837_);
  or (_10512_, _10511_, _03279_);
  or (_10513_, _10512_, _10509_);
  nor (_10514_, _01558_, \oc8051_golden_model_1.PC [0]);
  nor (_10515_, _10514_, _02841_);
  and (_10516_, _10515_, _10513_);
  or (_10517_, _10516_, _10499_);
  and (_10518_, _10517_, _04353_);
  nor (_10519_, _08723_, _03628_);
  and (_10520_, _10519_, _02856_);
  or (_10521_, _10520_, _01878_);
  or (_10522_, _10521_, _10518_);
  nand (_10523_, _06850_, _01878_);
  and (_10524_, _10523_, _02962_);
  and (_10525_, _10524_, _10522_);
  nand (_10526_, _10510_, _02862_);
  nor (_10527_, _10526_, _08724_);
  or (_10528_, _10527_, _10525_);
  and (_10529_, _10528_, _01565_);
  or (_10530_, _01565_, _01280_);
  nand (_10531_, _01989_, _10530_);
  or (_10532_, _10531_, _10529_);
  and (_10533_, _10532_, _10498_);
  or (_10534_, _10533_, _02871_);
  and (_10535_, _04952_, _03673_);
  nand (_10536_, _06849_, _02871_);
  or (_10537_, _10536_, _10535_);
  and (_10538_, _10537_, _10534_);
  or (_10539_, _10538_, _02870_);
  nor (_10540_, _08357_, _03628_);
  and (_10541_, _03628_, \oc8051_golden_model_1.PSW [7]);
  nor (_10542_, _10541_, _10540_);
  nand (_10543_, _10542_, _02870_);
  and (_10544_, _10543_, _04310_);
  and (_10545_, _10544_, _10539_);
  nand (_10546_, _01604_, \oc8051_golden_model_1.PC [0]);
  nand (_10547_, _02887_, _10546_);
  or (_10548_, _10547_, _10545_);
  and (_10549_, _10548_, _10497_);
  or (_10550_, _10549_, _02889_);
  or (_10551_, _04952_, _02890_);
  and (_10552_, _10551_, _02880_);
  and (_10553_, _10552_, _10550_);
  and (_10554_, _04307_, _03028_);
  not (_10555_, _10554_);
  and (_10556_, _04662_, \oc8051_golden_model_1.TH1 [0]);
  and (_10557_, _04667_, \oc8051_golden_model_1.DPH [0]);
  nor (_10558_, _10557_, _10556_);
  and (_10559_, _04675_, \oc8051_golden_model_1.P2INREG [0]);
  not (_10560_, _10559_);
  and (_10561_, _04681_, \oc8051_golden_model_1.TMOD [0]);
  and (_10562_, _04686_, \oc8051_golden_model_1.TL0 [0]);
  nor (_10563_, _10562_, _10561_);
  and (_10564_, _10563_, _10560_);
  and (_10565_, _04691_, \oc8051_golden_model_1.IE [0]);
  not (_10566_, _10565_);
  and (_10567_, _04697_, \oc8051_golden_model_1.SCON [0]);
  and (_10568_, _04699_, \oc8051_golden_model_1.SBUF [0]);
  nor (_10569_, _10568_, _10567_);
  and (_10570_, _10569_, _10566_);
  and (_10571_, _04703_, \oc8051_golden_model_1.P0INREG [0]);
  not (_10572_, _10571_);
  and (_10573_, _04706_, \oc8051_golden_model_1.P1INREG [0]);
  and (_10574_, _04710_, \oc8051_golden_model_1.P3INREG [0]);
  nor (_10575_, _10574_, _10573_);
  and (_10576_, _10575_, _10572_);
  and (_10577_, _10576_, _10570_);
  and (_10578_, _10577_, _10564_);
  and (_10579_, _10578_, _10558_);
  and (_10580_, _04717_, \oc8051_golden_model_1.TH0 [0]);
  and (_10581_, _04719_, \oc8051_golden_model_1.TL1 [0]);
  nor (_10582_, _10581_, _10580_);
  and (_10583_, _04722_, \oc8051_golden_model_1.TCON [0]);
  and (_10584_, _04726_, \oc8051_golden_model_1.PCON [0]);
  nor (_10585_, _10584_, _10583_);
  and (_10586_, _10585_, _10582_);
  and (_10587_, _04730_, \oc8051_golden_model_1.IP [0]);
  and (_10588_, _04734_, \oc8051_golden_model_1.ACC [0]);
  nor (_10589_, _10588_, _10587_);
  and (_10590_, _04737_, \oc8051_golden_model_1.PSW [0]);
  and (_10591_, _04739_, \oc8051_golden_model_1.B [0]);
  nor (_10592_, _10591_, _10590_);
  and (_10593_, _10592_, _10589_);
  and (_10594_, _04744_, \oc8051_golden_model_1.DPL [0]);
  and (_10595_, _04746_, \oc8051_golden_model_1.SP [0]);
  nor (_10596_, _10595_, _10594_);
  and (_10597_, _10596_, _10593_);
  and (_10598_, _10597_, _10586_);
  and (_10599_, _10598_, _10579_);
  and (_10600_, _10599_, _10555_);
  nor (_10601_, _10600_, _02880_);
  or (_10602_, _10601_, _04758_);
  or (_10603_, _10602_, _10553_);
  and (_10604_, _04758_, _02441_);
  nor (_10605_, _10604_, _01871_);
  and (_10606_, _10605_, _10603_);
  and (_10607_, _04562_, _01871_);
  or (_10608_, _10607_, _01638_);
  or (_10609_, _10608_, _10606_);
  and (_10610_, _01638_, _01280_);
  nor (_10611_, _10610_, _02914_);
  and (_10612_, _10611_, _10609_);
  nor (_10613_, _04106_, _04562_);
  nor (_10614_, _10495_, _10613_);
  nor (_10615_, _10614_, _02913_);
  nor (_10616_, _10615_, _02915_);
  or (_10617_, _10616_, _10612_);
  and (_10618_, _04106_, \oc8051_golden_model_1.ACC [0]);
  nor (_10619_, _04106_, \oc8051_golden_model_1.ACC [0]);
  nor (_10620_, _10619_, _10618_);
  or (_10621_, _10620_, _04775_);
  and (_10622_, _10621_, _02911_);
  and (_10623_, _10622_, _10617_);
  or (_10624_, _10623_, _10496_);
  and (_10625_, _10624_, _02909_);
  and (_10626_, _10618_, _02908_);
  or (_10627_, _10626_, _01632_);
  or (_10628_, _10627_, _10625_);
  and (_10629_, _01632_, _01280_);
  nor (_10630_, _10629_, _04789_);
  and (_10631_, _10630_, _10628_);
  nor (_10632_, _10613_, _04795_);
  or (_10633_, _10632_, _04794_);
  or (_10634_, _10633_, _10631_);
  nand (_10635_, _10619_, _04794_);
  and (_10636_, _10635_, _10634_);
  or (_10637_, _10636_, _01636_);
  nand (_10638_, _01641_, _01533_);
  nand (_10639_, _01636_, _01280_);
  and (_10640_, _10639_, _10638_);
  and (_10641_, _10640_, _10637_);
  nor (_10642_, _10638_, _03028_);
  or (_10643_, _10642_, _02935_);
  or (_10644_, _10643_, _10641_);
  nand (_10645_, _04952_, _02935_);
  and (_10646_, _10645_, _04814_);
  and (_10647_, _10646_, _10644_);
  nor (_10648_, _04106_, _04814_);
  or (_10649_, _10648_, _02058_);
  or (_10650_, _10649_, _10647_);
  and (_10651_, _10650_, _10494_);
  or (_10652_, _10651_, _01642_);
  and (_10653_, _01642_, _01280_);
  nor (_10654_, _10653_, _02941_);
  and (_10655_, _10654_, _10652_);
  and (_10656_, _10540_, _02941_);
  or (_10657_, _10656_, _05171_);
  or (_10658_, _10657_, _10655_);
  nand (_10659_, _05171_, _03028_);
  and (_10660_, _10659_, _05178_);
  and (_10661_, _10660_, _10658_);
  nor (_10662_, _04952_, _05178_);
  or (_10663_, _10662_, _01791_);
  or (_10664_, _10663_, _10661_);
  nand (_10665_, _04106_, _01791_);
  and (_10666_, _10665_, _03186_);
  and (_10667_, _10666_, _10664_);
  nor (_10668_, _03187_, _02956_);
  nor (_10669_, _10668_, _03189_);
  nor (_10670_, _03386_, _03187_);
  nor (_10671_, _10670_, _03540_);
  and (_10672_, _10671_, _03186_);
  and (_10673_, _10672_, _10669_);
  not (_10674_, _10673_);
  or (_10675_, _10674_, _10667_);
  or (_10676_, _10673_, \oc8051_golden_model_1.IRAM[0] [0]);
  not (_10677_, _03557_);
  not (_10678_, _03548_);
  and (_10679_, _03556_, _10678_);
  and (_10680_, _10679_, _10677_);
  and (_10681_, _10680_, _01865_);
  not (_10682_, _10681_);
  and (_10683_, _10682_, _10676_);
  and (_10684_, _10683_, _10675_);
  not (_10685_, _10030_);
  nor (_10686_, _10685_, _02058_);
  and (_10687_, _09969_, _02058_);
  or (_10688_, _10687_, _10686_);
  and (_10689_, _10688_, _10681_);
  or (_37199_, _10689_, _10684_);
  nor (_10690_, _05179_, _04953_);
  or (_10691_, _10690_, _05178_);
  nor (_10692_, _04057_, _02687_);
  and (_10693_, _10692_, _02910_);
  or (_10694_, _02887_, _02812_);
  nand (_10695_, _06838_, _02503_);
  nor (_10696_, _08698_, _03619_);
  or (_10697_, _10696_, _04353_);
  nor (_10698_, _04489_, _04107_);
  nor (_10699_, _10698_, _02816_);
  nor (_10700_, _05161_, _04372_);
  nand (_10701_, _10700_, _04380_);
  nor (_10702_, _01562_, \oc8051_golden_model_1.PC [1]);
  and (_10703_, _01562_, \oc8051_golden_model_1.ACC [1]);
  or (_10704_, _10703_, _10702_);
  nor (_10705_, _10704_, _04380_);
  nor (_10706_, _10705_, _02815_);
  and (_10707_, _10706_, _10701_);
  or (_10708_, _10707_, _02837_);
  or (_10709_, _10708_, _10699_);
  nand (_10710_, _08698_, _08275_);
  or (_10711_, _10710_, _04366_);
  and (_10712_, _10711_, _10709_);
  or (_10713_, _10712_, _03279_);
  nor (_10714_, _01558_, _01253_);
  nor (_10715_, _10714_, _02841_);
  and (_10716_, _10715_, _10713_);
  and (_10717_, _02841_, _02812_);
  or (_10718_, _10717_, _02856_);
  or (_10719_, _10718_, _10716_);
  and (_10720_, _10719_, _10697_);
  or (_10721_, _10720_, _01878_);
  nand (_10722_, _06838_, _01878_);
  and (_10723_, _10722_, _02962_);
  and (_10724_, _10723_, _10721_);
  not (_10725_, _08699_);
  and (_10726_, _10710_, _10725_);
  and (_10727_, _10726_, _02862_);
  or (_10728_, _10727_, _10724_);
  and (_10729_, _10728_, _01565_);
  or (_10730_, _01565_, \oc8051_golden_model_1.PC [1]);
  nand (_10731_, _01989_, _10730_);
  or (_10732_, _10731_, _10729_);
  and (_10733_, _10732_, _10695_);
  or (_10734_, _10733_, _02871_);
  and (_10735_, _04907_, _03673_);
  nand (_10736_, _06837_, _02871_);
  or (_10737_, _10736_, _10735_);
  and (_10738_, _10737_, _10734_);
  or (_10739_, _10738_, _02870_);
  nor (_10740_, _08298_, _03619_);
  and (_10741_, _03619_, \oc8051_golden_model_1.PSW [7]);
  nor (_10742_, _10741_, _10740_);
  nand (_10743_, _10742_, _02870_);
  and (_10744_, _10743_, _04310_);
  and (_10745_, _10744_, _10739_);
  nand (_10746_, _01604_, _01253_);
  nand (_10747_, _02887_, _10746_);
  or (_10748_, _10747_, _10745_);
  and (_10749_, _10748_, _10694_);
  or (_10750_, _10749_, _02889_);
  or (_10751_, _04907_, _02890_);
  and (_10752_, _10751_, _02880_);
  and (_10753_, _10752_, _10750_);
  nor (_10754_, _04560_, _02811_);
  and (_10755_, _04722_, \oc8051_golden_model_1.TCON [1]);
  not (_10756_, _10755_);
  and (_10757_, _04734_, \oc8051_golden_model_1.ACC [1]);
  and (_10758_, _04737_, \oc8051_golden_model_1.PSW [1]);
  nor (_10759_, _10758_, _10757_);
  and (_10760_, _10759_, _10756_);
  and (_10761_, _04717_, \oc8051_golden_model_1.TH0 [1]);
  not (_10762_, _10761_);
  and (_10763_, _04730_, \oc8051_golden_model_1.IP [1]);
  and (_10764_, _04739_, \oc8051_golden_model_1.B [1]);
  nor (_10765_, _10764_, _10763_);
  and (_10766_, _10765_, _10762_);
  and (_10767_, _04726_, \oc8051_golden_model_1.PCON [1]);
  and (_10768_, _04719_, \oc8051_golden_model_1.TL1 [1]);
  nor (_10769_, _10768_, _10767_);
  and (_10770_, _10769_, _10766_);
  and (_10771_, _10770_, _10760_);
  and (_10772_, _04686_, \oc8051_golden_model_1.TL0 [1]);
  and (_10773_, _04662_, \oc8051_golden_model_1.TH1 [1]);
  nor (_10774_, _10773_, _10772_);
  and (_10775_, _04667_, \oc8051_golden_model_1.DPH [1]);
  not (_10776_, _10775_);
  and (_10777_, _10776_, _10774_);
  and (_10778_, _04703_, \oc8051_golden_model_1.P0INREG [1]);
  not (_10779_, _10778_);
  and (_10780_, _04706_, \oc8051_golden_model_1.P1INREG [1]);
  and (_10781_, _04710_, \oc8051_golden_model_1.P3INREG [1]);
  nor (_10782_, _10781_, _10780_);
  and (_10783_, _10782_, _10779_);
  and (_10784_, _04681_, \oc8051_golden_model_1.TMOD [1]);
  and (_10785_, _04675_, \oc8051_golden_model_1.P2INREG [1]);
  nor (_10786_, _10785_, _10784_);
  and (_10787_, _10786_, _10783_);
  and (_10788_, _04691_, \oc8051_golden_model_1.IE [1]);
  not (_10789_, _10788_);
  and (_10790_, _04697_, \oc8051_golden_model_1.SCON [1]);
  and (_10791_, _04699_, \oc8051_golden_model_1.SBUF [1]);
  nor (_10792_, _10791_, _10790_);
  and (_10793_, _10792_, _10789_);
  and (_10794_, _04744_, \oc8051_golden_model_1.DPL [1]);
  and (_10795_, _04746_, \oc8051_golden_model_1.SP [1]);
  nor (_10796_, _10795_, _10794_);
  and (_10797_, _10796_, _10793_);
  and (_10798_, _10797_, _10787_);
  and (_10799_, _10798_, _10777_);
  and (_10800_, _10799_, _10771_);
  not (_10801_, _10800_);
  nor (_10802_, _10801_, _10754_);
  nor (_10803_, _10802_, _02880_);
  or (_10804_, _10803_, _04758_);
  or (_10805_, _10804_, _10753_);
  and (_10806_, _04758_, _01822_);
  nor (_10807_, _10806_, _01871_);
  and (_10808_, _10807_, _10805_);
  and (_10809_, _04683_, _01871_);
  or (_10810_, _10809_, _01638_);
  or (_10811_, _10810_, _10808_);
  and (_10812_, _01638_, \oc8051_golden_model_1.PC [1]);
  nor (_10813_, _10812_, _02914_);
  and (_10814_, _10813_, _10811_);
  and (_10815_, _04057_, _02687_);
  nor (_10816_, _10815_, _10692_);
  nor (_10817_, _10816_, _02913_);
  nor (_10818_, _10817_, _02915_);
  or (_10819_, _10818_, _10814_);
  nor (_10820_, _04057_, _01613_);
  and (_10821_, _04057_, _01613_);
  nor (_10822_, _10821_, _10820_);
  or (_10823_, _10822_, _04775_);
  and (_10824_, _10823_, _02911_);
  and (_10825_, _10824_, _10819_);
  or (_10826_, _10825_, _10693_);
  and (_10827_, _10826_, _02909_);
  and (_10828_, _10820_, _02908_);
  or (_10829_, _10828_, _01632_);
  or (_10830_, _10829_, _10827_);
  and (_10831_, _01632_, \oc8051_golden_model_1.PC [1]);
  nor (_10832_, _10831_, _04789_);
  and (_10833_, _10832_, _10830_);
  nor (_10834_, _10815_, _04795_);
  or (_10835_, _10834_, _04794_);
  or (_10836_, _10835_, _10833_);
  nand (_10837_, _10821_, _04794_);
  and (_10838_, _10837_, _04799_);
  and (_10839_, _10838_, _10836_);
  and (_10840_, _01636_, _01253_);
  not (_10841_, _10638_);
  or (_10842_, _10841_, _10840_);
  or (_10843_, _10842_, _10839_);
  nand (_10844_, _10700_, _10841_);
  and (_10845_, _10844_, _04815_);
  and (_10846_, _10845_, _10843_);
  nor (_10847_, _10690_, _04815_);
  or (_10848_, _10847_, _10846_);
  and (_10849_, _10848_, _04814_);
  nor (_10850_, _10698_, _04814_);
  or (_10851_, _10850_, _02058_);
  or (_10852_, _10851_, _10849_);
  nand (_10853_, _02058_, _01723_);
  and (_10854_, _10853_, _10453_);
  and (_10855_, _10854_, _10852_);
  and (_10856_, _01642_, _01253_);
  or (_10857_, _02941_, _10856_);
  or (_10858_, _10857_, _10855_);
  or (_10859_, _10740_, _02958_);
  and (_10860_, _10859_, _05172_);
  and (_10861_, _10860_, _10858_);
  and (_10862_, _10700_, _05171_);
  or (_10863_, _10862_, _02952_);
  or (_10864_, _10863_, _10861_);
  and (_10865_, _10864_, _10691_);
  or (_10866_, _10865_, _01791_);
  or (_10867_, _10698_, _03118_);
  and (_10868_, _10867_, _03186_);
  and (_10869_, _10868_, _10866_);
  or (_10870_, _10869_, _10674_);
  or (_10871_, _10673_, \oc8051_golden_model_1.IRAM[0] [1]);
  and (_10872_, _10871_, _10682_);
  and (_10873_, _10872_, _10870_);
  and (_10874_, _09912_, _02058_);
  and (_10875_, _10026_, _05195_);
  or (_10876_, _10875_, _10874_);
  and (_10877_, _10876_, _10681_);
  or (_37200_, _10877_, _10873_);
  nor (_10878_, _10673_, _03397_);
  or (_10879_, _05161_, _03456_);
  nor (_10880_, _05172_, _06733_);
  and (_10881_, _10880_, _10879_);
  not (_10882_, _05043_);
  and (_10883_, _04953_, _10882_);
  nor (_10884_, _04953_, _10882_);
  or (_10885_, _10884_, _10883_);
  and (_10886_, _10885_, _02935_);
  and (_10887_, _04372_, _03455_);
  nor (_10888_, _04372_, _03455_);
  or (_10889_, _10888_, _10887_);
  or (_10890_, _10889_, _04804_);
  nor (_10891_, _04155_, _02338_);
  and (_10892_, _10891_, _02910_);
  or (_10893_, _03456_, _02887_);
  nor (_10894_, _08687_, _03855_);
  or (_10895_, _10894_, _04353_);
  or (_10896_, _10889_, _04381_);
  nor (_10897_, _01562_, _01554_);
  and (_10898_, _01562_, \oc8051_golden_model_1.ACC [2]);
  or (_10899_, _10898_, _04380_);
  or (_10900_, _10899_, _10897_);
  and (_10901_, _10900_, _10896_);
  and (_10902_, _10901_, _02816_);
  and (_10903_, _04489_, _04155_);
  nor (_10904_, _04489_, _04155_);
  nor (_10905_, _10904_, _10903_);
  nor (_10906_, _10905_, _02816_);
  or (_10907_, _10906_, _10902_);
  and (_10908_, _10907_, _04366_);
  nand (_10909_, _08687_, _08250_);
  and (_10910_, _10909_, _02837_);
  or (_10911_, _10910_, _03279_);
  or (_10912_, _10911_, _10908_);
  nor (_10913_, _01558_, _01553_);
  nor (_10914_, _10913_, _02841_);
  and (_10915_, _10914_, _10912_);
  and (_10916_, _03456_, _02841_);
  or (_10917_, _10916_, _02856_);
  or (_10918_, _10917_, _10915_);
  and (_10919_, _10918_, _10895_);
  or (_10920_, _10919_, _01878_);
  nand (_10921_, _06816_, _01878_);
  and (_10922_, _10921_, _02962_);
  and (_10923_, _10922_, _10920_);
  not (_10924_, _08688_);
  and (_10925_, _10909_, _10924_);
  and (_10926_, _10925_, _02862_);
  or (_10927_, _10926_, _10923_);
  and (_10928_, _10927_, _01565_);
  or (_10929_, _01565_, _01554_);
  nand (_10930_, _01989_, _10929_);
  or (_10931_, _10930_, _10928_);
  nand (_10932_, _06816_, _02503_);
  and (_10933_, _10932_, _10931_);
  or (_10934_, _10933_, _02871_);
  and (_10935_, _05043_, _03673_);
  nand (_10936_, _06815_, _02871_);
  or (_10937_, _10936_, _10935_);
  and (_10938_, _10937_, _10934_);
  or (_10939_, _10938_, _02870_);
  nor (_10940_, _08273_, _03855_);
  and (_10941_, _03855_, \oc8051_golden_model_1.PSW [7]);
  nor (_10942_, _10941_, _10940_);
  nand (_10943_, _10942_, _02870_);
  and (_10944_, _10943_, _04310_);
  and (_10945_, _10944_, _10939_);
  nand (_10946_, _01604_, _01553_);
  nand (_10947_, _02887_, _10946_);
  or (_10948_, _10947_, _10945_);
  and (_10949_, _10948_, _10893_);
  or (_10950_, _10949_, _02889_);
  or (_10951_, _05043_, _02890_);
  and (_10952_, _10951_, _02880_);
  and (_10953_, _10952_, _10950_);
  nor (_10954_, _04560_, _03455_);
  not (_10955_, _10954_);
  and (_10956_, _04730_, \oc8051_golden_model_1.IP [2]);
  and (_10957_, _04734_, \oc8051_golden_model_1.ACC [2]);
  nor (_10958_, _10957_, _10956_);
  and (_10959_, _04737_, \oc8051_golden_model_1.PSW [2]);
  and (_10960_, _04739_, \oc8051_golden_model_1.B [2]);
  nor (_10961_, _10960_, _10959_);
  and (_10962_, _10961_, _10958_);
  and (_10963_, _04686_, \oc8051_golden_model_1.TL0 [2]);
  not (_10964_, _10963_);
  and (_10965_, _04706_, \oc8051_golden_model_1.P1INREG [2]);
  and (_10966_, _04710_, \oc8051_golden_model_1.P3INREG [2]);
  nor (_10967_, _10966_, _10965_);
  and (_10968_, _10967_, _10964_);
  and (_10969_, _04703_, \oc8051_golden_model_1.P0INREG [2]);
  and (_10970_, _04675_, \oc8051_golden_model_1.P2INREG [2]);
  nor (_10971_, _10970_, _10969_);
  and (_10972_, _10971_, _10968_);
  and (_10973_, _04746_, \oc8051_golden_model_1.SP [2]);
  not (_10974_, _10973_);
  and (_10975_, _04691_, \oc8051_golden_model_1.IE [2]);
  not (_10976_, _10975_);
  and (_10977_, _04697_, \oc8051_golden_model_1.SCON [2]);
  and (_10978_, _04699_, \oc8051_golden_model_1.SBUF [2]);
  nor (_10979_, _10978_, _10977_);
  and (_10980_, _10979_, _10976_);
  and (_10981_, _10980_, _10974_);
  and (_10982_, _10981_, _10972_);
  and (_10983_, _10982_, _10962_);
  and (_10984_, _04681_, \oc8051_golden_model_1.TMOD [2]);
  and (_10985_, _04662_, \oc8051_golden_model_1.TH1 [2]);
  nor (_10986_, _10985_, _10984_);
  and (_10987_, _04744_, \oc8051_golden_model_1.DPL [2]);
  and (_10988_, _04667_, \oc8051_golden_model_1.DPH [2]);
  nor (_10989_, _10988_, _10987_);
  and (_10990_, _10989_, _10986_);
  and (_10991_, _04722_, \oc8051_golden_model_1.TCON [2]);
  and (_10992_, _04717_, \oc8051_golden_model_1.TH0 [2]);
  nor (_10993_, _10992_, _10991_);
  and (_10994_, _04726_, \oc8051_golden_model_1.PCON [2]);
  and (_10995_, _04719_, \oc8051_golden_model_1.TL1 [2]);
  nor (_10996_, _10995_, _10994_);
  and (_10997_, _10996_, _10993_);
  and (_10998_, _10997_, _10990_);
  and (_10999_, _10998_, _10983_);
  and (_11000_, _10999_, _10955_);
  nor (_11001_, _11000_, _02880_);
  or (_11002_, _11001_, _04758_);
  or (_11003_, _11002_, _10953_);
  and (_11004_, _04758_, _02294_);
  nor (_11005_, _11004_, _01871_);
  and (_11006_, _11005_, _11003_);
  and (_11007_, _04724_, _01871_);
  or (_11008_, _11007_, _01638_);
  or (_11009_, _11008_, _11006_);
  and (_11010_, _01638_, _01554_);
  nor (_11011_, _11010_, _02914_);
  and (_11012_, _11011_, _11009_);
  and (_11013_, _04155_, _02338_);
  nor (_11014_, _11013_, _10891_);
  nor (_11015_, _11014_, _02913_);
  nor (_11016_, _11015_, _02915_);
  or (_11017_, _11016_, _11012_);
  nor (_11018_, _04155_, _06184_);
  and (_11019_, _04155_, _06184_);
  nor (_11020_, _11019_, _11018_);
  or (_11021_, _11020_, _04775_);
  and (_11022_, _11021_, _02911_);
  and (_11023_, _11022_, _11017_);
  or (_11024_, _11023_, _10892_);
  and (_11025_, _11024_, _02909_);
  and (_11026_, _11018_, _02908_);
  or (_11027_, _11026_, _01632_);
  or (_11028_, _11027_, _11025_);
  and (_11029_, _01632_, _01554_);
  nor (_11030_, _11029_, _04789_);
  and (_11031_, _11030_, _11028_);
  nor (_11032_, _11013_, _04795_);
  or (_11033_, _11032_, _04794_);
  or (_11034_, _11033_, _11031_);
  nand (_11035_, _11019_, _04794_);
  and (_11036_, _11035_, _04799_);
  and (_11037_, _11036_, _11034_);
  and (_11038_, _01978_, _01641_);
  or (_11039_, _02718_, _11038_);
  and (_11040_, _01636_, _01553_);
  and (_11041_, _01983_, _01641_);
  or (_11042_, _11041_, _11040_);
  or (_11043_, _11042_, _11039_);
  or (_11044_, _11043_, _11037_);
  and (_11045_, _11044_, _10890_);
  or (_11046_, _11045_, _02930_);
  or (_11047_, _10889_, _04807_);
  and (_11048_, _11047_, _04815_);
  and (_11049_, _11048_, _11046_);
  or (_11050_, _11049_, _10886_);
  and (_11051_, _11050_, _04814_);
  nor (_11052_, _10905_, _04814_);
  or (_11053_, _11052_, _02058_);
  or (_11054_, _11053_, _11051_);
  nand (_11055_, _09943_, _02058_);
  and (_11056_, _11055_, _10453_);
  and (_11057_, _11056_, _11054_);
  and (_11058_, _01642_, _01553_);
  or (_11059_, _02941_, _11058_);
  or (_11060_, _11059_, _11057_);
  or (_11061_, _10940_, _02958_);
  and (_11062_, _11061_, _05172_);
  and (_11063_, _11062_, _11060_);
  or (_11064_, _11063_, _10881_);
  and (_11065_, _11064_, _05178_);
  or (_11066_, _05179_, _05043_);
  nor (_11067_, _06572_, _05178_);
  and (_11068_, _11067_, _11066_);
  or (_11069_, _11068_, _01791_);
  or (_11070_, _11069_, _11065_);
  nor (_11071_, _04156_, _04107_);
  nor (_11072_, _11071_, _04157_);
  or (_11073_, _11072_, _03118_);
  and (_11074_, _11073_, _03186_);
  and (_11075_, _11074_, _11070_);
  and (_11076_, _11075_, _10673_);
  or (_11077_, _11076_, _10878_);
  and (_11078_, _11077_, _10682_);
  and (_11079_, _09906_, _02058_);
  not (_11080_, _10021_);
  nor (_11081_, _11080_, _02058_);
  or (_11082_, _11081_, _11079_);
  and (_11083_, _11082_, _10681_);
  or (_37201_, _11083_, _11078_);
  or (_11084_, _06733_, _06732_);
  nor (_11085_, _05172_, _05163_);
  and (_11086_, _11085_, _11084_);
  not (_11087_, _04998_);
  nor (_11088_, _10883_, _11087_);
  or (_11089_, _11088_, _05045_);
  and (_11090_, _11089_, _02935_);
  and (_11091_, _01682_, _01636_);
  nor (_11092_, _04013_, _01689_);
  and (_11093_, _04013_, _01689_);
  nor (_11094_, _11093_, _11092_);
  and (_11095_, _11094_, _02913_);
  nor (_11096_, _08746_, _03849_);
  or (_11097_, _11096_, _04353_);
  nand (_11098_, _08746_, _08386_);
  or (_11099_, _11098_, _04366_);
  nor (_11100_, _10903_, _04013_);
  nor (_11101_, _11100_, _04491_);
  nor (_11102_, _11101_, _02816_);
  nor (_11103_, _10887_, _03268_);
  or (_11104_, _11103_, _04374_);
  or (_11105_, _11104_, _04381_);
  nor (_11106_, _01683_, _01562_);
  and (_11107_, _01562_, \oc8051_golden_model_1.ACC [3]);
  or (_11108_, _11107_, _11106_);
  nor (_11109_, _11108_, _04380_);
  nor (_11110_, _11109_, _02815_);
  and (_11111_, _11110_, _11105_);
  or (_11112_, _11111_, _02837_);
  or (_11113_, _11112_, _11102_);
  and (_11114_, _11113_, _11099_);
  or (_11115_, _11114_, _03279_);
  nor (_11116_, _01682_, _01558_);
  nor (_11117_, _11116_, _02841_);
  and (_11118_, _11117_, _11115_);
  and (_11119_, _06732_, _02841_);
  or (_11120_, _11119_, _02856_);
  or (_11121_, _11120_, _11118_);
  and (_11122_, _11121_, _11097_);
  or (_11123_, _11122_, _01878_);
  nand (_11124_, _06804_, _01878_);
  and (_11125_, _11124_, _02962_);
  and (_11126_, _11125_, _11123_);
  not (_11127_, _08747_);
  and (_11128_, _11098_, _11127_);
  and (_11129_, _11128_, _02862_);
  or (_11130_, _11129_, _11126_);
  and (_11131_, _11130_, _01565_);
  or (_11132_, _01683_, _01565_);
  nand (_11133_, _01989_, _11132_);
  or (_11134_, _11133_, _11131_);
  nand (_11135_, _06804_, _02503_);
  and (_11136_, _11135_, _11134_);
  or (_11137_, _11136_, _02871_);
  and (_11138_, _04998_, _03673_);
  nand (_11139_, _06803_, _02871_);
  or (_11140_, _11139_, _11138_);
  and (_11141_, _11140_, _11137_);
  or (_11142_, _11141_, _02870_);
  and (_11143_, _03849_, \oc8051_golden_model_1.PSW [7]);
  nor (_11144_, _08409_, _03849_);
  nor (_11145_, _11144_, _11143_);
  nand (_11146_, _11145_, _02870_);
  and (_11147_, _11146_, _04310_);
  and (_11148_, _11147_, _11142_);
  nand (_11149_, _01682_, _01604_);
  nand (_11150_, _02887_, _11149_);
  or (_11151_, _11150_, _11148_);
  or (_11152_, _06732_, _02887_);
  and (_11153_, _11152_, _11151_);
  or (_11154_, _11153_, _02889_);
  or (_11155_, _04998_, _02890_);
  and (_11156_, _11155_, _02880_);
  and (_11157_, _11156_, _11154_);
  nor (_11158_, _04560_, _03268_);
  not (_11159_, _11158_);
  and (_11160_, _04734_, \oc8051_golden_model_1.ACC [3]);
  not (_11161_, _11160_);
  and (_11162_, _04681_, \oc8051_golden_model_1.TMOD [3]);
  and (_11163_, _04739_, \oc8051_golden_model_1.B [3]);
  nor (_11164_, _11163_, _11162_);
  and (_11165_, _11164_, _11161_);
  and (_11166_, _04662_, \oc8051_golden_model_1.TH1 [3]);
  not (_11167_, _11166_);
  and (_11168_, _04730_, \oc8051_golden_model_1.IP [3]);
  and (_11169_, _04737_, \oc8051_golden_model_1.PSW [3]);
  nor (_11170_, _11169_, _11168_);
  and (_11171_, _11170_, _11167_);
  and (_11172_, _04744_, \oc8051_golden_model_1.DPL [3]);
  and (_11173_, _04667_, \oc8051_golden_model_1.DPH [3]);
  nor (_11174_, _11173_, _11172_);
  and (_11175_, _11174_, _11171_);
  and (_11176_, _11175_, _11165_);
  and (_11177_, _04722_, \oc8051_golden_model_1.TCON [3]);
  and (_11178_, _04717_, \oc8051_golden_model_1.TH0 [3]);
  nor (_11179_, _11178_, _11177_);
  and (_11180_, _04726_, \oc8051_golden_model_1.PCON [3]);
  and (_11181_, _04719_, \oc8051_golden_model_1.TL1 [3]);
  nor (_11182_, _11181_, _11180_);
  and (_11183_, _11182_, _11179_);
  and (_11184_, _04675_, \oc8051_golden_model_1.P2INREG [3]);
  not (_11185_, _11184_);
  and (_11186_, _04706_, \oc8051_golden_model_1.P1INREG [3]);
  and (_11187_, _04710_, \oc8051_golden_model_1.P3INREG [3]);
  nor (_11188_, _11187_, _11186_);
  and (_11189_, _11188_, _11185_);
  and (_11190_, _04703_, \oc8051_golden_model_1.P0INREG [3]);
  and (_11191_, _04686_, \oc8051_golden_model_1.TL0 [3]);
  nor (_11192_, _11191_, _11190_);
  and (_11193_, _11192_, _11189_);
  and (_11194_, _04746_, \oc8051_golden_model_1.SP [3]);
  not (_11195_, _11194_);
  and (_11196_, _04691_, \oc8051_golden_model_1.IE [3]);
  not (_11197_, _11196_);
  and (_11198_, _04697_, \oc8051_golden_model_1.SCON [3]);
  and (_11199_, _04699_, \oc8051_golden_model_1.SBUF [3]);
  nor (_11200_, _11199_, _11198_);
  and (_11201_, _11200_, _11197_);
  and (_11202_, _11201_, _11195_);
  and (_11203_, _11202_, _11193_);
  and (_11204_, _11203_, _11183_);
  and (_11205_, _11204_, _11176_);
  and (_11206_, _11205_, _11159_);
  nor (_11207_, _11206_, _02880_);
  or (_11208_, _11207_, _04758_);
  or (_11209_, _11208_, _11157_);
  and (_11210_, _04758_, _01954_);
  nor (_11211_, _11210_, _01871_);
  and (_11212_, _11211_, _11209_);
  and (_11213_, _04678_, _01871_);
  or (_11214_, _11213_, _01638_);
  or (_11215_, _11214_, _11212_);
  nand (_11216_, _01683_, _01638_);
  and (_11217_, _11216_, _11215_);
  or (_11218_, _11217_, _02914_);
  not (_11219_, _02914_);
  and (_11220_, _04013_, _02159_);
  nor (_11221_, _04013_, _02159_);
  nor (_11222_, _11221_, _11220_);
  or (_11223_, _11222_, _11219_);
  and (_11224_, _11223_, _04775_);
  and (_11225_, _11224_, _11218_);
  or (_11226_, _11225_, _11095_);
  and (_11227_, _11226_, _02911_);
  and (_11228_, _11221_, _02910_);
  or (_11229_, _11228_, _11227_);
  and (_11230_, _11229_, _02909_);
  and (_11231_, _11092_, _02908_);
  or (_11232_, _11231_, _01632_);
  or (_11233_, _11232_, _11230_);
  and (_11234_, _01683_, _01632_);
  nor (_11235_, _11234_, _04789_);
  and (_11236_, _11235_, _11233_);
  nor (_11237_, _11220_, _04795_);
  or (_11238_, _11237_, _04794_);
  or (_11239_, _11238_, _11236_);
  nand (_11240_, _11093_, _04794_);
  and (_11241_, _11240_, _04799_);
  nand (_11242_, _11241_, _11239_);
  nand (_11243_, _11242_, _04804_);
  or (_11244_, _11243_, _11091_);
  or (_11245_, _11104_, _04804_);
  and (_11246_, _11245_, _11244_);
  or (_11247_, _11246_, _02930_);
  or (_11248_, _11104_, _04807_);
  and (_11249_, _11248_, _04815_);
  and (_11250_, _11249_, _11247_);
  or (_11251_, _11250_, _11090_);
  and (_11252_, _11251_, _04814_);
  nor (_11253_, _11101_, _04814_);
  or (_11254_, _11253_, _02058_);
  or (_11255_, _11254_, _11252_);
  nand (_11256_, _09938_, _02058_);
  and (_11257_, _11256_, _10453_);
  and (_11258_, _11257_, _11255_);
  and (_11259_, _01682_, _01642_);
  or (_11260_, _02941_, _11259_);
  or (_11261_, _11260_, _11258_);
  or (_11262_, _11144_, _02958_);
  and (_11263_, _11262_, _05172_);
  and (_11264_, _11263_, _11261_);
  or (_11265_, _11264_, _11086_);
  and (_11266_, _11265_, _05178_);
  or (_11267_, _06572_, _04998_);
  nor (_11268_, _05181_, _05178_);
  and (_11269_, _11268_, _11267_);
  or (_11270_, _11269_, _01791_);
  or (_11271_, _11270_, _11266_);
  nor (_11272_, _04157_, _04014_);
  nor (_11273_, _11272_, _04158_);
  or (_11274_, _11273_, _03118_);
  and (_11275_, _11274_, _03186_);
  and (_11276_, _11275_, _11271_);
  or (_11277_, _11276_, _10674_);
  or (_11278_, _10673_, \oc8051_golden_model_1.IRAM[0] [3]);
  and (_11279_, _11278_, _10682_);
  and (_11280_, _11279_, _11277_);
  not (_11281_, _10017_);
  nor (_11282_, _11281_, _02058_);
  and (_11283_, _09900_, _02058_);
  or (_11284_, _11283_, _11282_);
  and (_11285_, _11284_, _10681_);
  or (_37203_, _11285_, _11280_);
  not (_11286_, _05135_);
  and (_11287_, _05045_, _11286_);
  nor (_11288_, _05045_, _11286_);
  or (_11289_, _11288_, _11287_);
  and (_11290_, _11289_, _02935_);
  nor (_11291_, _04374_, _04211_);
  and (_11292_, _04374_, _04211_);
  or (_11293_, _11292_, _11291_);
  or (_11294_, _11293_, _04804_);
  nor (_11295_, _04657_, _04257_);
  and (_11296_, _11295_, _02910_);
  nor (_11297_, _08329_, _08301_);
  and (_11298_, _08301_, \oc8051_golden_model_1.PSW [7]);
  nor (_11299_, _11298_, _11297_);
  nor (_11300_, _11299_, _04311_);
  nor (_11301_, _08301_, _08710_);
  or (_11302_, _11301_, _04353_);
  nand (_11303_, _08302_, _08710_);
  or (_11304_, _11303_, _04366_);
  or (_11305_, _11293_, _04381_);
  and (_11306_, _01562_, \oc8051_golden_model_1.ACC [4]);
  nor (_11307_, _10049_, _01562_);
  or (_11308_, _11307_, _04380_);
  or (_11309_, _11308_, _11306_);
  and (_11310_, _11309_, _11305_);
  or (_11311_, _11310_, _01883_);
  or (_11312_, _05135_, _04394_);
  and (_11313_, _11312_, _11311_);
  or (_11314_, _11313_, _02815_);
  and (_11315_, _04491_, _04257_);
  nor (_11316_, _04491_, _04257_);
  nor (_11317_, _11316_, _11315_);
  nand (_11318_, _11317_, _02815_);
  and (_11319_, _11318_, _11314_);
  or (_11320_, _11319_, _02837_);
  and (_11321_, _11320_, _11304_);
  or (_11322_, _11321_, _03279_);
  nor (_11323_, _10048_, _01558_);
  nor (_11324_, _11323_, _02841_);
  and (_11325_, _11324_, _11322_);
  and (_11326_, _05160_, _02841_);
  or (_11327_, _11326_, _02856_);
  or (_11328_, _11327_, _11325_);
  and (_11329_, _11328_, _11302_);
  or (_11330_, _11329_, _01878_);
  nand (_11331_, _06884_, _01878_);
  and (_11332_, _11331_, _02962_);
  and (_11333_, _11332_, _11330_);
  not (_11334_, _08711_);
  and (_11335_, _11303_, _11334_);
  and (_11336_, _11335_, _02862_);
  or (_11337_, _11336_, _11333_);
  and (_11338_, _11337_, _01565_);
  or (_11339_, _10049_, _01565_);
  nand (_11340_, _11339_, _01989_);
  or (_11341_, _11340_, _11338_);
  nand (_11342_, _06884_, _02503_);
  and (_11343_, _11342_, _11341_);
  or (_11344_, _11343_, _02871_);
  and (_11345_, _05135_, _03673_);
  nand (_11346_, _06883_, _02871_);
  or (_11347_, _11346_, _11345_);
  and (_11348_, _11347_, _04311_);
  and (_11349_, _11348_, _11344_);
  or (_11350_, _11349_, _11300_);
  and (_11351_, _11350_, _04310_);
  nand (_11352_, _10048_, _01604_);
  nand (_11353_, _11352_, _02887_);
  or (_11354_, _11353_, _11351_);
  or (_11355_, _05160_, _02887_);
  and (_11356_, _11355_, _11354_);
  or (_11357_, _11356_, _02889_);
  or (_11358_, _05135_, _02890_);
  and (_11359_, _11358_, _02880_);
  and (_11360_, _11359_, _11357_);
  nor (_11361_, _04560_, _04211_);
  not (_11362_, _11361_);
  and (_11363_, _04662_, \oc8051_golden_model_1.TH1 [4]);
  and (_11364_, _04667_, \oc8051_golden_model_1.DPH [4]);
  nor (_11365_, _11364_, _11363_);
  and (_11366_, _04734_, \oc8051_golden_model_1.ACC [4]);
  and (_11367_, _04732_, _04708_);
  and (_11368_, _11367_, _04671_);
  and (_11369_, _11368_, \oc8051_golden_model_1.B [4]);
  nor (_11370_, _11369_, _11366_);
  and (_11371_, _04730_, \oc8051_golden_model_1.IP [4]);
  and (_11372_, _04737_, \oc8051_golden_model_1.PSW [4]);
  nor (_11373_, _11372_, _11371_);
  and (_11374_, _11373_, _11370_);
  and (_11375_, _04675_, \oc8051_golden_model_1.P2INREG [4]);
  not (_11376_, _11375_);
  and (_11377_, _04681_, \oc8051_golden_model_1.TMOD [4]);
  and (_11378_, _04686_, \oc8051_golden_model_1.TL0 [4]);
  nor (_11379_, _11378_, _11377_);
  and (_11380_, _11379_, _11376_);
  and (_11381_, _11380_, _11374_);
  and (_11382_, _11381_, _11365_);
  and (_11383_, _04717_, \oc8051_golden_model_1.TH0 [4]);
  and (_11384_, _04719_, \oc8051_golden_model_1.TL1 [4]);
  nor (_11385_, _11384_, _11383_);
  and (_11386_, _04722_, \oc8051_golden_model_1.TCON [4]);
  and (_11387_, _04726_, \oc8051_golden_model_1.PCON [4]);
  nor (_11388_, _11387_, _11386_);
  and (_11389_, _11388_, _11385_);
  and (_11390_, _04744_, \oc8051_golden_model_1.DPL [4]);
  not (_11391_, _11390_);
  and (_11392_, _04703_, \oc8051_golden_model_1.P0INREG [4]);
  not (_11393_, _11392_);
  and (_11394_, _04706_, \oc8051_golden_model_1.P1INREG [4]);
  and (_11395_, _04710_, \oc8051_golden_model_1.P3INREG [4]);
  nor (_11396_, _11395_, _11394_);
  and (_11397_, _11396_, _11393_);
  and (_11398_, _11397_, _11391_);
  and (_11399_, _04691_, \oc8051_golden_model_1.IE [4]);
  not (_11400_, _11399_);
  and (_11401_, _04697_, \oc8051_golden_model_1.SCON [4]);
  and (_11402_, _04699_, \oc8051_golden_model_1.SBUF [4]);
  nor (_11403_, _11402_, _11401_);
  and (_11404_, _11403_, _11400_);
  and (_11405_, _04746_, \oc8051_golden_model_1.SP [4]);
  not (_11406_, _11405_);
  and (_11407_, _11406_, _11404_);
  and (_11408_, _11407_, _11398_);
  and (_11409_, _11408_, _11389_);
  and (_11410_, _11409_, _11382_);
  and (_11411_, _11410_, _11362_);
  nor (_11412_, _11411_, _02880_);
  or (_11413_, _11412_, _04758_);
  or (_11414_, _11413_, _11360_);
  and (_11415_, _04758_, _01855_);
  nor (_11416_, _11415_, _01871_);
  and (_11417_, _11416_, _11414_);
  and (_11418_, _04694_, _01871_);
  or (_11419_, _11418_, _01638_);
  or (_11420_, _11419_, _11417_);
  and (_11421_, _10049_, _01638_);
  nor (_11422_, _11421_, _02914_);
  and (_11423_, _11422_, _11420_);
  and (_11424_, _04657_, _04257_);
  nor (_11425_, _11424_, _11295_);
  nor (_11426_, _11425_, _02913_);
  nor (_11427_, _11426_, _02915_);
  or (_11428_, _11427_, _11423_);
  nor (_11429_, _04257_, _06085_);
  and (_11430_, _04257_, _06085_);
  nor (_11431_, _11430_, _11429_);
  or (_11432_, _11431_, _04775_);
  and (_11433_, _11432_, _02911_);
  and (_11434_, _11433_, _11428_);
  or (_11435_, _11434_, _11296_);
  and (_11436_, _11435_, _02909_);
  and (_11437_, _11429_, _02908_);
  or (_11438_, _11437_, _01632_);
  or (_11439_, _11438_, _11436_);
  and (_11440_, _10049_, _01632_);
  nor (_11441_, _11440_, _04789_);
  and (_11442_, _11441_, _11439_);
  nor (_11443_, _11424_, _04795_);
  or (_11444_, _11443_, _04794_);
  or (_11445_, _11444_, _11442_);
  nand (_11446_, _11430_, _04794_);
  and (_11447_, _11446_, _04799_);
  and (_11448_, _11447_, _11445_);
  and (_11449_, _10048_, _01636_);
  or (_11450_, _11449_, _11041_);
  or (_11451_, _11450_, _11039_);
  or (_11452_, _11451_, _11448_);
  and (_11453_, _11452_, _11294_);
  or (_11454_, _11453_, _02930_);
  or (_11455_, _11293_, _04807_);
  and (_11456_, _11455_, _04815_);
  and (_11457_, _11456_, _11454_);
  or (_11458_, _11457_, _11290_);
  and (_11459_, _11458_, _04814_);
  nor (_11460_, _11317_, _04814_);
  or (_11461_, _11460_, _02058_);
  or (_11462_, _11461_, _11459_);
  or (_11463_, _09934_, _05195_);
  and (_11464_, _11463_, _10453_);
  and (_11465_, _11464_, _11462_);
  and (_11466_, _10048_, _01642_);
  or (_11467_, _11466_, _02941_);
  or (_11468_, _11467_, _11465_);
  or (_11469_, _11297_, _02958_);
  and (_11470_, _05154_, _03144_);
  and (_11471_, _11470_, _11469_);
  and (_11472_, _11471_, _11468_);
  nor (_11473_, _05181_, _05135_);
  nor (_11474_, _11473_, _06554_);
  and (_11475_, _11474_, _03143_);
  nor (_11476_, _05163_, _05160_);
  nor (_11477_, _11476_, _05164_);
  and (_11478_, _11477_, _05171_);
  or (_11479_, _11478_, _03121_);
  or (_11480_, _11479_, _11475_);
  or (_11481_, _11480_, _11472_);
  not (_11482_, _02645_);
  or (_11483_, _11474_, _11482_);
  and (_11484_, _11483_, _11481_);
  or (_11485_, _11484_, _01791_);
  nor (_11486_, _04258_, _04158_);
  nor (_11487_, _11486_, _04259_);
  or (_11488_, _11487_, _03118_);
  and (_11489_, _11488_, _03186_);
  and (_11490_, _11489_, _11485_);
  or (_11491_, _11490_, _10674_);
  or (_11492_, _10673_, \oc8051_golden_model_1.IRAM[0] [4]);
  and (_11493_, _11492_, _10682_);
  and (_11494_, _11493_, _11491_);
  and (_11495_, _10013_, _05195_);
  and (_11496_, _09895_, _02058_);
  or (_11497_, _11496_, _11495_);
  and (_11498_, _11497_, _10681_);
  or (_37204_, _11498_, _11494_);
  nor (_11499_, _05164_, _05159_);
  nor (_11500_, _11499_, _05165_);
  and (_11501_, _11500_, _05171_);
  nor (_11502_, _04626_, _03964_);
  and (_11503_, _11502_, _02910_);
  nor (_11504_, _08435_, _08411_);
  and (_11505_, _08411_, \oc8051_golden_model_1.PSW [7]);
  nor (_11506_, _11505_, _11504_);
  nor (_11507_, _11506_, _04311_);
  nor (_11508_, _08411_, _08757_);
  or (_11509_, _11508_, _04353_);
  nand (_11510_, _08412_, _08757_);
  or (_11511_, _11510_, _04366_);
  or (_11512_, _05090_, _04394_);
  nor (_11513_, _11292_, _03916_);
  or (_11514_, _11513_, _04375_);
  and (_11515_, _11514_, _04380_);
  or (_11516_, _10043_, _01562_);
  nand (_11517_, _01562_, _06079_);
  and (_11518_, _11517_, _11516_);
  and (_11519_, _11518_, _04381_);
  or (_11520_, _11519_, _01883_);
  or (_11521_, _11520_, _11515_);
  and (_11522_, _11521_, _11512_);
  or (_11523_, _11522_, _02815_);
  nor (_11524_, _11315_, _03964_);
  nor (_11525_, _11524_, _04492_);
  nand (_11526_, _11525_, _02815_);
  and (_11527_, _11526_, _11523_);
  or (_11528_, _11527_, _02837_);
  and (_11529_, _11528_, _11511_);
  or (_11530_, _11529_, _03279_);
  nor (_11531_, _10043_, _01558_);
  nor (_11532_, _11531_, _02841_);
  and (_11533_, _11532_, _11530_);
  and (_11534_, _05159_, _02841_);
  or (_11535_, _11534_, _02856_);
  or (_11536_, _11535_, _11533_);
  and (_11537_, _11536_, _11509_);
  or (_11538_, _11537_, _01878_);
  nand (_11539_, _06867_, _01878_);
  and (_11540_, _11539_, _02962_);
  and (_11541_, _11540_, _11538_);
  not (_11542_, _08758_);
  and (_11543_, _11510_, _11542_);
  and (_11544_, _11543_, _02862_);
  or (_11545_, _11544_, _11541_);
  and (_11546_, _11545_, _01565_);
  or (_11547_, _10044_, _01565_);
  nand (_11548_, _11547_, _01989_);
  or (_11549_, _11548_, _11546_);
  nand (_11550_, _06867_, _02503_);
  and (_11551_, _11550_, _11549_);
  or (_11552_, _11551_, _02871_);
  and (_11553_, _05090_, _03673_);
  nand (_11554_, _06866_, _02871_);
  or (_11555_, _11554_, _11553_);
  and (_11556_, _11555_, _04311_);
  and (_11557_, _11556_, _11552_);
  or (_11558_, _11557_, _11507_);
  and (_11559_, _11558_, _04310_);
  nand (_11560_, _10043_, _01604_);
  nand (_11561_, _11560_, _02887_);
  or (_11562_, _11561_, _11559_);
  or (_11563_, _05159_, _02887_);
  and (_11564_, _11563_, _11562_);
  or (_11565_, _11564_, _02889_);
  or (_11566_, _05090_, _02890_);
  and (_11567_, _11566_, _02880_);
  and (_11568_, _11567_, _11565_);
  nor (_11569_, _04560_, _03916_);
  not (_11570_, _11569_);
  and (_11571_, _04730_, \oc8051_golden_model_1.IP [5]);
  and (_11572_, _04739_, \oc8051_golden_model_1.B [5]);
  nor (_11573_, _11572_, _11571_);
  and (_11574_, _04734_, \oc8051_golden_model_1.ACC [5]);
  and (_11575_, _04737_, \oc8051_golden_model_1.PSW [5]);
  nor (_11576_, _11575_, _11574_);
  and (_11577_, _11576_, _11573_);
  and (_11578_, _04686_, \oc8051_golden_model_1.TL0 [5]);
  not (_11579_, _11578_);
  and (_11580_, _04706_, \oc8051_golden_model_1.P1INREG [5]);
  and (_11581_, _04710_, \oc8051_golden_model_1.P3INREG [5]);
  nor (_11582_, _11581_, _11580_);
  and (_11583_, _11582_, _11579_);
  and (_11584_, _04703_, \oc8051_golden_model_1.P0INREG [5]);
  and (_11585_, _04675_, \oc8051_golden_model_1.P2INREG [5]);
  nor (_11586_, _11585_, _11584_);
  and (_11587_, _11586_, _11583_);
  and (_11588_, _04746_, \oc8051_golden_model_1.SP [5]);
  not (_11589_, _11588_);
  and (_11590_, _04691_, \oc8051_golden_model_1.IE [5]);
  not (_11591_, _11590_);
  and (_11592_, _04697_, \oc8051_golden_model_1.SCON [5]);
  and (_11593_, _04699_, \oc8051_golden_model_1.SBUF [5]);
  nor (_11594_, _11593_, _11592_);
  and (_11595_, _11594_, _11591_);
  and (_11596_, _11595_, _11589_);
  and (_11597_, _11596_, _11587_);
  and (_11598_, _11597_, _11577_);
  and (_11599_, _04717_, \oc8051_golden_model_1.TH0 [5]);
  and (_11600_, _04719_, \oc8051_golden_model_1.TL1 [5]);
  nor (_11601_, _11600_, _11599_);
  and (_11602_, _04722_, \oc8051_golden_model_1.TCON [5]);
  and (_11603_, _04726_, \oc8051_golden_model_1.PCON [5]);
  nor (_11604_, _11603_, _11602_);
  and (_11605_, _11604_, _11601_);
  and (_11606_, _04681_, \oc8051_golden_model_1.TMOD [5]);
  and (_11607_, _04662_, \oc8051_golden_model_1.TH1 [5]);
  nor (_11608_, _11607_, _11606_);
  and (_11609_, _04744_, \oc8051_golden_model_1.DPL [5]);
  and (_11610_, _04667_, \oc8051_golden_model_1.DPH [5]);
  nor (_11611_, _11610_, _11609_);
  and (_11612_, _11611_, _11608_);
  and (_11613_, _11612_, _11605_);
  and (_11614_, _11613_, _11598_);
  and (_11615_, _11614_, _11570_);
  nor (_11616_, _11615_, _02880_);
  or (_11617_, _11616_, _04758_);
  or (_11618_, _11617_, _11568_);
  and (_11619_, _04758_, _02252_);
  nor (_11620_, _11619_, _01871_);
  and (_11621_, _11620_, _11618_);
  and (_11622_, _04672_, _01871_);
  or (_11623_, _11622_, _01638_);
  or (_11624_, _11623_, _11621_);
  and (_11625_, _10044_, _01638_);
  nor (_11626_, _11625_, _02914_);
  and (_11627_, _11626_, _11624_);
  and (_11628_, _04626_, _03964_);
  nor (_11629_, _11628_, _11502_);
  nor (_11630_, _11629_, _02913_);
  nor (_11631_, _11630_, _02915_);
  or (_11632_, _11631_, _11627_);
  nor (_11633_, _03964_, _06079_);
  and (_11634_, _03964_, _06079_);
  nor (_11635_, _11634_, _11633_);
  or (_11636_, _11635_, _04775_);
  and (_11637_, _11636_, _02911_);
  and (_11638_, _11637_, _11632_);
  or (_11639_, _11638_, _11503_);
  and (_11640_, _11639_, _02909_);
  and (_11641_, _11633_, _02908_);
  or (_11642_, _11641_, _01632_);
  or (_11643_, _11642_, _11640_);
  and (_11644_, _10044_, _01632_);
  nor (_11645_, _11644_, _04789_);
  and (_11646_, _11645_, _11643_);
  nor (_11647_, _11628_, _04795_);
  or (_11648_, _11647_, _04794_);
  or (_11649_, _11648_, _11646_);
  nand (_11650_, _11634_, _04794_);
  and (_11651_, _11650_, _04799_);
  and (_11652_, _11651_, _11649_);
  and (_11653_, _10043_, _01636_);
  or (_11654_, _11653_, _10841_);
  or (_11655_, _11654_, _11652_);
  or (_11656_, _11514_, _10638_);
  and (_11657_, _11656_, _04815_);
  and (_11658_, _11657_, _11655_);
  not (_11659_, _05090_);
  nor (_11660_, _11287_, _11659_);
  or (_11661_, _11660_, _05137_);
  and (_11662_, _11661_, _02935_);
  or (_11663_, _11662_, _11658_);
  and (_11664_, _11663_, _04814_);
  nor (_11665_, _11525_, _04814_);
  or (_11666_, _11665_, _02058_);
  or (_11667_, _11666_, _11664_);
  nand (_11668_, _09930_, _02058_);
  and (_11669_, _11668_, _10453_);
  and (_11670_, _11669_, _11667_);
  and (_11671_, _10043_, _01642_);
  or (_11672_, _11671_, _02941_);
  or (_11673_, _11672_, _11670_);
  or (_11674_, _11504_, _02958_);
  and (_11675_, _11674_, _05172_);
  and (_11676_, _11675_, _11673_);
  or (_11677_, _11676_, _11501_);
  and (_11678_, _11677_, _05178_);
  or (_11679_, _06554_, _05090_);
  nor (_11680_, _05183_, _05178_);
  and (_11681_, _11680_, _11679_);
  or (_11682_, _11681_, _01791_);
  or (_11683_, _11682_, _11678_);
  nor (_11684_, _04259_, _03965_);
  nor (_11685_, _11684_, _04260_);
  or (_11686_, _11685_, _03118_);
  and (_11687_, _11686_, _03186_);
  and (_11688_, _11687_, _11683_);
  or (_11689_, _11688_, _10674_);
  or (_11690_, _10673_, \oc8051_golden_model_1.IRAM[0] [5]);
  and (_11691_, _11690_, _10682_);
  and (_11692_, _11691_, _11689_);
  and (_11693_, _09890_, _02058_);
  not (_11694_, _10009_);
  nor (_11695_, _11694_, _02058_);
  or (_11696_, _11695_, _11693_);
  and (_11697_, _11696_, _10681_);
  or (_37206_, _11697_, _11692_);
  nor (_11698_, _05183_, _04861_);
  nor (_11699_, _11698_, _05184_);
  or (_11700_, _11699_, _05178_);
  nor (_11701_, _05137_, _04862_);
  or (_11702_, _11701_, _05138_);
  and (_11703_, _11702_, _02935_);
  nor (_11704_, _04375_, _03808_);
  or (_11705_, _11704_, _04376_);
  or (_11706_, _11705_, _04804_);
  nor (_11707_, _03862_, _06026_);
  and (_11708_, _03862_, _06026_);
  nor (_11709_, _11708_, _11707_);
  and (_11710_, _11709_, _02913_);
  nor (_11711_, _08383_, _08359_);
  and (_11712_, _08359_, \oc8051_golden_model_1.PSW [7]);
  nor (_11713_, _11712_, _11711_);
  nor (_11714_, _11713_, _04311_);
  nor (_11715_, _08359_, _08734_);
  or (_11716_, _11715_, _04353_);
  nand (_11717_, _08360_, _08734_);
  or (_11718_, _11717_, _04366_);
  or (_11719_, _11705_, _04381_);
  and (_11720_, _01562_, \oc8051_golden_model_1.ACC [6]);
  nor (_11721_, _10037_, _01562_);
  or (_11722_, _11721_, _11720_);
  or (_11723_, _11722_, _04380_);
  and (_11724_, _11723_, _11719_);
  or (_11725_, _11724_, _01883_);
  or (_11726_, _04861_, _04394_);
  and (_11727_, _11726_, _11725_);
  or (_11728_, _11727_, _02815_);
  nor (_11729_, _04492_, _03862_);
  nor (_11730_, _11729_, _04493_);
  nand (_11731_, _11730_, _02815_);
  and (_11732_, _11731_, _11728_);
  or (_11733_, _11732_, _02837_);
  and (_11734_, _11733_, _11718_);
  or (_11735_, _11734_, _03279_);
  nor (_11736_, _10036_, _01558_);
  nor (_11737_, _11736_, _02841_);
  and (_11738_, _11737_, _11735_);
  and (_11739_, _05158_, _02841_);
  or (_11740_, _11739_, _02856_);
  or (_11741_, _11740_, _11738_);
  and (_11742_, _11741_, _11716_);
  or (_11743_, _11742_, _01878_);
  nand (_11744_, _06791_, _01878_);
  and (_11745_, _11744_, _02962_);
  and (_11746_, _11745_, _11743_);
  not (_11747_, _08735_);
  and (_11748_, _11717_, _11747_);
  and (_11749_, _11748_, _02862_);
  or (_11750_, _11749_, _11746_);
  and (_11751_, _11750_, _01565_);
  or (_11752_, _10037_, _01565_);
  nand (_11753_, _11752_, _01989_);
  or (_11754_, _11753_, _11751_);
  nand (_11755_, _06791_, _02503_);
  and (_11756_, _11755_, _11754_);
  or (_11757_, _11756_, _02871_);
  and (_11758_, _04861_, _03673_);
  nand (_11759_, _06790_, _02871_);
  or (_11760_, _11759_, _11758_);
  and (_11761_, _11760_, _04311_);
  and (_11762_, _11761_, _11757_);
  or (_11763_, _11762_, _11714_);
  and (_11764_, _11763_, _04310_);
  nand (_11765_, _10036_, _01604_);
  nand (_11766_, _11765_, _02887_);
  or (_11767_, _11766_, _11764_);
  or (_11768_, _05158_, _02887_);
  and (_11769_, _11768_, _11767_);
  or (_11770_, _11769_, _02889_);
  or (_11771_, _04861_, _02890_);
  and (_11772_, _11771_, _02880_);
  and (_11773_, _11772_, _11770_);
  nor (_11774_, _04560_, _03808_);
  and (_11775_, _04662_, \oc8051_golden_model_1.TH1 [6]);
  and (_11776_, _04667_, \oc8051_golden_model_1.DPH [6]);
  nor (_11777_, _11776_, _11775_);
  and (_11778_, _04675_, \oc8051_golden_model_1.P2INREG [6]);
  not (_11779_, _11778_);
  and (_11780_, _04681_, \oc8051_golden_model_1.TMOD [6]);
  and (_11781_, _04686_, \oc8051_golden_model_1.TL0 [6]);
  nor (_11782_, _11781_, _11780_);
  and (_11783_, _11782_, _11779_);
  and (_11784_, _04691_, \oc8051_golden_model_1.IE [6]);
  not (_11785_, _11784_);
  and (_11786_, _04697_, \oc8051_golden_model_1.SCON [6]);
  and (_11787_, _04699_, \oc8051_golden_model_1.SBUF [6]);
  nor (_11788_, _11787_, _11786_);
  and (_11789_, _11788_, _11785_);
  and (_11790_, _04703_, \oc8051_golden_model_1.P0INREG [6]);
  not (_11791_, _11790_);
  and (_11792_, _04706_, \oc8051_golden_model_1.P1INREG [6]);
  and (_11793_, _04710_, \oc8051_golden_model_1.P3INREG [6]);
  nor (_11794_, _11793_, _11792_);
  and (_11795_, _11794_, _11791_);
  and (_11796_, _11795_, _11789_);
  and (_11797_, _11796_, _11783_);
  and (_11798_, _11797_, _11777_);
  and (_11799_, _04717_, \oc8051_golden_model_1.TH0 [6]);
  and (_11800_, _04719_, \oc8051_golden_model_1.TL1 [6]);
  nor (_11801_, _11800_, _11799_);
  and (_11802_, _04722_, \oc8051_golden_model_1.TCON [6]);
  and (_11803_, _04726_, \oc8051_golden_model_1.PCON [6]);
  nor (_11804_, _11803_, _11802_);
  and (_11805_, _11804_, _11801_);
  and (_11806_, _04730_, \oc8051_golden_model_1.IP [6]);
  and (_11807_, _04739_, \oc8051_golden_model_1.B [6]);
  nor (_11808_, _11807_, _11806_);
  and (_11809_, _04734_, \oc8051_golden_model_1.ACC [6]);
  and (_11810_, _04737_, \oc8051_golden_model_1.PSW [6]);
  nor (_11811_, _11810_, _11809_);
  and (_11812_, _11811_, _11808_);
  and (_11813_, _04744_, \oc8051_golden_model_1.DPL [6]);
  and (_11814_, _04746_, \oc8051_golden_model_1.SP [6]);
  nor (_11815_, _11814_, _11813_);
  and (_11816_, _11815_, _11812_);
  and (_11817_, _11816_, _11805_);
  and (_11818_, _11817_, _11798_);
  not (_11819_, _11818_);
  nor (_11820_, _11819_, _11774_);
  nor (_11821_, _11820_, _02880_);
  or (_11822_, _11821_, _04758_);
  or (_11823_, _11822_, _11773_);
  and (_11824_, _04758_, _01922_);
  nor (_11825_, _11824_, _01871_);
  and (_11826_, _11825_, _11823_);
  and (_11827_, _09920_, _01871_);
  or (_11828_, _11827_, _01638_);
  or (_11829_, _11828_, _11826_);
  and (_11830_, _10037_, _01638_);
  nor (_11831_, _11830_, _02914_);
  and (_11832_, _11831_, _11829_);
  and (_11833_, _04594_, _03862_);
  nor (_11834_, _04594_, _03862_);
  nor (_11835_, _11834_, _11833_);
  and (_11836_, _11835_, _02914_);
  or (_11837_, _11836_, _11832_);
  and (_11838_, _11837_, _04775_);
  or (_11839_, _11838_, _11710_);
  and (_11840_, _11839_, _02911_);
  and (_11841_, _11834_, _02910_);
  or (_11842_, _11841_, _11840_);
  and (_11843_, _11842_, _02909_);
  and (_11844_, _11707_, _02908_);
  or (_11845_, _11844_, _01632_);
  or (_11846_, _11845_, _11843_);
  and (_11847_, _10037_, _01632_);
  nor (_11848_, _11847_, _04789_);
  and (_11849_, _11848_, _11846_);
  nor (_11850_, _11833_, _04795_);
  or (_11851_, _11850_, _04794_);
  or (_11852_, _11851_, _11849_);
  nand (_11853_, _11708_, _04794_);
  and (_11854_, _11853_, _04799_);
  and (_11855_, _11854_, _11852_);
  and (_11856_, _10036_, _01636_);
  or (_11857_, _11856_, _11041_);
  or (_11858_, _11857_, _11039_);
  or (_11859_, _11858_, _11855_);
  and (_11860_, _11859_, _11706_);
  or (_11861_, _11860_, _02930_);
  or (_11862_, _11705_, _04807_);
  and (_11863_, _11862_, _04815_);
  and (_11864_, _11863_, _11861_);
  or (_11865_, _11864_, _11703_);
  and (_11866_, _11865_, _04814_);
  nor (_11867_, _11730_, _04814_);
  or (_11868_, _11867_, _02058_);
  or (_11869_, _11868_, _11866_);
  or (_11870_, _09923_, _05195_);
  and (_11871_, _11870_, _10453_);
  and (_11872_, _11871_, _11869_);
  and (_11873_, _10036_, _01642_);
  or (_11874_, _11873_, _02941_);
  or (_11875_, _11874_, _11872_);
  or (_11876_, _11711_, _02958_);
  and (_11877_, _11876_, _05172_);
  and (_11878_, _11877_, _11875_);
  or (_11879_, _05165_, _05158_);
  and (_11880_, _11879_, _05171_);
  and (_11881_, _11880_, _05166_);
  or (_11882_, _11881_, _02952_);
  or (_11883_, _11882_, _11878_);
  and (_11884_, _11883_, _11700_);
  or (_11885_, _11884_, _01791_);
  nor (_11886_, _04260_, _03863_);
  nor (_11887_, _11886_, _04261_);
  or (_11888_, _11887_, _03118_);
  and (_11889_, _11888_, _03186_);
  and (_11890_, _11889_, _11885_);
  or (_11891_, _11890_, _10674_);
  or (_11892_, _10673_, \oc8051_golden_model_1.IRAM[0] [6]);
  and (_11893_, _11892_, _10682_);
  and (_11894_, _11893_, _11891_);
  not (_11895_, _10001_);
  nor (_11896_, _11895_, _02058_);
  and (_11897_, _09879_, _02058_);
  or (_11898_, _11897_, _11896_);
  and (_11899_, _11898_, _10681_);
  or (_37207_, _11899_, _11894_);
  or (_11900_, _10674_, _05191_);
  or (_11901_, _10673_, \oc8051_golden_model_1.IRAM[0] [7]);
  and (_11902_, _11901_, _10682_);
  and (_11903_, _11902_, _11900_);
  and (_11904_, _10681_, _05230_);
  or (_37208_, _11904_, _11903_);
  and (_11905_, _10688_, _03556_);
  and (_11906_, _10680_, _03272_);
  not (_11907_, _11906_);
  or (_11908_, _11907_, _11905_);
  and (_11909_, _03189_, _02956_);
  and (_11910_, _11909_, _10671_);
  and (_11911_, _11910_, _10667_);
  nor (_11912_, _11910_, _02977_);
  or (_11913_, _11912_, _11906_);
  or (_11914_, _11913_, _11911_);
  and (_37211_, _11914_, _11908_);
  not (_11915_, _11910_);
  or (_11916_, _11915_, _10869_);
  or (_11917_, _11910_, \oc8051_golden_model_1.IRAM[1] [1]);
  and (_11918_, _11917_, _11907_);
  and (_11919_, _11918_, _11916_);
  and (_11920_, _10876_, _03556_);
  and (_11921_, _11920_, _11906_);
  or (_37213_, _11921_, _11919_);
  nor (_11922_, _11910_, _03399_);
  and (_11923_, _11910_, _11075_);
  or (_11924_, _11923_, _11922_);
  and (_11925_, _11924_, _11907_);
  and (_11926_, _11082_, _03556_);
  and (_11927_, _11926_, _11906_);
  or (_37214_, _11927_, _11925_);
  or (_11928_, _11915_, _11276_);
  or (_11929_, _11910_, \oc8051_golden_model_1.IRAM[1] [3]);
  and (_11930_, _11929_, _11907_);
  and (_11931_, _11930_, _11928_);
  and (_11932_, _11284_, _03556_);
  and (_11933_, _11932_, _11906_);
  or (_37215_, _11933_, _11931_);
  or (_11934_, _11915_, _11490_);
  or (_11935_, _11910_, \oc8051_golden_model_1.IRAM[1] [4]);
  and (_11936_, _11935_, _11907_);
  and (_11937_, _11936_, _11934_);
  and (_11938_, _11497_, _03556_);
  and (_11939_, _11938_, _11906_);
  or (_37216_, _11939_, _11937_);
  or (_11940_, _11915_, _11688_);
  or (_11941_, _11910_, \oc8051_golden_model_1.IRAM[1] [5]);
  and (_11942_, _11941_, _11907_);
  and (_11943_, _11942_, _11940_);
  and (_11944_, _11696_, _03556_);
  and (_11945_, _11944_, _11906_);
  or (_37217_, _11945_, _11943_);
  or (_11946_, _11915_, _11890_);
  or (_11947_, _11910_, \oc8051_golden_model_1.IRAM[1] [6]);
  and (_11948_, _11947_, _11907_);
  and (_11949_, _11948_, _11946_);
  and (_11950_, _11898_, _03556_);
  and (_11951_, _11950_, _11906_);
  or (_37219_, _11951_, _11949_);
  or (_11952_, _11915_, _05192_);
  or (_11953_, _11910_, \oc8051_golden_model_1.IRAM[1] [7]);
  and (_11954_, _11953_, _11907_);
  and (_11955_, _11954_, _11952_);
  and (_11956_, _11906_, _05231_);
  or (_37220_, _11956_, _11955_);
  and (_11957_, _10668_, _03106_);
  and (_11958_, _11957_, _10671_);
  not (_11959_, _11958_);
  or (_11960_, _11959_, _10667_);
  or (_11961_, _11958_, \oc8051_golden_model_1.IRAM[2] [0]);
  and (_11962_, _10680_, _04395_);
  not (_11963_, _11962_);
  and (_11964_, _11963_, _11961_);
  and (_11965_, _11964_, _11960_);
  and (_11966_, _11962_, _10688_);
  or (_37223_, _11966_, _11965_);
  or (_11967_, _11959_, _10869_);
  or (_11968_, _11958_, \oc8051_golden_model_1.IRAM[2] [1]);
  and (_11969_, _11968_, _11963_);
  and (_11970_, _11969_, _11967_);
  and (_11971_, _11962_, _10876_);
  or (_37224_, _11971_, _11970_);
  nor (_11972_, _11958_, _03405_);
  and (_11973_, _11958_, _11075_);
  or (_11974_, _11973_, _11972_);
  and (_11975_, _11974_, _11963_);
  and (_11976_, _11962_, _11082_);
  or (_37226_, _11976_, _11975_);
  or (_11977_, _11959_, _11276_);
  or (_11978_, _11958_, \oc8051_golden_model_1.IRAM[2] [3]);
  and (_11979_, _11978_, _11963_);
  and (_11980_, _11979_, _11977_);
  and (_11981_, _11962_, _11284_);
  or (_37227_, _11981_, _11980_);
  or (_11982_, _11959_, _11490_);
  or (_11983_, _11958_, \oc8051_golden_model_1.IRAM[2] [4]);
  and (_11984_, _11983_, _11963_);
  and (_11985_, _11984_, _11982_);
  and (_11986_, _11962_, _11497_);
  or (_37228_, _11986_, _11985_);
  or (_11987_, _11959_, _11688_);
  or (_11988_, _11958_, \oc8051_golden_model_1.IRAM[2] [5]);
  and (_11989_, _11988_, _11963_);
  and (_11990_, _11989_, _11987_);
  and (_11991_, _11962_, _11696_);
  or (_37229_, _11991_, _11990_);
  or (_11992_, _11959_, _11890_);
  or (_11993_, _11958_, \oc8051_golden_model_1.IRAM[2] [6]);
  and (_11994_, _11993_, _11963_);
  and (_11995_, _11994_, _11992_);
  and (_11996_, _11962_, _11898_);
  or (_37230_, _11996_, _11995_);
  or (_11997_, _11959_, _05192_);
  or (_11998_, _11958_, \oc8051_golden_model_1.IRAM[2] [7]);
  and (_11999_, _11998_, _11963_);
  and (_12000_, _11999_, _11997_);
  and (_12001_, _11962_, _05230_);
  or (_37232_, _12001_, _12000_);
  and (_12002_, _10671_, _03190_);
  or (_12003_, _12002_, \oc8051_golden_model_1.IRAM[3] [0]);
  and (_12004_, _10680_, _01863_);
  not (_12005_, _12004_);
  and (_12006_, _12005_, _12003_);
  not (_12007_, _12002_);
  or (_12008_, _12007_, _10667_);
  and (_12009_, _12008_, _12006_);
  and (_12010_, _12004_, _11905_);
  or (_37235_, _12010_, _12009_);
  or (_12011_, _12002_, \oc8051_golden_model_1.IRAM[3] [1]);
  and (_12012_, _12011_, _12005_);
  or (_12013_, _12007_, _10869_);
  and (_12014_, _12013_, _12012_);
  and (_12015_, _12004_, _11920_);
  or (_37236_, _12015_, _12014_);
  nor (_12016_, _12002_, _03403_);
  and (_12017_, _12002_, _11075_);
  or (_12018_, _12017_, _12016_);
  and (_12019_, _12018_, _12005_);
  and (_12020_, _12004_, _11926_);
  or (_37237_, _12020_, _12019_);
  or (_12021_, _12002_, \oc8051_golden_model_1.IRAM[3] [3]);
  and (_12022_, _12021_, _12005_);
  or (_12023_, _12007_, _11276_);
  and (_12024_, _12023_, _12022_);
  and (_12025_, _12004_, _11932_);
  or (_37238_, _12025_, _12024_);
  or (_12026_, _12002_, \oc8051_golden_model_1.IRAM[3] [4]);
  and (_12027_, _12026_, _12005_);
  or (_12028_, _12007_, _11490_);
  and (_12029_, _12028_, _12027_);
  and (_12030_, _12004_, _11938_);
  or (_37239_, _12030_, _12029_);
  or (_12031_, _12002_, \oc8051_golden_model_1.IRAM[3] [5]);
  and (_12032_, _12031_, _12005_);
  or (_12033_, _12007_, _11688_);
  and (_12034_, _12033_, _12032_);
  and (_12035_, _12004_, _11944_);
  or (_37240_, _12035_, _12034_);
  or (_12036_, _12002_, \oc8051_golden_model_1.IRAM[3] [6]);
  and (_12037_, _12036_, _12005_);
  or (_12038_, _12007_, _11890_);
  and (_12039_, _12038_, _12037_);
  and (_12040_, _12004_, _11950_);
  or (_37242_, _12040_, _12039_);
  or (_12041_, _12002_, \oc8051_golden_model_1.IRAM[3] [7]);
  and (_12042_, _12041_, _12005_);
  or (_12043_, _12007_, _05192_);
  and (_12044_, _12043_, _12042_);
  and (_12045_, _12004_, _05231_);
  or (_37243_, _12045_, _12044_);
  and (_12046_, _03540_, _03386_);
  and (_12047_, _12046_, _10669_);
  and (_12048_, _12047_, _10667_);
  nor (_12049_, _12047_, _02995_);
  or (_12050_, _12049_, _12048_);
  nor (_12051_, _03555_, _01864_);
  and (_12052_, _12051_, _38087_);
  and (_12053_, _12052_, _37580_);
  nor (_12054_, _03555_, \oc8051_golden_model_1.SP [1]);
  and (_12055_, _12054_, _38087_);
  and (_12056_, _12055_, _37580_);
  or (_12057_, _12056_, _12053_);
  nor (_12058_, _03555_, _10678_);
  and (_12059_, _12058_, _38087_);
  and (_12060_, _12059_, _37580_);
  not (_12061_, _03552_);
  nor (_12062_, _03555_, _12061_);
  and (_12063_, _12062_, _38087_);
  and (_12064_, _12063_, _37580_);
  not (_12065_, _12064_);
  nand (_12066_, _12065_, _12060_);
  or (_12067_, _12066_, _12057_);
  and (_12068_, _12067_, _12050_);
  and (_12069_, _03556_, _03548_);
  and (_12070_, _12069_, _12061_);
  and (_12071_, _12070_, _01865_);
  and (_12072_, _12071_, _11905_);
  or (_37247_, _12072_, _12068_);
  not (_12073_, _12047_);
  or (_12074_, _12073_, _10869_);
  not (_12075_, _12071_);
  or (_12076_, _12047_, \oc8051_golden_model_1.IRAM[4] [1]);
  and (_12077_, _12076_, _12075_);
  and (_12078_, _12077_, _12074_);
  and (_12079_, _12071_, _11920_);
  or (_37248_, _12079_, _12078_);
  or (_12080_, _12073_, _11075_);
  or (_12081_, _12047_, \oc8051_golden_model_1.IRAM[4] [2]);
  and (_12082_, _12081_, _12075_);
  and (_12083_, _12082_, _12080_);
  and (_12084_, _12071_, _11926_);
  or (_37250_, _12084_, _12083_);
  or (_12085_, _12073_, _11276_);
  or (_12086_, _12047_, \oc8051_golden_model_1.IRAM[4] [3]);
  and (_12087_, _12086_, _12075_);
  and (_12088_, _12087_, _12085_);
  and (_12089_, _12071_, _11932_);
  or (_37251_, _12089_, _12088_);
  or (_12090_, _12073_, _11490_);
  or (_12091_, _12047_, \oc8051_golden_model_1.IRAM[4] [4]);
  and (_12092_, _12091_, _12075_);
  and (_12093_, _12092_, _12090_);
  and (_12094_, _12071_, _11938_);
  or (_37252_, _12094_, _12093_);
  or (_12095_, _12073_, _11688_);
  or (_12096_, _12047_, \oc8051_golden_model_1.IRAM[4] [5]);
  and (_12097_, _12096_, _12075_);
  and (_12098_, _12097_, _12095_);
  and (_12099_, _12071_, _11944_);
  or (_37253_, _12099_, _12098_);
  or (_12100_, _12073_, _11890_);
  or (_12101_, _12047_, \oc8051_golden_model_1.IRAM[4] [6]);
  and (_12102_, _12101_, _12075_);
  and (_12103_, _12102_, _12100_);
  and (_12104_, _12071_, _11950_);
  or (_37254_, _12104_, _12103_);
  or (_12105_, _12073_, _05192_);
  or (_12106_, _12047_, \oc8051_golden_model_1.IRAM[4] [7]);
  and (_12107_, _12106_, _12075_);
  and (_12108_, _12107_, _12105_);
  and (_12109_, _12071_, _05231_);
  or (_37255_, _12109_, _12108_);
  and (_12110_, _12046_, _11909_);
  not (_12111_, _12110_);
  or (_12112_, _12111_, _10667_);
  and (_12113_, _12070_, _03272_);
  not (_12114_, _12113_);
  or (_12115_, _12110_, \oc8051_golden_model_1.IRAM[5] [0]);
  and (_12116_, _12115_, _12114_);
  and (_12117_, _12116_, _12112_);
  and (_12118_, _12113_, _11905_);
  or (_37258_, _12118_, _12117_);
  or (_12119_, _12111_, _10869_);
  or (_12120_, _12110_, \oc8051_golden_model_1.IRAM[5] [1]);
  and (_12121_, _12120_, _12114_);
  and (_12122_, _12121_, _12119_);
  and (_12123_, _12113_, _11920_);
  or (_37259_, _12123_, _12122_);
  or (_12124_, _12111_, _11075_);
  or (_12125_, _12110_, \oc8051_golden_model_1.IRAM[5] [2]);
  and (_12126_, _12125_, _12114_);
  and (_12127_, _12126_, _12124_);
  and (_12128_, _12113_, _11926_);
  or (_37261_, _12128_, _12127_);
  or (_12129_, _12111_, _11276_);
  or (_12130_, _12110_, \oc8051_golden_model_1.IRAM[5] [3]);
  and (_12131_, _12130_, _12114_);
  and (_12132_, _12131_, _12129_);
  and (_12133_, _12113_, _11932_);
  or (_37262_, _12133_, _12132_);
  or (_12134_, _12111_, _11490_);
  or (_12135_, _12110_, \oc8051_golden_model_1.IRAM[5] [4]);
  and (_12136_, _12135_, _12114_);
  and (_12137_, _12136_, _12134_);
  and (_12138_, _12113_, _11938_);
  or (_37263_, _12138_, _12137_);
  or (_12139_, _12111_, _11688_);
  or (_12140_, _12110_, \oc8051_golden_model_1.IRAM[5] [5]);
  and (_12141_, _12140_, _12114_);
  and (_12142_, _12141_, _12139_);
  and (_12143_, _12113_, _11944_);
  or (_37264_, _12143_, _12142_);
  or (_12144_, _12111_, _11890_);
  or (_12145_, _12110_, \oc8051_golden_model_1.IRAM[5] [6]);
  and (_12146_, _12145_, _12114_);
  and (_12147_, _12146_, _12144_);
  and (_12148_, _12113_, _11950_);
  or (_37265_, _12148_, _12147_);
  or (_12149_, _12111_, _05192_);
  or (_12150_, _12110_, \oc8051_golden_model_1.IRAM[5] [7]);
  and (_12151_, _12150_, _12114_);
  and (_12152_, _12151_, _12149_);
  and (_12153_, _12113_, _05231_);
  or (_37267_, _12153_, _12152_);
  and (_12154_, _12046_, _11957_);
  not (_12155_, _12154_);
  or (_12156_, _12155_, _10667_);
  and (_12157_, _12070_, _04395_);
  not (_12158_, _12157_);
  or (_12159_, _12154_, \oc8051_golden_model_1.IRAM[6] [0]);
  and (_12160_, _12159_, _12158_);
  and (_12161_, _12160_, _12156_);
  and (_12162_, _12157_, _11905_);
  or (_37269_, _12162_, _12161_);
  or (_12163_, _12155_, _10869_);
  or (_12164_, _12154_, \oc8051_golden_model_1.IRAM[6] [1]);
  and (_12165_, _12164_, _12158_);
  and (_12166_, _12165_, _12163_);
  and (_12167_, _12157_, _11920_);
  or (_37271_, _12167_, _12166_);
  or (_12168_, _12155_, _11075_);
  or (_12169_, _12154_, \oc8051_golden_model_1.IRAM[6] [2]);
  and (_12170_, _12169_, _12158_);
  and (_12171_, _12170_, _12168_);
  and (_12172_, _12157_, _11926_);
  or (_37272_, _12172_, _12171_);
  or (_12173_, _12155_, _11276_);
  or (_12174_, _12154_, \oc8051_golden_model_1.IRAM[6] [3]);
  and (_12175_, _12174_, _12158_);
  and (_12176_, _12175_, _12173_);
  and (_12177_, _12157_, _11932_);
  or (_37273_, _12177_, _12176_);
  or (_12178_, _12155_, _11490_);
  or (_12179_, _12154_, \oc8051_golden_model_1.IRAM[6] [4]);
  and (_12180_, _12179_, _12158_);
  and (_12181_, _12180_, _12178_);
  and (_12182_, _12157_, _11938_);
  or (_37274_, _12182_, _12181_);
  or (_12183_, _12155_, _11688_);
  or (_12184_, _12154_, \oc8051_golden_model_1.IRAM[6] [5]);
  and (_12185_, _12184_, _12158_);
  and (_12186_, _12185_, _12183_);
  and (_12187_, _12157_, _11944_);
  or (_37275_, _12187_, _12186_);
  or (_12188_, _12155_, _11890_);
  or (_12189_, _12154_, \oc8051_golden_model_1.IRAM[6] [6]);
  and (_12190_, _12189_, _12158_);
  and (_12191_, _12190_, _12188_);
  and (_12192_, _12157_, _11950_);
  or (_37277_, _12192_, _12191_);
  or (_12193_, _12155_, _05192_);
  or (_12194_, _12154_, \oc8051_golden_model_1.IRAM[6] [7]);
  and (_12195_, _12194_, _12158_);
  and (_12196_, _12195_, _12193_);
  and (_12197_, _12157_, _05231_);
  or (_37278_, _12197_, _12196_);
  and (_12198_, _12070_, _01863_);
  not (_12199_, _12198_);
  or (_12200_, _12199_, _11905_);
  and (_12201_, _12046_, _03190_);
  and (_12202_, _12201_, _10667_);
  nor (_12203_, _12201_, _02989_);
  or (_12204_, _12203_, _12198_);
  or (_12205_, _12204_, _12202_);
  and (_37281_, _12205_, _12200_);
  or (_12206_, _12201_, \oc8051_golden_model_1.IRAM[7] [1]);
  and (_12207_, _12206_, _12199_);
  not (_12208_, _12201_);
  or (_12209_, _12208_, _10869_);
  and (_12210_, _12209_, _12207_);
  and (_12211_, _12198_, _11920_);
  or (_37283_, _12211_, _12210_);
  nor (_12212_, _12201_, _03411_);
  and (_12213_, _12201_, _11075_);
  or (_12214_, _12213_, _12212_);
  and (_12215_, _12214_, _12199_);
  and (_12216_, _12198_, _11926_);
  or (_37284_, _12216_, _12215_);
  or (_12217_, _12201_, \oc8051_golden_model_1.IRAM[7] [3]);
  and (_12218_, _12217_, _12199_);
  or (_12219_, _12208_, _11276_);
  and (_12220_, _12219_, _12218_);
  and (_12221_, _12198_, _11932_);
  or (_37285_, _12221_, _12220_);
  or (_12222_, _12201_, \oc8051_golden_model_1.IRAM[7] [4]);
  and (_12223_, _12222_, _12199_);
  or (_12224_, _12208_, _11490_);
  and (_12225_, _12224_, _12223_);
  and (_12226_, _12198_, _11938_);
  or (_37286_, _12226_, _12225_);
  or (_12227_, _12201_, \oc8051_golden_model_1.IRAM[7] [5]);
  and (_12228_, _12227_, _12199_);
  or (_12229_, _12208_, _11688_);
  and (_12230_, _12229_, _12228_);
  and (_12231_, _12198_, _11944_);
  or (_37287_, _12231_, _12230_);
  or (_12232_, _12201_, \oc8051_golden_model_1.IRAM[7] [6]);
  and (_12233_, _12232_, _12199_);
  or (_12234_, _12208_, _11890_);
  and (_12235_, _12234_, _12233_);
  and (_12236_, _12198_, _11950_);
  or (_37288_, _12236_, _12235_);
  or (_12237_, _12208_, _05192_);
  or (_12238_, _12201_, \oc8051_golden_model_1.IRAM[7] [7]);
  and (_12239_, _12238_, _12199_);
  and (_12240_, _12239_, _12237_);
  and (_12241_, _12198_, _05231_);
  or (_37289_, _12241_, _12240_);
  and (_12242_, _03557_, _03546_);
  not (_12243_, _12242_);
  or (_12244_, _12243_, _11905_);
  and (_12245_, _10670_, _03539_);
  and (_12246_, _12245_, _10669_);
  and (_12247_, _12246_, _10667_);
  nor (_12248_, _12246_, _03009_);
  or (_12249_, _12248_, _12242_);
  or (_12250_, _12249_, _12247_);
  and (_37293_, _12250_, _12244_);
  or (_12251_, _12243_, _11920_);
  and (_12252_, _12246_, _10869_);
  nor (_12253_, _12246_, _02788_);
  or (_12254_, _12253_, _12242_);
  or (_12255_, _12254_, _12252_);
  and (_37294_, _12255_, _12251_);
  nor (_12256_, _12246_, _03432_);
  and (_12257_, _12246_, _11075_);
  or (_12258_, _12257_, _12256_);
  and (_12259_, _12258_, _12243_);
  and (_12260_, _12242_, _11926_);
  or (_37296_, _12260_, _12259_);
  not (_12261_, _12246_);
  or (_12262_, _12261_, _11276_);
  or (_12263_, _12246_, \oc8051_golden_model_1.IRAM[8] [3]);
  and (_12264_, _12263_, _12243_);
  and (_12265_, _12264_, _12262_);
  and (_12266_, _12242_, _11932_);
  or (_37297_, _12266_, _12265_);
  or (_12268_, _12261_, _11490_);
  or (_12270_, _12246_, \oc8051_golden_model_1.IRAM[8] [4]);
  and (_12271_, _12270_, _12243_);
  and (_12273_, _12271_, _12268_);
  and (_12274_, _12242_, _11938_);
  or (_37298_, _12274_, _12273_);
  or (_12276_, _12261_, _11688_);
  or (_12278_, _12246_, \oc8051_golden_model_1.IRAM[8] [5]);
  and (_12279_, _12278_, _12243_);
  and (_12281_, _12279_, _12276_);
  and (_12282_, _12242_, _11944_);
  or (_37299_, _12282_, _12281_);
  or (_12284_, _12261_, _11890_);
  or (_12286_, _12246_, \oc8051_golden_model_1.IRAM[8] [6]);
  and (_12287_, _12286_, _12243_);
  and (_12289_, _12287_, _12284_);
  and (_12290_, _12242_, _11950_);
  or (_37300_, _12290_, _12289_);
  or (_12292_, _12261_, _05192_);
  or (_12294_, _12246_, \oc8051_golden_model_1.IRAM[8] [7]);
  and (_12295_, _12294_, _12243_);
  and (_12297_, _12295_, _12292_);
  and (_12298_, _12242_, _05231_);
  or (_37302_, _12298_, _12297_);
  and (_12300_, _12245_, _11909_);
  not (_12301_, _12300_);
  or (_12302_, _12301_, _10667_);
  and (_12303_, _03557_, _10678_);
  and (_12304_, _12303_, _03272_);
  not (_12305_, _12304_);
  or (_12306_, _12300_, \oc8051_golden_model_1.IRAM[9] [0]);
  and (_12307_, _12306_, _12305_);
  and (_12308_, _12307_, _12302_);
  and (_12309_, _12304_, _11905_);
  or (_37304_, _12309_, _12308_);
  or (_12310_, _12301_, _10869_);
  or (_12311_, _12300_, \oc8051_golden_model_1.IRAM[9] [1]);
  and (_12312_, _12311_, _12305_);
  and (_12313_, _12312_, _12310_);
  and (_12314_, _12304_, _11920_);
  or (_37305_, _12314_, _12313_);
  or (_12315_, _12301_, _11075_);
  and (_12316_, _03557_, _03273_);
  not (_12317_, _12316_);
  or (_12318_, _12300_, \oc8051_golden_model_1.IRAM[9] [2]);
  and (_12319_, _12318_, _12317_);
  and (_12320_, _12319_, _12315_);
  and (_12321_, _12316_, _11926_);
  or (_37307_, _12321_, _12320_);
  or (_12322_, _12301_, _11276_);
  or (_12323_, _12300_, \oc8051_golden_model_1.IRAM[9] [3]);
  and (_12324_, _12323_, _12317_);
  and (_12325_, _12324_, _12322_);
  and (_12326_, _12316_, _11932_);
  or (_37308_, _12326_, _12325_);
  or (_12327_, _12301_, _11490_);
  or (_12328_, _12300_, \oc8051_golden_model_1.IRAM[9] [4]);
  and (_12329_, _12328_, _12317_);
  and (_12330_, _12329_, _12327_);
  and (_12331_, _12316_, _11938_);
  or (_37309_, _12331_, _12330_);
  or (_12332_, _12301_, _11688_);
  or (_12333_, _12300_, \oc8051_golden_model_1.IRAM[9] [5]);
  and (_12334_, _12333_, _12317_);
  and (_12335_, _12334_, _12332_);
  and (_12336_, _12316_, _11944_);
  or (_37310_, _12336_, _12335_);
  or (_12337_, _12301_, _11890_);
  or (_12338_, _12300_, \oc8051_golden_model_1.IRAM[9] [6]);
  and (_12339_, _12338_, _12317_);
  and (_12340_, _12339_, _12337_);
  and (_12342_, _12316_, _11950_);
  or (_37311_, _12342_, _12340_);
  or (_12344_, _12301_, _05192_);
  or (_12346_, _12300_, \oc8051_golden_model_1.IRAM[9] [7]);
  and (_12347_, _12346_, _12317_);
  and (_12349_, _12347_, _12344_);
  and (_12350_, _12316_, _05231_);
  or (_37313_, _12350_, _12349_);
  and (_12352_, _12245_, _11957_);
  not (_12354_, _12352_);
  or (_12355_, _12354_, _10667_);
  and (_12357_, _12303_, _04395_);
  not (_12358_, _12357_);
  or (_12360_, _12352_, \oc8051_golden_model_1.IRAM[10] [0]);
  and (_12361_, _12360_, _12358_);
  and (_12363_, _12361_, _12355_);
  and (_12364_, _12357_, _11905_);
  or (_37316_, _12364_, _12363_);
  or (_12366_, _12354_, _10869_);
  nand (_12368_, _04396_, _03557_);
  or (_12369_, _12352_, \oc8051_golden_model_1.IRAM[10] [1]);
  and (_12371_, _12369_, _12368_);
  and (_12372_, _12371_, _12366_);
  and (_12373_, _12357_, _11920_);
  or (_37317_, _12373_, _12372_);
  or (_12374_, _12354_, _11075_);
  or (_12375_, _12352_, \oc8051_golden_model_1.IRAM[10] [2]);
  and (_12376_, _12375_, _12358_);
  and (_12377_, _12376_, _12374_);
  and (_12378_, _12357_, _11926_);
  or (_37318_, _12378_, _12377_);
  or (_12379_, _12354_, _11276_);
  or (_12380_, _12352_, \oc8051_golden_model_1.IRAM[10] [3]);
  and (_12381_, _12380_, _12368_);
  and (_12382_, _12381_, _12379_);
  and (_12383_, _12357_, _11932_);
  or (_37319_, _12383_, _12382_);
  or (_12384_, _12354_, _11490_);
  or (_12385_, _12352_, \oc8051_golden_model_1.IRAM[10] [4]);
  and (_12386_, _12385_, _12368_);
  and (_12387_, _12386_, _12384_);
  and (_12388_, _12357_, _11938_);
  or (_37320_, _12388_, _12387_);
  or (_12389_, _12354_, _11688_);
  or (_12390_, _12352_, \oc8051_golden_model_1.IRAM[10] [5]);
  and (_12391_, _12390_, _12368_);
  and (_12392_, _12391_, _12389_);
  and (_12393_, _12357_, _11944_);
  or (_37321_, _12393_, _12392_);
  or (_12394_, _12354_, _11890_);
  or (_12395_, _12352_, \oc8051_golden_model_1.IRAM[10] [6]);
  and (_12396_, _12395_, _12368_);
  and (_12397_, _12396_, _12394_);
  and (_12398_, _12357_, _11950_);
  or (_37323_, _12398_, _12397_);
  nand (_12399_, _12352_, _05192_);
  or (_12400_, _12352_, _03594_);
  and (_12401_, _12400_, _12368_);
  nand (_12402_, _12401_, _12399_);
  or (_12403_, _12358_, _05231_);
  and (_37324_, _12403_, _12402_);
  not (_12404_, _03106_);
  and (_12405_, _10668_, _12404_);
  and (_12406_, _12245_, _12405_);
  not (_12407_, _12406_);
  or (_12408_, _12407_, _10667_);
  and (_12409_, _12303_, _01863_);
  not (_12410_, _12409_);
  or (_12411_, _12406_, \oc8051_golden_model_1.IRAM[11] [0]);
  and (_12412_, _12411_, _12410_);
  and (_12413_, _12412_, _12408_);
  and (_12414_, _12409_, _11905_);
  or (_37327_, _12414_, _12413_);
  or (_12415_, _12407_, _10869_);
  or (_12416_, _12406_, \oc8051_golden_model_1.IRAM[11] [1]);
  and (_12417_, _12416_, _12410_);
  and (_12418_, _12417_, _12415_);
  and (_12419_, _12409_, _11920_);
  or (_37329_, _12419_, _12418_);
  and (_12420_, _12245_, _03190_);
  or (_12421_, _12420_, \oc8051_golden_model_1.IRAM[11] [2]);
  and (_12422_, _12421_, _12410_);
  not (_12423_, _12420_);
  or (_12424_, _12423_, _11075_);
  and (_12425_, _12424_, _12422_);
  and (_12426_, _12409_, _11926_);
  or (_37330_, _12426_, _12425_);
  or (_12427_, _12420_, \oc8051_golden_model_1.IRAM[11] [3]);
  and (_12428_, _12427_, _12410_);
  or (_12429_, _12423_, _11276_);
  and (_12430_, _12429_, _12428_);
  and (_12431_, _12409_, _11932_);
  or (_37331_, _12431_, _12430_);
  or (_12432_, _12420_, \oc8051_golden_model_1.IRAM[11] [4]);
  and (_12433_, _12432_, _12410_);
  or (_12434_, _12423_, _11490_);
  and (_12435_, _12434_, _12433_);
  and (_12436_, _12409_, _11938_);
  or (_37332_, _12436_, _12435_);
  or (_12437_, _12420_, \oc8051_golden_model_1.IRAM[11] [5]);
  and (_12438_, _12437_, _12410_);
  or (_12439_, _12423_, _11688_);
  and (_12440_, _12439_, _12438_);
  and (_12441_, _12409_, _11944_);
  or (_37333_, _12441_, _12440_);
  or (_12442_, _12420_, \oc8051_golden_model_1.IRAM[11] [6]);
  and (_12443_, _12442_, _12410_);
  or (_12444_, _12423_, _11890_);
  and (_12445_, _12444_, _12443_);
  and (_12446_, _12409_, _11950_);
  or (_37335_, _12446_, _12445_);
  or (_12447_, _12420_, \oc8051_golden_model_1.IRAM[11] [7]);
  and (_12448_, _12447_, _12410_);
  or (_12449_, _12423_, _05192_);
  and (_12450_, _12449_, _12448_);
  and (_12451_, _12409_, _05231_);
  or (_37336_, _12451_, _12450_);
  and (_12452_, _10669_, _03542_);
  or (_12453_, _12452_, \oc8051_golden_model_1.IRAM[12] [0]);
  and (_12454_, _03558_, _01865_);
  not (_12455_, _12454_);
  and (_12456_, _12455_, _12453_);
  not (_12457_, _12452_);
  or (_12458_, _12457_, _10667_);
  and (_12459_, _12458_, _12456_);
  and (_12460_, _12454_, _11905_);
  or (_37339_, _12460_, _12459_);
  and (_12461_, _12069_, _03552_);
  nand (_12462_, _12461_, _01865_);
  or (_12463_, _12462_, _11920_);
  and (_12464_, _12452_, _10869_);
  or (_12465_, _12452_, _02801_);
  nand (_12466_, _12465_, _12462_);
  or (_12467_, _12466_, _12464_);
  and (_37340_, _12467_, _12463_);
  nor (_12468_, _12452_, _03445_);
  and (_12469_, _12452_, _11075_);
  or (_12470_, _12469_, _12468_);
  and (_12471_, _12470_, _12462_);
  and (_12472_, _12454_, _11926_);
  or (_37341_, _12472_, _12471_);
  or (_12473_, _12452_, \oc8051_golden_model_1.IRAM[12] [3]);
  and (_12474_, _12473_, _12455_);
  or (_12475_, _12457_, _11276_);
  and (_12476_, _12475_, _12474_);
  and (_12477_, _12454_, _11932_);
  or (_37342_, _12477_, _12476_);
  or (_12478_, _12452_, \oc8051_golden_model_1.IRAM[12] [4]);
  and (_12479_, _12478_, _12455_);
  or (_12480_, _12457_, _11490_);
  and (_12481_, _12480_, _12479_);
  and (_12482_, _12454_, _11938_);
  or (_37344_, _12482_, _12481_);
  or (_12483_, _12452_, \oc8051_golden_model_1.IRAM[12] [5]);
  and (_12484_, _12483_, _12455_);
  or (_12485_, _12457_, _11688_);
  and (_12486_, _12485_, _12484_);
  and (_12487_, _12454_, _11944_);
  or (_37345_, _12487_, _12486_);
  or (_12488_, _12452_, \oc8051_golden_model_1.IRAM[12] [6]);
  and (_12489_, _12488_, _12455_);
  or (_12490_, _12457_, _11890_);
  and (_12491_, _12490_, _12489_);
  and (_12492_, _12454_, _11950_);
  or (_37346_, _12492_, _12491_);
  or (_12493_, _12452_, \oc8051_golden_model_1.IRAM[12] [7]);
  and (_12494_, _12493_, _12455_);
  or (_12495_, _12457_, _05192_);
  and (_12496_, _12495_, _12494_);
  and (_12497_, _12454_, _05231_);
  or (_37347_, _12497_, _12496_);
  and (_12498_, _11909_, _03542_);
  not (_12499_, _12498_);
  or (_12500_, _12499_, _10667_);
  or (_12501_, _12498_, \oc8051_golden_model_1.IRAM[13] [0]);
  and (_12502_, _12461_, _03272_);
  not (_12503_, _12502_);
  and (_12504_, _12503_, _12501_);
  and (_12505_, _12504_, _12500_);
  and (_12506_, _12502_, _11905_);
  or (_37351_, _12506_, _12505_);
  or (_12507_, _12503_, _11920_);
  and (_12508_, _12498_, _10869_);
  nor (_12509_, _12498_, _02803_);
  or (_12510_, _12509_, _12502_);
  or (_12511_, _12510_, _12508_);
  and (_37352_, _12511_, _12507_);
  nor (_12512_, _12498_, _03447_);
  and (_12513_, _12498_, _11075_);
  or (_12514_, _12513_, _12512_);
  and (_12515_, _12514_, _12503_);
  and (_12516_, _03558_, _03272_);
  and (_12517_, _12516_, _11926_);
  or (_37353_, _12517_, _12515_);
  not (_12518_, _12516_);
  or (_12519_, _12498_, \oc8051_golden_model_1.IRAM[13] [3]);
  and (_12520_, _12519_, _12518_);
  or (_12521_, _12499_, _11276_);
  and (_12522_, _12521_, _12520_);
  and (_12523_, _12516_, _11932_);
  or (_37354_, _12523_, _12522_);
  or (_12524_, _12498_, \oc8051_golden_model_1.IRAM[13] [4]);
  and (_12525_, _12524_, _12518_);
  or (_12526_, _12499_, _11490_);
  and (_12527_, _12526_, _12525_);
  and (_12528_, _12516_, _11938_);
  or (_37355_, _12528_, _12527_);
  or (_12529_, _12498_, \oc8051_golden_model_1.IRAM[13] [5]);
  and (_12530_, _12529_, _12518_);
  or (_12531_, _12499_, _11688_);
  and (_12532_, _12531_, _12530_);
  and (_12533_, _12516_, _11944_);
  or (_37356_, _12533_, _12532_);
  or (_12534_, _12498_, \oc8051_golden_model_1.IRAM[13] [6]);
  and (_12535_, _12534_, _12518_);
  or (_12536_, _12499_, _11890_);
  and (_12537_, _12536_, _12535_);
  and (_12538_, _12516_, _11950_);
  or (_37357_, _12538_, _12537_);
  or (_12539_, _12498_, \oc8051_golden_model_1.IRAM[13] [7]);
  and (_12540_, _12539_, _12518_);
  or (_12541_, _12499_, _05192_);
  and (_12542_, _12541_, _12540_);
  and (_12543_, _12516_, _05231_);
  or (_37358_, _12543_, _12542_);
  and (_12544_, _11957_, _03542_);
  or (_12545_, _12544_, \oc8051_golden_model_1.IRAM[14] [0]);
  and (_12546_, _04395_, _03558_);
  not (_12547_, _12546_);
  and (_12548_, _12547_, _12545_);
  not (_12549_, _12544_);
  or (_12550_, _12549_, _10667_);
  and (_12551_, _12550_, _12548_);
  and (_12552_, _12546_, _11905_);
  or (_37362_, _12552_, _12551_);
  nand (_12553_, _04395_, _12461_);
  or (_12554_, _12553_, _11920_);
  and (_12555_, _12544_, _10869_);
  or (_12556_, _12544_, _02797_);
  nand (_12557_, _12556_, _12553_);
  or (_12558_, _12557_, _12555_);
  and (_37363_, _12558_, _12554_);
  nor (_12559_, _12544_, _03441_);
  and (_12560_, _12544_, _11075_);
  or (_12561_, _12560_, _12559_);
  and (_12562_, _12561_, _12553_);
  and (_12563_, _12546_, _11926_);
  or (_37364_, _12563_, _12562_);
  or (_12564_, _12544_, \oc8051_golden_model_1.IRAM[14] [3]);
  and (_12565_, _12564_, _12547_);
  or (_12566_, _12549_, _11276_);
  and (_12567_, _12566_, _12565_);
  and (_12568_, _12546_, _11932_);
  or (_37366_, _12568_, _12567_);
  or (_12569_, _12544_, \oc8051_golden_model_1.IRAM[14] [4]);
  and (_12570_, _12569_, _12547_);
  or (_12571_, _12549_, _11490_);
  and (_12572_, _12571_, _12570_);
  and (_12573_, _12546_, _11938_);
  or (_37367_, _12573_, _12572_);
  or (_12574_, _12544_, \oc8051_golden_model_1.IRAM[14] [5]);
  and (_12575_, _12574_, _12547_);
  or (_12576_, _12549_, _11688_);
  and (_12577_, _12576_, _12575_);
  and (_12578_, _12546_, _11944_);
  or (_37368_, _12578_, _12577_);
  or (_12579_, _12544_, \oc8051_golden_model_1.IRAM[14] [6]);
  and (_12580_, _12579_, _12547_);
  or (_12581_, _12549_, _11890_);
  and (_12582_, _12581_, _12580_);
  and (_12583_, _12546_, _11950_);
  or (_37369_, _12583_, _12582_);
  or (_12584_, _12544_, \oc8051_golden_model_1.IRAM[14] [7]);
  and (_12585_, _12584_, _12547_);
  or (_12586_, _12549_, _05192_);
  and (_12587_, _12586_, _12585_);
  and (_12588_, _12546_, _05231_);
  or (_37370_, _12588_, _12587_);
  or (_12589_, _03543_, \oc8051_golden_model_1.IRAM[15] [0]);
  and (_12590_, _12589_, _03560_);
  or (_12591_, _10667_, _03562_);
  and (_12592_, _12591_, _12590_);
  and (_12593_, _11905_, _03559_);
  or (_37373_, _12593_, _12592_);
  nand (_12594_, _12461_, _01863_);
  or (_12595_, _11920_, _12594_);
  and (_12596_, _10869_, _03543_);
  or (_12597_, _03543_, _02795_);
  nand (_12598_, _12597_, _12594_);
  or (_12599_, _12598_, _12596_);
  and (_37374_, _12599_, _12595_);
  nor (_12600_, _03543_, _03439_);
  and (_12601_, _11075_, _03543_);
  or (_12602_, _12601_, _12600_);
  and (_12603_, _12602_, _12594_);
  and (_12604_, _11926_, _03559_);
  or (_37375_, _12604_, _12603_);
  or (_12605_, _03543_, \oc8051_golden_model_1.IRAM[15] [3]);
  and (_12606_, _12605_, _03560_);
  or (_12607_, _11276_, _03562_);
  and (_12608_, _12607_, _12606_);
  and (_12609_, _11932_, _03559_);
  or (_37377_, _12609_, _12608_);
  or (_12610_, _03543_, \oc8051_golden_model_1.IRAM[15] [4]);
  and (_12611_, _12610_, _03560_);
  or (_12612_, _11490_, _03562_);
  and (_12613_, _12612_, _12611_);
  and (_12614_, _11938_, _03559_);
  or (_37378_, _12614_, _12613_);
  or (_12615_, _03543_, \oc8051_golden_model_1.IRAM[15] [5]);
  and (_12616_, _12615_, _03560_);
  or (_12617_, _11688_, _03562_);
  and (_12618_, _12617_, _12616_);
  and (_12619_, _11944_, _03559_);
  or (_37379_, _12619_, _12618_);
  or (_12620_, _03543_, \oc8051_golden_model_1.IRAM[15] [6]);
  and (_12621_, _12620_, _03560_);
  or (_12622_, _11890_, _03562_);
  and (_12623_, _12622_, _12621_);
  and (_12624_, _11950_, _03559_);
  or (_37380_, _12624_, _12623_);
  nor (_12625_, _38087_, _06020_);
  nor (_12626_, _03683_, _06020_);
  and (_12627_, _10620_, _03683_);
  or (_12628_, _12627_, _12626_);
  and (_12629_, _12628_, _02167_);
  and (_12630_, _03683_, _04562_);
  or (_12631_, _12630_, _12626_);
  or (_12632_, _12631_, _01870_);
  and (_12633_, _03683_, _03028_);
  or (_12634_, _12633_, _12626_);
  or (_12635_, _12634_, _05249_);
  nor (_12636_, _04106_, _05239_);
  or (_12637_, _12636_, _12626_);
  or (_12638_, _12637_, _02814_);
  and (_12639_, _03683_, \oc8051_golden_model_1.ACC [0]);
  or (_12640_, _12639_, _12626_);
  and (_12641_, _12640_, _02817_);
  nor (_12642_, _02817_, _06020_);
  or (_12643_, _12642_, _02001_);
  or (_12644_, _12643_, _12641_);
  and (_12645_, _12644_, _02024_);
  and (_12646_, _12645_, _12638_);
  and (_12647_, _10510_, _04318_);
  nor (_12648_, _04318_, _06020_);
  or (_12649_, _12648_, _12647_);
  and (_12650_, _12649_, _02007_);
  or (_12651_, _12650_, _12646_);
  and (_12652_, _12651_, _02840_);
  and (_12653_, _12634_, _01999_);
  or (_12654_, _12653_, _02006_);
  or (_12655_, _12654_, _12652_);
  or (_12656_, _12640_, _02021_);
  and (_12657_, _12656_, _02025_);
  and (_12658_, _12657_, _12655_);
  and (_12659_, _12626_, _01997_);
  or (_12660_, _12659_, _01991_);
  or (_12661_, _12660_, _12658_);
  or (_12662_, _12637_, _02861_);
  and (_12663_, _12662_, _12661_);
  or (_12664_, _12663_, _05279_);
  nor (_12665_, _05942_, _05938_);
  nor (_12666_, _12665_, _05944_);
  or (_12667_, _12666_, _05285_);
  and (_12668_, _12667_, _02408_);
  and (_12669_, _12668_, _12664_);
  nor (_12670_, _10542_, _05995_);
  or (_12671_, _12670_, _12648_);
  and (_12672_, _12671_, _01875_);
  or (_12673_, _12672_, _05994_);
  or (_12674_, _12673_, _12669_);
  and (_12675_, _12674_, _12635_);
  or (_12676_, _12675_, _02528_);
  and (_12677_, _04952_, _03683_);
  or (_12678_, _12626_, _02888_);
  or (_12679_, _12678_, _12677_);
  and (_12680_, _12679_, _12676_);
  or (_12681_, _12680_, _01602_);
  nor (_12682_, _10600_, _05239_);
  or (_12683_, _12626_, _02043_);
  or (_12684_, _12683_, _12682_);
  and (_12685_, _12684_, _06355_);
  and (_12686_, _12685_, _12681_);
  nand (_12687_, _06353_, _01710_);
  or (_12688_, _06347_, _06322_);
  or (_12689_, _06353_, _12688_);
  and (_12690_, _12689_, _06008_);
  and (_12691_, _12690_, _12687_);
  or (_12692_, _12691_, _01869_);
  or (_12693_, _12692_, _12686_);
  and (_12694_, _12693_, _12632_);
  or (_12695_, _12694_, _02079_);
  and (_12696_, _10614_, _03683_);
  or (_12697_, _12626_, _02166_);
  or (_12698_, _12697_, _12696_);
  and (_12699_, _12698_, _02912_);
  and (_12700_, _12699_, _12695_);
  or (_12701_, _12700_, _12629_);
  and (_12702_, _12701_, _02176_);
  nand (_12703_, _12631_, _02072_);
  nor (_12704_, _12703_, _12636_);
  or (_12705_, _12704_, _12702_);
  and (_12706_, _12705_, _02907_);
  or (_12707_, _12626_, _04106_);
  and (_12708_, _12640_, _02177_);
  and (_12709_, _12708_, _12707_);
  or (_12710_, _12709_, _02071_);
  or (_12711_, _12710_, _12706_);
  nor (_12712_, _10613_, _05239_);
  or (_12713_, _12626_, _04788_);
  or (_12714_, _12713_, _12712_);
  and (_12715_, _12714_, _04793_);
  and (_12716_, _12715_, _12711_);
  nor (_12717_, _10619_, _05239_);
  or (_12718_, _12717_, _12626_);
  and (_12719_, _12718_, _02173_);
  or (_12720_, _12719_, _02201_);
  or (_12721_, _12720_, _12716_);
  or (_12722_, _12637_, _02303_);
  and (_12723_, _12722_, _01887_);
  and (_12724_, _12723_, _12721_);
  and (_12725_, _12626_, _01860_);
  or (_12726_, _12725_, _01537_);
  or (_12727_, _12726_, _12724_);
  or (_12728_, _12637_, _01538_);
  and (_12729_, _12728_, _38087_);
  and (_12730_, _12729_, _12727_);
  or (_12731_, _12730_, _12625_);
  and (_40184_, _12731_, _37580_);
  nor (_12732_, _38087_, _06014_);
  nor (_12733_, _04318_, _06014_);
  and (_12734_, _10696_, _04318_);
  or (_12735_, _12734_, _12733_);
  and (_12736_, _12735_, _01997_);
  nor (_12737_, _03683_, _06014_);
  nor (_12738_, _05239_, _02811_);
  or (_12739_, _12738_, _12737_);
  or (_12740_, _12739_, _02840_);
  or (_12741_, _03683_, \oc8051_golden_model_1.B [1]);
  and (_12742_, _10698_, _03683_);
  not (_12743_, _12742_);
  and (_12744_, _12743_, _12741_);
  or (_12745_, _12744_, _02814_);
  nand (_12746_, _03683_, _01613_);
  and (_12747_, _12746_, _12741_);
  and (_12748_, _12747_, _02817_);
  nor (_12749_, _02817_, _06014_);
  or (_12750_, _12749_, _02001_);
  or (_12751_, _12750_, _12748_);
  and (_12752_, _12751_, _02024_);
  and (_12753_, _12752_, _12745_);
  and (_12754_, _10710_, _04318_);
  or (_12755_, _12754_, _12733_);
  and (_12756_, _12755_, _02007_);
  or (_12757_, _12756_, _01999_);
  or (_12758_, _12757_, _12753_);
  and (_12759_, _12758_, _12740_);
  or (_12760_, _12759_, _02006_);
  or (_12761_, _12747_, _02021_);
  and (_12762_, _12761_, _02025_);
  and (_12763_, _12762_, _12760_);
  or (_12764_, _12763_, _12736_);
  and (_12765_, _12764_, _02861_);
  and (_12766_, _12754_, _10725_);
  or (_12767_, _12766_, _12733_);
  and (_12768_, _12767_, _01991_);
  or (_12769_, _12768_, _05279_);
  or (_12770_, _12769_, _12765_);
  nor (_12771_, _05948_, _05834_);
  nor (_12772_, _12771_, _05950_);
  or (_12773_, _12772_, _05285_);
  and (_12774_, _12773_, _02408_);
  and (_12775_, _12774_, _12770_);
  nor (_12776_, _10742_, _05995_);
  or (_12777_, _12776_, _12733_);
  and (_12778_, _12777_, _01875_);
  or (_12779_, _12778_, _05994_);
  or (_12780_, _12779_, _12775_);
  or (_12781_, _12739_, _05249_);
  and (_12782_, _12781_, _12780_);
  or (_12783_, _12782_, _02528_);
  and (_12784_, _04907_, _03683_);
  or (_12785_, _12737_, _02888_);
  or (_12786_, _12785_, _12784_);
  and (_12787_, _12786_, _02043_);
  and (_12788_, _12787_, _12783_);
  nand (_12789_, _10802_, _03683_);
  and (_12790_, _12741_, _01602_);
  and (_12791_, _12790_, _12789_);
  or (_12792_, _12791_, _06008_);
  or (_12793_, _12792_, _12788_);
  nor (_12794_, _06348_, _06346_);
  or (_12795_, _12794_, _06349_);
  nor (_12796_, _12795_, _06353_);
  and (_12797_, _06353_, _06319_);
  or (_12798_, _12797_, _12796_);
  or (_12799_, _12798_, _06355_);
  and (_12800_, _12799_, _01870_);
  and (_12801_, _12800_, _12793_);
  nand (_12802_, _03683_, _02687_);
  and (_12803_, _12802_, _01869_);
  and (_12804_, _12803_, _12741_);
  or (_12805_, _12804_, _12801_);
  and (_12806_, _12805_, _02166_);
  or (_12807_, _10816_, _05239_);
  and (_12808_, _12741_, _02079_);
  and (_12809_, _12808_, _12807_);
  or (_12810_, _12809_, _12806_);
  and (_12811_, _12810_, _02912_);
  or (_12812_, _10822_, _05239_);
  and (_12813_, _12741_, _02167_);
  and (_12814_, _12813_, _12812_);
  or (_12815_, _12814_, _12811_);
  and (_12816_, _12815_, _02176_);
  or (_12817_, _10692_, _05239_);
  and (_12818_, _12741_, _02072_);
  and (_12819_, _12818_, _12817_);
  or (_12820_, _12819_, _12816_);
  and (_12821_, _12820_, _02907_);
  or (_12822_, _12737_, _04058_);
  and (_12823_, _12747_, _02177_);
  and (_12824_, _12823_, _12822_);
  or (_12825_, _12824_, _12821_);
  and (_12826_, _12825_, _02174_);
  or (_12827_, _12746_, _04058_);
  and (_12828_, _12741_, _02173_);
  and (_12829_, _12828_, _12827_);
  or (_12830_, _12829_, _02201_);
  or (_12831_, _12802_, _04058_);
  and (_12832_, _12741_, _02071_);
  and (_12833_, _12832_, _12831_);
  or (_12834_, _12833_, _12830_);
  or (_12835_, _12834_, _12826_);
  or (_12836_, _12744_, _02303_);
  and (_12837_, _12836_, _01887_);
  and (_12838_, _12837_, _12835_);
  and (_12839_, _12735_, _01860_);
  or (_12840_, _12839_, _01537_);
  or (_12841_, _12840_, _12838_);
  or (_12842_, _12737_, _01538_);
  or (_12843_, _12842_, _12742_);
  and (_12844_, _12843_, _38087_);
  and (_12845_, _12844_, _12841_);
  or (_12846_, _12845_, _12732_);
  and (_40185_, _12846_, _37580_);
  nor (_12847_, _38087_, _06068_);
  nor (_12848_, _03683_, _06068_);
  and (_12849_, _11020_, _03683_);
  or (_12850_, _12849_, _12848_);
  and (_12851_, _12850_, _02167_);
  and (_12852_, _03683_, _04724_);
  or (_12853_, _12852_, _12848_);
  or (_12854_, _12853_, _01870_);
  nor (_12855_, _05239_, _03455_);
  or (_12856_, _12855_, _12848_);
  or (_12857_, _12856_, _05249_);
  and (_12858_, _10909_, _04318_);
  and (_12859_, _12858_, _10924_);
  nor (_12860_, _04318_, _06068_);
  or (_12861_, _12860_, _02861_);
  or (_12862_, _12861_, _12859_);
  or (_12863_, _12856_, _02840_);
  nor (_12864_, _10905_, _05239_);
  or (_12865_, _12864_, _12848_);
  or (_12866_, _12865_, _02814_);
  and (_12867_, _03683_, \oc8051_golden_model_1.ACC [2]);
  or (_12868_, _12867_, _12848_);
  and (_12869_, _12868_, _02817_);
  nor (_12870_, _02817_, _06068_);
  or (_12871_, _12870_, _02001_);
  or (_12872_, _12871_, _12869_);
  and (_12873_, _12872_, _02024_);
  and (_12874_, _12873_, _12866_);
  or (_12875_, _12860_, _12858_);
  and (_12876_, _12875_, _02007_);
  or (_12877_, _12876_, _01999_);
  or (_12878_, _12877_, _12874_);
  and (_12879_, _12878_, _12863_);
  or (_12880_, _12879_, _02006_);
  or (_12881_, _12868_, _02021_);
  and (_12882_, _12881_, _02025_);
  and (_12883_, _12882_, _12880_);
  and (_12884_, _10894_, _04318_);
  or (_12885_, _12884_, _12860_);
  and (_12886_, _12885_, _01997_);
  or (_12887_, _12886_, _01991_);
  or (_12888_, _12887_, _12883_);
  and (_12889_, _12888_, _12862_);
  or (_12890_, _12889_, _05279_);
  or (_12891_, _05952_, _05744_);
  and (_12892_, _12891_, _05954_);
  or (_12893_, _12892_, _05285_);
  and (_12894_, _12893_, _02408_);
  and (_12895_, _12894_, _12890_);
  nor (_12896_, _10942_, _05995_);
  or (_12897_, _12896_, _12860_);
  and (_12898_, _12897_, _01875_);
  or (_12899_, _12898_, _05994_);
  or (_12900_, _12899_, _12895_);
  and (_12901_, _12900_, _12857_);
  or (_12902_, _12901_, _02528_);
  and (_12903_, _05043_, _03683_);
  or (_12904_, _12848_, _02888_);
  or (_12905_, _12904_, _12903_);
  and (_12906_, _12905_, _12902_);
  or (_12907_, _12906_, _01602_);
  nor (_12908_, _11000_, _05239_);
  or (_12909_, _12848_, _02043_);
  or (_12910_, _12909_, _12908_);
  and (_12911_, _12910_, _06355_);
  and (_12912_, _12911_, _12907_);
  nand (_12913_, _06353_, _06309_);
  nor (_12914_, _06349_, _06320_);
  not (_12915_, _12914_);
  and (_12916_, _12915_, _06312_);
  nor (_12917_, _12915_, _06312_);
  nor (_12918_, _12917_, _12916_);
  or (_12919_, _12918_, _06353_);
  and (_12920_, _12919_, _06008_);
  and (_12921_, _12920_, _12913_);
  or (_12922_, _12921_, _01869_);
  or (_12923_, _12922_, _12912_);
  and (_12924_, _12923_, _12854_);
  or (_12925_, _12924_, _02079_);
  and (_12926_, _11014_, _03683_);
  or (_12927_, _12848_, _02166_);
  or (_12928_, _12927_, _12926_);
  and (_12929_, _12928_, _02912_);
  and (_12930_, _12929_, _12925_);
  or (_12931_, _12930_, _12851_);
  and (_12932_, _12931_, _02176_);
  or (_12933_, _12848_, _04156_);
  and (_12934_, _12853_, _02072_);
  and (_12935_, _12934_, _12933_);
  or (_12936_, _12935_, _12932_);
  and (_12937_, _12936_, _02907_);
  and (_12938_, _12868_, _02177_);
  and (_12939_, _12938_, _12933_);
  or (_12940_, _12939_, _02071_);
  or (_12941_, _12940_, _12937_);
  nor (_12942_, _11013_, _05239_);
  or (_12943_, _12848_, _04788_);
  or (_12944_, _12943_, _12942_);
  and (_12945_, _12944_, _04793_);
  and (_12946_, _12945_, _12941_);
  nor (_12947_, _11019_, _05239_);
  or (_12948_, _12947_, _12848_);
  and (_12949_, _12948_, _02173_);
  or (_12950_, _12949_, _02201_);
  or (_12951_, _12950_, _12946_);
  or (_12952_, _12865_, _02303_);
  and (_12953_, _12952_, _01887_);
  and (_12954_, _12953_, _12951_);
  and (_12955_, _12885_, _01860_);
  or (_12956_, _12955_, _01537_);
  or (_12957_, _12956_, _12954_);
  and (_12958_, _11072_, _03683_);
  or (_12959_, _12848_, _01538_);
  or (_12960_, _12959_, _12958_);
  and (_12961_, _12960_, _38087_);
  and (_12962_, _12961_, _12957_);
  or (_12963_, _12962_, _12847_);
  and (_40186_, _12963_, _37580_);
  nor (_12964_, _38087_, _06096_);
  nor (_12965_, _03683_, _06096_);
  and (_12966_, _11094_, _03683_);
  or (_12967_, _12966_, _12965_);
  and (_12968_, _12967_, _02167_);
  and (_12969_, _03683_, _04678_);
  or (_12970_, _12969_, _12965_);
  or (_12971_, _12970_, _01870_);
  nor (_12972_, _11206_, _05239_);
  or (_12973_, _12972_, _12965_);
  and (_12974_, _12973_, _01602_);
  nor (_12975_, _04318_, _06096_);
  and (_12976_, _11098_, _04318_);
  or (_12977_, _12976_, _12975_);
  or (_12978_, _12975_, _11127_);
  and (_12979_, _12978_, _12977_);
  or (_12980_, _12979_, _02861_);
  nor (_12981_, _11101_, _05239_);
  or (_12982_, _12981_, _12965_);
  or (_12983_, _12982_, _02814_);
  and (_12984_, _03683_, \oc8051_golden_model_1.ACC [3]);
  or (_12985_, _12984_, _12965_);
  and (_12986_, _12985_, _02817_);
  nor (_12987_, _02817_, _06096_);
  or (_12988_, _12987_, _02001_);
  or (_12989_, _12988_, _12986_);
  and (_12990_, _12989_, _02024_);
  and (_12991_, _12990_, _12983_);
  and (_12992_, _12977_, _02007_);
  or (_12993_, _12992_, _01999_);
  or (_12994_, _12993_, _12991_);
  nor (_12995_, _05239_, _03268_);
  or (_12996_, _12995_, _12965_);
  or (_12997_, _12996_, _02840_);
  and (_12998_, _12997_, _12994_);
  or (_12999_, _12998_, _02006_);
  or (_13000_, _12985_, _02021_);
  and (_13001_, _13000_, _02025_);
  and (_13002_, _13001_, _12999_);
  and (_13003_, _11096_, _04318_);
  or (_13004_, _13003_, _12975_);
  and (_13005_, _13004_, _01997_);
  or (_13006_, _13005_, _01991_);
  or (_13007_, _13006_, _13002_);
  and (_13008_, _13007_, _12980_);
  or (_13009_, _13008_, _05279_);
  nor (_13010_, _05958_, _05638_);
  nor (_13011_, _13010_, _05960_);
  or (_13012_, _13011_, _05285_);
  and (_13013_, _13012_, _02408_);
  and (_13014_, _13013_, _13009_);
  nor (_13015_, _11145_, _05995_);
  or (_13016_, _13015_, _12975_);
  and (_13017_, _13016_, _01875_);
  or (_13018_, _13017_, _05994_);
  or (_13019_, _13018_, _13014_);
  or (_13020_, _12996_, _05249_);
  and (_13021_, _13020_, _13019_);
  or (_13022_, _13021_, _02528_);
  and (_13023_, _04998_, _03683_);
  or (_13024_, _12965_, _02888_);
  or (_13025_, _13024_, _13023_);
  and (_13026_, _13025_, _02043_);
  and (_13027_, _13026_, _13022_);
  or (_13028_, _13027_, _12974_);
  and (_13029_, _13028_, _06355_);
  nor (_13030_, _12916_, _06311_);
  nor (_13031_, _13030_, _06304_);
  and (_13032_, _13030_, _06304_);
  or (_13033_, _13032_, _13031_);
  or (_13034_, _13033_, _06353_);
  not (_13035_, _06353_);
  or (_13036_, _13035_, _06301_);
  and (_13037_, _13036_, _06008_);
  and (_13038_, _13037_, _13034_);
  or (_13039_, _13038_, _01869_);
  or (_13040_, _13039_, _13029_);
  and (_13041_, _13040_, _12971_);
  or (_13042_, _13041_, _02079_);
  and (_13043_, _11222_, _03683_);
  or (_13044_, _12965_, _02166_);
  or (_13045_, _13044_, _13043_);
  and (_13046_, _13045_, _02912_);
  and (_13047_, _13046_, _13042_);
  or (_13048_, _13047_, _12968_);
  and (_13049_, _13048_, _02176_);
  or (_13050_, _12965_, _04014_);
  and (_13051_, _12970_, _02072_);
  and (_13052_, _13051_, _13050_);
  or (_13053_, _13052_, _13049_);
  and (_13054_, _13053_, _02907_);
  and (_13055_, _12985_, _02177_);
  and (_13056_, _13055_, _13050_);
  or (_13057_, _13056_, _02071_);
  or (_13058_, _13057_, _13054_);
  nor (_13059_, _11220_, _05239_);
  or (_13060_, _12965_, _04788_);
  or (_13061_, _13060_, _13059_);
  and (_13062_, _13061_, _04793_);
  and (_13063_, _13062_, _13058_);
  nor (_13064_, _11093_, _05239_);
  or (_13065_, _13064_, _12965_);
  and (_13066_, _13065_, _02173_);
  or (_13067_, _13066_, _02201_);
  or (_13068_, _13067_, _13063_);
  or (_13069_, _12982_, _02303_);
  and (_13070_, _13069_, _01887_);
  and (_13071_, _13070_, _13068_);
  and (_13072_, _13004_, _01860_);
  or (_13073_, _13072_, _01537_);
  or (_13074_, _13073_, _13071_);
  and (_13075_, _11273_, _03683_);
  or (_13076_, _12965_, _01538_);
  or (_13077_, _13076_, _13075_);
  and (_13078_, _13077_, _38087_);
  and (_13079_, _13078_, _13074_);
  or (_13080_, _13079_, _12964_);
  and (_40187_, _13080_, _37580_);
  nor (_13081_, _38087_, _06151_);
  nor (_13082_, _03683_, _06151_);
  and (_13083_, _11431_, _03683_);
  or (_13084_, _13083_, _13082_);
  and (_13085_, _13084_, _02167_);
  and (_13086_, _04694_, _03683_);
  or (_13087_, _13086_, _13082_);
  or (_13088_, _13087_, _01870_);
  nor (_13089_, _11411_, _05239_);
  or (_13090_, _13089_, _13082_);
  and (_13091_, _13090_, _01602_);
  nor (_13092_, _04211_, _05239_);
  or (_13093_, _13092_, _13082_);
  or (_13094_, _13093_, _05249_);
  nor (_13095_, _04318_, _06151_);
  and (_13096_, _11301_, _04318_);
  or (_13097_, _13096_, _13095_);
  and (_13098_, _13097_, _01997_);
  nor (_13099_, _11317_, _05239_);
  or (_13100_, _13099_, _13082_);
  or (_13101_, _13100_, _02814_);
  and (_13102_, _03683_, \oc8051_golden_model_1.ACC [4]);
  or (_13103_, _13102_, _13082_);
  and (_13104_, _13103_, _02817_);
  nor (_13105_, _02817_, _06151_);
  or (_13106_, _13105_, _02001_);
  or (_13107_, _13106_, _13104_);
  and (_13108_, _13107_, _02024_);
  and (_13109_, _13108_, _13101_);
  and (_13110_, _11303_, _04318_);
  or (_13111_, _13110_, _13095_);
  and (_13112_, _13111_, _02007_);
  or (_13113_, _13112_, _01999_);
  or (_13114_, _13113_, _13109_);
  or (_13115_, _13093_, _02840_);
  and (_13116_, _13115_, _13114_);
  or (_13117_, _13116_, _02006_);
  or (_13118_, _13103_, _02021_);
  and (_13119_, _13118_, _02025_);
  and (_13120_, _13119_, _13117_);
  or (_13121_, _13120_, _13098_);
  and (_13122_, _13121_, _02861_);
  or (_13123_, _13095_, _11334_);
  and (_13124_, _13123_, _01991_);
  and (_13125_, _13124_, _13111_);
  or (_13126_, _13125_, _05279_);
  or (_13127_, _13126_, _13122_);
  or (_13128_, _05966_, _05962_);
  and (_13129_, _13128_, _05968_);
  or (_13130_, _13129_, _05285_);
  and (_13131_, _13130_, _02408_);
  and (_13132_, _13131_, _13127_);
  nor (_13133_, _11299_, _05995_);
  or (_13134_, _13133_, _13095_);
  and (_13135_, _13134_, _01875_);
  or (_13136_, _13135_, _05994_);
  or (_13137_, _13136_, _13132_);
  and (_13138_, _13137_, _13094_);
  or (_13139_, _13138_, _02528_);
  and (_13140_, _05135_, _03683_);
  or (_13141_, _13082_, _02888_);
  or (_13142_, _13141_, _13140_);
  and (_13143_, _13142_, _02043_);
  and (_13144_, _13143_, _13139_);
  or (_13145_, _13144_, _13091_);
  and (_13146_, _13145_, _06355_);
  or (_13147_, _13035_, _06293_);
  nor (_13148_, _13030_, _06302_);
  or (_13149_, _13148_, _06303_);
  nand (_13150_, _13149_, _06340_);
  or (_13151_, _13149_, _06340_);
  and (_13152_, _13151_, _13150_);
  or (_13153_, _13152_, _06353_);
  and (_13154_, _13153_, _06008_);
  and (_13155_, _13154_, _13147_);
  or (_13156_, _13155_, _01869_);
  or (_13157_, _13156_, _13146_);
  and (_13158_, _13157_, _13088_);
  or (_13159_, _13158_, _02079_);
  and (_13160_, _11425_, _03683_);
  or (_13161_, _13082_, _02166_);
  or (_13162_, _13161_, _13160_);
  and (_13163_, _13162_, _02912_);
  and (_13164_, _13163_, _13159_);
  or (_13165_, _13164_, _13085_);
  and (_13166_, _13165_, _02176_);
  or (_13167_, _13082_, _04258_);
  and (_13168_, _13087_, _02072_);
  and (_13169_, _13168_, _13167_);
  or (_13170_, _13169_, _13166_);
  and (_13171_, _13170_, _02907_);
  and (_13172_, _13103_, _02177_);
  and (_13173_, _13172_, _13167_);
  or (_13174_, _13173_, _02071_);
  or (_13175_, _13174_, _13171_);
  nor (_13176_, _11424_, _05239_);
  or (_13177_, _13082_, _04788_);
  or (_13178_, _13177_, _13176_);
  and (_13179_, _13178_, _04793_);
  and (_13180_, _13179_, _13175_);
  nor (_13181_, _11430_, _05239_);
  or (_13182_, _13181_, _13082_);
  and (_13183_, _13182_, _02173_);
  or (_13184_, _13183_, _02201_);
  or (_13185_, _13184_, _13180_);
  or (_13186_, _13100_, _02303_);
  and (_13187_, _13186_, _01887_);
  and (_13188_, _13187_, _13185_);
  and (_13189_, _13097_, _01860_);
  or (_13190_, _13189_, _01537_);
  or (_13191_, _13190_, _13188_);
  and (_13192_, _11487_, _03683_);
  or (_13193_, _13082_, _01538_);
  or (_13194_, _13193_, _13192_);
  and (_13195_, _13194_, _38087_);
  and (_13196_, _13195_, _13191_);
  or (_13197_, _13196_, _13081_);
  and (_40188_, _13197_, _37580_);
  nor (_13198_, _38087_, _06140_);
  nor (_13199_, _03683_, _06140_);
  and (_13200_, _11635_, _03683_);
  or (_13201_, _13200_, _13199_);
  and (_13202_, _13201_, _02167_);
  and (_13203_, _04672_, _03683_);
  or (_13204_, _13203_, _13199_);
  or (_13205_, _13204_, _01870_);
  nor (_13206_, _11615_, _05239_);
  or (_13207_, _13206_, _13199_);
  and (_13208_, _13207_, _01602_);
  nor (_13209_, _03916_, _05239_);
  or (_13210_, _13209_, _13199_);
  or (_13211_, _13210_, _05249_);
  nor (_13212_, _04318_, _06140_);
  and (_13213_, _11508_, _04318_);
  or (_13214_, _13213_, _13212_);
  and (_13215_, _13214_, _01997_);
  nor (_13216_, _11525_, _05239_);
  or (_13217_, _13216_, _13199_);
  or (_13218_, _13217_, _02814_);
  and (_13219_, _03683_, \oc8051_golden_model_1.ACC [5]);
  or (_13220_, _13219_, _13199_);
  and (_13221_, _13220_, _02817_);
  nor (_13222_, _02817_, _06140_);
  or (_13223_, _13222_, _02001_);
  or (_13224_, _13223_, _13221_);
  and (_13225_, _13224_, _02024_);
  and (_13226_, _13225_, _13218_);
  and (_13227_, _11510_, _04318_);
  or (_13228_, _13227_, _13212_);
  and (_13229_, _13228_, _02007_);
  or (_13230_, _13229_, _01999_);
  or (_13231_, _13230_, _13226_);
  or (_13232_, _13210_, _02840_);
  and (_13233_, _13232_, _13231_);
  or (_13234_, _13233_, _02006_);
  or (_13235_, _13220_, _02021_);
  and (_13236_, _13235_, _02025_);
  and (_13237_, _13236_, _13234_);
  or (_13238_, _13237_, _13215_);
  and (_13239_, _13238_, _02861_);
  or (_13240_, _13212_, _11542_);
  and (_13241_, _13240_, _01991_);
  and (_13242_, _13241_, _13228_);
  or (_13243_, _13242_, _05279_);
  or (_13244_, _13243_, _13239_);
  or (_13245_, _05490_, _05489_);
  not (_13246_, _13245_);
  nor (_13247_, _13246_, _05970_);
  and (_13248_, _13246_, _05970_);
  or (_13249_, _13248_, _13247_);
  or (_13250_, _13249_, _05285_);
  and (_13251_, _13250_, _02408_);
  and (_13252_, _13251_, _13244_);
  nor (_13253_, _11506_, _05995_);
  or (_13254_, _13253_, _13212_);
  and (_13255_, _13254_, _01875_);
  or (_13256_, _13255_, _05994_);
  or (_13257_, _13256_, _13252_);
  and (_13258_, _13257_, _13211_);
  or (_13259_, _13258_, _02528_);
  and (_13260_, _05090_, _03683_);
  or (_13261_, _13199_, _02888_);
  or (_13262_, _13261_, _13260_);
  and (_13263_, _13262_, _02043_);
  and (_13264_, _13263_, _13259_);
  or (_13265_, _13264_, _13208_);
  and (_13266_, _13265_, _06355_);
  or (_13267_, _13035_, _06285_);
  not (_13268_, _06331_);
  and (_13269_, _13150_, _13268_);
  nor (_13270_, _13269_, _06341_);
  and (_13271_, _13269_, _06341_);
  or (_13272_, _13271_, _13270_);
  or (_13273_, _13272_, _06353_);
  and (_13274_, _13273_, _06008_);
  and (_13275_, _13274_, _13267_);
  or (_13276_, _13275_, _01869_);
  or (_13277_, _13276_, _13266_);
  and (_13278_, _13277_, _13205_);
  or (_13279_, _13278_, _02079_);
  and (_13280_, _11629_, _03683_);
  or (_13281_, _13199_, _02166_);
  or (_13282_, _13281_, _13280_);
  and (_13283_, _13282_, _02912_);
  and (_13284_, _13283_, _13279_);
  or (_13285_, _13284_, _13202_);
  and (_13286_, _13285_, _02176_);
  or (_13287_, _13199_, _03965_);
  and (_13288_, _13204_, _02072_);
  and (_13289_, _13288_, _13287_);
  or (_13290_, _13289_, _13286_);
  and (_13291_, _13290_, _02907_);
  and (_13292_, _13220_, _02177_);
  and (_13293_, _13292_, _13287_);
  or (_13294_, _13293_, _02071_);
  or (_13295_, _13294_, _13291_);
  nor (_13296_, _11628_, _05239_);
  or (_13297_, _13199_, _04788_);
  or (_13298_, _13297_, _13296_);
  and (_13299_, _13298_, _04793_);
  and (_13300_, _13299_, _13295_);
  nor (_13301_, _11634_, _05239_);
  or (_13302_, _13301_, _13199_);
  and (_13303_, _13302_, _02173_);
  or (_13304_, _13303_, _02201_);
  or (_13305_, _13304_, _13300_);
  or (_13306_, _13217_, _02303_);
  and (_13307_, _13306_, _01887_);
  and (_13308_, _13307_, _13305_);
  and (_13309_, _13214_, _01860_);
  or (_13310_, _13309_, _01537_);
  or (_13311_, _13310_, _13308_);
  and (_13312_, _11685_, _03683_);
  or (_13313_, _13199_, _01538_);
  or (_13314_, _13313_, _13312_);
  and (_13315_, _13314_, _38087_);
  and (_13316_, _13315_, _13311_);
  or (_13317_, _13316_, _13198_);
  and (_40189_, _13317_, _37580_);
  nor (_13318_, _38087_, _06270_);
  nor (_13319_, _03683_, _06270_);
  and (_13320_, _11709_, _03683_);
  or (_13321_, _13320_, _13319_);
  and (_13322_, _13321_, _02167_);
  and (_13323_, _09920_, _03683_);
  or (_13324_, _13323_, _13319_);
  or (_13325_, _13324_, _01870_);
  nor (_13326_, _11820_, _05239_);
  or (_13327_, _13326_, _13319_);
  and (_13328_, _13327_, _01602_);
  nor (_13329_, _03808_, _05239_);
  or (_13330_, _13329_, _13319_);
  or (_13331_, _13330_, _05249_);
  nor (_13332_, _04318_, _06270_);
  and (_13333_, _11715_, _04318_);
  or (_13334_, _13333_, _13332_);
  and (_13335_, _13334_, _01997_);
  nor (_13336_, _11730_, _05239_);
  or (_13337_, _13336_, _13319_);
  or (_13338_, _13337_, _02814_);
  and (_13339_, _03683_, \oc8051_golden_model_1.ACC [6]);
  or (_13340_, _13339_, _13319_);
  and (_13341_, _13340_, _02817_);
  nor (_13342_, _02817_, _06270_);
  or (_13343_, _13342_, _02001_);
  or (_13344_, _13343_, _13341_);
  and (_13345_, _13344_, _02024_);
  and (_13346_, _13345_, _13338_);
  and (_13347_, _11717_, _04318_);
  or (_13348_, _13347_, _13332_);
  and (_13349_, _13348_, _02007_);
  or (_13350_, _13349_, _01999_);
  or (_13351_, _13350_, _13346_);
  or (_13352_, _13330_, _02840_);
  and (_13353_, _13352_, _13351_);
  or (_13354_, _13353_, _02006_);
  or (_13355_, _13340_, _02021_);
  and (_13356_, _13355_, _02025_);
  and (_13357_, _13356_, _13354_);
  or (_13358_, _13357_, _13335_);
  and (_13359_, _13358_, _02861_);
  or (_13360_, _13332_, _11747_);
  and (_13361_, _13360_, _01991_);
  and (_13362_, _13361_, _13348_);
  or (_13363_, _13362_, _05279_);
  or (_13364_, _13363_, _13359_);
  nor (_13365_, _05982_, _05974_);
  nor (_13366_, _13365_, _05984_);
  or (_13367_, _13366_, _05285_);
  and (_13368_, _13367_, _02408_);
  and (_13369_, _13368_, _13364_);
  nor (_13370_, _11713_, _05995_);
  or (_13371_, _13370_, _13332_);
  and (_13372_, _13371_, _01875_);
  or (_13373_, _13372_, _05994_);
  or (_13374_, _13373_, _13369_);
  and (_13375_, _13374_, _13331_);
  or (_13376_, _13375_, _02528_);
  and (_13377_, _04861_, _03683_);
  or (_13378_, _13319_, _02888_);
  or (_13379_, _13378_, _13377_);
  and (_13380_, _13379_, _02043_);
  and (_13381_, _13380_, _13376_);
  or (_13382_, _13381_, _13328_);
  and (_13383_, _13382_, _06355_);
  or (_13384_, _13035_, _06276_);
  nor (_13385_, _13269_, _06286_);
  or (_13386_, _13385_, _06287_);
  or (_13387_, _13386_, _06343_);
  nand (_13388_, _13386_, _06343_);
  and (_13389_, _13388_, _13387_);
  or (_13390_, _13389_, _06353_);
  and (_13391_, _13390_, _06008_);
  and (_13392_, _13391_, _13384_);
  or (_13393_, _13392_, _01869_);
  or (_13394_, _13393_, _13383_);
  and (_13395_, _13394_, _13325_);
  or (_13396_, _13395_, _02079_);
  and (_13397_, _11835_, _03683_);
  or (_13398_, _13319_, _02166_);
  or (_13399_, _13398_, _13397_);
  and (_13400_, _13399_, _02912_);
  and (_13401_, _13400_, _13396_);
  or (_13402_, _13401_, _13322_);
  and (_13403_, _13402_, _02176_);
  or (_13404_, _13319_, _03863_);
  and (_13405_, _13324_, _02072_);
  and (_13406_, _13405_, _13404_);
  or (_13407_, _13406_, _13403_);
  and (_13408_, _13407_, _02907_);
  and (_13409_, _13340_, _02177_);
  and (_13410_, _13409_, _13404_);
  or (_13411_, _13410_, _02071_);
  or (_13412_, _13411_, _13408_);
  nor (_13413_, _11833_, _05239_);
  or (_13414_, _13319_, _04788_);
  or (_13415_, _13414_, _13413_);
  and (_13416_, _13415_, _04793_);
  and (_13417_, _13416_, _13412_);
  nor (_13418_, _11708_, _05239_);
  or (_13419_, _13418_, _13319_);
  and (_13420_, _13419_, _02173_);
  or (_13421_, _13420_, _02201_);
  or (_13422_, _13421_, _13417_);
  or (_13423_, _13337_, _02303_);
  and (_13424_, _13423_, _01887_);
  and (_13425_, _13424_, _13422_);
  and (_13426_, _13334_, _01860_);
  or (_13427_, _13426_, _01537_);
  or (_13428_, _13427_, _13425_);
  and (_13429_, _11887_, _03683_);
  or (_13430_, _13319_, _01538_);
  or (_13431_, _13430_, _13429_);
  and (_13432_, _13431_, _38087_);
  and (_13433_, _13432_, _13428_);
  or (_13434_, _13433_, _13318_);
  and (_40190_, _13434_, _37580_);
  nor (_13435_, _38087_, _01710_);
  nand (_13436_, _07304_, _04776_);
  nor (_13437_, _06591_, _01710_);
  nor (_13438_, _13437_, _06592_);
  nand (_13439_, _07114_, _13438_);
  and (_13440_, _03042_, _01710_);
  nand (_13441_, _07051_, _13440_);
  not (_13442_, _06433_);
  not (_13443_, _02345_);
  and (_13444_, _01972_, _01631_);
  not (_13445_, _13444_);
  and (_13446_, _06454_, _01631_);
  or (_13447_, _13446_, _02689_);
  nor (_13448_, _13447_, _02696_);
  and (_13449_, _13448_, _13445_);
  and (_13450_, _13449_, _13443_);
  nor (_13451_, _13450_, _13442_);
  nor (_13452_, _03680_, _01710_);
  and (_13453_, _03680_, _03028_);
  nor (_13454_, _13453_, _13452_);
  nand (_13455_, _13454_, _05994_);
  or (_13456_, _06613_, _03028_);
  nor (_13457_, _06620_, _01883_);
  or (_13458_, _13457_, _04952_);
  nor (_13459_, _06850_, _06618_);
  and (_13460_, _06623_, _03028_);
  not (_13461_, _06623_);
  and (_13462_, _06625_, _01710_);
  nor (_13463_, _06625_, _01710_);
  or (_13464_, _13463_, _06620_);
  or (_13465_, _13464_, _13462_);
  and (_13466_, _13465_, _13461_);
  or (_13467_, _13466_, _13460_);
  and (_13468_, _13467_, _06618_);
  or (_13469_, _13468_, _13459_);
  and (_13470_, _13469_, _10136_);
  or (_13471_, _13470_, _01883_);
  and (_13472_, _13471_, _02814_);
  and (_13473_, _13472_, _13458_);
  nor (_13474_, _04106_, _06472_);
  nor (_13475_, _13474_, _13452_);
  nor (_13476_, _13475_, _02814_);
  or (_13477_, _13476_, _02007_);
  or (_13478_, _13477_, _13473_);
  nor (_13479_, _04326_, _01710_);
  and (_13480_, _10510_, _04326_);
  nor (_13481_, _13480_, _13479_);
  nand (_13482_, _13481_, _02007_);
  and (_13483_, _13482_, _02840_);
  and (_13484_, _13483_, _13478_);
  nor (_13485_, _13454_, _02840_);
  or (_13486_, _13485_, _06614_);
  or (_13487_, _13486_, _13484_);
  and (_13488_, _13487_, _13456_);
  or (_13489_, _13488_, _02850_);
  or (_13490_, _04952_, _06675_);
  and (_13491_, _13490_, _02021_);
  and (_13492_, _13491_, _13489_);
  nor (_13493_, _06850_, _02021_);
  or (_13494_, _13493_, _06679_);
  or (_13495_, _13494_, _13492_);
  nand (_13496_, _06679_, _06085_);
  and (_13497_, _13496_, _13495_);
  or (_13498_, _13497_, _01997_);
  or (_13499_, _13452_, _02025_);
  and (_13500_, _13499_, _02861_);
  and (_13501_, _13500_, _13498_);
  nor (_13502_, _13475_, _02861_);
  or (_13503_, _13502_, _05279_);
  or (_13504_, _13503_, _13501_);
  not (_13505_, _05900_);
  nand (_13506_, _13505_, _05279_);
  and (_13507_, _13506_, _13504_);
  or (_13508_, _13507_, _06699_);
  nor (_13509_, _06752_, _01710_);
  nor (_13510_, _13509_, _06753_);
  nand (_13511_, _13510_, _06699_);
  and (_13512_, _13511_, _08245_);
  and (_13513_, _13512_, _13508_);
  nor (_13514_, _08245_, _13438_);
  or (_13515_, _13514_, _01963_);
  or (_13516_, _13515_, _13513_);
  nor (_13517_, _06931_, _01710_);
  nor (_13518_, _13517_, _06932_);
  nand (_13519_, _13518_, _01963_);
  and (_13520_, _13519_, _13516_);
  or (_13521_, _13520_, _06476_);
  and (_13522_, _06526_, _01710_);
  or (_13523_, _13522_, _07186_);
  nand (_13524_, _13523_, _06476_);
  and (_13525_, _13524_, _13521_);
  or (_13526_, _13525_, _01549_);
  nand (_13527_, _02441_, _01549_);
  and (_13528_, _13527_, _02408_);
  and (_13529_, _13528_, _13526_);
  nor (_13530_, _10542_, _06958_);
  nor (_13531_, _13530_, _13479_);
  nor (_13532_, _13531_, _02408_);
  or (_13533_, _13532_, _05994_);
  or (_13534_, _13533_, _13529_);
  and (_13535_, _13534_, _13455_);
  or (_13536_, _13535_, _02528_);
  and (_13537_, _04952_, _03680_);
  nor (_13538_, _13537_, _13452_);
  nand (_13539_, _13538_, _02528_);
  and (_13540_, _13539_, _02043_);
  and (_13541_, _13540_, _13536_);
  nor (_13542_, _10600_, _06472_);
  nor (_13543_, _13542_, _13452_);
  nor (_13544_, _13543_, _02043_);
  or (_13545_, _13544_, _06008_);
  or (_13546_, _13545_, _13541_);
  nand (_13547_, _06353_, _06008_);
  and (_13548_, _13547_, _13546_);
  and (_13549_, _13548_, _01609_);
  nor (_13550_, _02441_, _01609_);
  or (_13551_, _13550_, _01869_);
  or (_13552_, _13551_, _13549_);
  and (_13553_, _03680_, _04562_);
  nor (_13554_, _13553_, _13452_);
  nand (_13555_, _13554_, _01869_);
  and (_13556_, _13555_, _06985_);
  and (_13557_, _13556_, _13552_);
  nor (_13558_, _06985_, _02441_);
  or (_13559_, _13558_, _06990_);
  or (_13560_, _13559_, _13557_);
  nor (_13561_, _13440_, _06433_);
  nand (_13562_, _06994_, _13561_);
  nand (_13563_, _13562_, _06996_);
  and (_13564_, _13563_, _13560_);
  or (_13565_, _06999_, _13561_);
  and (_13566_, _13565_, _07002_);
  or (_13567_, _13566_, _13564_);
  not (_13568_, _13561_);
  nand (_13569_, _06999_, _13568_);
  and (_13570_, _13569_, _07006_);
  and (_13571_, _13570_, _13567_);
  nor (_13572_, _04952_, \oc8051_golden_model_1.ACC [0]);
  nor (_13573_, _07234_, _13572_);
  and (_13574_, _13573_, _02579_);
  or (_13575_, _13574_, _02168_);
  or (_13576_, _13575_, _13571_);
  or (_13577_, _10620_, _07014_);
  and (_13578_, _13577_, _07013_);
  and (_13579_, _13578_, _13576_);
  and (_13580_, _07012_, _08661_);
  or (_13581_, _13580_, _02079_);
  or (_13582_, _13581_, _13579_);
  and (_13583_, _10614_, _03680_);
  nor (_13584_, _13583_, _13452_);
  nand (_13585_, _13584_, _02079_);
  and (_13586_, _13585_, _02912_);
  and (_13587_, _13586_, _13582_);
  and (_13588_, _13452_, _02167_);
  or (_13589_, _13588_, _02390_);
  or (_13590_, _13589_, _13587_);
  or (_13591_, _06433_, _02344_);
  and (_13592_, _13591_, _13450_);
  and (_13593_, _13592_, _13590_);
  nor (_13594_, _13593_, _13451_);
  nor (_13595_, _13594_, _07031_);
  and (_13596_, _07031_, _07234_);
  or (_13597_, _13596_, _02178_);
  or (_13598_, _13597_, _13595_);
  or (_13599_, _10618_, _07035_);
  and (_13600_, _13599_, _07046_);
  and (_13601_, _13600_, _13598_);
  and (_13602_, _07040_, _07323_);
  or (_13603_, _13602_, _13601_);
  and (_13604_, _13603_, _02176_);
  nor (_13605_, _13554_, _13474_);
  and (_13606_, _13605_, _02072_);
  or (_13607_, _13606_, _07051_);
  or (_13608_, _13607_, _13604_);
  and (_13609_, _13608_, _13441_);
  or (_13610_, _13609_, _07055_);
  nand (_13611_, _07055_, _13440_);
  and (_13612_, _13611_, _07060_);
  and (_13613_, _13612_, _13610_);
  nor (_13614_, _13440_, _07060_);
  or (_13615_, _13614_, _06462_);
  or (_13616_, _13615_, _13613_);
  nand (_13617_, _13572_, _06462_);
  and (_13618_, _13617_, _02172_);
  and (_13619_, _13618_, _13616_);
  nor (_13620_, _10619_, _02172_);
  or (_13621_, _13620_, _07069_);
  or (_13622_, _13621_, _13619_);
  nand (_13623_, _07069_, _08660_);
  and (_13624_, _13623_, _13622_);
  or (_13625_, _13624_, _02071_);
  nor (_13626_, _10613_, _06472_);
  nor (_13627_, _13626_, _13452_);
  nand (_13628_, _13627_, _02071_);
  and (_13629_, _13628_, _07084_);
  and (_13630_, _13629_, _13625_);
  nor (_13631_, _07083_, _13510_);
  nor (_13632_, _07081_, _13510_);
  or (_13633_, _13632_, _07114_);
  or (_13634_, _13633_, _13631_);
  or (_13635_, _13634_, _13630_);
  and (_13636_, _13635_, _13439_);
  or (_13637_, _13636_, _02164_);
  nand (_13638_, _13518_, _02164_);
  and (_13639_, _13638_, _07177_);
  and (_13640_, _13639_, _13637_);
  nor (_13641_, _07177_, _13523_);
  or (_13642_, _13641_, _07175_);
  or (_13643_, _13642_, _13640_);
  nand (_13644_, _07175_, _06518_);
  and (_13645_, _13644_, _06451_);
  and (_13646_, _13645_, _06457_);
  and (_13647_, _13646_, _13643_);
  and (_13648_, _13561_, _06459_);
  or (_13649_, _13648_, _07210_);
  or (_13650_, _13649_, _13647_);
  or (_13651_, _07212_, _13573_);
  and (_13652_, _13651_, _13650_);
  or (_13653_, _13652_, _01890_);
  nand (_13654_, _08622_, _01890_);
  and (_13655_, _13654_, _07256_);
  and (_13656_, _13655_, _13653_);
  and (_13657_, _07253_, _08661_);
  or (_13658_, _13657_, _07304_);
  or (_13659_, _13658_, _13656_);
  and (_13660_, _13659_, _13436_);
  or (_13661_, _13660_, _02201_);
  nand (_13662_, _13475_, _02201_);
  and (_13663_, _13662_, _07346_);
  and (_13664_, _13663_, _13661_);
  nor (_13665_, _07350_, _01710_);
  nor (_13666_, _13665_, _10442_);
  or (_13667_, _13666_, _13664_);
  nand (_13668_, _07350_, _01613_);
  and (_13669_, _13668_, _01887_);
  and (_13670_, _13669_, _13667_);
  and (_13671_, _13452_, _01860_);
  or (_13672_, _13671_, _01537_);
  or (_13673_, _13672_, _13670_);
  nand (_13674_, _13475_, _01537_);
  and (_13675_, _13674_, _07368_);
  and (_13676_, _13675_, _13673_);
  and (_13677_, _07367_, _01710_);
  or (_13678_, _13677_, _07374_);
  or (_13679_, _13678_, _13676_);
  nand (_13680_, _07374_, _01613_);
  and (_13681_, _13680_, _38087_);
  and (_13682_, _13681_, _13679_);
  or (_13683_, _13682_, _13435_);
  and (_40192_, _13683_, _37580_);
  nor (_13684_, _38087_, _01613_);
  nand (_13685_, _07304_, _01710_);
  nand (_13686_, _07069_, _07321_);
  nor (_13687_, _03680_, _01613_);
  and (_13688_, _10692_, _03680_);
  nor (_13689_, _13688_, _13687_);
  nor (_13690_, _13689_, _02176_);
  or (_13691_, _06429_, _13445_);
  and (_13692_, _10816_, _03680_);
  nor (_13693_, _13692_, _13687_);
  nand (_13694_, _13693_, _02079_);
  nor (_13695_, _06472_, _02811_);
  nor (_13696_, _13695_, _13687_);
  nand (_13697_, _13696_, _05994_);
  and (_13698_, \oc8051_golden_model_1.PSW [7], _01710_);
  and (_13699_, _06518_, \oc8051_golden_model_1.ACC [0]);
  nor (_13700_, _06850_, _13699_);
  nor (_13701_, _13700_, _13698_);
  and (_13702_, _13701_, _07283_);
  nor (_13703_, _13701_, _07283_);
  or (_13704_, _13703_, _13702_);
  nand (_13705_, _13704_, _01963_);
  and (_13706_, _13705_, _06777_);
  nand (_13707_, _06614_, _02811_);
  nor (_13708_, _06838_, _06618_);
  nor (_13709_, _13461_, _02811_);
  and (_13710_, _06625_, _01613_);
  nor (_13711_, _06625_, _01613_);
  or (_13712_, _13711_, _06620_);
  or (_13713_, _13712_, _13710_);
  and (_13714_, _13713_, _13461_);
  or (_13715_, _13714_, _13709_);
  and (_13716_, _13715_, _06618_);
  or (_13717_, _13716_, _13708_);
  and (_13718_, _13717_, _10136_);
  or (_13719_, _13718_, _01883_);
  or (_13720_, _13457_, _04907_);
  and (_13721_, _13720_, _13719_);
  or (_13722_, _13721_, _02001_);
  nor (_13723_, _03680_, \oc8051_golden_model_1.ACC [1]);
  and (_13724_, _10698_, _03680_);
  nor (_13725_, _13724_, _13723_);
  or (_13726_, _13725_, _02814_);
  and (_13727_, _13726_, _13722_);
  or (_13728_, _13727_, _06636_);
  nor (_13729_, _06644_, \oc8051_golden_model_1.PSW [6]);
  nor (_13730_, _13729_, \oc8051_golden_model_1.ACC [1]);
  and (_13731_, _13729_, \oc8051_golden_model_1.ACC [1]);
  nor (_13732_, _13731_, _13730_);
  nand (_13733_, _13732_, _06636_);
  and (_13734_, _13733_, _02008_);
  and (_13735_, _13734_, _13728_);
  nor (_13736_, _04326_, _01613_);
  and (_13737_, _10710_, _04326_);
  nor (_13738_, _13737_, _13736_);
  nor (_13739_, _13738_, _02024_);
  nor (_13740_, _13696_, _02840_);
  or (_13741_, _13740_, _06614_);
  or (_13742_, _13741_, _13739_);
  or (_13743_, _13742_, _13735_);
  and (_13744_, _13743_, _13707_);
  or (_13745_, _13744_, _02850_);
  or (_13746_, _04907_, _06675_);
  and (_13747_, _13746_, _02021_);
  and (_13748_, _13747_, _13745_);
  nor (_13749_, _06838_, _02021_);
  or (_13750_, _13749_, _06679_);
  or (_13751_, _13750_, _13748_);
  nand (_13752_, _06679_, _06079_);
  and (_13753_, _13752_, _13751_);
  or (_13754_, _13753_, _01997_);
  and (_13755_, _10696_, _04326_);
  nor (_13756_, _13755_, _13736_);
  nand (_13757_, _13756_, _01997_);
  and (_13758_, _13757_, _02861_);
  and (_13759_, _13758_, _13754_);
  and (_13760_, _13737_, _10725_);
  nor (_13761_, _13760_, _13736_);
  nor (_13762_, _13761_, _02861_);
  or (_13763_, _13762_, _05279_);
  or (_13764_, _13763_, _13759_);
  and (_13765_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [0]);
  nor (_13766_, _13765_, _06315_);
  nor (_13767_, _13766_, _05902_);
  or (_13768_, _13767_, _05285_);
  and (_13769_, _13768_, _13764_);
  or (_13770_, _13769_, _06699_);
  not (_13771_, _13699_);
  and (_13772_, _13771_, _03028_);
  nor (_13773_, _13772_, _13698_);
  and (_13774_, _13773_, _06432_);
  nor (_13775_, _13773_, _06432_);
  or (_13776_, _13775_, _13774_);
  or (_13777_, _13776_, _06700_);
  and (_13778_, _13777_, _08245_);
  and (_13779_, _13778_, _13770_);
  and (_13780_, _13771_, _04952_);
  nor (_13781_, _13780_, _13698_);
  and (_13782_, _13781_, _07233_);
  nor (_13783_, _13781_, _07233_);
  or (_13784_, _13783_, _13782_);
  and (_13785_, _06609_, _13784_);
  or (_13786_, _13785_, _01963_);
  or (_13787_, _13786_, _13779_);
  and (_13788_, _13787_, _13706_);
  nor (_13789_, _13699_, _02441_);
  nor (_13790_, _13789_, _13698_);
  and (_13791_, _13790_, _07322_);
  nor (_13792_, _13790_, _07322_);
  nor (_13793_, _13792_, _13791_);
  nor (_13794_, _13793_, _06777_);
  or (_13795_, _13794_, _01549_);
  or (_13796_, _13795_, _13788_);
  nand (_13797_, _01822_, _01549_);
  and (_13798_, _13797_, _02408_);
  and (_13799_, _13798_, _13796_);
  nor (_13800_, _10742_, _06958_);
  nor (_13801_, _13800_, _13736_);
  nor (_13802_, _13801_, _02408_);
  or (_13803_, _13802_, _05994_);
  or (_13804_, _13803_, _13799_);
  and (_13805_, _13804_, _13697_);
  or (_13806_, _13805_, _02528_);
  and (_13807_, _04907_, _03680_);
  nor (_13808_, _13807_, _13687_);
  nand (_13809_, _13808_, _02528_);
  and (_13810_, _13809_, _02043_);
  and (_13811_, _13810_, _13806_);
  nor (_13812_, _10802_, _06472_);
  nor (_13813_, _13812_, _13687_);
  nor (_13814_, _13813_, _02043_);
  or (_13815_, _13814_, _06008_);
  or (_13816_, _13815_, _13811_);
  nand (_13817_, _06263_, _06008_);
  and (_13818_, _13817_, _13816_);
  and (_13819_, _13818_, _01609_);
  nor (_13820_, _01822_, _01609_);
  or (_13821_, _13820_, _01869_);
  or (_13822_, _13821_, _13819_);
  and (_13823_, _03680_, _02687_);
  nor (_13824_, _13823_, _13723_);
  or (_13825_, _13824_, _01870_);
  and (_13826_, _13825_, _06985_);
  and (_13827_, _13826_, _13822_);
  not (_13828_, _10326_);
  nor (_13829_, _06985_, _01822_);
  or (_13830_, _13829_, _13828_);
  or (_13831_, _13830_, _13827_);
  nor (_13832_, _10326_, _06432_);
  nor (_13833_, _13832_, _02579_);
  and (_13834_, _13833_, _13831_);
  and (_13835_, _07233_, _02579_);
  or (_13836_, _13835_, _02168_);
  or (_13837_, _13836_, _13834_);
  or (_13838_, _10822_, _07014_);
  and (_13839_, _13838_, _07013_);
  and (_13840_, _13839_, _13837_);
  and (_13841_, _07012_, _07322_);
  or (_13842_, _13841_, _02079_);
  or (_13843_, _13842_, _13840_);
  and (_13844_, _13843_, _13694_);
  or (_13845_, _13844_, _02167_);
  and (_13846_, _13448_, _02344_);
  or (_13847_, _13687_, _02912_);
  and (_13848_, _13847_, _13846_);
  and (_13849_, _13848_, _13845_);
  or (_13850_, _06429_, _13444_);
  and (_13851_, _13850_, _07026_);
  or (_13852_, _13851_, _13849_);
  and (_13853_, _13852_, _13691_);
  or (_13854_, _13853_, _07031_);
  or (_13855_, _07036_, _07231_);
  and (_13856_, _13855_, _07035_);
  and (_13857_, _13856_, _13854_);
  or (_13858_, _10820_, _07040_);
  and (_13859_, _13858_, _07042_);
  or (_13860_, _13859_, _13857_);
  or (_13861_, _07046_, _07320_);
  and (_13862_, _13861_, _02176_);
  and (_13863_, _13862_, _13860_);
  or (_13864_, _13863_, _13690_);
  and (_13865_, _13864_, _09859_);
  nor (_13866_, _03122_, _02595_);
  nor (_13867_, _09859_, _06430_);
  or (_13868_, _13867_, _13866_);
  or (_13869_, _13868_, _13865_);
  nand (_13870_, _13866_, _06430_);
  and (_13871_, _13870_, _07060_);
  and (_13872_, _13871_, _13869_);
  nor (_13873_, _06430_, _07060_);
  or (_13874_, _13873_, _06462_);
  or (_13875_, _13874_, _13872_);
  nand (_13876_, _07232_, _06462_);
  and (_13877_, _13876_, _02172_);
  and (_13878_, _13877_, _13875_);
  nand (_13879_, _10821_, _07070_);
  and (_13880_, _13879_, _09854_);
  or (_13881_, _13880_, _13878_);
  and (_13882_, _13881_, _13686_);
  or (_13883_, _13882_, _02071_);
  nor (_13884_, _10815_, _06472_);
  or (_13885_, _13884_, _13687_);
  or (_13886_, _13885_, _04788_);
  and (_13887_, _13886_, _07084_);
  and (_13888_, _13887_, _13883_);
  and (_13889_, _07096_, _07094_);
  nor (_13890_, _13889_, _07097_);
  or (_13891_, _13890_, _07114_);
  and (_13892_, _13891_, _10385_);
  or (_13893_, _13892_, _13888_);
  and (_13894_, _07125_, _07123_);
  nor (_13895_, _13894_, _07126_);
  or (_13896_, _13895_, _07116_);
  and (_13897_, _13896_, _13893_);
  or (_13898_, _13897_, _02164_);
  and (_13899_, _07155_, _07153_);
  nor (_13900_, _13899_, _07156_);
  or (_13901_, _13900_, _02165_);
  and (_13902_, _13901_, _07177_);
  and (_13903_, _13902_, _13898_);
  and (_13904_, _07187_, _07185_);
  nor (_13905_, _13904_, _07188_);
  and (_13906_, _13905_, _07144_);
  or (_13907_, _13906_, _07175_);
  or (_13908_, _13907_, _13903_);
  nand (_13909_, _07175_, _01710_);
  and (_13910_, _13909_, _06458_);
  and (_13911_, _13910_, _13908_);
  or (_13912_, _06433_, _06432_);
  nor (_13913_, _06458_, _06434_);
  and (_13914_, _13913_, _13912_);
  or (_13915_, _13914_, _13911_);
  and (_13916_, _13915_, _07212_);
  or (_13917_, _07234_, _07233_);
  nor (_13918_, _07235_, _07212_);
  and (_13919_, _13918_, _13917_);
  or (_13920_, _13919_, _01890_);
  or (_13921_, _13920_, _13916_);
  and (_13922_, _07285_, _07283_);
  nor (_13923_, _13922_, _07286_);
  or (_13924_, _13923_, _01891_);
  and (_13925_, _13924_, _07256_);
  and (_13926_, _13925_, _13921_);
  nor (_13927_, _07323_, _07322_);
  nor (_13928_, _13927_, _07324_);
  and (_13929_, _13928_, _07253_);
  or (_13930_, _13929_, _07304_);
  or (_13931_, _13930_, _13926_);
  and (_13932_, _13931_, _13685_);
  or (_13933_, _13932_, _02201_);
  or (_13934_, _13725_, _02303_);
  and (_13935_, _13934_, _07346_);
  and (_13936_, _13935_, _13933_);
  nor (_13937_, _07375_, _07351_);
  and (_13938_, _13937_, _08922_);
  nor (_13939_, _13938_, _10442_);
  or (_13940_, _13939_, _13936_);
  nand (_13941_, _07350_, _06184_);
  and (_13942_, _13941_, _01887_);
  and (_13943_, _13942_, _13940_);
  nor (_13944_, _13756_, _01887_);
  or (_13945_, _13944_, _01537_);
  or (_13946_, _13945_, _13943_);
  nor (_13947_, _13724_, _13687_);
  nand (_13948_, _13947_, _01537_);
  and (_13949_, _13948_, _07368_);
  and (_13950_, _13949_, _13946_);
  and (_13951_, _13937_, _07367_);
  or (_13952_, _13951_, _07374_);
  or (_13953_, _13952_, _13950_);
  nand (_13954_, _07374_, _06184_);
  and (_13955_, _13954_, _38087_);
  and (_13956_, _13955_, _13953_);
  or (_13957_, _13956_, _13684_);
  and (_40193_, _13957_, _37580_);
  nor (_13958_, _38087_, _06184_);
  nand (_13959_, _07304_, _01613_);
  and (_13960_, _07127_, _06583_);
  nor (_13961_, _13960_, _07128_);
  or (_13962_, _13961_, _07116_);
  nand (_13963_, _07069_, _07317_);
  not (_13964_, _09856_);
  nand (_13965_, _13964_, _06426_);
  nor (_13966_, _03680_, _06184_);
  and (_13967_, _11014_, _03680_);
  nor (_13968_, _13967_, _13966_);
  nand (_13969_, _13968_, _02079_);
  nor (_13970_, _06472_, _03455_);
  nor (_13971_, _13970_, _13966_);
  nand (_13972_, _13971_, _05994_);
  nor (_13973_, _04907_, _01613_);
  and (_13974_, _04952_, _01710_);
  nor (_13975_, _13974_, _07233_);
  nor (_13976_, _13975_, _13973_);
  nor (_13977_, _07229_, _13976_);
  and (_13978_, _07229_, _13976_);
  nor (_13979_, _13978_, _13977_);
  nor (_13980_, _13573_, _07233_);
  not (_13981_, _13980_);
  or (_13982_, _13981_, _13979_);
  and (_13983_, _13982_, \oc8051_golden_model_1.PSW [7]);
  nor (_13984_, _13979_, \oc8051_golden_model_1.PSW [7]);
  or (_13985_, _13984_, _13983_);
  nand (_13986_, _13981_, _13979_);
  and (_13987_, _13986_, _13985_);
  nand (_13988_, _13987_, _06609_);
  nand (_13989_, _06614_, _03455_);
  nor (_13990_, _06816_, _06618_);
  nor (_13991_, _13461_, _03455_);
  and (_13992_, _06625_, _06184_);
  nor (_13993_, _06625_, _06184_);
  or (_13994_, _13993_, _06620_);
  or (_13995_, _13994_, _13992_);
  and (_13996_, _13995_, _13461_);
  or (_13997_, _13996_, _13991_);
  and (_13998_, _13997_, _06618_);
  or (_13999_, _13998_, _13990_);
  and (_14000_, _13999_, _10136_);
  or (_14001_, _14000_, _01883_);
  or (_14002_, _13457_, _05043_);
  and (_14003_, _14002_, _14001_);
  or (_14004_, _14003_, _02001_);
  nor (_14005_, _10905_, _06472_);
  nor (_14006_, _14005_, _13966_);
  nand (_14007_, _14006_, _02001_);
  and (_14008_, _14007_, _14004_);
  or (_14009_, _14008_, _06636_);
  nand (_14010_, _13729_, \oc8051_golden_model_1.ACC [2]);
  and (_14011_, \oc8051_golden_model_1.ACC [2], \oc8051_golden_model_1.ACC [1]);
  nor (_14012_, _14011_, _06643_);
  or (_14013_, _14012_, _13729_);
  and (_14014_, _14013_, _14010_);
  nand (_14015_, _14014_, _06636_);
  and (_14016_, _14015_, _02008_);
  and (_14017_, _14016_, _14009_);
  nor (_14018_, _04326_, _06184_);
  and (_14019_, _10909_, _04326_);
  nor (_14020_, _14019_, _14018_);
  nor (_14021_, _14020_, _02024_);
  nor (_14022_, _13971_, _02840_);
  or (_14023_, _14022_, _06614_);
  or (_14024_, _14023_, _14021_);
  or (_14025_, _14024_, _14017_);
  and (_14026_, _14025_, _13989_);
  or (_14027_, _14026_, _02850_);
  or (_14028_, _05043_, _06675_);
  and (_14029_, _14028_, _02021_);
  and (_14030_, _14029_, _14027_);
  nor (_14031_, _06816_, _02021_);
  or (_14032_, _14031_, _06679_);
  or (_14033_, _14032_, _14030_);
  nand (_14034_, _06679_, _06026_);
  and (_14035_, _14034_, _14033_);
  or (_14036_, _14035_, _01997_);
  and (_14037_, _10894_, _04326_);
  nor (_14038_, _14037_, _14018_);
  nand (_14039_, _14038_, _01997_);
  and (_14040_, _14039_, _02861_);
  and (_14041_, _14040_, _14036_);
  and (_14042_, _14019_, _10924_);
  nor (_14043_, _14042_, _14018_);
  nor (_14044_, _14043_, _02861_);
  or (_14045_, _14044_, _05279_);
  or (_14046_, _14045_, _14041_);
  nor (_14047_, _05906_, _05902_);
  nor (_14048_, _14047_, _05908_);
  or (_14049_, _14048_, _05285_);
  and (_14050_, _14049_, _06700_);
  and (_14051_, _14050_, _14046_);
  and (_14052_, _02811_, \oc8051_golden_model_1.ACC [1]);
  and (_14053_, _03028_, _01710_);
  nor (_14054_, _14053_, _06432_);
  nor (_14055_, _14054_, _14052_);
  nor (_14056_, _14055_, _06427_);
  and (_14057_, _14055_, _06427_);
  nor (_14058_, _14057_, _14056_);
  nor (_14059_, _13561_, _06432_);
  not (_14060_, _14059_);
  or (_14061_, _14060_, _14058_);
  and (_14062_, _14061_, \oc8051_golden_model_1.PSW [7]);
  nor (_14063_, _14058_, \oc8051_golden_model_1.PSW [7]);
  or (_14064_, _14063_, _14062_);
  nand (_14065_, _14060_, _14058_);
  and (_14066_, _14065_, _14064_);
  nor (_14067_, _14066_, _06700_);
  or (_14068_, _14067_, _06609_);
  or (_14069_, _14068_, _14051_);
  and (_14070_, _14069_, _13988_);
  or (_14071_, _14070_, _01963_);
  nor (_14072_, _08621_, _07281_);
  or (_14073_, _14072_, _07282_);
  and (_14074_, _07279_, _14073_);
  nor (_14075_, _07279_, _14073_);
  nor (_14076_, _14075_, _14074_);
  and (_14077_, _08623_, \oc8051_golden_model_1.PSW [7]);
  not (_14078_, _14077_);
  nor (_14079_, _14078_, _14076_);
  and (_14080_, _14078_, _14076_);
  nor (_14081_, _14080_, _14079_);
  nand (_14082_, _14081_, _01963_);
  and (_14083_, _14082_, _06777_);
  and (_14084_, _14083_, _14071_);
  nor (_14085_, _02441_, \oc8051_golden_model_1.ACC [0]);
  nor (_14086_, _14085_, _07322_);
  nor (_14087_, _14086_, _08632_);
  nor (_14088_, _07318_, _14087_);
  and (_14089_, _07318_, _14087_);
  nor (_14090_, _14089_, _14088_);
  not (_14091_, _08662_);
  or (_14092_, _14091_, _14090_);
  and (_14093_, _14092_, \oc8051_golden_model_1.PSW [7]);
  nor (_14094_, _14090_, \oc8051_golden_model_1.PSW [7]);
  or (_14095_, _14094_, _14093_);
  nand (_14096_, _14091_, _14090_);
  and (_14097_, _14096_, _14095_);
  nor (_14098_, _14097_, _06777_);
  or (_14099_, _14098_, _01549_);
  or (_14100_, _14099_, _14084_);
  nand (_14101_, _02294_, _01549_);
  and (_14102_, _14101_, _02408_);
  and (_14103_, _14102_, _14100_);
  nor (_14104_, _10942_, _06958_);
  nor (_14105_, _14104_, _14018_);
  nor (_14106_, _14105_, _02408_);
  or (_14107_, _14106_, _05994_);
  or (_14108_, _14107_, _14103_);
  and (_14109_, _14108_, _13972_);
  or (_14110_, _14109_, _02528_);
  and (_14111_, _05043_, _03680_);
  nor (_14112_, _14111_, _13966_);
  nand (_14113_, _14112_, _02528_);
  and (_14114_, _14113_, _02043_);
  and (_14115_, _14114_, _14110_);
  nor (_14116_, _11000_, _06472_);
  nor (_14117_, _14116_, _13966_);
  nor (_14118_, _14117_, _02043_);
  or (_14119_, _14118_, _06008_);
  or (_14120_, _14119_, _14115_);
  or (_14121_, _06198_, _06355_);
  and (_14122_, _14121_, _14120_);
  and (_14123_, _14122_, _01609_);
  nor (_14124_, _02294_, _01609_);
  or (_14125_, _14124_, _01869_);
  or (_14126_, _14125_, _14123_);
  and (_14127_, _03680_, _04724_);
  nor (_14128_, _14127_, _13966_);
  nand (_14129_, _14128_, _01869_);
  and (_14130_, _14129_, _06985_);
  and (_14131_, _14130_, _14126_);
  nor (_14132_, _06985_, _02294_);
  or (_14133_, _14132_, _06990_);
  or (_14134_, _14133_, _14131_);
  nand (_14135_, _06994_, _06427_);
  nand (_14136_, _14135_, _06996_);
  and (_14137_, _14136_, _14134_);
  or (_14138_, _06999_, _06427_);
  and (_14139_, _14138_, _07002_);
  or (_14140_, _14139_, _14137_);
  and (_14141_, _02047_, _01644_);
  not (_14142_, _14141_);
  nand (_14143_, _06999_, _06428_);
  and (_14144_, _14143_, _14142_);
  and (_14145_, _14144_, _14140_);
  or (_14146_, _07229_, _01434_);
  and (_14147_, _14146_, _02579_);
  or (_14148_, _14147_, _14145_);
  and (_14149_, _02053_, _01644_);
  not (_14150_, _14149_);
  or (_14151_, _07229_, _14150_);
  and (_14152_, _14151_, _14148_);
  or (_14153_, _14152_, _02168_);
  or (_14154_, _11020_, _07014_);
  and (_14155_, _14154_, _07013_);
  and (_14156_, _14155_, _14153_);
  and (_14157_, _07012_, _07318_);
  or (_14158_, _14157_, _02079_);
  or (_14159_, _14158_, _14156_);
  and (_14160_, _14159_, _13969_);
  or (_14161_, _14160_, _02167_);
  or (_14162_, _13966_, _02912_);
  and (_14163_, _14162_, _09864_);
  and (_14164_, _14163_, _14161_);
  and (_14165_, _07031_, _07227_);
  and (_14166_, _06425_, _07026_);
  or (_14167_, _14166_, _02178_);
  or (_14168_, _14167_, _14165_);
  or (_14169_, _14168_, _14164_);
  or (_14170_, _11018_, _07035_);
  and (_14171_, _14170_, _14169_);
  or (_14172_, _14171_, _07040_);
  or (_14173_, _07046_, _07316_);
  and (_14174_, _14173_, _02176_);
  and (_14175_, _14174_, _14172_);
  or (_14176_, _14128_, _11019_);
  nor (_14177_, _14176_, _02176_);
  or (_14178_, _14177_, _09858_);
  or (_14179_, _14178_, _14175_);
  not (_14180_, _06426_);
  and (_14181_, _14180_, _02730_);
  or (_14182_, _14181_, _09860_);
  and (_14183_, _14182_, _14179_);
  and (_14184_, _01971_, _01647_);
  nand (_14185_, _09856_, _06426_);
  and (_14186_, _14185_, _14184_);
  or (_14187_, _14186_, _14183_);
  and (_14188_, _14187_, _13965_);
  or (_14189_, _14188_, _06462_);
  nand (_14190_, _07228_, _06462_);
  and (_14191_, _14190_, _02172_);
  and (_14192_, _14191_, _14189_);
  nand (_14193_, _11019_, _07070_);
  and (_14194_, _14193_, _09854_);
  or (_14195_, _14194_, _14192_);
  and (_14196_, _14195_, _13963_);
  or (_14197_, _14196_, _02071_);
  nor (_14198_, _11013_, _06472_);
  nor (_14199_, _14198_, _13966_);
  nand (_14200_, _14199_, _02071_);
  and (_14201_, _14200_, _07084_);
  and (_14202_, _14201_, _14197_);
  and (_14203_, _07098_, _06744_);
  nor (_14204_, _14203_, _07099_);
  and (_14205_, _14204_, _07085_);
  or (_14206_, _14205_, _07114_);
  or (_14207_, _14206_, _14202_);
  and (_14208_, _14207_, _13962_);
  or (_14209_, _14208_, _02164_);
  and (_14210_, _07157_, _06924_);
  nor (_14211_, _14210_, _07158_);
  or (_14212_, _14211_, _02165_);
  and (_14213_, _14212_, _07177_);
  and (_14214_, _14213_, _14209_);
  and (_14215_, _07189_, _06516_);
  nor (_14216_, _14215_, _07190_);
  and (_14217_, _14216_, _07144_);
  or (_14218_, _14217_, _07175_);
  or (_14219_, _14218_, _14214_);
  nand (_14220_, _07175_, _01613_);
  and (_14221_, _14220_, _06458_);
  and (_14222_, _14221_, _14219_);
  and (_14223_, _06435_, _06428_);
  nor (_14224_, _14223_, _06436_);
  and (_14225_, _14224_, _06459_);
  or (_14226_, _14225_, _14222_);
  and (_14227_, _14226_, _07212_);
  and (_14228_, _07236_, _07230_);
  nor (_14229_, _14228_, _07237_);
  and (_14230_, _14229_, _07210_);
  or (_14231_, _14230_, _01890_);
  or (_14232_, _14231_, _14227_);
  and (_14233_, _07287_, _07279_);
  nor (_14234_, _14233_, _07288_);
  or (_14235_, _14234_, _01891_);
  and (_14236_, _14235_, _07256_);
  and (_14237_, _14236_, _14232_);
  and (_14238_, _07325_, _07319_);
  nor (_14239_, _14238_, _07326_);
  and (_14240_, _14239_, _07253_);
  or (_14241_, _14240_, _07304_);
  or (_14242_, _14241_, _14237_);
  and (_14243_, _14242_, _13959_);
  or (_14244_, _14243_, _02201_);
  nand (_14245_, _14006_, _02201_);
  and (_14246_, _14245_, _07346_);
  and (_14247_, _14246_, _14244_);
  and (_14248_, _06643_, _01710_);
  nor (_14249_, _07351_, _06184_);
  or (_14250_, _14249_, _14248_);
  nor (_14251_, _14250_, _07350_);
  nor (_14252_, _14251_, _10442_);
  or (_14253_, _14252_, _14247_);
  nand (_14254_, _07350_, _01689_);
  and (_14255_, _14254_, _01887_);
  and (_14256_, _14255_, _14253_);
  nor (_14257_, _14038_, _01887_);
  or (_14258_, _14257_, _01537_);
  or (_14259_, _14258_, _14256_);
  and (_14260_, _11072_, _03680_);
  nor (_14261_, _14260_, _13966_);
  nand (_14262_, _14261_, _01537_);
  and (_14263_, _14262_, _07368_);
  and (_14264_, _14263_, _14259_);
  and (_14265_, _07375_, \oc8051_golden_model_1.ACC [2]);
  nor (_14266_, _07375_, \oc8051_golden_model_1.ACC [2]);
  nor (_14267_, _14266_, _14265_);
  nor (_14268_, _14267_, _07374_);
  nor (_14269_, _14268_, _10465_);
  or (_14270_, _14269_, _14264_);
  nand (_14271_, _07374_, _01689_);
  and (_14272_, _14271_, _38087_);
  and (_14273_, _14272_, _14270_);
  or (_14274_, _14273_, _13958_);
  and (_40194_, _14274_, _37580_);
  nor (_14275_, _38087_, _01689_);
  nor (_14276_, _06421_, _06423_);
  nor (_14277_, _14276_, _06437_);
  and (_14278_, _14276_, _06437_);
  nor (_14279_, _14278_, _14277_);
  nand (_14280_, _14279_, _06459_);
  nor (_14281_, _03680_, _01689_);
  nor (_14282_, _11220_, _06472_);
  nor (_14283_, _14282_, _14281_);
  nor (_14284_, _14283_, _04788_);
  and (_14285_, _11222_, _03680_);
  nor (_14286_, _14285_, _14281_);
  nand (_14287_, _14286_, _02079_);
  nor (_14288_, _07225_, _07223_);
  or (_14289_, _14288_, _07006_);
  nor (_14290_, _06472_, _03268_);
  nor (_14291_, _14290_, _14281_);
  nand (_14292_, _14291_, _05994_);
  nor (_14293_, _05043_, _06184_);
  nor (_14294_, _13977_, _14293_);
  and (_14295_, _14288_, _14294_);
  nor (_14296_, _14288_, _14294_);
  or (_14297_, _14296_, _14295_);
  nor (_14298_, _14297_, _06518_);
  and (_14299_, _14297_, _06518_);
  nor (_14300_, _14299_, _14298_);
  and (_14301_, _14300_, _13983_);
  nor (_14302_, _14300_, _13983_);
  nor (_14303_, _14302_, _14301_);
  or (_14304_, _14303_, _08245_);
  nor (_14305_, _04326_, _01689_);
  and (_14306_, _11098_, _04326_);
  and (_14307_, _14306_, _11127_);
  nor (_14308_, _14307_, _14305_);
  nor (_14309_, _14308_, _02861_);
  nand (_14310_, _06614_, _03268_);
  nor (_14311_, _11101_, _06472_);
  nor (_14312_, _14311_, _14281_);
  nor (_14313_, _14312_, _02814_);
  or (_14314_, _13457_, _04998_);
  nor (_14315_, _06804_, _06618_);
  nor (_14316_, _13461_, _03268_);
  and (_14317_, _06625_, _01689_);
  nor (_14318_, _06625_, _01689_);
  or (_14319_, _14318_, _06620_);
  or (_14320_, _14319_, _14317_);
  and (_14321_, _14320_, _13461_);
  or (_14322_, _14321_, _14316_);
  and (_14323_, _14322_, _06618_);
  or (_14324_, _14323_, _14315_);
  and (_14325_, _14324_, _10136_);
  or (_14326_, _14325_, _01883_);
  and (_14327_, _14326_, _02814_);
  and (_14328_, _14327_, _14314_);
  or (_14329_, _14328_, _14313_);
  and (_14330_, _14329_, _06642_);
  not (_14331_, \oc8051_golden_model_1.PSW [6]);
  nor (_14332_, _06643_, _14331_);
  nor (_14333_, _14332_, \oc8051_golden_model_1.ACC [3]);
  nor (_14334_, _14333_, _06644_);
  and (_14335_, _14334_, _06636_);
  or (_14336_, _14335_, _02007_);
  or (_14337_, _14336_, _14330_);
  nor (_14338_, _14306_, _14305_);
  nand (_14339_, _14338_, _02007_);
  and (_14340_, _14339_, _02840_);
  and (_14341_, _14340_, _14337_);
  nor (_14342_, _14291_, _02840_);
  or (_14343_, _14342_, _06614_);
  or (_14344_, _14343_, _14341_);
  and (_14345_, _14344_, _14310_);
  or (_14346_, _14345_, _02850_);
  or (_14347_, _04998_, _06675_);
  and (_14348_, _14347_, _02021_);
  and (_14349_, _14348_, _14346_);
  nor (_14350_, _06804_, _02021_);
  or (_14351_, _14350_, _06679_);
  or (_14352_, _14351_, _14349_);
  nand (_14353_, _06679_, _04776_);
  and (_14354_, _14353_, _14352_);
  or (_14355_, _14354_, _01997_);
  and (_14356_, _11096_, _04326_);
  nor (_14357_, _14356_, _14305_);
  nand (_14358_, _14357_, _01997_);
  and (_14359_, _14358_, _02861_);
  and (_14360_, _14359_, _14355_);
  or (_14361_, _14360_, _14309_);
  and (_14362_, _14361_, _05285_);
  nor (_14363_, _05912_, _05908_);
  nor (_14364_, _14363_, _05914_);
  nand (_14365_, _14364_, _05279_);
  nand (_14366_, _14365_, _08771_);
  or (_14367_, _14366_, _14362_);
  and (_14368_, _03455_, \oc8051_golden_model_1.ACC [2]);
  nor (_14369_, _14056_, _14368_);
  nor (_14370_, _14369_, _14276_);
  and (_14371_, _14369_, _14276_);
  nor (_14372_, _14371_, _14370_);
  and (_14373_, _14372_, \oc8051_golden_model_1.PSW [7]);
  nor (_14374_, _14372_, \oc8051_golden_model_1.PSW [7]);
  nor (_14375_, _14374_, _14373_);
  and (_14376_, _14375_, _14062_);
  nor (_14377_, _14375_, _14062_);
  or (_14378_, _14377_, _14376_);
  nand (_14379_, _14378_, _08772_);
  and (_14380_, _14379_, _08778_);
  and (_14381_, _14380_, _14367_);
  nor (_14382_, _14378_, _08778_);
  or (_14383_, _14382_, _06609_);
  or (_14384_, _14383_, _14381_);
  and (_14385_, _14384_, _14304_);
  or (_14386_, _14385_, _01963_);
  nor (_14387_, _14074_, _07277_);
  nor (_14388_, _08596_, _14387_);
  and (_14389_, _08596_, _14387_);
  or (_14390_, _14389_, _14388_);
  not (_14391_, _14079_);
  nor (_14392_, _14391_, _14390_);
  and (_14393_, _14391_, _14390_);
  nor (_14394_, _14393_, _14392_);
  nand (_14395_, _14394_, _01963_);
  and (_14396_, _14395_, _06777_);
  and (_14397_, _14396_, _14386_);
  and (_14398_, _02294_, \oc8051_golden_model_1.ACC [2]);
  nor (_14399_, _14088_, _14398_);
  nor (_14400_, _08629_, _14399_);
  and (_14401_, _08629_, _14399_);
  nor (_14402_, _14401_, _14400_);
  and (_14403_, _14402_, \oc8051_golden_model_1.PSW [7]);
  nor (_14404_, _14402_, \oc8051_golden_model_1.PSW [7]);
  nor (_14405_, _14404_, _14403_);
  and (_14406_, _14405_, _14093_);
  nor (_14407_, _14405_, _14093_);
  or (_14408_, _14407_, _14406_);
  nor (_14409_, _14408_, _06777_);
  or (_14410_, _14409_, _01549_);
  or (_14411_, _14410_, _14397_);
  nand (_14412_, _01954_, _01549_);
  and (_14413_, _14412_, _02408_);
  and (_14414_, _14413_, _14411_);
  nor (_14415_, _11145_, _06958_);
  nor (_14416_, _14415_, _14305_);
  nor (_14417_, _14416_, _02408_);
  or (_14418_, _14417_, _05994_);
  or (_14419_, _14418_, _14414_);
  and (_14420_, _14419_, _14292_);
  or (_14421_, _14420_, _02528_);
  and (_14422_, _04998_, _03680_);
  nor (_14423_, _14422_, _14281_);
  nand (_14424_, _14423_, _02528_);
  and (_14425_, _14424_, _02043_);
  and (_14426_, _14425_, _14421_);
  nor (_14427_, _11206_, _06472_);
  nor (_14428_, _14427_, _14281_);
  nor (_14429_, _14428_, _02043_);
  or (_14430_, _14429_, _06008_);
  or (_14431_, _14430_, _14426_);
  or (_14432_, _06146_, _06355_);
  and (_14433_, _14432_, _14431_);
  and (_14434_, _14433_, _01609_);
  nor (_14435_, _01954_, _01609_);
  or (_14436_, _14435_, _01869_);
  or (_14437_, _14436_, _14434_);
  and (_14438_, _03680_, _04678_);
  nor (_14439_, _14438_, _14281_);
  nand (_14440_, _14439_, _01869_);
  and (_14441_, _14440_, _06985_);
  and (_14442_, _14441_, _14437_);
  and (_14443_, _02062_, _01644_);
  nor (_14444_, _06985_, _01954_);
  or (_14445_, _14444_, _14443_);
  or (_14446_, _14445_, _14442_);
  not (_14447_, _14443_);
  or (_14448_, _14276_, _14447_);
  and (_14449_, _14448_, _14446_);
  and (_14450_, _02351_, _01434_);
  not (_14451_, _14450_);
  and (_14452_, _02074_, _01644_);
  nor (_14453_, _06999_, _14452_);
  and (_14454_, _14453_, _14451_);
  and (_14455_, _14454_, _06994_);
  and (_14456_, _14455_, _14449_);
  not (_14457_, _14455_);
  and (_14458_, _14457_, _14276_);
  or (_14459_, _14458_, _02579_);
  or (_14460_, _14459_, _14456_);
  and (_14461_, _14460_, _14289_);
  or (_14462_, _14461_, _02168_);
  or (_14463_, _11094_, _07014_);
  and (_14464_, _14463_, _07013_);
  and (_14465_, _14464_, _14462_);
  and (_14466_, _07012_, _08629_);
  or (_14467_, _14466_, _02079_);
  or (_14468_, _14467_, _14465_);
  and (_14469_, _14468_, _14287_);
  or (_14470_, _14469_, _02167_);
  or (_14471_, _14281_, _02912_);
  and (_14472_, _14471_, _13846_);
  and (_14473_, _14472_, _14470_);
  or (_14474_, _06423_, _13444_);
  and (_14475_, _14474_, _07026_);
  or (_14476_, _14475_, _14473_);
  or (_14477_, _06423_, _13445_);
  and (_14478_, _14477_, _07036_);
  and (_14479_, _14478_, _14476_);
  and (_14480_, _07031_, _07225_);
  or (_14481_, _14480_, _02178_);
  or (_14482_, _14481_, _14479_);
  or (_14483_, _11092_, _07035_);
  and (_14484_, _14483_, _07046_);
  and (_14485_, _14484_, _14482_);
  and (_14486_, _07040_, _07314_);
  or (_14487_, _14486_, _14485_);
  and (_14488_, _14487_, _02176_);
  or (_14489_, _14439_, _11093_);
  nor (_14490_, _14489_, _02176_);
  or (_14491_, _14490_, _07051_);
  or (_14492_, _14491_, _14488_);
  nand (_14493_, _07051_, _06421_);
  nor (_14494_, _13964_, _02594_);
  and (_14495_, _14494_, _14493_);
  and (_14496_, _14495_, _14492_);
  nor (_14497_, _14494_, _06421_);
  or (_14498_, _14497_, _06462_);
  or (_14499_, _14498_, _14496_);
  nand (_14500_, _07223_, _06462_);
  and (_14501_, _14500_, _02172_);
  and (_14502_, _14501_, _14499_);
  nand (_14503_, _11093_, _07070_);
  and (_14504_, _14503_, _09854_);
  or (_14505_, _14504_, _14502_);
  nand (_14506_, _07069_, _07315_);
  and (_14507_, _14506_, _04788_);
  and (_14508_, _14507_, _14505_);
  or (_14509_, _14508_, _14284_);
  and (_14510_, _14509_, _07084_);
  and (_14511_, _07100_, _06739_);
  nor (_14512_, _14511_, _07101_);
  and (_14513_, _14512_, _07085_);
  or (_14514_, _14513_, _07114_);
  or (_14515_, _14514_, _14510_);
  and (_14516_, _07129_, _06578_);
  nor (_14517_, _14516_, _07130_);
  or (_14518_, _14517_, _07116_);
  and (_14519_, _14518_, _02165_);
  and (_14520_, _14519_, _14515_);
  and (_14521_, _07159_, _06922_);
  nor (_14522_, _14521_, _07160_);
  or (_14523_, _14522_, _07144_);
  and (_14524_, _14523_, _07146_);
  or (_14525_, _14524_, _14520_);
  and (_14526_, _07191_, _06511_);
  nor (_14527_, _14526_, _07192_);
  or (_14528_, _14527_, _07177_);
  and (_14529_, _14528_, _07176_);
  and (_14530_, _14529_, _14525_);
  nand (_14531_, _07175_, \oc8051_golden_model_1.ACC [2]);
  nand (_14532_, _14531_, _06458_);
  or (_14533_, _14532_, _14530_);
  and (_14534_, _14533_, _14280_);
  or (_14535_, _14534_, _07210_);
  nor (_14536_, _07238_, _14288_);
  and (_14537_, _07238_, _14288_);
  nor (_14538_, _14537_, _14536_);
  nand (_14539_, _14538_, _07210_);
  and (_14540_, _14539_, _01891_);
  and (_14541_, _14540_, _14535_);
  nor (_14542_, _07289_, _08596_);
  and (_14543_, _07289_, _08596_);
  nor (_14544_, _14543_, _14542_);
  or (_14545_, _14544_, _07253_);
  and (_14546_, _14545_, _07255_);
  or (_14547_, _14546_, _14541_);
  nor (_14548_, _07327_, _08629_);
  and (_14549_, _07327_, _08629_);
  nor (_14550_, _14549_, _14548_);
  nand (_14551_, _14550_, _07253_);
  and (_14552_, _14551_, _07305_);
  and (_14553_, _14552_, _14547_);
  and (_14554_, _07304_, \oc8051_golden_model_1.ACC [2]);
  or (_14555_, _14554_, _02201_);
  or (_14556_, _14555_, _14553_);
  nand (_14557_, _14312_, _02201_);
  and (_14558_, _14557_, _07346_);
  and (_14559_, _14558_, _14556_);
  nor (_14560_, _14248_, _01689_);
  or (_14561_, _14560_, _07352_);
  and (_14562_, _14561_, _07345_);
  or (_14563_, _14562_, _07350_);
  or (_14564_, _14563_, _14559_);
  nand (_14565_, _07350_, _06085_);
  and (_14566_, _14565_, _01887_);
  and (_14567_, _14566_, _14564_);
  nor (_14568_, _14357_, _01887_);
  or (_14569_, _14568_, _01537_);
  or (_14570_, _14569_, _14567_);
  and (_14571_, _11273_, _03680_);
  nor (_14572_, _14571_, _14281_);
  nand (_14573_, _14572_, _01537_);
  and (_14574_, _14573_, _07368_);
  and (_14575_, _14574_, _14570_);
  or (_14576_, _14265_, \oc8051_golden_model_1.ACC [3]);
  and (_14577_, _14576_, _07376_);
  and (_14578_, _14577_, _07367_);
  or (_14579_, _14578_, _07374_);
  or (_14580_, _14579_, _14575_);
  nand (_14581_, _07374_, _06085_);
  and (_14582_, _14581_, _38087_);
  and (_14583_, _14582_, _14580_);
  or (_14584_, _14583_, _14275_);
  and (_40195_, _14584_, _37580_);
  nor (_14585_, _38087_, _06085_);
  nand (_14586_, _07304_, _01689_);
  nor (_14587_, _07193_, _06505_);
  nor (_14588_, _14587_, _07194_);
  or (_14589_, _14588_, _07177_);
  nand (_14590_, _07069_, _07312_);
  and (_14591_, _01647_, _01533_);
  nand (_14592_, _14591_, _06418_);
  or (_14593_, _07036_, _07220_);
  nor (_14594_, _03680_, _06085_);
  and (_14595_, _11425_, _03680_);
  nor (_14596_, _14595_, _14594_);
  nand (_14597_, _14596_, _02079_);
  nor (_14598_, _04211_, _06472_);
  nor (_14599_, _14598_, _14594_);
  nand (_14600_, _14599_, _05994_);
  or (_14601_, _14406_, _14403_);
  or (_14602_, _14399_, _08638_);
  and (_14603_, _14602_, _08637_);
  nor (_14604_, _07313_, _14603_);
  and (_14605_, _07313_, _14603_);
  nor (_14606_, _14605_, _14604_);
  and (_14607_, _14606_, \oc8051_golden_model_1.PSW [7]);
  nor (_14608_, _14606_, \oc8051_golden_model_1.PSW [7]);
  nor (_14609_, _14608_, _14607_);
  and (_14610_, _14609_, _14601_);
  nor (_14611_, _14609_, _14601_);
  nor (_14612_, _14611_, _14610_);
  or (_14613_, _14612_, _06777_);
  nand (_14614_, _06614_, _04211_);
  nor (_14615_, _06884_, _06618_);
  or (_14616_, _05135_, _06621_);
  nor (_14617_, _13461_, _04211_);
  and (_14618_, _06625_, _06085_);
  nor (_14619_, _06625_, _06085_);
  or (_14620_, _14619_, _06620_);
  or (_14621_, _14620_, _14618_);
  and (_14622_, _14621_, _13461_);
  or (_14623_, _14622_, _14617_);
  and (_14624_, _14623_, _06618_);
  and (_14625_, _14624_, _14616_);
  or (_14626_, _14625_, _14615_);
  and (_14627_, _14626_, _06617_);
  nor (_14628_, _11317_, _06472_);
  nor (_14629_, _14628_, _14594_);
  nor (_14630_, _14629_, _02814_);
  or (_14631_, _14630_, _06636_);
  or (_14632_, _14631_, _14627_);
  nor (_14633_, _06644_, \oc8051_golden_model_1.ACC [4]);
  nor (_14634_, _14633_, _06650_);
  not (_14635_, _14634_);
  nand (_14636_, _14635_, _06636_);
  and (_14637_, _14636_, _02008_);
  and (_14638_, _14637_, _14632_);
  nor (_14639_, _04326_, _06085_);
  and (_14640_, _11303_, _04326_);
  nor (_14641_, _14640_, _14639_);
  nor (_14642_, _14641_, _02024_);
  nor (_14643_, _14599_, _02840_);
  or (_14644_, _14643_, _06614_);
  or (_14645_, _14644_, _14642_);
  or (_14646_, _14645_, _14638_);
  and (_14647_, _14646_, _14614_);
  or (_14648_, _14647_, _02850_);
  or (_14649_, _05135_, _06675_);
  and (_14650_, _14649_, _02021_);
  and (_14651_, _14650_, _14648_);
  nor (_14652_, _06884_, _02021_);
  or (_14653_, _14652_, _06679_);
  or (_14654_, _14653_, _14651_);
  nand (_14655_, _06679_, _01710_);
  and (_14656_, _14655_, _14654_);
  or (_14657_, _14656_, _01997_);
  and (_14658_, _11301_, _04326_);
  nor (_14659_, _14658_, _14639_);
  nand (_14660_, _14659_, _01997_);
  and (_14661_, _14660_, _02861_);
  and (_14662_, _14661_, _14657_);
  and (_14663_, _14640_, _11334_);
  nor (_14664_, _14663_, _14639_);
  nor (_14665_, _14664_, _02861_);
  or (_14666_, _14665_, _05279_);
  or (_14667_, _14666_, _14662_);
  nor (_14668_, _05918_, _05914_);
  nor (_14669_, _14668_, _05920_);
  or (_14670_, _14669_, _05285_);
  and (_14671_, _14670_, _14667_);
  or (_14672_, _14671_, _06699_);
  or (_14673_, _14376_, _14373_);
  nor (_14674_, _03268_, \oc8051_golden_model_1.ACC [3]);
  nand (_14675_, _03268_, \oc8051_golden_model_1.ACC [3]);
  and (_14676_, _14369_, _14675_);
  or (_14677_, _14676_, _14674_);
  nor (_14678_, _14677_, _06419_);
  and (_14679_, _14677_, _06419_);
  nor (_14680_, _14679_, _14678_);
  and (_14681_, _14680_, \oc8051_golden_model_1.PSW [7]);
  nor (_14682_, _14680_, \oc8051_golden_model_1.PSW [7]);
  nor (_14683_, _14682_, _14681_);
  and (_14684_, _14683_, _14673_);
  nor (_14685_, _14683_, _14673_);
  nor (_14686_, _14685_, _14684_);
  or (_14687_, _14686_, _06700_);
  and (_14688_, _14687_, _08245_);
  and (_14689_, _14688_, _14672_);
  or (_14690_, _14301_, _14298_);
  and (_14691_, _04998_, _01689_);
  or (_14692_, _04998_, _01689_);
  and (_14693_, _14692_, _14294_);
  or (_14694_, _14693_, _14691_);
  nor (_14695_, _07222_, _14694_);
  and (_14696_, _07222_, _14694_);
  nor (_14697_, _14696_, _14695_);
  and (_14698_, _14697_, \oc8051_golden_model_1.PSW [7]);
  nor (_14699_, _14697_, \oc8051_golden_model_1.PSW [7]);
  nor (_14700_, _14699_, _14698_);
  and (_14701_, _14700_, _14690_);
  nor (_14702_, _14700_, _14690_);
  nor (_14703_, _14702_, _14701_);
  and (_14704_, _14703_, _06609_);
  or (_14705_, _14704_, _01963_);
  or (_14706_, _14705_, _14689_);
  or (_14707_, _14387_, _08594_);
  and (_14708_, _14707_, _08603_);
  nor (_14709_, _07273_, _14708_);
  and (_14710_, _07273_, _14708_);
  nor (_14711_, _14710_, _14709_);
  or (_14712_, _14392_, _14711_);
  nand (_14713_, _14392_, _14711_);
  and (_14714_, _14713_, _14712_);
  or (_14715_, _14714_, _02036_);
  and (_14716_, _14715_, _14706_);
  or (_14717_, _14716_, _06476_);
  and (_14718_, _14717_, _14613_);
  or (_14719_, _14718_, _01549_);
  nand (_14720_, _01855_, _01549_);
  and (_14721_, _14720_, _02408_);
  and (_14722_, _14721_, _14719_);
  nor (_14723_, _11299_, _06958_);
  nor (_14724_, _14723_, _14639_);
  nor (_14725_, _14724_, _02408_);
  or (_14726_, _14725_, _05994_);
  or (_14727_, _14726_, _14722_);
  and (_14728_, _14727_, _14600_);
  or (_14729_, _14728_, _02528_);
  and (_14730_, _05135_, _03680_);
  nor (_14731_, _14730_, _14594_);
  nand (_14732_, _14731_, _02528_);
  and (_14733_, _14732_, _02043_);
  and (_14734_, _14733_, _14729_);
  nor (_14735_, _11411_, _06472_);
  nor (_14736_, _14735_, _14594_);
  nor (_14737_, _14736_, _02043_);
  or (_14738_, _14737_, _06008_);
  or (_14739_, _14738_, _14734_);
  or (_14740_, _06092_, _06355_);
  and (_14741_, _14740_, _14739_);
  and (_14742_, _14741_, _01609_);
  nor (_14743_, _01855_, _01609_);
  or (_14744_, _14743_, _01869_);
  or (_14745_, _14744_, _14742_);
  and (_14746_, _04694_, _03680_);
  nor (_14747_, _14746_, _14594_);
  nand (_14748_, _14747_, _01869_);
  and (_14749_, _14748_, _06985_);
  and (_14750_, _14749_, _14745_);
  nor (_14751_, _06985_, _01855_);
  or (_14752_, _14751_, _02351_);
  or (_14753_, _14752_, _14750_);
  or (_14754_, _06419_, _02352_);
  nor (_14755_, _14452_, _06993_);
  not (_14756_, _14755_);
  nor (_14757_, _03122_, _02371_);
  nor (_14758_, _14757_, _14756_);
  and (_14759_, _14758_, _14754_);
  and (_14760_, _14759_, _14753_);
  and (_14761_, _01972_, _01644_);
  not (_14762_, _14758_);
  and (_14763_, _14762_, _06419_);
  or (_14764_, _14763_, _14761_);
  or (_14765_, _14764_, _14760_);
  not (_14766_, _14761_);
  or (_14767_, _06419_, _14766_);
  and (_14768_, _14767_, _07006_);
  and (_14769_, _14768_, _14765_);
  and (_14770_, _07222_, _02579_);
  or (_14771_, _14770_, _02168_);
  or (_14772_, _14771_, _14769_);
  or (_14773_, _11431_, _07014_);
  and (_14774_, _14773_, _07013_);
  and (_14775_, _14774_, _14772_);
  and (_14776_, _07012_, _07313_);
  or (_14777_, _14776_, _02079_);
  or (_14778_, _14777_, _14775_);
  and (_14779_, _14778_, _14597_);
  or (_14780_, _14779_, _02167_);
  or (_14781_, _14594_, _02912_);
  and (_14782_, _14781_, _07027_);
  and (_14783_, _14782_, _14780_);
  and (_14784_, _06417_, _07026_);
  or (_14785_, _14784_, _07031_);
  or (_14786_, _14785_, _14783_);
  and (_14787_, _14786_, _14593_);
  or (_14788_, _14787_, _02178_);
  or (_14789_, _11429_, _07035_);
  and (_14790_, _14789_, _07046_);
  and (_14791_, _14790_, _14788_);
  and (_14792_, _07040_, _07311_);
  or (_14793_, _14792_, _14791_);
  and (_14794_, _14793_, _02176_);
  or (_14795_, _14747_, _11430_);
  nor (_14796_, _14795_, _02176_);
  or (_14797_, _14796_, _14591_);
  or (_14798_, _14797_, _14794_);
  and (_14799_, _14798_, _14592_);
  or (_14800_, _14799_, _06462_);
  nand (_14801_, _07221_, _06462_);
  and (_14802_, _14801_, _02172_);
  and (_14803_, _14802_, _14800_);
  nand (_14804_, _11430_, _07070_);
  and (_14805_, _14804_, _09854_);
  or (_14806_, _14805_, _14803_);
  and (_14807_, _14806_, _14590_);
  or (_14808_, _14807_, _02071_);
  nor (_14809_, _11424_, _06472_);
  nor (_14810_, _14809_, _14594_);
  nand (_14811_, _14810_, _02071_);
  and (_14812_, _14811_, _07084_);
  and (_14813_, _14812_, _14808_);
  nor (_14814_, _07102_, _06730_);
  nor (_14815_, _14814_, _07103_);
  or (_14816_, _14815_, _07114_);
  and (_14817_, _14816_, _10385_);
  or (_14818_, _14817_, _14813_);
  nor (_14819_, _07131_, _06570_);
  nor (_14820_, _14819_, _07132_);
  or (_14821_, _14820_, _07116_);
  and (_14822_, _14821_, _02165_);
  and (_14823_, _14822_, _14818_);
  nor (_14824_, _07161_, _06911_);
  nor (_14825_, _14824_, _07162_);
  or (_14826_, _14825_, _07144_);
  and (_14827_, _14826_, _07146_);
  or (_14828_, _14827_, _14823_);
  and (_14829_, _14828_, _14589_);
  or (_14830_, _14829_, _07175_);
  nand (_14831_, _07175_, _01689_);
  and (_14832_, _14831_, _06458_);
  and (_14833_, _14832_, _14830_);
  nor (_14834_, _06439_, _06419_);
  nor (_14835_, _14834_, _06440_);
  and (_14836_, _14835_, _06459_);
  or (_14837_, _14836_, _14833_);
  and (_14838_, _14837_, _07212_);
  nor (_14839_, _07240_, _07222_);
  nor (_14840_, _14839_, _07241_);
  and (_14841_, _14840_, _07210_);
  or (_14842_, _14841_, _01890_);
  or (_14843_, _14842_, _14838_);
  nor (_14844_, _07291_, _07273_);
  nor (_14845_, _14844_, _07292_);
  or (_14846_, _14845_, _01891_);
  and (_14847_, _14846_, _07256_);
  and (_14848_, _14847_, _14843_);
  nor (_14849_, _07329_, _07313_);
  nor (_14850_, _14849_, _07330_);
  and (_14851_, _14850_, _07253_);
  or (_14852_, _14851_, _07304_);
  or (_14853_, _14852_, _14848_);
  and (_14854_, _14853_, _14586_);
  or (_14855_, _14854_, _02201_);
  nand (_14856_, _14629_, _02201_);
  and (_14857_, _14856_, _07346_);
  and (_14858_, _14857_, _14855_);
  and (_14859_, _07352_, _06085_);
  nor (_14860_, _07352_, _06085_);
  nor (_14861_, _14860_, _14859_);
  not (_14862_, _14861_);
  and (_14863_, _14862_, _07345_);
  or (_14864_, _14863_, _07350_);
  or (_14865_, _14864_, _14858_);
  nand (_14866_, _07350_, _06079_);
  and (_14867_, _14866_, _01887_);
  and (_14868_, _14867_, _14865_);
  nor (_14869_, _14659_, _01887_);
  or (_14870_, _14869_, _01537_);
  or (_14871_, _14870_, _14868_);
  and (_14872_, _11487_, _03680_);
  nor (_14873_, _14872_, _14594_);
  nand (_14874_, _14873_, _01537_);
  and (_14875_, _14874_, _07368_);
  and (_14876_, _14875_, _14871_);
  and (_14877_, _07376_, _06085_);
  nor (_14878_, _14877_, _07377_);
  and (_14879_, _14878_, _07367_);
  or (_14880_, _14879_, _07374_);
  or (_14881_, _14880_, _14876_);
  nand (_14882_, _07374_, _06079_);
  and (_14883_, _14882_, _38087_);
  and (_14884_, _14883_, _14881_);
  or (_14885_, _14884_, _14585_);
  and (_40196_, _14885_, _37580_);
  nor (_14886_, _38087_, _06079_);
  and (_14887_, _02049_, _01652_);
  nor (_14888_, _03680_, _06079_);
  nor (_14889_, _11628_, _06472_);
  nor (_14890_, _14889_, _14888_);
  nor (_14891_, _14890_, _04788_);
  or (_14892_, _07036_, _07216_);
  and (_14893_, _11629_, _03680_);
  nor (_14894_, _14893_, _14888_);
  nand (_14895_, _14894_, _02079_);
  and (_14896_, _07218_, _14141_);
  and (_14897_, _06415_, _14761_);
  and (_14898_, _06454_, _01644_);
  and (_14899_, _01975_, _01644_);
  and (_14900_, _06415_, _02351_);
  nor (_14901_, _06985_, _02252_);
  nor (_14902_, _03916_, _06472_);
  nor (_14903_, _14902_, _14888_);
  nand (_14904_, _14903_, _05994_);
  and (_14905_, _01855_, \oc8051_golden_model_1.ACC [4]);
  nor (_14906_, _14604_, _14905_);
  nor (_14907_, _08643_, _14906_);
  and (_14908_, _08643_, _14906_);
  nor (_14909_, _14908_, _14907_);
  and (_14910_, _14909_, \oc8051_golden_model_1.PSW [7]);
  nor (_14911_, _14909_, \oc8051_golden_model_1.PSW [7]);
  nor (_14912_, _14911_, _14910_);
  nor (_14913_, _14610_, _14607_);
  not (_14914_, _14913_);
  and (_14915_, _14914_, _14912_);
  nor (_14916_, _14914_, _14912_);
  nor (_14917_, _14916_, _14915_);
  or (_14918_, _14917_, _06777_);
  nor (_14919_, _05135_, _06085_);
  nor (_14920_, _14695_, _14919_);
  nor (_14921_, _07218_, _14920_);
  and (_14922_, _07218_, _14920_);
  nor (_14923_, _14922_, _14921_);
  and (_14924_, _14923_, \oc8051_golden_model_1.PSW [7]);
  nor (_14925_, _14923_, \oc8051_golden_model_1.PSW [7]);
  nor (_14926_, _14925_, _14924_);
  nor (_14927_, _14701_, _14698_);
  not (_14928_, _14927_);
  and (_14929_, _14928_, _14926_);
  nor (_14930_, _14928_, _14926_);
  nor (_14931_, _14930_, _14929_);
  and (_14932_, _14931_, _06609_);
  nor (_14933_, _04326_, _06079_);
  and (_14934_, _11510_, _04326_);
  and (_14935_, _14934_, _11542_);
  nor (_14936_, _14935_, _14933_);
  nor (_14937_, _14936_, _02861_);
  nand (_14938_, _06614_, _03916_);
  nor (_14939_, _06867_, _06618_);
  or (_14940_, _05090_, _06621_);
  nor (_14941_, _13461_, _03916_);
  and (_14942_, _06625_, _06079_);
  nor (_14943_, _06625_, _06079_);
  or (_14944_, _14943_, _06620_);
  or (_14945_, _14944_, _14942_);
  and (_14946_, _14945_, _13461_);
  or (_14947_, _14946_, _14941_);
  and (_14948_, _14947_, _06618_);
  and (_14949_, _14948_, _14940_);
  or (_14950_, _14949_, _14939_);
  and (_14951_, _14950_, _06617_);
  nor (_14952_, _11525_, _06472_);
  nor (_14953_, _14952_, _14888_);
  nor (_14954_, _14953_, _02814_);
  or (_14955_, _14954_, _06636_);
  or (_14956_, _14955_, _14951_);
  and (_14957_, _08514_, _06652_);
  nor (_14958_, _08514_, _06652_);
  nor (_14959_, _14958_, _14957_);
  nand (_14960_, _14959_, _06636_);
  and (_14961_, _14960_, _02008_);
  and (_14962_, _14961_, _14956_);
  nor (_14963_, _14934_, _14933_);
  nor (_14964_, _14963_, _02024_);
  nor (_14965_, _14903_, _02840_);
  or (_14966_, _14965_, _06614_);
  or (_14967_, _14966_, _14964_);
  or (_14968_, _14967_, _14962_);
  and (_14969_, _14968_, _14938_);
  or (_14970_, _14969_, _02850_);
  or (_14971_, _05090_, _06675_);
  and (_14972_, _14971_, _02021_);
  and (_14973_, _14972_, _14970_);
  nor (_14974_, _06867_, _02021_);
  or (_14975_, _14974_, _06679_);
  or (_14976_, _14975_, _14973_);
  nand (_14977_, _06679_, _01613_);
  and (_14978_, _14977_, _14976_);
  or (_14979_, _14978_, _01997_);
  and (_14980_, _11508_, _04326_);
  nor (_14981_, _14980_, _14933_);
  nand (_14982_, _14981_, _01997_);
  and (_14983_, _14982_, _02861_);
  and (_14984_, _14983_, _14979_);
  or (_14985_, _14984_, _14937_);
  and (_14986_, _14985_, _05285_);
  nor (_14987_, _05924_, _05920_);
  nor (_14988_, _14987_, _05926_);
  and (_14989_, _14988_, _05279_);
  or (_14990_, _14989_, _06699_);
  or (_14991_, _14990_, _14986_);
  and (_14992_, _04211_, \oc8051_golden_model_1.ACC [4]);
  nor (_14993_, _14678_, _14992_);
  nor (_14994_, _14993_, _06415_);
  and (_14995_, _14993_, _06415_);
  nor (_14996_, _14995_, _14994_);
  and (_14997_, _14996_, \oc8051_golden_model_1.PSW [7]);
  nor (_14998_, _14996_, \oc8051_golden_model_1.PSW [7]);
  nor (_14999_, _14998_, _14997_);
  nor (_15000_, _14684_, _14681_);
  not (_15001_, _15000_);
  and (_15002_, _15001_, _14999_);
  nor (_15003_, _15001_, _14999_);
  nor (_15004_, _15003_, _15002_);
  or (_15005_, _15004_, _06700_);
  and (_15006_, _15005_, _08245_);
  and (_15007_, _15006_, _14991_);
  or (_15008_, _15007_, _14932_);
  and (_15009_, _15008_, _02036_);
  not (_15010_, _08624_);
  nor (_15011_, _15010_, _14711_);
  nor (_15012_, _15011_, _06518_);
  not (_15013_, _15012_);
  nor (_15014_, _14709_, _07270_);
  nor (_15015_, _07268_, _15014_);
  and (_15016_, _07268_, _15014_);
  or (_15017_, _15016_, _15015_);
  and (_15018_, _15017_, _06518_);
  nor (_15019_, _15017_, _06518_);
  nor (_15020_, _15019_, _15018_);
  and (_15021_, _15020_, _15013_);
  nor (_15022_, _15020_, _15013_);
  nor (_15023_, _15022_, _15021_);
  and (_15024_, _15023_, _01963_);
  or (_15025_, _15024_, _06476_);
  or (_15026_, _15025_, _15009_);
  and (_15027_, _15026_, _14918_);
  or (_15028_, _15027_, _01549_);
  nand (_15029_, _02252_, _01549_);
  and (_15030_, _15029_, _02408_);
  and (_15031_, _15030_, _15028_);
  nor (_15032_, _11506_, _06958_);
  nor (_15033_, _15032_, _14933_);
  nor (_15034_, _15033_, _02408_);
  or (_15035_, _15034_, _05994_);
  or (_15036_, _15035_, _15031_);
  and (_15037_, _15036_, _14904_);
  or (_15038_, _15037_, _02528_);
  and (_15039_, _05090_, _03680_);
  nor (_15040_, _15039_, _14888_);
  nand (_15041_, _15040_, _02528_);
  and (_15042_, _15041_, _02043_);
  and (_15043_, _15042_, _15038_);
  nor (_15044_, _11615_, _06472_);
  nor (_15045_, _15044_, _14888_);
  nor (_15046_, _15045_, _02043_);
  or (_15047_, _15046_, _06008_);
  or (_15048_, _15047_, _15043_);
  or (_15049_, _06059_, _06355_);
  and (_15050_, _15049_, _15048_);
  and (_15051_, _15050_, _01609_);
  nor (_15052_, _02252_, _01609_);
  or (_15053_, _15052_, _01869_);
  or (_15054_, _15053_, _15051_);
  and (_15055_, _04672_, _03680_);
  nor (_15056_, _15055_, _14888_);
  nand (_15057_, _15056_, _01869_);
  and (_15058_, _15057_, _06985_);
  and (_15059_, _15058_, _15054_);
  or (_15060_, _15059_, _14901_);
  and (_15061_, _15060_, _02352_);
  nor (_15062_, _15061_, _14900_);
  nor (_15063_, _15062_, _14452_);
  and (_15064_, _06415_, _14452_);
  nor (_15065_, _15064_, _15063_);
  nor (_15066_, _15065_, _10322_);
  and (_15067_, _10322_, _06415_);
  nor (_15068_, _15067_, _15066_);
  nor (_15069_, _15068_, _14899_);
  and (_15070_, _06415_, _14899_);
  or (_15071_, _15070_, _15069_);
  or (_15072_, _15071_, _14898_);
  nand (_15073_, _14898_, _06416_);
  and (_15074_, _15073_, _14766_);
  and (_15075_, _15074_, _15072_);
  or (_15076_, _15075_, _14897_);
  and (_15077_, _15076_, _14142_);
  or (_15078_, _15077_, _14896_);
  and (_15079_, _15078_, _14150_);
  and (_15080_, _07218_, _02580_);
  or (_15081_, _15080_, _02168_);
  or (_15082_, _15081_, _15079_);
  or (_15083_, _11635_, _07014_);
  and (_15084_, _15083_, _07013_);
  and (_15085_, _15084_, _15082_);
  and (_15086_, _07012_, _08643_);
  or (_15087_, _15086_, _02079_);
  or (_15088_, _15087_, _15085_);
  and (_15089_, _15088_, _14895_);
  or (_15090_, _15089_, _02167_);
  or (_15091_, _14888_, _02912_);
  and (_15092_, _15091_, _07027_);
  and (_15093_, _15092_, _15090_);
  and (_15094_, _06413_, _07026_);
  or (_15095_, _15094_, _07031_);
  or (_15096_, _15095_, _15093_);
  and (_15097_, _15096_, _14892_);
  or (_15098_, _15097_, _02178_);
  or (_15099_, _11633_, _07035_);
  and (_15100_, _15099_, _07046_);
  and (_15101_, _15100_, _15098_);
  and (_15102_, _07040_, _07309_);
  or (_15103_, _15102_, _15101_);
  and (_15104_, _15103_, _02176_);
  or (_15105_, _15056_, _11634_);
  nor (_15106_, _15105_, _02176_);
  or (_15107_, _15106_, _14591_);
  or (_15108_, _15107_, _15104_);
  nand (_15109_, _14591_, _06414_);
  and (_15110_, _15109_, _15108_);
  or (_15111_, _15110_, _06462_);
  nand (_15112_, _07217_, _06462_);
  and (_15113_, _15112_, _02172_);
  and (_15114_, _15113_, _15111_);
  nand (_15115_, _11634_, _07070_);
  and (_15116_, _15115_, _09854_);
  or (_15117_, _15116_, _15114_);
  nand (_15118_, _07069_, _07310_);
  and (_15119_, _15118_, _04788_);
  and (_15120_, _15119_, _15117_);
  or (_15121_, _15120_, _14891_);
  and (_15122_, _15121_, _07084_);
  and (_15123_, _07104_, _06727_);
  nor (_15124_, _15123_, _07105_);
  and (_15125_, _15124_, _07085_);
  or (_15126_, _15125_, _07114_);
  or (_15127_, _15126_, _15122_);
  and (_15128_, _07133_, _06567_);
  nor (_15129_, _15128_, _07134_);
  or (_15130_, _15129_, _07116_);
  and (_15131_, _15130_, _02165_);
  and (_15132_, _15131_, _15127_);
  and (_15133_, _07164_, _06905_);
  nor (_15134_, _15133_, _07165_);
  or (_15135_, _15134_, _07144_);
  and (_15136_, _15135_, _07146_);
  or (_15137_, _15136_, _15132_);
  and (_15138_, _07195_, _06502_);
  nor (_15139_, _15138_, _07196_);
  or (_15140_, _15139_, _07177_);
  and (_15141_, _15140_, _07176_);
  and (_15142_, _15141_, _15137_);
  nor (_15143_, _06453_, _02693_);
  nand (_15144_, _07175_, \oc8051_golden_model_1.ACC [4]);
  nand (_15145_, _15144_, _15143_);
  or (_15146_, _15145_, _15142_);
  and (_15147_, _06441_, _06416_);
  nor (_15148_, _15147_, _06443_);
  or (_15149_, _15148_, _15143_);
  nand (_15150_, _15149_, _15146_);
  nor (_15151_, _15150_, _14887_);
  and (_15152_, _15148_, _14887_);
  or (_15153_, _15152_, _07210_);
  or (_15154_, _15153_, _15151_);
  and (_15155_, _07242_, _07219_);
  nor (_15156_, _15155_, _07243_);
  or (_15157_, _15156_, _07212_);
  and (_15158_, _15157_, _01891_);
  and (_15159_, _15158_, _15154_);
  and (_15160_, _07293_, _07268_);
  nor (_15161_, _15160_, _07294_);
  or (_15162_, _15161_, _07253_);
  and (_15163_, _15162_, _07255_);
  or (_15164_, _15163_, _15159_);
  not (_15165_, _08643_);
  nor (_15166_, _07331_, _15165_);
  and (_15167_, _07331_, _15165_);
  nor (_15168_, _15167_, _15166_);
  or (_15169_, _15168_, _07256_);
  and (_15170_, _15169_, _07305_);
  and (_15171_, _15170_, _15164_);
  and (_15172_, _07304_, \oc8051_golden_model_1.ACC [4]);
  or (_15173_, _15172_, _02201_);
  or (_15174_, _15173_, _15171_);
  nand (_15175_, _14953_, _02201_);
  and (_15176_, _15175_, _07346_);
  and (_15177_, _15176_, _15174_);
  nor (_15178_, _14859_, _06079_);
  or (_15179_, _15178_, _07353_);
  and (_15180_, _15179_, _07345_);
  or (_15181_, _15180_, _07350_);
  or (_15182_, _15181_, _15177_);
  nand (_15183_, _07350_, _06026_);
  and (_15184_, _15183_, _01887_);
  and (_15185_, _15184_, _15182_);
  nor (_15186_, _14981_, _01887_);
  or (_15187_, _15186_, _01537_);
  or (_15188_, _15187_, _15185_);
  and (_15189_, _11685_, _03680_);
  nor (_15190_, _15189_, _14888_);
  nand (_15191_, _15190_, _01537_);
  and (_15192_, _15191_, _07368_);
  and (_15193_, _15192_, _15188_);
  nor (_15194_, _07377_, \oc8051_golden_model_1.ACC [5]);
  nor (_15195_, _15194_, _07378_);
  and (_15196_, _15195_, _07367_);
  or (_15197_, _15196_, _07374_);
  or (_15198_, _15197_, _15193_);
  nand (_15199_, _07374_, _06026_);
  and (_15200_, _15199_, _38087_);
  and (_15201_, _15200_, _15198_);
  or (_15202_, _15201_, _14886_);
  and (_40197_, _15202_, _37580_);
  nor (_15203_, _38087_, _06026_);
  nand (_15204_, _07304_, _06079_);
  nand (_15205_, _07069_, _07307_);
  nand (_15206_, _09858_, _06411_);
  nand (_15207_, _06410_, _07026_);
  nor (_15208_, _03680_, _06026_);
  and (_15209_, _11835_, _03680_);
  nor (_15210_, _15209_, _15208_);
  and (_15211_, _15210_, _02079_);
  nor (_15212_, _07215_, _07006_);
  and (_15213_, _14757_, _06412_);
  not (_15214_, _06412_);
  nand (_15215_, _06990_, _15214_);
  nor (_15216_, _03808_, _06472_);
  nor (_15217_, _15216_, _15208_);
  nand (_15218_, _15217_, _05994_);
  or (_15219_, _15014_, _07266_);
  and (_15220_, _15219_, _08612_);
  nor (_15221_, _15220_, _07264_);
  and (_15222_, _15220_, _07264_);
  nor (_15223_, _15222_, _15221_);
  nor (_15224_, _15012_, _15017_);
  nor (_15225_, _15018_, _15224_);
  nor (_15226_, _15225_, _06518_);
  nand (_15227_, _15226_, _15223_);
  or (_15228_, _15226_, _15223_);
  and (_15229_, _15228_, _15227_);
  or (_15230_, _15229_, _02036_);
  and (_15231_, _15230_, _06777_);
  or (_15232_, _05090_, _06079_);
  and (_15233_, _05090_, _06079_);
  or (_15234_, _14920_, _15233_);
  and (_15235_, _15234_, _15232_);
  nor (_15236_, _15235_, _07215_);
  and (_15237_, _15235_, _07215_);
  nor (_15238_, _15237_, _15236_);
  nor (_15239_, _14929_, _14924_);
  and (_15240_, _15239_, \oc8051_golden_model_1.PSW [7]);
  nor (_15241_, _15240_, _15238_);
  and (_15242_, _15240_, _15238_);
  nor (_15243_, _15242_, _15241_);
  and (_15244_, _15243_, _06609_);
  nand (_15245_, _03916_, \oc8051_golden_model_1.ACC [5]);
  nor (_15246_, _03916_, \oc8051_golden_model_1.ACC [5]);
  or (_15247_, _14993_, _15246_);
  and (_15248_, _15247_, _15245_);
  nor (_15249_, _15248_, _06412_);
  and (_15250_, _15248_, _06412_);
  nor (_15251_, _15250_, _15249_);
  nor (_15252_, _15002_, _14997_);
  and (_15253_, _15252_, \oc8051_golden_model_1.PSW [7]);
  nor (_15254_, _15253_, _15251_);
  and (_15255_, _15253_, _15251_);
  nor (_15256_, _15255_, _15254_);
  and (_15257_, _15256_, _06699_);
  nand (_15258_, _06614_, _03808_);
  nor (_15259_, _06791_, _06618_);
  or (_15260_, _04861_, _06621_);
  nor (_15261_, _13461_, _03808_);
  and (_15262_, _06625_, _06026_);
  nor (_15263_, _06625_, _06026_);
  or (_15264_, _15263_, _06620_);
  or (_15265_, _15264_, _15262_);
  and (_15266_, _15265_, _13461_);
  or (_15267_, _15266_, _15261_);
  and (_15268_, _15267_, _06618_);
  and (_15269_, _15268_, _15260_);
  or (_15270_, _15269_, _15259_);
  and (_15271_, _15270_, _06617_);
  nor (_15272_, _11730_, _06472_);
  nor (_15273_, _15272_, _15208_);
  nor (_15274_, _15273_, _02814_);
  or (_15275_, _15274_, _06636_);
  or (_15276_, _15275_, _15271_);
  not (_15277_, _06654_);
  nor (_15278_, _14958_, _15277_);
  and (_15279_, _08513_, _06655_);
  nor (_15280_, _15279_, _15278_);
  nand (_15281_, _15280_, _06636_);
  and (_15282_, _15281_, _02008_);
  and (_15283_, _15282_, _15276_);
  nor (_15284_, _04326_, _06026_);
  and (_15285_, _11717_, _04326_);
  nor (_15286_, _15285_, _15284_);
  nor (_15287_, _15286_, _02024_);
  nor (_15288_, _15217_, _02840_);
  or (_15289_, _15288_, _06614_);
  or (_15290_, _15289_, _15287_);
  or (_15291_, _15290_, _15283_);
  and (_15292_, _15291_, _15258_);
  or (_15293_, _15292_, _02850_);
  or (_15294_, _04861_, _06675_);
  and (_15295_, _15294_, _02021_);
  and (_15296_, _15295_, _15293_);
  nor (_15297_, _06791_, _02021_);
  or (_15298_, _15297_, _06679_);
  or (_15299_, _15298_, _15296_);
  nand (_15300_, _06679_, _06184_);
  and (_15301_, _15300_, _15299_);
  or (_15302_, _15301_, _01997_);
  and (_15303_, _11715_, _04326_);
  nor (_15304_, _15303_, _15284_);
  nand (_15305_, _15304_, _01997_);
  and (_15306_, _15305_, _02861_);
  and (_15307_, _15306_, _15302_);
  and (_15308_, _15285_, _11747_);
  nor (_15309_, _15308_, _15284_);
  nor (_15310_, _15309_, _02861_);
  or (_15311_, _15310_, _05279_);
  or (_15312_, _15311_, _15307_);
  nor (_15313_, _05930_, _05926_);
  nor (_15314_, _15313_, _05932_);
  or (_15315_, _15314_, _05285_);
  and (_15316_, _15315_, _06700_);
  and (_15317_, _15316_, _15312_);
  or (_15318_, _15317_, _15257_);
  and (_15319_, _15318_, _08245_);
  or (_15320_, _15319_, _01963_);
  or (_15321_, _15320_, _15244_);
  and (_15322_, _15321_, _15231_);
  or (_15323_, _14906_, _08649_);
  and (_15324_, _15323_, _08648_);
  nor (_15325_, _15324_, _07308_);
  and (_15326_, _15324_, _07308_);
  nor (_15327_, _15326_, _15325_);
  nor (_15328_, _14915_, _14910_);
  and (_15329_, _15328_, \oc8051_golden_model_1.PSW [7]);
  nor (_15330_, _15329_, _15327_);
  and (_15331_, _15329_, _15327_);
  nor (_15332_, _15331_, _15330_);
  and (_15333_, _15332_, _06476_);
  or (_15334_, _15333_, _01549_);
  or (_15335_, _15334_, _15322_);
  nand (_15336_, _01922_, _01549_);
  and (_15337_, _15336_, _02408_);
  and (_15338_, _15337_, _15335_);
  nor (_15339_, _11713_, _06958_);
  nor (_15340_, _15339_, _15284_);
  nor (_15341_, _15340_, _02408_);
  or (_15342_, _15341_, _05994_);
  or (_15343_, _15342_, _15338_);
  and (_15344_, _15343_, _15218_);
  or (_15345_, _15344_, _02528_);
  and (_15346_, _04861_, _03680_);
  nor (_15347_, _15346_, _15208_);
  nand (_15348_, _15347_, _02528_);
  and (_15349_, _15348_, _02043_);
  and (_15350_, _15349_, _15345_);
  nor (_15351_, _11820_, _06472_);
  nor (_15352_, _15351_, _15208_);
  nor (_15353_, _15352_, _02043_);
  or (_15354_, _15353_, _06008_);
  or (_15355_, _15354_, _15350_);
  not (_15356_, _06027_);
  and (_15357_, _06032_, _15356_);
  or (_15358_, _15357_, _06355_);
  and (_15359_, _15358_, _15355_);
  and (_15360_, _15359_, _01609_);
  nor (_15361_, _01922_, _01609_);
  or (_15362_, _15361_, _01869_);
  or (_15363_, _15362_, _15360_);
  and (_15364_, _09920_, _03680_);
  nor (_15365_, _15364_, _15208_);
  nand (_15366_, _15365_, _01869_);
  and (_15367_, _15366_, _06985_);
  and (_15368_, _15367_, _15363_);
  nor (_15369_, _06985_, _01922_);
  or (_15370_, _15369_, _06990_);
  or (_15371_, _15370_, _15368_);
  and (_15372_, _15371_, _15215_);
  or (_15373_, _15372_, _06993_);
  and (_15374_, _15214_, _06993_);
  nor (_15375_, _15374_, _14757_);
  and (_15376_, _15375_, _15373_);
  or (_15377_, _15376_, _15213_);
  nand (_15378_, _15377_, _14766_);
  nand (_15379_, _06412_, _14761_);
  and (_15380_, _15379_, _07006_);
  and (_15381_, _15380_, _15378_);
  or (_15382_, _15381_, _15212_);
  and (_15383_, _15382_, _07014_);
  nor (_15384_, _11709_, _07014_);
  or (_15385_, _15384_, _07012_);
  or (_15386_, _15385_, _15383_);
  nand (_15387_, _07012_, _07308_);
  and (_15388_, _15387_, _02166_);
  and (_15389_, _15388_, _15386_);
  or (_15390_, _15389_, _15211_);
  and (_15391_, _15390_, _02912_);
  nor (_15392_, _15208_, _02912_);
  or (_15393_, _15392_, _07026_);
  or (_15394_, _15393_, _15391_);
  and (_15395_, _15394_, _15207_);
  nor (_15396_, _15395_, _07031_);
  and (_15397_, _07031_, _07213_);
  or (_15398_, _15397_, _02178_);
  or (_15399_, _15398_, _15396_);
  or (_15400_, _11707_, _07035_);
  and (_15401_, _15400_, _07046_);
  and (_15402_, _15401_, _15399_);
  and (_15403_, _07040_, _07306_);
  or (_15404_, _15403_, _15402_);
  and (_15405_, _15404_, _02176_);
  or (_15406_, _15365_, _11708_);
  nor (_15407_, _15406_, _02176_);
  or (_15408_, _15407_, _09858_);
  or (_15409_, _15408_, _15405_);
  and (_15410_, _15409_, _15206_);
  or (_15411_, _15410_, _13866_);
  or (_15412_, _06411_, _01858_);
  nand (_15413_, _15412_, _14184_);
  and (_15414_, _15413_, _15411_);
  nor (_15415_, _06411_, _07060_);
  or (_15416_, _15415_, _06462_);
  or (_15417_, _15416_, _15414_);
  nand (_15418_, _07214_, _06462_);
  and (_15419_, _15418_, _02172_);
  and (_15420_, _15419_, _15417_);
  nand (_15421_, _11708_, _07070_);
  and (_15422_, _15421_, _09854_);
  or (_15423_, _15422_, _15420_);
  and (_15424_, _15423_, _15205_);
  or (_15425_, _15424_, _02071_);
  nor (_15426_, _11833_, _06472_);
  nor (_15427_, _15426_, _15208_);
  nand (_15428_, _15427_, _02071_);
  and (_15429_, _15428_, _07084_);
  and (_15430_, _15429_, _15425_);
  nor (_15431_, _07106_, _06764_);
  nor (_15432_, _15431_, _07107_);
  and (_15433_, _15432_, _07085_);
  or (_15434_, _15433_, _07114_);
  or (_15435_, _15434_, _15430_);
  nor (_15436_, _07135_, _06603_);
  nor (_15437_, _15436_, _07136_);
  or (_15438_, _15437_, _07116_);
  and (_15439_, _15438_, _15435_);
  or (_15440_, _15439_, _02164_);
  nor (_15441_, _07166_, _06944_);
  nor (_15442_, _15441_, _07167_);
  or (_15443_, _15442_, _02165_);
  and (_15444_, _15443_, _07177_);
  and (_15445_, _15444_, _15440_);
  and (_15446_, _07197_, _07179_);
  nor (_15447_, _15446_, _07198_);
  and (_15448_, _15447_, _07144_);
  or (_15449_, _15448_, _07175_);
  or (_15450_, _15449_, _15445_);
  nand (_15451_, _07175_, _06079_);
  and (_15452_, _15451_, _06458_);
  and (_15453_, _15452_, _15450_);
  nor (_15454_, _06444_, _06412_);
  nor (_15455_, _15454_, _06445_);
  and (_15456_, _15455_, _06459_);
  or (_15457_, _15456_, _07210_);
  or (_15458_, _15457_, _15453_);
  nor (_15459_, _07244_, _07215_);
  nor (_15460_, _15459_, _07245_);
  or (_15461_, _15460_, _07212_);
  and (_15462_, _15461_, _15458_);
  or (_15463_, _15462_, _01890_);
  nor (_15464_, _07295_, _07264_);
  nor (_15465_, _15464_, _07296_);
  or (_15466_, _15465_, _01891_);
  and (_15467_, _15466_, _07256_);
  and (_15468_, _15467_, _15463_);
  nor (_15469_, _07333_, _07308_);
  nor (_15470_, _15469_, _07334_);
  and (_15471_, _15470_, _07253_);
  or (_15472_, _15471_, _07304_);
  or (_15473_, _15472_, _15468_);
  and (_15474_, _15473_, _15204_);
  or (_15475_, _15474_, _02201_);
  nand (_15476_, _15273_, _02201_);
  and (_15477_, _15476_, _07346_);
  and (_15478_, _15477_, _15475_);
  nor (_15479_, _07353_, _06026_);
  or (_15480_, _15479_, _07354_);
  nor (_15481_, _15480_, _07350_);
  nor (_15482_, _15481_, _10442_);
  or (_15483_, _15482_, _15478_);
  nand (_15484_, _07350_, _04776_);
  and (_15485_, _15484_, _01887_);
  and (_15486_, _15485_, _15483_);
  nor (_15487_, _15304_, _01887_);
  or (_15488_, _15487_, _01537_);
  or (_15489_, _15488_, _15486_);
  and (_15490_, _11887_, _03680_);
  nor (_15491_, _15490_, _15208_);
  nand (_15492_, _15491_, _01537_);
  and (_15493_, _15492_, _07368_);
  and (_15494_, _15493_, _15489_);
  nor (_15495_, _07378_, \oc8051_golden_model_1.ACC [6]);
  nor (_15496_, _15495_, _07379_);
  and (_15497_, _15496_, _07367_);
  or (_15498_, _15497_, _07374_);
  or (_15499_, _15498_, _15494_);
  nand (_15500_, _07374_, _04776_);
  and (_15501_, _15500_, _38087_);
  and (_15502_, _15501_, _15499_);
  or (_15503_, _15502_, _15203_);
  and (_40199_, _15503_, _37580_);
  not (_15504_, \oc8051_golden_model_1.DPL [0]);
  nor (_15505_, _38087_, _15504_);
  nor (_15506_, _03856_, _15504_);
  and (_15507_, _03856_, _03028_);
  or (_15508_, _15507_, _15506_);
  or (_15509_, _15508_, _05249_);
  and (_15510_, _03748_, \oc8051_golden_model_1.ACC [0]);
  or (_15511_, _15510_, _15506_);
  or (_15512_, _15511_, _02021_);
  nor (_15513_, _04106_, _07397_);
  or (_15514_, _15513_, _15506_);
  or (_15515_, _15514_, _02814_);
  and (_15516_, _15511_, _02817_);
  nor (_15517_, _02817_, _15504_);
  or (_15518_, _15517_, _02001_);
  or (_15519_, _15518_, _15516_);
  and (_15520_, _15519_, _02840_);
  and (_15521_, _15520_, _15515_);
  and (_15522_, _15508_, _01999_);
  or (_15523_, _15522_, _02006_);
  or (_15524_, _15523_, _15521_);
  and (_15525_, _15524_, _15512_);
  or (_15526_, _15525_, _07416_);
  nand (_15527_, _07416_, \oc8051_golden_model_1.DPL [0]);
  and (_15528_, _15527_, _07401_);
  and (_15529_, _15528_, _15526_);
  nor (_15530_, _02568_, _07401_);
  or (_15531_, _15530_, _05994_);
  or (_15532_, _15531_, _15529_);
  and (_15533_, _15532_, _15509_);
  or (_15534_, _15533_, _02528_);
  or (_15535_, _15506_, _02888_);
  and (_15536_, _04952_, _03748_);
  or (_15537_, _15536_, _15535_);
  and (_15538_, _15537_, _15534_);
  or (_15539_, _15538_, _01602_);
  nor (_15540_, _10600_, _07443_);
  or (_15541_, _15540_, _15506_);
  or (_15542_, _15541_, _02043_);
  and (_15543_, _15542_, _01870_);
  and (_15544_, _15543_, _15539_);
  and (_15545_, _03748_, _04562_);
  or (_15546_, _15545_, _15506_);
  and (_15547_, _15546_, _01869_);
  or (_15548_, _15547_, _02079_);
  or (_15549_, _15548_, _15544_);
  and (_15550_, _10614_, _03748_);
  or (_15551_, _15550_, _15506_);
  or (_15552_, _15551_, _02166_);
  and (_15553_, _15552_, _15549_);
  or (_15555_, _15553_, _02167_);
  and (_15556_, _10620_, _03856_);
  or (_15557_, _15506_, _02912_);
  or (_15558_, _15557_, _15556_);
  and (_15559_, _15558_, _02176_);
  and (_15560_, _15559_, _15555_);
  nand (_15561_, _15546_, _02072_);
  nor (_15562_, _15561_, _15513_);
  or (_15563_, _15562_, _15560_);
  and (_15564_, _15563_, _02907_);
  or (_15566_, _15506_, _04106_);
  and (_15567_, _15511_, _02177_);
  and (_15568_, _15567_, _15566_);
  or (_15569_, _15568_, _02071_);
  or (_15570_, _15569_, _15564_);
  nor (_15571_, _10613_, _07397_);
  or (_15572_, _15506_, _04788_);
  or (_15573_, _15572_, _15571_);
  and (_15574_, _15573_, _04793_);
  and (_15575_, _15574_, _15570_);
  not (_15577_, _02743_);
  nor (_15578_, _10619_, _07397_);
  or (_15579_, _15578_, _15506_);
  and (_15580_, _15579_, _02173_);
  or (_15581_, _15580_, _15577_);
  or (_15582_, _15581_, _15575_);
  or (_15583_, _15514_, _02743_);
  and (_15584_, _15583_, _38087_);
  and (_15585_, _15584_, _15582_);
  or (_15586_, _15585_, _15505_);
  and (_40200_, _15586_, _37580_);
  and (_15587_, _38088_, \oc8051_golden_model_1.DPL [1]);
  or (_15588_, _10822_, _07397_);
  or (_15589_, _03856_, \oc8051_golden_model_1.DPL [1]);
  and (_15590_, _15589_, _02167_);
  and (_15591_, _15590_, _15588_);
  nor (_15592_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.DPL [0]);
  nor (_15593_, _15592_, _07421_);
  and (_15594_, _15593_, _07416_);
  and (_15595_, _10698_, _03856_);
  not (_15598_, _15595_);
  and (_15599_, _15598_, _15589_);
  or (_15600_, _15599_, _02814_);
  nand (_15601_, _03856_, _01613_);
  and (_15602_, _15601_, _15589_);
  and (_15603_, _15602_, _02817_);
  and (_15604_, _02818_, \oc8051_golden_model_1.DPL [1]);
  or (_15605_, _15604_, _02001_);
  or (_15606_, _15605_, _15603_);
  and (_15607_, _15606_, _02840_);
  and (_15609_, _15607_, _15600_);
  and (_15610_, _07397_, \oc8051_golden_model_1.DPL [1]);
  nor (_15611_, _07397_, _02811_);
  or (_15612_, _15611_, _15610_);
  and (_15613_, _15612_, _01999_);
  or (_15614_, _15613_, _02006_);
  or (_15615_, _15614_, _15609_);
  or (_15616_, _15602_, _02021_);
  and (_15617_, _15616_, _07417_);
  and (_15618_, _15617_, _15615_);
  or (_15620_, _15618_, _15594_);
  and (_15621_, _15620_, _07401_);
  nor (_15622_, _02687_, _07401_);
  or (_15623_, _15622_, _05994_);
  or (_15624_, _15623_, _15621_);
  or (_15625_, _15612_, _05249_);
  and (_15626_, _15625_, _15624_);
  or (_15627_, _15626_, _02528_);
  and (_15628_, _04907_, _03748_);
  or (_15629_, _15610_, _02888_);
  or (_15631_, _15629_, _15628_);
  and (_15632_, _15631_, _02043_);
  and (_15633_, _15632_, _15627_);
  and (_15634_, _15589_, _01602_);
  nand (_15635_, _10802_, _03856_);
  and (_15636_, _15635_, _15634_);
  or (_15637_, _15636_, _15633_);
  and (_15638_, _15637_, _01870_);
  and (_15639_, _15589_, _01869_);
  nand (_15640_, _03856_, _02687_);
  and (_15642_, _15640_, _15639_);
  or (_15643_, _15642_, _15638_);
  and (_15644_, _15643_, _02166_);
  or (_15645_, _10816_, _07397_);
  and (_15646_, _15589_, _02079_);
  and (_15647_, _15646_, _15645_);
  or (_15648_, _15647_, _15644_);
  and (_15649_, _15648_, _02912_);
  or (_15650_, _15649_, _15591_);
  and (_15651_, _15650_, _02176_);
  or (_15653_, _10692_, _07397_);
  and (_15654_, _15589_, _02072_);
  and (_15655_, _15654_, _15653_);
  or (_15656_, _15655_, _15651_);
  and (_15657_, _15656_, _02907_);
  or (_15658_, _15610_, _04058_);
  and (_15659_, _15602_, _02177_);
  and (_15660_, _15659_, _15658_);
  or (_15661_, _15660_, _15657_);
  and (_15662_, _15661_, _02174_);
  or (_15664_, _15601_, _04058_);
  and (_15665_, _15589_, _02173_);
  and (_15666_, _15665_, _15664_);
  or (_15667_, _15666_, _02201_);
  or (_15668_, _15640_, _04058_);
  and (_15669_, _15589_, _02071_);
  and (_15670_, _15669_, _15668_);
  or (_15671_, _15670_, _15667_);
  or (_15672_, _15671_, _15662_);
  or (_15673_, _15599_, _02303_);
  and (_15675_, _15673_, _15672_);
  or (_15676_, _15675_, _01537_);
  or (_15677_, _15610_, _01538_);
  or (_15678_, _15677_, _15595_);
  and (_15679_, _15678_, _38087_);
  and (_15680_, _15679_, _15676_);
  or (_15681_, _15680_, _15587_);
  and (_40201_, _15681_, _37580_);
  and (_15682_, _38088_, \oc8051_golden_model_1.DPL [2]);
  and (_15683_, _07397_, \oc8051_golden_model_1.DPL [2]);
  nor (_15685_, _11019_, _07397_);
  or (_15686_, _15685_, _15683_);
  and (_15687_, _15686_, _02173_);
  or (_15688_, _15683_, _04156_);
  and (_15689_, _03748_, _04724_);
  or (_15690_, _15689_, _15683_);
  and (_15691_, _15690_, _02072_);
  and (_15692_, _15691_, _15688_);
  and (_15693_, _11020_, _03856_);
  or (_15694_, _15693_, _15683_);
  and (_15696_, _15694_, _02167_);
  nor (_15697_, _07397_, _03455_);
  or (_15698_, _15697_, _15683_);
  or (_15699_, _15698_, _05249_);
  nor (_15700_, _07421_, \oc8051_golden_model_1.DPL [2]);
  nor (_15701_, _15700_, _07422_);
  and (_15702_, _15701_, _07416_);
  nor (_15703_, _10905_, _07397_);
  or (_15704_, _15703_, _15683_);
  or (_15705_, _15704_, _02814_);
  and (_15707_, _03748_, \oc8051_golden_model_1.ACC [2]);
  or (_15708_, _15707_, _15683_);
  and (_15709_, _15708_, _02817_);
  and (_15710_, _02818_, \oc8051_golden_model_1.DPL [2]);
  or (_15711_, _15710_, _02001_);
  or (_15712_, _15711_, _15709_);
  and (_15713_, _15712_, _02840_);
  and (_15714_, _15713_, _15705_);
  and (_15715_, _15698_, _01999_);
  or (_15716_, _15715_, _02006_);
  or (_15718_, _15716_, _15714_);
  or (_15719_, _15708_, _02021_);
  and (_15720_, _15719_, _07417_);
  and (_15721_, _15720_, _15718_);
  or (_15722_, _15721_, _15702_);
  and (_15723_, _15722_, _07401_);
  nor (_15724_, _02338_, _07401_);
  or (_15725_, _15724_, _05994_);
  or (_15726_, _15725_, _15723_);
  and (_15727_, _15726_, _15699_);
  or (_15729_, _15727_, _02528_);
  or (_15730_, _15683_, _02888_);
  and (_15731_, _05043_, _03748_);
  or (_15732_, _15731_, _15730_);
  and (_15733_, _15732_, _02043_);
  and (_15734_, _15733_, _15729_);
  nor (_15735_, _11000_, _07443_);
  or (_15736_, _15735_, _15683_);
  and (_15737_, _15736_, _01602_);
  or (_15738_, _15737_, _01869_);
  or (_15740_, _15738_, _15734_);
  or (_15741_, _15690_, _01870_);
  and (_15742_, _15741_, _15740_);
  or (_15743_, _15742_, _02079_);
  and (_15744_, _11014_, _03856_);
  or (_15745_, _15683_, _02166_);
  or (_15746_, _15745_, _15744_);
  and (_15747_, _15746_, _02912_);
  and (_15748_, _15747_, _15743_);
  or (_15749_, _15748_, _15696_);
  and (_15751_, _15749_, _02176_);
  or (_15752_, _15751_, _15692_);
  and (_15753_, _15752_, _02907_);
  and (_15754_, _15708_, _02177_);
  and (_15755_, _15754_, _15688_);
  or (_15756_, _15755_, _02071_);
  or (_15757_, _15756_, _15753_);
  nor (_15758_, _11013_, _07397_);
  or (_15759_, _15683_, _04788_);
  or (_15760_, _15759_, _15758_);
  and (_15762_, _15760_, _04793_);
  and (_15763_, _15762_, _15757_);
  or (_15764_, _15763_, _15687_);
  and (_15765_, _15764_, _02303_);
  and (_15766_, _15704_, _02201_);
  or (_15767_, _15766_, _01537_);
  or (_15768_, _15767_, _15765_);
  and (_15769_, _11072_, _03856_);
  or (_15770_, _15683_, _01538_);
  or (_15771_, _15770_, _15769_);
  and (_15773_, _15771_, _38087_);
  and (_15774_, _15773_, _15768_);
  or (_15775_, _15774_, _15682_);
  and (_40203_, _15775_, _37580_);
  or (_15776_, _38087_, \oc8051_golden_model_1.DPL [3]);
  and (_15777_, _15776_, _37580_);
  and (_15778_, _07397_, \oc8051_golden_model_1.DPL [3]);
  and (_15779_, _11094_, _03856_);
  or (_15780_, _15779_, _15778_);
  and (_15781_, _15780_, _02167_);
  nor (_15783_, _07397_, _03268_);
  or (_15784_, _15783_, _15778_);
  or (_15785_, _15784_, _05249_);
  nor (_15786_, _07422_, \oc8051_golden_model_1.DPL [3]);
  nor (_15787_, _15786_, _07423_);
  and (_15788_, _15787_, _07416_);
  nor (_15789_, _11101_, _07397_);
  or (_15790_, _15789_, _15778_);
  or (_15791_, _15790_, _02814_);
  and (_15792_, _03748_, \oc8051_golden_model_1.ACC [3]);
  or (_15794_, _15792_, _15778_);
  and (_15795_, _15794_, _02817_);
  and (_15796_, _02818_, \oc8051_golden_model_1.DPL [3]);
  or (_15797_, _15796_, _02001_);
  or (_15798_, _15797_, _15795_);
  and (_15799_, _15798_, _02840_);
  and (_15800_, _15799_, _15791_);
  and (_15801_, _15784_, _01999_);
  or (_15802_, _15801_, _02006_);
  or (_15803_, _15802_, _15800_);
  or (_15805_, _15794_, _02021_);
  and (_15806_, _15805_, _07417_);
  and (_15807_, _15806_, _15803_);
  or (_15808_, _15807_, _15788_);
  and (_15809_, _15808_, _07401_);
  nor (_15810_, _02159_, _07401_);
  or (_15811_, _15810_, _05994_);
  or (_15812_, _15811_, _15809_);
  and (_15813_, _15812_, _15785_);
  or (_15814_, _15813_, _02528_);
  or (_15816_, _15778_, _02888_);
  and (_15817_, _04998_, _03748_);
  or (_15818_, _15817_, _15816_);
  and (_15819_, _15818_, _02043_);
  and (_15820_, _15819_, _15814_);
  nor (_15821_, _11206_, _07443_);
  or (_15822_, _15821_, _15778_);
  and (_15823_, _15822_, _01602_);
  or (_15824_, _15823_, _01869_);
  or (_15825_, _15824_, _15820_);
  and (_15827_, _03748_, _04678_);
  or (_15828_, _15827_, _15778_);
  or (_15829_, _15828_, _01870_);
  and (_15830_, _15829_, _15825_);
  or (_15831_, _15830_, _02079_);
  and (_15832_, _11222_, _03856_);
  or (_15833_, _15778_, _02166_);
  or (_15834_, _15833_, _15832_);
  and (_15835_, _15834_, _02912_);
  and (_15836_, _15835_, _15831_);
  or (_15838_, _15836_, _15781_);
  and (_15839_, _15838_, _02176_);
  or (_15840_, _15778_, _04014_);
  and (_15841_, _15828_, _02072_);
  and (_15842_, _15841_, _15840_);
  or (_15843_, _15842_, _15839_);
  and (_15844_, _15843_, _02907_);
  and (_15845_, _15794_, _02177_);
  and (_15846_, _15845_, _15840_);
  or (_15847_, _15846_, _02071_);
  or (_15849_, _15847_, _15844_);
  nor (_15850_, _11220_, _07397_);
  or (_15851_, _15778_, _04788_);
  or (_15852_, _15851_, _15850_);
  and (_15853_, _15852_, _04793_);
  and (_15854_, _15853_, _15849_);
  nor (_15855_, _11093_, _07397_);
  or (_15856_, _15855_, _15778_);
  and (_15857_, _15856_, _02173_);
  or (_15858_, _15857_, _02201_);
  or (_15860_, _15858_, _15854_);
  or (_15861_, _15790_, _02303_);
  and (_15862_, _15861_, _01538_);
  and (_15863_, _15862_, _15860_);
  and (_15864_, _11273_, _03856_);
  or (_15865_, _15864_, _15778_);
  and (_15866_, _15865_, _01537_);
  or (_15867_, _15866_, _38088_);
  or (_15868_, _15867_, _15863_);
  and (_40204_, _15868_, _15777_);
  or (_15870_, _38087_, \oc8051_golden_model_1.DPL [4]);
  and (_15871_, _15870_, _37580_);
  and (_15872_, _07397_, \oc8051_golden_model_1.DPL [4]);
  and (_15873_, _11431_, _03856_);
  or (_15874_, _15873_, _15872_);
  and (_15875_, _15874_, _02167_);
  nor (_15876_, _04211_, _07397_);
  or (_15877_, _15876_, _15872_);
  or (_15878_, _15877_, _05249_);
  nor (_15879_, _11317_, _07397_);
  or (_15881_, _15879_, _15872_);
  or (_15882_, _15881_, _02814_);
  and (_15883_, _03748_, \oc8051_golden_model_1.ACC [4]);
  or (_15884_, _15883_, _15872_);
  and (_15885_, _15884_, _02817_);
  and (_15886_, _02818_, \oc8051_golden_model_1.DPL [4]);
  or (_15887_, _15886_, _02001_);
  or (_15888_, _15887_, _15885_);
  and (_15889_, _15888_, _02840_);
  and (_15890_, _15889_, _15882_);
  and (_15892_, _15877_, _01999_);
  or (_15893_, _15892_, _02006_);
  or (_15894_, _15893_, _15890_);
  or (_15895_, _15884_, _02021_);
  and (_15896_, _15895_, _07417_);
  and (_15897_, _15896_, _15894_);
  nor (_15898_, _07423_, \oc8051_golden_model_1.DPL [4]);
  nor (_15899_, _15898_, _07424_);
  and (_15900_, _15899_, _07416_);
  or (_15901_, _15900_, _15897_);
  and (_15903_, _15901_, _07401_);
  nor (_15904_, _04657_, _07401_);
  or (_15905_, _15904_, _05994_);
  or (_15906_, _15905_, _15903_);
  and (_15907_, _15906_, _15878_);
  or (_15908_, _15907_, _02528_);
  or (_15909_, _15872_, _02888_);
  and (_15910_, _05135_, _03748_);
  or (_15911_, _15910_, _15909_);
  and (_15912_, _15911_, _02043_);
  and (_15914_, _15912_, _15908_);
  nor (_15915_, _11411_, _07443_);
  or (_15916_, _15915_, _15872_);
  and (_15917_, _15916_, _01602_);
  or (_15918_, _15917_, _01869_);
  or (_15919_, _15918_, _15914_);
  and (_15920_, _04694_, _03748_);
  or (_15921_, _15920_, _15872_);
  or (_15922_, _15921_, _01870_);
  and (_15923_, _15922_, _15919_);
  or (_15925_, _15923_, _02079_);
  and (_15926_, _11425_, _03856_);
  or (_15927_, _15872_, _02166_);
  or (_15928_, _15927_, _15926_);
  and (_15929_, _15928_, _02912_);
  and (_15930_, _15929_, _15925_);
  or (_15931_, _15930_, _15875_);
  and (_15932_, _15931_, _02176_);
  or (_15933_, _15872_, _04258_);
  and (_15934_, _15921_, _02072_);
  and (_15936_, _15934_, _15933_);
  or (_15937_, _15936_, _15932_);
  and (_15938_, _15937_, _02907_);
  and (_15939_, _15884_, _02177_);
  and (_15940_, _15939_, _15933_);
  or (_15941_, _15940_, _02071_);
  or (_15942_, _15941_, _15938_);
  nor (_15943_, _11424_, _07397_);
  or (_15944_, _15872_, _04788_);
  or (_15945_, _15944_, _15943_);
  and (_15947_, _15945_, _04793_);
  and (_15948_, _15947_, _15942_);
  nor (_15949_, _11430_, _07397_);
  or (_15950_, _15949_, _15872_);
  and (_15951_, _15950_, _02173_);
  or (_15952_, _15951_, _02201_);
  or (_15953_, _15952_, _15948_);
  or (_15954_, _15881_, _02303_);
  and (_15955_, _15954_, _01538_);
  and (_15956_, _15955_, _15953_);
  and (_15958_, _11487_, _03856_);
  or (_15959_, _15958_, _15872_);
  and (_15960_, _15959_, _01537_);
  or (_15961_, _15960_, _38088_);
  or (_15962_, _15961_, _15956_);
  and (_40205_, _15962_, _15871_);
  or (_15963_, _38087_, \oc8051_golden_model_1.DPL [5]);
  and (_15964_, _15963_, _37580_);
  and (_15965_, _07397_, \oc8051_golden_model_1.DPL [5]);
  and (_15966_, _11635_, _03856_);
  or (_15968_, _15966_, _15965_);
  and (_15969_, _15968_, _02167_);
  nor (_15970_, _03916_, _07397_);
  or (_15971_, _15970_, _15965_);
  or (_15972_, _15971_, _05249_);
  nor (_15973_, _11525_, _07397_);
  or (_15974_, _15973_, _15965_);
  or (_15975_, _15974_, _02814_);
  and (_15976_, _03748_, \oc8051_golden_model_1.ACC [5]);
  or (_15977_, _15976_, _15965_);
  and (_15979_, _15977_, _02817_);
  and (_15980_, _02818_, \oc8051_golden_model_1.DPL [5]);
  or (_15981_, _15980_, _02001_);
  or (_15982_, _15981_, _15979_);
  and (_15983_, _15982_, _02840_);
  and (_15984_, _15983_, _15975_);
  and (_15985_, _15971_, _01999_);
  or (_15986_, _15985_, _02006_);
  or (_15987_, _15986_, _15984_);
  or (_15988_, _15977_, _02021_);
  and (_15990_, _15988_, _07417_);
  and (_15991_, _15990_, _15987_);
  nor (_15992_, _07424_, \oc8051_golden_model_1.DPL [5]);
  nor (_15993_, _15992_, _07425_);
  and (_15994_, _15993_, _07416_);
  or (_15995_, _15994_, _15991_);
  and (_15996_, _15995_, _07401_);
  nor (_15997_, _04626_, _07401_);
  or (_15998_, _15997_, _05994_);
  or (_15999_, _15998_, _15996_);
  and (_16001_, _15999_, _15972_);
  or (_16002_, _16001_, _02528_);
  or (_16003_, _15965_, _02888_);
  and (_16004_, _05090_, _03748_);
  or (_16005_, _16004_, _16003_);
  and (_16006_, _16005_, _02043_);
  and (_16007_, _16006_, _16002_);
  nor (_16008_, _11615_, _07443_);
  or (_16009_, _16008_, _15965_);
  and (_16010_, _16009_, _01602_);
  or (_16012_, _16010_, _01869_);
  or (_16013_, _16012_, _16007_);
  and (_16014_, _04672_, _03748_);
  or (_16015_, _16014_, _15965_);
  or (_16016_, _16015_, _01870_);
  and (_16017_, _16016_, _16013_);
  or (_16018_, _16017_, _02079_);
  and (_16019_, _11629_, _03856_);
  or (_16020_, _15965_, _02166_);
  or (_16021_, _16020_, _16019_);
  and (_16023_, _16021_, _02912_);
  and (_16024_, _16023_, _16018_);
  or (_16025_, _16024_, _15969_);
  and (_16026_, _16025_, _02176_);
  or (_16027_, _15965_, _03965_);
  and (_16028_, _16015_, _02072_);
  and (_16029_, _16028_, _16027_);
  or (_16030_, _16029_, _16026_);
  and (_16031_, _16030_, _02907_);
  and (_16032_, _15977_, _02177_);
  and (_16033_, _16032_, _16027_);
  or (_16034_, _16033_, _02071_);
  or (_16035_, _16034_, _16031_);
  nor (_16036_, _11628_, _07397_);
  or (_16037_, _15965_, _04788_);
  or (_16038_, _16037_, _16036_);
  and (_16039_, _16038_, _04793_);
  and (_16040_, _16039_, _16035_);
  nor (_16041_, _11634_, _07397_);
  or (_16042_, _16041_, _15965_);
  and (_16045_, _16042_, _02173_);
  or (_16046_, _16045_, _02201_);
  or (_16047_, _16046_, _16040_);
  or (_16048_, _15974_, _02303_);
  and (_16049_, _16048_, _01538_);
  and (_16050_, _16049_, _16047_);
  and (_16051_, _11685_, _03856_);
  or (_16052_, _16051_, _15965_);
  and (_16053_, _16052_, _01537_);
  or (_16054_, _16053_, _38088_);
  or (_16056_, _16054_, _16050_);
  and (_40206_, _16056_, _15964_);
  or (_16057_, _38087_, \oc8051_golden_model_1.DPL [6]);
  and (_16058_, _16057_, _37580_);
  and (_16059_, _07397_, \oc8051_golden_model_1.DPL [6]);
  and (_16060_, _11709_, _03856_);
  or (_16061_, _16060_, _16059_);
  and (_16062_, _16061_, _02167_);
  nor (_16063_, _03808_, _07397_);
  or (_16064_, _16063_, _16059_);
  or (_16066_, _16064_, _05249_);
  nor (_16067_, _11730_, _07397_);
  or (_16068_, _16067_, _16059_);
  or (_16069_, _16068_, _02814_);
  and (_16070_, _03748_, \oc8051_golden_model_1.ACC [6]);
  or (_16071_, _16070_, _16059_);
  and (_16072_, _16071_, _02817_);
  and (_16073_, _02818_, \oc8051_golden_model_1.DPL [6]);
  or (_16074_, _16073_, _02001_);
  or (_16075_, _16074_, _16072_);
  and (_16077_, _16075_, _02840_);
  and (_16078_, _16077_, _16069_);
  and (_16079_, _16064_, _01999_);
  or (_16080_, _16079_, _02006_);
  or (_16081_, _16080_, _16078_);
  or (_16082_, _16071_, _02021_);
  and (_16083_, _16082_, _07417_);
  and (_16084_, _16083_, _16081_);
  nor (_16085_, _07425_, \oc8051_golden_model_1.DPL [6]);
  nor (_16086_, _16085_, _07426_);
  and (_16088_, _16086_, _07416_);
  or (_16089_, _16088_, _16084_);
  and (_16090_, _16089_, _07401_);
  nor (_16091_, _04594_, _07401_);
  or (_16092_, _16091_, _05994_);
  or (_16093_, _16092_, _16090_);
  and (_16094_, _16093_, _16066_);
  or (_16095_, _16094_, _02528_);
  or (_16096_, _16059_, _02888_);
  and (_16097_, _04861_, _03748_);
  or (_16099_, _16097_, _16096_);
  and (_16100_, _16099_, _02043_);
  and (_16101_, _16100_, _16095_);
  nor (_16102_, _11820_, _07443_);
  or (_16103_, _16102_, _16059_);
  and (_16104_, _16103_, _01602_);
  or (_16105_, _16104_, _01869_);
  or (_16106_, _16105_, _16101_);
  and (_16107_, _09920_, _03748_);
  or (_16108_, _16107_, _16059_);
  or (_16110_, _16108_, _01870_);
  and (_16111_, _16110_, _16106_);
  or (_16112_, _16111_, _02079_);
  and (_16113_, _11835_, _03856_);
  or (_16114_, _16059_, _02166_);
  or (_16115_, _16114_, _16113_);
  and (_16116_, _16115_, _02912_);
  and (_16117_, _16116_, _16112_);
  or (_16118_, _16117_, _16062_);
  and (_16119_, _16118_, _02176_);
  or (_16121_, _16059_, _03863_);
  and (_16122_, _16108_, _02072_);
  and (_16123_, _16122_, _16121_);
  or (_16124_, _16123_, _16119_);
  and (_16125_, _16124_, _02907_);
  and (_16126_, _16071_, _02177_);
  and (_16127_, _16126_, _16121_);
  or (_16128_, _16127_, _02071_);
  or (_16129_, _16128_, _16125_);
  nor (_16130_, _11833_, _07397_);
  or (_16132_, _16059_, _04788_);
  or (_16133_, _16132_, _16130_);
  and (_16134_, _16133_, _04793_);
  and (_16135_, _16134_, _16129_);
  nor (_16136_, _11708_, _07397_);
  or (_16137_, _16136_, _16059_);
  and (_16138_, _16137_, _02173_);
  or (_16139_, _16138_, _02201_);
  or (_16140_, _16139_, _16135_);
  or (_16141_, _16068_, _02303_);
  and (_16143_, _16141_, _01538_);
  and (_16144_, _16143_, _16140_);
  and (_16145_, _11887_, _03856_);
  or (_16146_, _16145_, _16059_);
  and (_16147_, _16146_, _01537_);
  or (_16148_, _16147_, _38088_);
  or (_16149_, _16148_, _16144_);
  and (_40207_, _16149_, _16058_);
  and (_16150_, _38088_, \oc8051_golden_model_1.DPH [0]);
  nor (_16151_, _07428_, \oc8051_golden_model_1.DPH [0]);
  nor (_16153_, _16151_, _07517_);
  and (_16154_, _16153_, _07416_);
  and (_16155_, _07495_, \oc8051_golden_model_1.DPH [0]);
  nor (_16156_, _04106_, _07495_);
  or (_16157_, _16156_, _16155_);
  or (_16158_, _16157_, _02814_);
  and (_16159_, _03741_, \oc8051_golden_model_1.ACC [0]);
  or (_16160_, _16159_, _16155_);
  and (_16161_, _16160_, _02817_);
  and (_16162_, _02818_, \oc8051_golden_model_1.DPH [0]);
  or (_16164_, _16162_, _02001_);
  or (_16165_, _16164_, _16161_);
  and (_16166_, _16165_, _02840_);
  and (_16167_, _16166_, _16158_);
  and (_16168_, _03850_, _03028_);
  or (_16169_, _16168_, _16155_);
  and (_16170_, _16169_, _01999_);
  or (_16171_, _16170_, _02006_);
  or (_16172_, _16171_, _16167_);
  or (_16173_, _16160_, _02021_);
  and (_16175_, _16173_, _07417_);
  and (_16176_, _16175_, _16172_);
  or (_16177_, _16176_, _16154_);
  and (_16178_, _16177_, _07401_);
  nor (_16179_, _02441_, _07401_);
  or (_16180_, _16179_, _05994_);
  or (_16181_, _16180_, _16178_);
  or (_16182_, _16169_, _05249_);
  and (_16183_, _16182_, _16181_);
  or (_16184_, _16183_, _02528_);
  and (_16186_, _04952_, _03741_);
  or (_16187_, _16155_, _02888_);
  or (_16188_, _16187_, _16186_);
  and (_16189_, _16188_, _16184_);
  or (_16190_, _16189_, _01602_);
  nor (_16191_, _10600_, _07540_);
  or (_16192_, _16191_, _16155_);
  or (_16193_, _16192_, _02043_);
  and (_16194_, _16193_, _01870_);
  and (_16195_, _16194_, _16190_);
  and (_16197_, _03741_, _04562_);
  or (_16198_, _16197_, _16155_);
  and (_16199_, _16198_, _01869_);
  or (_16200_, _16199_, _02079_);
  or (_16201_, _16200_, _16195_);
  and (_16202_, _10614_, _03741_);
  or (_16203_, _16202_, _16155_);
  or (_16204_, _16203_, _02166_);
  and (_16205_, _16204_, _16201_);
  or (_16206_, _16205_, _02167_);
  and (_16208_, _10620_, _03850_);
  or (_16209_, _16155_, _02912_);
  or (_16210_, _16209_, _16208_);
  and (_16211_, _16210_, _02176_);
  and (_16212_, _16211_, _16206_);
  nand (_16213_, _16198_, _02072_);
  nor (_16214_, _16213_, _16156_);
  or (_16215_, _16214_, _16212_);
  and (_16216_, _16215_, _02907_);
  or (_16217_, _16155_, _04106_);
  and (_16219_, _16160_, _02177_);
  and (_16220_, _16219_, _16217_);
  or (_16221_, _16220_, _02071_);
  or (_16222_, _16221_, _16216_);
  nor (_16223_, _10613_, _07495_);
  or (_16224_, _16155_, _04788_);
  or (_16225_, _16224_, _16223_);
  and (_16226_, _16225_, _04793_);
  and (_16227_, _16226_, _16222_);
  nor (_16228_, _10619_, _07495_);
  or (_16230_, _16228_, _16155_);
  and (_16231_, _16230_, _02173_);
  or (_16232_, _16231_, _15577_);
  or (_16233_, _16232_, _16227_);
  or (_16234_, _16157_, _02743_);
  and (_16235_, _16234_, _38087_);
  and (_16236_, _16235_, _16233_);
  or (_16237_, _16236_, _16150_);
  and (_40209_, _16237_, _37580_);
  and (_16238_, _38088_, \oc8051_golden_model_1.DPH [1]);
  or (_16240_, _10822_, _07495_);
  or (_16241_, _03850_, \oc8051_golden_model_1.DPH [1]);
  and (_16242_, _16241_, _02167_);
  and (_16243_, _16242_, _16240_);
  or (_16244_, _07517_, \oc8051_golden_model_1.DPH [1]);
  and (_16245_, _16244_, _07518_);
  and (_16246_, _16245_, _07416_);
  and (_16247_, _10698_, _03850_);
  not (_16248_, _16247_);
  and (_16249_, _16248_, _16241_);
  or (_16251_, _16249_, _02814_);
  nand (_16252_, _03850_, _01613_);
  and (_16253_, _16252_, _16241_);
  and (_16254_, _16253_, _02817_);
  and (_16255_, _02818_, \oc8051_golden_model_1.DPH [1]);
  or (_16256_, _16255_, _02001_);
  or (_16257_, _16256_, _16254_);
  and (_16258_, _16257_, _02840_);
  and (_16259_, _16258_, _16251_);
  and (_16260_, _07495_, \oc8051_golden_model_1.DPH [1]);
  nor (_16262_, _07495_, _02811_);
  or (_16263_, _16262_, _16260_);
  and (_16264_, _16263_, _01999_);
  or (_16265_, _16264_, _02006_);
  or (_16266_, _16265_, _16259_);
  or (_16267_, _16253_, _02021_);
  and (_16268_, _16267_, _07417_);
  and (_16269_, _16268_, _16266_);
  or (_16270_, _16269_, _16246_);
  and (_16271_, _16270_, _07401_);
  nor (_16273_, _07401_, _01822_);
  or (_16274_, _16273_, _05994_);
  or (_16275_, _16274_, _16271_);
  or (_16276_, _16263_, _05249_);
  and (_16277_, _16276_, _16275_);
  or (_16278_, _16277_, _02528_);
  and (_16279_, _04907_, _03741_);
  or (_16280_, _16260_, _02888_);
  or (_16281_, _16280_, _16279_);
  and (_16282_, _16281_, _02043_);
  and (_16284_, _16282_, _16278_);
  and (_16285_, _16241_, _01602_);
  nand (_16286_, _10802_, _03850_);
  and (_16287_, _16286_, _16285_);
  or (_16288_, _16287_, _16284_);
  and (_16289_, _16288_, _01870_);
  and (_16290_, _16241_, _01869_);
  nand (_16291_, _03850_, _02687_);
  and (_16292_, _16291_, _16290_);
  or (_16293_, _16292_, _16289_);
  and (_16295_, _16293_, _02166_);
  or (_16296_, _10816_, _07495_);
  and (_16297_, _16241_, _02079_);
  and (_16298_, _16297_, _16296_);
  or (_16299_, _16298_, _16295_);
  and (_16300_, _16299_, _02912_);
  or (_16301_, _16300_, _16243_);
  and (_16302_, _16301_, _02176_);
  or (_16303_, _10692_, _07495_);
  and (_16304_, _16241_, _02072_);
  and (_16306_, _16304_, _16303_);
  or (_16307_, _16306_, _16302_);
  and (_16308_, _16307_, _02907_);
  or (_16309_, _16260_, _04058_);
  and (_16310_, _16253_, _02177_);
  and (_16311_, _16310_, _16309_);
  or (_16312_, _16311_, _16308_);
  and (_16313_, _16312_, _02174_);
  or (_16314_, _16252_, _04058_);
  and (_16315_, _16241_, _02173_);
  and (_16317_, _16315_, _16314_);
  or (_16318_, _16317_, _02201_);
  or (_16319_, _16291_, _04058_);
  and (_16320_, _16241_, _02071_);
  and (_16321_, _16320_, _16319_);
  or (_16322_, _16321_, _16318_);
  or (_16323_, _16322_, _16313_);
  or (_16324_, _16249_, _02303_);
  and (_16325_, _16324_, _16323_);
  or (_16326_, _16325_, _01537_);
  or (_16328_, _16260_, _01538_);
  or (_16329_, _16328_, _16247_);
  and (_16330_, _16329_, _38087_);
  and (_16331_, _16330_, _16326_);
  or (_16332_, _16331_, _16238_);
  and (_40210_, _16332_, _37580_);
  nor (_16333_, _38087_, _07516_);
  nor (_16334_, _03850_, _07516_);
  nor (_16335_, _11019_, _07495_);
  or (_16336_, _16335_, _16334_);
  and (_16338_, _16336_, _02173_);
  and (_16339_, _11020_, _03850_);
  or (_16340_, _16339_, _16334_);
  and (_16341_, _16340_, _02167_);
  nor (_16342_, _07495_, _03455_);
  or (_16343_, _16342_, _16334_);
  or (_16344_, _16343_, _05249_);
  or (_16345_, _16343_, _02840_);
  nor (_16346_, _10905_, _07495_);
  or (_16347_, _16346_, _16334_);
  and (_16349_, _16347_, _02001_);
  nor (_16350_, _02817_, _07516_);
  and (_16351_, _03741_, \oc8051_golden_model_1.ACC [2]);
  or (_16352_, _16351_, _16334_);
  and (_16353_, _16352_, _02817_);
  or (_16354_, _16353_, _16350_);
  and (_16355_, _16354_, _02814_);
  or (_16356_, _16355_, _01999_);
  or (_16357_, _16356_, _16349_);
  and (_16358_, _16357_, _16345_);
  or (_16360_, _16358_, _02006_);
  or (_16361_, _16352_, _02021_);
  and (_16362_, _16361_, _07417_);
  and (_16363_, _16362_, _16360_);
  nand (_16364_, _07518_, _07516_);
  nor (_16365_, _07519_, _07417_);
  and (_16366_, _16365_, _16364_);
  or (_16367_, _16366_, _16363_);
  and (_16368_, _16367_, _07401_);
  nor (_16369_, _02294_, _07401_);
  or (_16371_, _16369_, _05994_);
  or (_16372_, _16371_, _16368_);
  and (_16373_, _16372_, _16344_);
  or (_16374_, _16373_, _02528_);
  or (_16375_, _16334_, _02888_);
  and (_16376_, _05043_, _03741_);
  or (_16377_, _16376_, _16375_);
  and (_16378_, _16377_, _02043_);
  and (_16379_, _16378_, _16374_);
  nor (_16380_, _11000_, _07540_);
  or (_16382_, _16380_, _16334_);
  and (_16383_, _16382_, _01602_);
  or (_16384_, _16383_, _01869_);
  or (_16385_, _16384_, _16379_);
  and (_16386_, _03741_, _04724_);
  or (_16387_, _16386_, _16334_);
  or (_16388_, _16387_, _01870_);
  and (_16389_, _16388_, _16385_);
  or (_16390_, _16389_, _02079_);
  and (_16391_, _11014_, _03850_);
  or (_16393_, _16334_, _02166_);
  or (_16394_, _16393_, _16391_);
  and (_16395_, _16394_, _02912_);
  and (_16396_, _16395_, _16390_);
  or (_16397_, _16396_, _16341_);
  and (_16398_, _16397_, _02176_);
  or (_16399_, _16334_, _04156_);
  and (_16400_, _16387_, _02072_);
  and (_16401_, _16400_, _16399_);
  or (_16402_, _16401_, _16398_);
  and (_16404_, _16402_, _02907_);
  and (_16405_, _16352_, _02177_);
  and (_16406_, _16405_, _16399_);
  or (_16407_, _16406_, _02071_);
  or (_16408_, _16407_, _16404_);
  nor (_16409_, _11013_, _07495_);
  or (_16410_, _16334_, _04788_);
  or (_16411_, _16410_, _16409_);
  and (_16412_, _16411_, _04793_);
  and (_16413_, _16412_, _16408_);
  or (_16415_, _16413_, _16338_);
  and (_16416_, _16415_, _02303_);
  and (_16417_, _16347_, _02201_);
  or (_16418_, _16417_, _01537_);
  or (_16419_, _16418_, _16416_);
  and (_16420_, _11072_, _03850_);
  or (_16421_, _16334_, _01538_);
  or (_16422_, _16421_, _16420_);
  and (_16423_, _16422_, _38087_);
  and (_16424_, _16423_, _16419_);
  or (_16426_, _16424_, _16333_);
  and (_40211_, _16426_, _37580_);
  or (_16427_, _38087_, \oc8051_golden_model_1.DPH [3]);
  and (_16428_, _16427_, _37580_);
  and (_16429_, _07495_, \oc8051_golden_model_1.DPH [3]);
  and (_16430_, _11094_, _03850_);
  or (_16431_, _16430_, _16429_);
  and (_16432_, _16431_, _02167_);
  nor (_16433_, _07495_, _03268_);
  or (_16434_, _16433_, _16429_);
  or (_16436_, _16434_, _05249_);
  or (_16437_, _07519_, \oc8051_golden_model_1.DPH [3]);
  nor (_16438_, _07520_, _07417_);
  and (_16439_, _16438_, _16437_);
  nor (_16440_, _11101_, _07495_);
  or (_16441_, _16440_, _16429_);
  or (_16442_, _16441_, _02814_);
  and (_16443_, _03741_, \oc8051_golden_model_1.ACC [3]);
  or (_16444_, _16443_, _16429_);
  and (_16445_, _16444_, _02817_);
  and (_16447_, _02818_, \oc8051_golden_model_1.DPH [3]);
  or (_16448_, _16447_, _02001_);
  or (_16449_, _16448_, _16445_);
  and (_16450_, _16449_, _02840_);
  and (_16451_, _16450_, _16442_);
  and (_16452_, _16434_, _01999_);
  or (_16453_, _16452_, _02006_);
  or (_16454_, _16453_, _16451_);
  or (_16455_, _16444_, _02021_);
  and (_16456_, _16455_, _07417_);
  and (_16458_, _16456_, _16454_);
  or (_16459_, _16458_, _16439_);
  and (_16460_, _16459_, _07401_);
  nor (_16461_, _07401_, _01954_);
  or (_16462_, _16461_, _05994_);
  or (_16463_, _16462_, _16460_);
  and (_16464_, _16463_, _16436_);
  or (_16465_, _16464_, _02528_);
  or (_16466_, _16429_, _02888_);
  and (_16467_, _04998_, _03741_);
  or (_16469_, _16467_, _16466_);
  and (_16470_, _16469_, _02043_);
  and (_16471_, _16470_, _16465_);
  nor (_16472_, _11206_, _07540_);
  or (_16473_, _16472_, _16429_);
  and (_16474_, _16473_, _01602_);
  or (_16475_, _16474_, _01869_);
  or (_16476_, _16475_, _16471_);
  and (_16477_, _03741_, _04678_);
  or (_16478_, _16477_, _16429_);
  or (_16480_, _16478_, _01870_);
  and (_16481_, _16480_, _16476_);
  or (_16482_, _16481_, _02079_);
  and (_16483_, _11222_, _03850_);
  or (_16484_, _16429_, _02166_);
  or (_16485_, _16484_, _16483_);
  and (_16486_, _16485_, _02912_);
  and (_16487_, _16486_, _16482_);
  or (_16488_, _16487_, _16432_);
  and (_16489_, _16488_, _02176_);
  or (_16491_, _16429_, _04014_);
  and (_16492_, _16478_, _02072_);
  and (_16493_, _16492_, _16491_);
  or (_16494_, _16493_, _16489_);
  and (_16495_, _16494_, _02907_);
  and (_16496_, _16444_, _02177_);
  and (_16497_, _16496_, _16491_);
  or (_16498_, _16497_, _02071_);
  or (_16499_, _16498_, _16495_);
  nor (_16500_, _11220_, _07495_);
  or (_16502_, _16429_, _04788_);
  or (_16503_, _16502_, _16500_);
  and (_16504_, _16503_, _04793_);
  and (_16505_, _16504_, _16499_);
  nor (_16506_, _11093_, _07495_);
  or (_16507_, _16506_, _16429_);
  and (_16508_, _16507_, _02173_);
  or (_16509_, _16508_, _02201_);
  or (_16510_, _16509_, _16505_);
  or (_16511_, _16441_, _02303_);
  and (_16513_, _16511_, _01538_);
  and (_16514_, _16513_, _16510_);
  and (_16515_, _11273_, _03850_);
  or (_16516_, _16515_, _16429_);
  and (_16517_, _16516_, _01537_);
  or (_16518_, _16517_, _38088_);
  or (_16519_, _16518_, _16514_);
  and (_40212_, _16519_, _16428_);
  or (_16520_, _38087_, \oc8051_golden_model_1.DPH [4]);
  and (_16521_, _16520_, _37580_);
  and (_16523_, _07495_, \oc8051_golden_model_1.DPH [4]);
  and (_16524_, _11431_, _03850_);
  or (_16525_, _16524_, _16523_);
  and (_16526_, _16525_, _02167_);
  nor (_16527_, _04211_, _07495_);
  or (_16528_, _16527_, _16523_);
  or (_16529_, _16528_, _05249_);
  nor (_16530_, _11317_, _07495_);
  or (_16531_, _16530_, _16523_);
  or (_16532_, _16531_, _02814_);
  and (_16534_, _03741_, \oc8051_golden_model_1.ACC [4]);
  or (_16535_, _16534_, _16523_);
  and (_16536_, _16535_, _02817_);
  and (_16537_, _02818_, \oc8051_golden_model_1.DPH [4]);
  or (_16538_, _16537_, _02001_);
  or (_16539_, _16538_, _16536_);
  and (_16540_, _16539_, _02840_);
  and (_16541_, _16540_, _16532_);
  and (_16542_, _16528_, _01999_);
  or (_16543_, _16542_, _02006_);
  or (_16545_, _16543_, _16541_);
  or (_16546_, _16535_, _02021_);
  and (_16547_, _16546_, _07417_);
  and (_16548_, _16547_, _16545_);
  or (_16549_, _07520_, \oc8051_golden_model_1.DPH [4]);
  nor (_16550_, _07521_, _07417_);
  and (_16551_, _16550_, _16549_);
  or (_16552_, _16551_, _16548_);
  and (_16553_, _16552_, _07401_);
  nor (_16554_, _07401_, _01855_);
  or (_16556_, _16554_, _05994_);
  or (_16557_, _16556_, _16553_);
  and (_16558_, _16557_, _16529_);
  or (_16559_, _16558_, _02528_);
  or (_16560_, _16523_, _02888_);
  and (_16561_, _05135_, _03741_);
  or (_16562_, _16561_, _16560_);
  and (_16563_, _16562_, _02043_);
  and (_16564_, _16563_, _16559_);
  nor (_16565_, _11411_, _07540_);
  or (_16567_, _16565_, _16523_);
  and (_16568_, _16567_, _01602_);
  or (_16569_, _16568_, _01869_);
  or (_16570_, _16569_, _16564_);
  and (_16571_, _04694_, _03741_);
  or (_16572_, _16571_, _16523_);
  or (_16573_, _16572_, _01870_);
  and (_16574_, _16573_, _16570_);
  or (_16575_, _16574_, _02079_);
  and (_16576_, _11425_, _03850_);
  or (_16578_, _16523_, _02166_);
  or (_16579_, _16578_, _16576_);
  and (_16580_, _16579_, _02912_);
  and (_16581_, _16580_, _16575_);
  or (_16582_, _16581_, _16526_);
  and (_16583_, _16582_, _02176_);
  or (_16584_, _16523_, _04258_);
  and (_16585_, _16572_, _02072_);
  and (_16586_, _16585_, _16584_);
  or (_16587_, _16586_, _16583_);
  and (_16589_, _16587_, _02907_);
  and (_16590_, _16535_, _02177_);
  and (_16591_, _16590_, _16584_);
  or (_16592_, _16591_, _02071_);
  or (_16593_, _16592_, _16589_);
  nor (_16594_, _11424_, _07495_);
  or (_16595_, _16523_, _04788_);
  or (_16596_, _16595_, _16594_);
  and (_16597_, _16596_, _04793_);
  and (_16598_, _16597_, _16593_);
  nor (_16600_, _11430_, _07495_);
  or (_16601_, _16600_, _16523_);
  and (_16602_, _16601_, _02173_);
  or (_16603_, _16602_, _02201_);
  or (_16604_, _16603_, _16598_);
  or (_16605_, _16531_, _02303_);
  and (_16606_, _16605_, _01538_);
  and (_16607_, _16606_, _16604_);
  and (_16608_, _11487_, _03850_);
  or (_16609_, _16608_, _16523_);
  and (_16611_, _16609_, _01537_);
  or (_16612_, _16611_, _38088_);
  or (_16613_, _16612_, _16607_);
  and (_40213_, _16613_, _16521_);
  or (_16614_, _38087_, \oc8051_golden_model_1.DPH [5]);
  and (_16615_, _16614_, _37580_);
  and (_16616_, _07495_, \oc8051_golden_model_1.DPH [5]);
  and (_16617_, _11635_, _03850_);
  or (_16618_, _16617_, _16616_);
  and (_16619_, _16618_, _02167_);
  nor (_16621_, _03916_, _07495_);
  or (_16622_, _16621_, _16616_);
  or (_16623_, _16622_, _05249_);
  nor (_16624_, _11525_, _07495_);
  or (_16625_, _16624_, _16616_);
  or (_16626_, _16625_, _02814_);
  and (_16627_, _03741_, \oc8051_golden_model_1.ACC [5]);
  or (_16628_, _16627_, _16616_);
  and (_16629_, _16628_, _02817_);
  and (_16630_, _02818_, \oc8051_golden_model_1.DPH [5]);
  or (_16632_, _16630_, _02001_);
  or (_16633_, _16632_, _16629_);
  and (_16634_, _16633_, _02840_);
  and (_16635_, _16634_, _16626_);
  and (_16636_, _16622_, _01999_);
  or (_16637_, _16636_, _02006_);
  or (_16638_, _16637_, _16635_);
  or (_16639_, _16628_, _02021_);
  and (_16640_, _16639_, _07417_);
  and (_16641_, _16640_, _16638_);
  or (_16643_, _07521_, \oc8051_golden_model_1.DPH [5]);
  nor (_16644_, _07522_, _07417_);
  and (_16645_, _16644_, _16643_);
  or (_16646_, _16645_, _16641_);
  and (_16647_, _16646_, _07401_);
  nor (_16648_, _02252_, _07401_);
  or (_16649_, _16648_, _05994_);
  or (_16650_, _16649_, _16647_);
  and (_16651_, _16650_, _16623_);
  or (_16652_, _16651_, _02528_);
  or (_16654_, _16616_, _02888_);
  and (_16655_, _05090_, _03741_);
  or (_16656_, _16655_, _16654_);
  and (_16657_, _16656_, _02043_);
  and (_16658_, _16657_, _16652_);
  nor (_16659_, _11615_, _07540_);
  or (_16660_, _16659_, _16616_);
  and (_16661_, _16660_, _01602_);
  or (_16662_, _16661_, _01869_);
  or (_16663_, _16662_, _16658_);
  and (_16664_, _04672_, _03741_);
  or (_16665_, _16664_, _16616_);
  or (_16666_, _16665_, _01870_);
  and (_16667_, _16666_, _16663_);
  or (_16668_, _16667_, _02079_);
  and (_16669_, _11629_, _03850_);
  or (_16670_, _16616_, _02166_);
  or (_16671_, _16670_, _16669_);
  and (_16672_, _16671_, _02912_);
  and (_16673_, _16672_, _16668_);
  or (_16676_, _16673_, _16619_);
  and (_16677_, _16676_, _02176_);
  or (_16678_, _16616_, _03965_);
  and (_16679_, _16665_, _02072_);
  and (_16680_, _16679_, _16678_);
  or (_16681_, _16680_, _16677_);
  and (_16682_, _16681_, _02907_);
  and (_16683_, _16628_, _02177_);
  and (_16684_, _16683_, _16678_);
  or (_16685_, _16684_, _02071_);
  or (_16687_, _16685_, _16682_);
  nor (_16688_, _11628_, _07495_);
  or (_16689_, _16616_, _04788_);
  or (_16690_, _16689_, _16688_);
  and (_16691_, _16690_, _04793_);
  and (_16692_, _16691_, _16687_);
  nor (_16693_, _11634_, _07495_);
  or (_16694_, _16693_, _16616_);
  and (_16695_, _16694_, _02173_);
  or (_16696_, _16695_, _02201_);
  or (_16698_, _16696_, _16692_);
  or (_16699_, _16625_, _02303_);
  and (_16700_, _16699_, _01538_);
  and (_16701_, _16700_, _16698_);
  and (_16702_, _11685_, _03850_);
  or (_16703_, _16702_, _16616_);
  and (_16704_, _16703_, _01537_);
  or (_16705_, _16704_, _38088_);
  or (_16706_, _16705_, _16701_);
  and (_40214_, _16706_, _16615_);
  or (_16708_, _38087_, \oc8051_golden_model_1.DPH [6]);
  and (_16709_, _16708_, _37580_);
  nor (_16710_, _03850_, _10272_);
  and (_16711_, _11709_, _03850_);
  or (_16712_, _16711_, _16710_);
  and (_16713_, _16712_, _02167_);
  nor (_16714_, _03808_, _07495_);
  or (_16715_, _16714_, _16710_);
  or (_16716_, _16715_, _05249_);
  nor (_16717_, _11730_, _07495_);
  or (_16719_, _16717_, _16710_);
  or (_16720_, _16719_, _02814_);
  and (_16721_, _03741_, \oc8051_golden_model_1.ACC [6]);
  or (_16722_, _16721_, _16710_);
  and (_16723_, _16722_, _02817_);
  nor (_16724_, _02817_, _10272_);
  or (_16725_, _16724_, _02001_);
  or (_16726_, _16725_, _16723_);
  and (_16727_, _16726_, _02840_);
  and (_16728_, _16727_, _16720_);
  and (_16730_, _16715_, _01999_);
  or (_16731_, _16730_, _02006_);
  or (_16732_, _16731_, _16728_);
  or (_16733_, _16722_, _02021_);
  and (_16734_, _16733_, _07417_);
  and (_16735_, _16734_, _16732_);
  or (_16736_, _07522_, \oc8051_golden_model_1.DPH [6]);
  nor (_16737_, _07523_, _07417_);
  and (_16738_, _16737_, _16736_);
  or (_16739_, _16738_, _16735_);
  and (_16741_, _16739_, _07401_);
  nor (_16742_, _07401_, _01922_);
  or (_16743_, _16742_, _05994_);
  or (_16744_, _16743_, _16741_);
  and (_16745_, _16744_, _16716_);
  or (_16746_, _16745_, _02528_);
  or (_16747_, _16710_, _02888_);
  and (_16748_, _04861_, _03741_);
  or (_16749_, _16748_, _16747_);
  and (_16750_, _16749_, _02043_);
  and (_16752_, _16750_, _16746_);
  nor (_16753_, _11820_, _07540_);
  or (_16754_, _16753_, _16710_);
  and (_16755_, _16754_, _01602_);
  or (_16756_, _16755_, _01869_);
  or (_16757_, _16756_, _16752_);
  and (_16758_, _09920_, _03741_);
  or (_16759_, _16758_, _16710_);
  or (_16760_, _16759_, _01870_);
  and (_16761_, _16760_, _16757_);
  or (_16763_, _16761_, _02079_);
  and (_16764_, _11835_, _03850_);
  or (_16765_, _16710_, _02166_);
  or (_16766_, _16765_, _16764_);
  and (_16767_, _16766_, _02912_);
  and (_16768_, _16767_, _16763_);
  or (_16769_, _16768_, _16713_);
  and (_16770_, _16769_, _02176_);
  or (_16771_, _16710_, _03863_);
  and (_16772_, _16759_, _02072_);
  and (_16774_, _16772_, _16771_);
  or (_16775_, _16774_, _16770_);
  and (_16776_, _16775_, _02907_);
  and (_16777_, _16722_, _02177_);
  and (_16778_, _16777_, _16771_);
  or (_16779_, _16778_, _02071_);
  or (_16780_, _16779_, _16776_);
  nor (_16781_, _11833_, _07495_);
  or (_16782_, _16710_, _04788_);
  or (_16783_, _16782_, _16781_);
  and (_16785_, _16783_, _04793_);
  and (_16786_, _16785_, _16780_);
  nor (_16787_, _11708_, _07495_);
  or (_16788_, _16787_, _16710_);
  and (_16789_, _16788_, _02173_);
  or (_16790_, _16789_, _02201_);
  or (_16791_, _16790_, _16786_);
  or (_16792_, _16719_, _02303_);
  and (_16793_, _16792_, _01538_);
  and (_16794_, _16793_, _16791_);
  and (_16796_, _11887_, _03850_);
  or (_16797_, _16796_, _16710_);
  and (_16798_, _16797_, _01537_);
  or (_16799_, _16798_, _38088_);
  or (_16800_, _16799_, _16794_);
  and (_40215_, _16800_, _16709_);
  and (_16801_, _38088_, \oc8051_golden_model_1.IE [0]);
  and (_16802_, _07586_, \oc8051_golden_model_1.IE [0]);
  and (_16803_, _10620_, _03633_);
  or (_16804_, _16803_, _16802_);
  and (_16806_, _16804_, _02167_);
  and (_16807_, _03633_, _03028_);
  or (_16808_, _16807_, _16802_);
  or (_16809_, _16808_, _05249_);
  nor (_16810_, _04106_, _07586_);
  or (_16811_, _16810_, _16802_);
  or (_16812_, _16811_, _02814_);
  and (_16813_, _03633_, \oc8051_golden_model_1.ACC [0]);
  or (_16814_, _16813_, _16802_);
  and (_16815_, _16814_, _02817_);
  and (_16817_, _02818_, \oc8051_golden_model_1.IE [0]);
  or (_16818_, _16817_, _02001_);
  or (_16819_, _16818_, _16815_);
  and (_16820_, _16819_, _02024_);
  and (_16821_, _16820_, _16812_);
  and (_16822_, _07594_, \oc8051_golden_model_1.IE [0]);
  and (_16823_, _10510_, _04333_);
  or (_16824_, _16823_, _16822_);
  and (_16825_, _16824_, _02007_);
  or (_16826_, _16825_, _16821_);
  and (_16828_, _16826_, _02840_);
  and (_16829_, _16808_, _01999_);
  or (_16830_, _16829_, _02006_);
  or (_16831_, _16830_, _16828_);
  or (_16832_, _16814_, _02021_);
  and (_16833_, _16832_, _02025_);
  and (_16834_, _16833_, _16831_);
  and (_16835_, _16802_, _01997_);
  or (_16836_, _16835_, _01991_);
  or (_16837_, _16836_, _16834_);
  or (_16839_, _16811_, _02861_);
  and (_16840_, _16839_, _02408_);
  and (_16841_, _16840_, _16837_);
  nor (_16842_, _10542_, _07594_);
  or (_16843_, _16842_, _16822_);
  and (_16844_, _16843_, _01875_);
  or (_16845_, _16844_, _05994_);
  or (_16846_, _16845_, _16841_);
  and (_16847_, _16846_, _16809_);
  or (_16848_, _16847_, _02528_);
  and (_16850_, _04952_, _03633_);
  or (_16851_, _16802_, _02888_);
  or (_16852_, _16851_, _16850_);
  and (_16853_, _16852_, _02043_);
  and (_16854_, _16853_, _16848_);
  nor (_16855_, _10600_, _07586_);
  or (_16856_, _16855_, _16802_);
  and (_16857_, _16856_, _01602_);
  or (_16858_, _16857_, _01869_);
  or (_16859_, _16858_, _16854_);
  and (_16861_, _03633_, _04562_);
  or (_16862_, _16861_, _16802_);
  or (_16863_, _16862_, _01870_);
  and (_16864_, _16863_, _16859_);
  or (_16865_, _16864_, _02079_);
  and (_16866_, _10614_, _03633_);
  or (_16867_, _16802_, _02166_);
  or (_16868_, _16867_, _16866_);
  and (_16869_, _16868_, _02912_);
  and (_16870_, _16869_, _16865_);
  or (_16872_, _16870_, _16806_);
  and (_16873_, _16872_, _02176_);
  nand (_16874_, _16862_, _02072_);
  nor (_16875_, _16874_, _16810_);
  or (_16876_, _16875_, _16873_);
  and (_16877_, _16876_, _02907_);
  or (_16878_, _16802_, _04106_);
  and (_16879_, _16814_, _02177_);
  and (_16880_, _16879_, _16878_);
  or (_16881_, _16880_, _02071_);
  or (_16883_, _16881_, _16877_);
  nor (_16884_, _10613_, _07586_);
  or (_16885_, _16802_, _04788_);
  or (_16886_, _16885_, _16884_);
  and (_16887_, _16886_, _04793_);
  and (_16888_, _16887_, _16883_);
  nor (_16889_, _10619_, _07586_);
  or (_16890_, _16889_, _16802_);
  and (_16891_, _16890_, _02173_);
  or (_16892_, _16891_, _02201_);
  or (_16894_, _16892_, _16888_);
  or (_16895_, _16811_, _02303_);
  and (_16896_, _16895_, _01887_);
  and (_16897_, _16896_, _16894_);
  and (_16898_, _16802_, _01860_);
  or (_16899_, _16898_, _01537_);
  or (_16900_, _16899_, _16897_);
  or (_16901_, _16811_, _01538_);
  and (_16902_, _16901_, _38087_);
  and (_16903_, _16902_, _16900_);
  or (_16905_, _16903_, _16801_);
  and (_40217_, _16905_, _37580_);
  and (_16906_, _38088_, \oc8051_golden_model_1.IE [1]);
  and (_16907_, _07586_, \oc8051_golden_model_1.IE [1]);
  nor (_16908_, _07586_, _02811_);
  or (_16909_, _16908_, _16907_);
  or (_16910_, _16909_, _02840_);
  or (_16911_, _03633_, \oc8051_golden_model_1.IE [1]);
  and (_16912_, _10698_, _03633_);
  not (_16913_, _16912_);
  and (_16915_, _16913_, _16911_);
  or (_16916_, _16915_, _02814_);
  nand (_16917_, _03633_, _01613_);
  and (_16918_, _16917_, _16911_);
  and (_16919_, _16918_, _02817_);
  and (_16920_, _02818_, \oc8051_golden_model_1.IE [1]);
  or (_16921_, _16920_, _02001_);
  or (_16922_, _16921_, _16919_);
  and (_16923_, _16922_, _02024_);
  and (_16924_, _16923_, _16916_);
  and (_16926_, _07594_, \oc8051_golden_model_1.IE [1]);
  and (_16927_, _10710_, _04333_);
  or (_16928_, _16927_, _16926_);
  and (_16929_, _16928_, _02007_);
  or (_16930_, _16929_, _01999_);
  or (_16931_, _16930_, _16924_);
  and (_16932_, _16931_, _16910_);
  or (_16933_, _16932_, _02006_);
  or (_16934_, _16918_, _02021_);
  and (_16935_, _16934_, _02025_);
  and (_16937_, _16935_, _16933_);
  and (_16938_, _10696_, _04333_);
  or (_16939_, _16938_, _16926_);
  and (_16940_, _16939_, _01997_);
  or (_16941_, _16940_, _01991_);
  or (_16942_, _16941_, _16937_);
  and (_16943_, _16927_, _10725_);
  or (_16944_, _16926_, _02861_);
  or (_16945_, _16944_, _16943_);
  and (_16946_, _16945_, _16942_);
  and (_16948_, _16946_, _02408_);
  nor (_16949_, _10742_, _07594_);
  or (_16950_, _16926_, _16949_);
  and (_16951_, _16950_, _01875_);
  or (_16952_, _16951_, _05994_);
  or (_16953_, _16952_, _16948_);
  or (_16954_, _16909_, _05249_);
  and (_16955_, _16954_, _16953_);
  or (_16956_, _16955_, _02528_);
  and (_16957_, _04907_, _03633_);
  or (_16959_, _16907_, _02888_);
  or (_16960_, _16959_, _16957_);
  and (_16961_, _16960_, _02043_);
  and (_16962_, _16961_, _16956_);
  nor (_16963_, _10802_, _07586_);
  or (_16964_, _16963_, _16907_);
  and (_16965_, _16964_, _01602_);
  or (_16966_, _16965_, _16962_);
  and (_16967_, _16966_, _01870_);
  nand (_16968_, _03633_, _02687_);
  and (_16970_, _16911_, _01869_);
  and (_16971_, _16970_, _16968_);
  or (_16972_, _16971_, _16967_);
  and (_16973_, _16972_, _02166_);
  or (_16974_, _10816_, _07586_);
  and (_16975_, _16911_, _02079_);
  and (_16976_, _16975_, _16974_);
  or (_16977_, _16976_, _16973_);
  and (_16978_, _16977_, _02912_);
  or (_16979_, _10822_, _07586_);
  and (_16981_, _16911_, _02167_);
  and (_16982_, _16981_, _16979_);
  or (_16983_, _16982_, _16978_);
  and (_16984_, _16983_, _02176_);
  or (_16985_, _10692_, _07586_);
  and (_16986_, _16911_, _02072_);
  and (_16987_, _16986_, _16985_);
  or (_16988_, _16987_, _16984_);
  and (_16989_, _16988_, _02907_);
  or (_16990_, _16907_, _04058_);
  and (_16992_, _16918_, _02177_);
  and (_16993_, _16992_, _16990_);
  or (_16994_, _16993_, _16989_);
  and (_16995_, _16994_, _02174_);
  or (_16996_, _16917_, _04058_);
  and (_16997_, _16911_, _02173_);
  and (_16998_, _16997_, _16996_);
  or (_16999_, _16998_, _02201_);
  or (_17000_, _16968_, _04058_);
  and (_17001_, _16911_, _02071_);
  and (_17003_, _17001_, _17000_);
  or (_17004_, _17003_, _16999_);
  or (_17005_, _17004_, _16995_);
  or (_17006_, _16915_, _02303_);
  and (_17007_, _17006_, _01887_);
  and (_17008_, _17007_, _17005_);
  and (_17009_, _16939_, _01860_);
  or (_17010_, _17009_, _01537_);
  or (_17011_, _17010_, _17008_);
  or (_17012_, _16907_, _01538_);
  or (_17014_, _17012_, _16912_);
  and (_17015_, _17014_, _38087_);
  and (_17016_, _17015_, _17011_);
  or (_17017_, _17016_, _16906_);
  and (_40218_, _17017_, _37580_);
  and (_17018_, _38088_, \oc8051_golden_model_1.IE [2]);
  and (_17019_, _07586_, \oc8051_golden_model_1.IE [2]);
  and (_17020_, _11020_, _03633_);
  or (_17021_, _17020_, _17019_);
  and (_17022_, _17021_, _02167_);
  nor (_17024_, _07586_, _03455_);
  or (_17025_, _17024_, _17019_);
  or (_17026_, _17025_, _05249_);
  or (_17027_, _17025_, _02840_);
  nor (_17028_, _10905_, _07586_);
  or (_17029_, _17028_, _17019_);
  or (_17030_, _17029_, _02814_);
  and (_17031_, _03633_, \oc8051_golden_model_1.ACC [2]);
  or (_17032_, _17031_, _17019_);
  and (_17033_, _17032_, _02817_);
  and (_17035_, _02818_, \oc8051_golden_model_1.IE [2]);
  or (_17036_, _17035_, _02001_);
  or (_17037_, _17036_, _17033_);
  and (_17038_, _17037_, _02024_);
  and (_17039_, _17038_, _17030_);
  and (_17040_, _07594_, \oc8051_golden_model_1.IE [2]);
  and (_17041_, _10909_, _04333_);
  or (_17042_, _17041_, _17040_);
  and (_17043_, _17042_, _02007_);
  or (_17044_, _17043_, _01999_);
  or (_17045_, _17044_, _17039_);
  and (_17046_, _17045_, _17027_);
  or (_17047_, _17046_, _02006_);
  or (_17048_, _17032_, _02021_);
  and (_17049_, _17048_, _02025_);
  and (_17050_, _17049_, _17047_);
  and (_17051_, _10894_, _04333_);
  or (_17052_, _17051_, _17040_);
  and (_17053_, _17052_, _01997_);
  or (_17054_, _17053_, _01991_);
  or (_17057_, _17054_, _17050_);
  and (_17058_, _17041_, _10924_);
  or (_17059_, _17040_, _02861_);
  or (_17060_, _17059_, _17058_);
  and (_17061_, _17060_, _02408_);
  and (_17062_, _17061_, _17057_);
  nor (_17063_, _10942_, _07594_);
  or (_17064_, _17063_, _17040_);
  and (_17065_, _17064_, _01875_);
  or (_17066_, _17065_, _05994_);
  or (_17068_, _17066_, _17062_);
  and (_17069_, _17068_, _17026_);
  or (_17070_, _17069_, _02528_);
  and (_17071_, _05043_, _03633_);
  or (_17072_, _17019_, _02888_);
  or (_17073_, _17072_, _17071_);
  and (_17074_, _17073_, _02043_);
  and (_17075_, _17074_, _17070_);
  nor (_17076_, _11000_, _07586_);
  or (_17077_, _17076_, _17019_);
  and (_17079_, _17077_, _01602_);
  or (_17080_, _17079_, _01869_);
  or (_17081_, _17080_, _17075_);
  and (_17082_, _03633_, _04724_);
  or (_17083_, _17082_, _17019_);
  or (_17084_, _17083_, _01870_);
  and (_17085_, _17084_, _17081_);
  or (_17086_, _17085_, _02079_);
  and (_17087_, _11014_, _03633_);
  or (_17088_, _17019_, _02166_);
  or (_17090_, _17088_, _17087_);
  and (_17091_, _17090_, _02912_);
  and (_17092_, _17091_, _17086_);
  or (_17093_, _17092_, _17022_);
  and (_17094_, _17093_, _02176_);
  or (_17095_, _17019_, _04156_);
  and (_17096_, _17083_, _02072_);
  and (_17097_, _17096_, _17095_);
  or (_17098_, _17097_, _17094_);
  and (_17099_, _17098_, _02907_);
  and (_17101_, _17032_, _02177_);
  and (_17102_, _17101_, _17095_);
  or (_17103_, _17102_, _02071_);
  or (_17104_, _17103_, _17099_);
  nor (_17105_, _11013_, _07586_);
  or (_17106_, _17019_, _04788_);
  or (_17107_, _17106_, _17105_);
  and (_17108_, _17107_, _04793_);
  and (_17109_, _17108_, _17104_);
  nor (_17110_, _11019_, _07586_);
  or (_17112_, _17110_, _17019_);
  and (_17113_, _17112_, _02173_);
  or (_17114_, _17113_, _02201_);
  or (_17115_, _17114_, _17109_);
  or (_17116_, _17029_, _02303_);
  and (_17117_, _17116_, _01887_);
  and (_17118_, _17117_, _17115_);
  and (_17119_, _17052_, _01860_);
  or (_17120_, _17119_, _01537_);
  or (_17121_, _17120_, _17118_);
  and (_17123_, _11072_, _03633_);
  or (_17124_, _17019_, _01538_);
  or (_17125_, _17124_, _17123_);
  and (_17126_, _17125_, _38087_);
  and (_17127_, _17126_, _17121_);
  or (_17128_, _17127_, _17018_);
  and (_40219_, _17128_, _37580_);
  and (_17129_, _38088_, \oc8051_golden_model_1.IE [3]);
  and (_17130_, _07586_, \oc8051_golden_model_1.IE [3]);
  and (_17131_, _11094_, _03633_);
  or (_17133_, _17131_, _17130_);
  and (_17134_, _17133_, _02167_);
  nor (_17135_, _07586_, _03268_);
  or (_17136_, _17135_, _17130_);
  or (_17137_, _17136_, _05249_);
  nor (_17138_, _11101_, _07586_);
  or (_17139_, _17138_, _17130_);
  or (_17140_, _17139_, _02814_);
  and (_17141_, _03633_, \oc8051_golden_model_1.ACC [3]);
  or (_17142_, _17141_, _17130_);
  and (_17144_, _17142_, _02817_);
  and (_17145_, _02818_, \oc8051_golden_model_1.IE [3]);
  or (_17146_, _17145_, _02001_);
  or (_17147_, _17146_, _17144_);
  and (_17148_, _17147_, _02024_);
  and (_17149_, _17148_, _17140_);
  and (_17150_, _07594_, \oc8051_golden_model_1.IE [3]);
  and (_17151_, _11098_, _04333_);
  or (_17152_, _17151_, _17150_);
  and (_17153_, _17152_, _02007_);
  or (_17155_, _17153_, _01999_);
  or (_17156_, _17155_, _17149_);
  or (_17157_, _17136_, _02840_);
  and (_17158_, _17157_, _17156_);
  or (_17159_, _17158_, _02006_);
  or (_17160_, _17142_, _02021_);
  and (_17161_, _17160_, _02025_);
  and (_17162_, _17161_, _17159_);
  and (_17163_, _11096_, _04333_);
  or (_17164_, _17163_, _17150_);
  and (_17166_, _17164_, _01997_);
  or (_17167_, _17166_, _01991_);
  or (_17168_, _17167_, _17162_);
  or (_17169_, _17150_, _11127_);
  and (_17170_, _17169_, _17152_);
  or (_17171_, _17170_, _02861_);
  and (_17172_, _17171_, _02408_);
  and (_17173_, _17172_, _17168_);
  nor (_17174_, _11145_, _07594_);
  or (_17175_, _17174_, _17150_);
  and (_17177_, _17175_, _01875_);
  or (_17178_, _17177_, _05994_);
  or (_17179_, _17178_, _17173_);
  and (_17180_, _17179_, _17137_);
  or (_17181_, _17180_, _02528_);
  and (_17182_, _04998_, _03633_);
  or (_17183_, _17130_, _02888_);
  or (_17184_, _17183_, _17182_);
  and (_17185_, _17184_, _02043_);
  and (_17186_, _17185_, _17181_);
  nor (_17188_, _11206_, _07586_);
  or (_17189_, _17188_, _17130_);
  and (_17190_, _17189_, _01602_);
  or (_17191_, _17190_, _01869_);
  or (_17192_, _17191_, _17186_);
  and (_17193_, _03633_, _04678_);
  or (_17194_, _17193_, _17130_);
  or (_17195_, _17194_, _01870_);
  and (_17196_, _17195_, _17192_);
  or (_17197_, _17196_, _02079_);
  and (_17199_, _11222_, _03633_);
  or (_17200_, _17130_, _02166_);
  or (_17201_, _17200_, _17199_);
  and (_17202_, _17201_, _02912_);
  and (_17203_, _17202_, _17197_);
  or (_17204_, _17203_, _17134_);
  and (_17205_, _17204_, _02176_);
  or (_17206_, _17130_, _04014_);
  and (_17207_, _17194_, _02072_);
  and (_17208_, _17207_, _17206_);
  or (_17210_, _17208_, _17205_);
  and (_17211_, _17210_, _02907_);
  and (_17212_, _17142_, _02177_);
  and (_17213_, _17212_, _17206_);
  or (_17214_, _17213_, _02071_);
  or (_17215_, _17214_, _17211_);
  nor (_17216_, _11220_, _07586_);
  or (_17217_, _17130_, _04788_);
  or (_17218_, _17217_, _17216_);
  and (_17219_, _17218_, _04793_);
  and (_17221_, _17219_, _17215_);
  nor (_17222_, _11093_, _07586_);
  or (_17223_, _17222_, _17130_);
  and (_17224_, _17223_, _02173_);
  or (_17225_, _17224_, _02201_);
  or (_17226_, _17225_, _17221_);
  or (_17227_, _17139_, _02303_);
  and (_17228_, _17227_, _01887_);
  and (_17229_, _17228_, _17226_);
  and (_17230_, _17164_, _01860_);
  or (_17232_, _17230_, _01537_);
  or (_17233_, _17232_, _17229_);
  and (_17234_, _11273_, _03633_);
  or (_17235_, _17130_, _01538_);
  or (_17236_, _17235_, _17234_);
  and (_17237_, _17236_, _38087_);
  and (_17238_, _17237_, _17233_);
  or (_17239_, _17238_, _17129_);
  and (_40220_, _17239_, _37580_);
  and (_17240_, _38088_, \oc8051_golden_model_1.IE [4]);
  and (_17242_, _07586_, \oc8051_golden_model_1.IE [4]);
  and (_17243_, _11431_, _03633_);
  or (_17244_, _17243_, _17242_);
  and (_17245_, _17244_, _02167_);
  nor (_17246_, _04211_, _07586_);
  or (_17247_, _17246_, _17242_);
  or (_17248_, _17247_, _05249_);
  and (_17249_, _07594_, \oc8051_golden_model_1.IE [4]);
  and (_17250_, _11301_, _04333_);
  or (_17251_, _17250_, _17249_);
  and (_17252_, _17251_, _01997_);
  nor (_17253_, _11317_, _07586_);
  or (_17254_, _17253_, _17242_);
  or (_17255_, _17254_, _02814_);
  and (_17256_, _03633_, \oc8051_golden_model_1.ACC [4]);
  or (_17257_, _17256_, _17242_);
  and (_17258_, _17257_, _02817_);
  and (_17259_, _02818_, \oc8051_golden_model_1.IE [4]);
  or (_17260_, _17259_, _02001_);
  or (_17261_, _17260_, _17258_);
  and (_17263_, _17261_, _02024_);
  and (_17264_, _17263_, _17255_);
  and (_17265_, _11303_, _04333_);
  or (_17266_, _17265_, _17249_);
  and (_17267_, _17266_, _02007_);
  or (_17268_, _17267_, _01999_);
  or (_17269_, _17268_, _17264_);
  or (_17270_, _17247_, _02840_);
  and (_17271_, _17270_, _17269_);
  or (_17272_, _17271_, _02006_);
  or (_17274_, _17257_, _02021_);
  and (_17275_, _17274_, _02025_);
  and (_17276_, _17275_, _17272_);
  or (_17277_, _17276_, _17252_);
  and (_17278_, _17277_, _02861_);
  or (_17279_, _17249_, _11334_);
  and (_17280_, _17279_, _01991_);
  and (_17281_, _17280_, _17266_);
  or (_17282_, _17281_, _17278_);
  and (_17283_, _17282_, _02408_);
  nor (_17285_, _11299_, _07594_);
  or (_17286_, _17285_, _17249_);
  and (_17287_, _17286_, _01875_);
  or (_17288_, _17287_, _05994_);
  or (_17289_, _17288_, _17283_);
  and (_17290_, _17289_, _17248_);
  or (_17291_, _17290_, _02528_);
  and (_17292_, _05135_, _03633_);
  or (_17293_, _17242_, _02888_);
  or (_17294_, _17293_, _17292_);
  and (_17296_, _17294_, _02043_);
  and (_17297_, _17296_, _17291_);
  nor (_17298_, _11411_, _07586_);
  or (_17299_, _17298_, _17242_);
  and (_17300_, _17299_, _01602_);
  or (_17301_, _17300_, _01869_);
  or (_17302_, _17301_, _17297_);
  and (_17303_, _04694_, _03633_);
  or (_17304_, _17303_, _17242_);
  or (_17305_, _17304_, _01870_);
  and (_17307_, _17305_, _17302_);
  or (_17308_, _17307_, _02079_);
  and (_17309_, _11425_, _03633_);
  or (_17310_, _17242_, _02166_);
  or (_17311_, _17310_, _17309_);
  and (_17312_, _17311_, _02912_);
  and (_17313_, _17312_, _17308_);
  or (_17314_, _17313_, _17245_);
  and (_17315_, _17314_, _02176_);
  or (_17316_, _17242_, _04258_);
  and (_17318_, _17304_, _02072_);
  and (_17319_, _17318_, _17316_);
  or (_17320_, _17319_, _17315_);
  and (_17321_, _17320_, _02907_);
  and (_17322_, _17257_, _02177_);
  and (_17323_, _17322_, _17316_);
  or (_17324_, _17323_, _02071_);
  or (_17325_, _17324_, _17321_);
  nor (_17326_, _11424_, _07586_);
  or (_17327_, _17242_, _04788_);
  or (_17329_, _17327_, _17326_);
  and (_17330_, _17329_, _04793_);
  and (_17331_, _17330_, _17325_);
  nor (_17332_, _11430_, _07586_);
  or (_17333_, _17332_, _17242_);
  and (_17334_, _17333_, _02173_);
  or (_17335_, _17334_, _02201_);
  or (_17336_, _17335_, _17331_);
  or (_17337_, _17254_, _02303_);
  and (_17338_, _17337_, _01887_);
  and (_17340_, _17338_, _17336_);
  and (_17341_, _17251_, _01860_);
  or (_17342_, _17341_, _01537_);
  or (_17343_, _17342_, _17340_);
  and (_17344_, _11487_, _03633_);
  or (_17345_, _17242_, _01538_);
  or (_17346_, _17345_, _17344_);
  and (_17347_, _17346_, _38087_);
  and (_17348_, _17347_, _17343_);
  or (_17349_, _17348_, _17240_);
  and (_40222_, _17349_, _37580_);
  and (_17351_, _38088_, \oc8051_golden_model_1.IE [5]);
  and (_17352_, _07586_, \oc8051_golden_model_1.IE [5]);
  and (_17353_, _11635_, _03633_);
  or (_17354_, _17353_, _17352_);
  and (_17355_, _17354_, _02167_);
  nor (_17356_, _11525_, _07586_);
  or (_17357_, _17356_, _17352_);
  or (_17358_, _17357_, _02814_);
  and (_17359_, _03633_, \oc8051_golden_model_1.ACC [5]);
  or (_17361_, _17359_, _17352_);
  and (_17362_, _17361_, _02817_);
  and (_17363_, _02818_, \oc8051_golden_model_1.IE [5]);
  or (_17364_, _17363_, _02001_);
  or (_17365_, _17364_, _17362_);
  and (_17366_, _17365_, _02024_);
  and (_17367_, _17366_, _17358_);
  and (_17368_, _07594_, \oc8051_golden_model_1.IE [5]);
  and (_17369_, _11510_, _04333_);
  or (_17370_, _17369_, _17368_);
  and (_17372_, _17370_, _02007_);
  or (_17373_, _17372_, _01999_);
  or (_17374_, _17373_, _17367_);
  nor (_17375_, _03916_, _07586_);
  or (_17376_, _17375_, _17352_);
  or (_17377_, _17376_, _02840_);
  and (_17378_, _17377_, _17374_);
  or (_17379_, _17378_, _02006_);
  or (_17380_, _17361_, _02021_);
  and (_17381_, _17380_, _02025_);
  and (_17383_, _17381_, _17379_);
  and (_17384_, _11508_, _04333_);
  or (_17385_, _17384_, _17368_);
  and (_17386_, _17385_, _01997_);
  or (_17387_, _17386_, _01991_);
  or (_17388_, _17387_, _17383_);
  or (_17389_, _17368_, _11542_);
  and (_17390_, _17389_, _17370_);
  or (_17391_, _17390_, _02861_);
  and (_17392_, _17391_, _02408_);
  and (_17393_, _17392_, _17388_);
  nor (_17394_, _11506_, _07594_);
  or (_17395_, _17394_, _17368_);
  and (_17396_, _17395_, _01875_);
  or (_17397_, _17396_, _05994_);
  or (_17398_, _17397_, _17393_);
  or (_17399_, _17376_, _05249_);
  and (_17400_, _17399_, _17398_);
  or (_17401_, _17400_, _02528_);
  and (_17402_, _05090_, _03633_);
  or (_17404_, _17352_, _02888_);
  or (_17405_, _17404_, _17402_);
  and (_17406_, _17405_, _02043_);
  and (_17407_, _17406_, _17401_);
  nor (_17408_, _11615_, _07586_);
  or (_17409_, _17408_, _17352_);
  and (_17410_, _17409_, _01602_);
  or (_17411_, _17410_, _01869_);
  or (_17412_, _17411_, _17407_);
  and (_17413_, _04672_, _03633_);
  or (_17415_, _17413_, _17352_);
  or (_17416_, _17415_, _01870_);
  and (_17417_, _17416_, _17412_);
  or (_17418_, _17417_, _02079_);
  and (_17419_, _11629_, _03633_);
  or (_17420_, _17352_, _02166_);
  or (_17421_, _17420_, _17419_);
  and (_17422_, _17421_, _02912_);
  and (_17423_, _17422_, _17418_);
  or (_17424_, _17423_, _17355_);
  and (_17426_, _17424_, _02176_);
  or (_17427_, _17352_, _03965_);
  and (_17428_, _17415_, _02072_);
  and (_17429_, _17428_, _17427_);
  or (_17430_, _17429_, _17426_);
  and (_17431_, _17430_, _02907_);
  and (_17432_, _17361_, _02177_);
  and (_17433_, _17432_, _17427_);
  or (_17434_, _17433_, _02071_);
  or (_17435_, _17434_, _17431_);
  nor (_17437_, _11628_, _07586_);
  or (_17438_, _17352_, _04788_);
  or (_17439_, _17438_, _17437_);
  and (_17440_, _17439_, _04793_);
  and (_17441_, _17440_, _17435_);
  nor (_17442_, _11634_, _07586_);
  or (_17443_, _17442_, _17352_);
  and (_17444_, _17443_, _02173_);
  or (_17445_, _17444_, _02201_);
  or (_17446_, _17445_, _17441_);
  or (_17448_, _17357_, _02303_);
  and (_17449_, _17448_, _01887_);
  and (_17450_, _17449_, _17446_);
  and (_17451_, _17385_, _01860_);
  or (_17452_, _17451_, _01537_);
  or (_17453_, _17452_, _17450_);
  and (_17454_, _11685_, _03633_);
  or (_17455_, _17352_, _01538_);
  or (_17456_, _17455_, _17454_);
  and (_17457_, _17456_, _38087_);
  and (_17458_, _17457_, _17453_);
  or (_17459_, _17458_, _17351_);
  and (_40223_, _17459_, _37580_);
  and (_17460_, _38088_, \oc8051_golden_model_1.IE [6]);
  and (_17461_, _07586_, \oc8051_golden_model_1.IE [6]);
  and (_17462_, _11709_, _03633_);
  or (_17463_, _17462_, _17461_);
  and (_17464_, _17463_, _02167_);
  nor (_17465_, _11730_, _07586_);
  or (_17466_, _17465_, _17461_);
  or (_17469_, _17466_, _02814_);
  and (_17470_, _03633_, \oc8051_golden_model_1.ACC [6]);
  or (_17471_, _17470_, _17461_);
  and (_17472_, _17471_, _02817_);
  and (_17473_, _02818_, \oc8051_golden_model_1.IE [6]);
  or (_17474_, _17473_, _02001_);
  or (_17475_, _17474_, _17472_);
  and (_17476_, _17475_, _02024_);
  and (_17477_, _17476_, _17469_);
  and (_17478_, _07594_, \oc8051_golden_model_1.IE [6]);
  and (_17480_, _11717_, _04333_);
  or (_17481_, _17480_, _17478_);
  and (_17482_, _17481_, _02007_);
  or (_17483_, _17482_, _01999_);
  or (_17484_, _17483_, _17477_);
  nor (_17485_, _03808_, _07586_);
  or (_17486_, _17485_, _17461_);
  or (_17487_, _17486_, _02840_);
  and (_17488_, _17487_, _17484_);
  or (_17489_, _17488_, _02006_);
  or (_17491_, _17471_, _02021_);
  and (_17492_, _17491_, _02025_);
  and (_17493_, _17492_, _17489_);
  and (_17494_, _11715_, _04333_);
  or (_17495_, _17494_, _17478_);
  and (_17496_, _17495_, _01997_);
  or (_17497_, _17496_, _01991_);
  or (_17498_, _17497_, _17493_);
  or (_17499_, _17478_, _11747_);
  and (_17500_, _17499_, _17481_);
  or (_17502_, _17500_, _02861_);
  and (_17503_, _17502_, _02408_);
  and (_17504_, _17503_, _17498_);
  nor (_17505_, _11713_, _07594_);
  or (_17506_, _17505_, _17478_);
  and (_17507_, _17506_, _01875_);
  or (_17508_, _17507_, _05994_);
  or (_17509_, _17508_, _17504_);
  or (_17510_, _17486_, _05249_);
  and (_17511_, _17510_, _17509_);
  or (_17513_, _17511_, _02528_);
  and (_17514_, _04861_, _03633_);
  or (_17515_, _17461_, _02888_);
  or (_17516_, _17515_, _17514_);
  and (_17517_, _17516_, _02043_);
  and (_17518_, _17517_, _17513_);
  nor (_17519_, _11820_, _07586_);
  or (_17520_, _17519_, _17461_);
  and (_17521_, _17520_, _01602_);
  or (_17522_, _17521_, _01869_);
  or (_17524_, _17522_, _17518_);
  and (_17525_, _09920_, _03633_);
  or (_17526_, _17525_, _17461_);
  or (_17527_, _17526_, _01870_);
  and (_17528_, _17527_, _17524_);
  or (_17529_, _17528_, _02079_);
  and (_17530_, _11835_, _03633_);
  or (_17531_, _17461_, _02166_);
  or (_17532_, _17531_, _17530_);
  and (_17533_, _17532_, _02912_);
  and (_17535_, _17533_, _17529_);
  or (_17536_, _17535_, _17464_);
  and (_17537_, _17536_, _02176_);
  or (_17538_, _17461_, _03863_);
  and (_17539_, _17526_, _02072_);
  and (_17540_, _17539_, _17538_);
  or (_17541_, _17540_, _17537_);
  and (_17542_, _17541_, _02907_);
  and (_17543_, _17471_, _02177_);
  and (_17544_, _17543_, _17538_);
  or (_17546_, _17544_, _02071_);
  or (_17547_, _17546_, _17542_);
  nor (_17548_, _11833_, _07586_);
  or (_17549_, _17461_, _04788_);
  or (_17550_, _17549_, _17548_);
  and (_17551_, _17550_, _04793_);
  and (_17552_, _17551_, _17547_);
  nor (_17553_, _11708_, _07586_);
  or (_17554_, _17553_, _17461_);
  and (_17555_, _17554_, _02173_);
  or (_17557_, _17555_, _02201_);
  or (_17558_, _17557_, _17552_);
  or (_17559_, _17466_, _02303_);
  and (_17560_, _17559_, _01887_);
  and (_17561_, _17560_, _17558_);
  and (_17562_, _17495_, _01860_);
  or (_17563_, _17562_, _01537_);
  or (_17564_, _17563_, _17561_);
  and (_17565_, _11887_, _03633_);
  or (_17566_, _17461_, _01538_);
  or (_17568_, _17566_, _17565_);
  and (_17569_, _17568_, _38087_);
  and (_17570_, _17569_, _17564_);
  or (_17571_, _17570_, _17460_);
  and (_40224_, _17571_, _37580_);
  and (_17572_, _38088_, \oc8051_golden_model_1.IP [0]);
  nor (_17573_, _04106_, _07689_);
  and (_17574_, _07689_, \oc8051_golden_model_1.IP [0]);
  and (_17575_, _03670_, _04562_);
  or (_17576_, _17575_, _17574_);
  nand (_17578_, _17576_, _02072_);
  nor (_17579_, _17578_, _17573_);
  and (_17580_, _10620_, _03670_);
  or (_17581_, _17580_, _17574_);
  and (_17582_, _17581_, _02167_);
  and (_17583_, _03670_, _03028_);
  or (_17584_, _17583_, _17574_);
  or (_17585_, _17584_, _05249_);
  or (_17586_, _17574_, _17573_);
  and (_17587_, _17586_, _02001_);
  and (_17588_, _02818_, \oc8051_golden_model_1.IP [0]);
  and (_17589_, _03670_, \oc8051_golden_model_1.ACC [0]);
  or (_17590_, _17589_, _17574_);
  and (_17591_, _17590_, _02817_);
  or (_17592_, _17591_, _17588_);
  and (_17593_, _17592_, _02814_);
  or (_17594_, _17593_, _02007_);
  or (_17595_, _17594_, _17587_);
  and (_17596_, _10510_, _04324_);
  and (_17597_, _07697_, \oc8051_golden_model_1.IP [0]);
  or (_17599_, _17597_, _02024_);
  or (_17600_, _17599_, _17596_);
  and (_17601_, _17600_, _02840_);
  and (_17602_, _17601_, _17595_);
  and (_17603_, _17584_, _01999_);
  or (_17604_, _17603_, _02006_);
  or (_17605_, _17604_, _17602_);
  or (_17606_, _17590_, _02021_);
  and (_17607_, _17606_, _02025_);
  and (_17608_, _17607_, _17605_);
  and (_17610_, _17574_, _01997_);
  or (_17611_, _17610_, _01991_);
  or (_17612_, _17611_, _17608_);
  or (_17613_, _17586_, _02861_);
  and (_17614_, _17613_, _02408_);
  and (_17615_, _17614_, _17612_);
  nor (_17616_, _10542_, _07697_);
  or (_17617_, _17616_, _17597_);
  and (_17618_, _17617_, _01875_);
  or (_17619_, _17618_, _05994_);
  or (_17621_, _17619_, _17615_);
  and (_17622_, _17621_, _17585_);
  or (_17623_, _17622_, _02528_);
  and (_17624_, _04952_, _03670_);
  or (_17625_, _17574_, _02888_);
  or (_17626_, _17625_, _17624_);
  and (_17627_, _17626_, _17623_);
  or (_17628_, _17627_, _01602_);
  nor (_17629_, _10600_, _07689_);
  or (_17630_, _17574_, _02043_);
  or (_17632_, _17630_, _17629_);
  and (_17633_, _17632_, _01870_);
  and (_17634_, _17633_, _17628_);
  and (_17635_, _17576_, _01869_);
  or (_17636_, _17635_, _02079_);
  or (_17637_, _17636_, _17634_);
  and (_17638_, _10614_, _03670_);
  or (_17639_, _17574_, _02166_);
  or (_17640_, _17639_, _17638_);
  and (_17641_, _17640_, _02912_);
  and (_17643_, _17641_, _17637_);
  or (_17644_, _17643_, _17582_);
  and (_17645_, _17644_, _02176_);
  or (_17646_, _17645_, _17579_);
  and (_17647_, _17646_, _02907_);
  or (_17648_, _17574_, _04106_);
  and (_17649_, _17590_, _02177_);
  and (_17650_, _17649_, _17648_);
  or (_17651_, _17650_, _02071_);
  or (_17652_, _17651_, _17647_);
  nor (_17654_, _10613_, _07689_);
  or (_17655_, _17574_, _04788_);
  or (_17656_, _17655_, _17654_);
  and (_17657_, _17656_, _04793_);
  and (_17658_, _17657_, _17652_);
  nor (_17659_, _10619_, _07689_);
  or (_17660_, _17659_, _17574_);
  and (_17661_, _17660_, _02173_);
  or (_17662_, _17661_, _02201_);
  or (_17663_, _17662_, _17658_);
  or (_17665_, _17586_, _02303_);
  and (_17666_, _17665_, _01887_);
  and (_17667_, _17666_, _17663_);
  and (_17668_, _17574_, _01860_);
  or (_17669_, _17668_, _01537_);
  or (_17670_, _17669_, _17667_);
  or (_17671_, _17586_, _01538_);
  and (_17672_, _17671_, _38087_);
  and (_17673_, _17672_, _17670_);
  or (_17674_, _17673_, _17572_);
  and (_40225_, _17674_, _37580_);
  and (_17676_, _38088_, \oc8051_golden_model_1.IP [1]);
  and (_17677_, _07689_, \oc8051_golden_model_1.IP [1]);
  nor (_17678_, _07689_, _02811_);
  or (_17679_, _17678_, _17677_);
  or (_17680_, _17679_, _02840_);
  or (_17681_, _03670_, \oc8051_golden_model_1.IP [1]);
  and (_17682_, _10698_, _03670_);
  not (_17683_, _17682_);
  and (_17684_, _17683_, _17681_);
  or (_17686_, _17684_, _02814_);
  nand (_17687_, _03670_, _01613_);
  and (_17688_, _17687_, _17681_);
  and (_17689_, _17688_, _02817_);
  and (_17690_, _02818_, \oc8051_golden_model_1.IP [1]);
  or (_17691_, _17690_, _02001_);
  or (_17692_, _17691_, _17689_);
  and (_17693_, _17692_, _02024_);
  and (_17694_, _17693_, _17686_);
  and (_17695_, _07697_, \oc8051_golden_model_1.IP [1]);
  and (_17697_, _10710_, _04324_);
  or (_17698_, _17697_, _17695_);
  and (_17699_, _17698_, _02007_);
  or (_17700_, _17699_, _01999_);
  or (_17701_, _17700_, _17694_);
  and (_17702_, _17701_, _17680_);
  or (_17703_, _17702_, _02006_);
  or (_17704_, _17688_, _02021_);
  and (_17705_, _17704_, _02025_);
  and (_17706_, _17705_, _17703_);
  and (_17708_, _10696_, _04324_);
  or (_17709_, _17708_, _17695_);
  and (_17710_, _17709_, _01997_);
  or (_17711_, _17710_, _01991_);
  or (_17712_, _17711_, _17706_);
  and (_17713_, _17697_, _10725_);
  or (_17714_, _17695_, _02861_);
  or (_17715_, _17714_, _17713_);
  and (_17716_, _17715_, _17712_);
  and (_17717_, _17716_, _02408_);
  nor (_17719_, _10742_, _07697_);
  or (_17720_, _17695_, _17719_);
  and (_17721_, _17720_, _01875_);
  or (_17722_, _17721_, _05994_);
  or (_17723_, _17722_, _17717_);
  or (_17724_, _17679_, _05249_);
  and (_17725_, _17724_, _17723_);
  or (_17726_, _17725_, _02528_);
  and (_17727_, _04907_, _03670_);
  or (_17728_, _17677_, _02888_);
  or (_17730_, _17728_, _17727_);
  and (_17731_, _17730_, _02043_);
  and (_17732_, _17731_, _17726_);
  nor (_17733_, _10802_, _07689_);
  or (_17734_, _17733_, _17677_);
  and (_17735_, _17734_, _01602_);
  or (_17736_, _17735_, _17732_);
  and (_17737_, _17736_, _01870_);
  nand (_17738_, _03670_, _02687_);
  and (_17739_, _17681_, _01869_);
  and (_17741_, _17739_, _17738_);
  or (_17742_, _17741_, _17737_);
  and (_17743_, _17742_, _02166_);
  or (_17744_, _10816_, _07689_);
  and (_17745_, _17681_, _02079_);
  and (_17746_, _17745_, _17744_);
  or (_17747_, _17746_, _17743_);
  and (_17748_, _17747_, _02912_);
  or (_17749_, _10822_, _07689_);
  and (_17750_, _17681_, _02167_);
  and (_17752_, _17750_, _17749_);
  or (_17753_, _17752_, _17748_);
  and (_17754_, _17753_, _02176_);
  or (_17755_, _10692_, _07689_);
  and (_17756_, _17681_, _02072_);
  and (_17757_, _17756_, _17755_);
  or (_17758_, _17757_, _17754_);
  and (_17759_, _17758_, _02907_);
  or (_17760_, _17677_, _04058_);
  and (_17761_, _17688_, _02177_);
  and (_17763_, _17761_, _17760_);
  or (_17764_, _17763_, _17759_);
  and (_17765_, _17764_, _02174_);
  or (_17766_, _17687_, _04058_);
  and (_17767_, _17681_, _02173_);
  and (_17768_, _17767_, _17766_);
  or (_17769_, _17768_, _02201_);
  or (_17770_, _17738_, _04058_);
  and (_17771_, _17681_, _02071_);
  and (_17772_, _17771_, _17770_);
  or (_17774_, _17772_, _17769_);
  or (_17775_, _17774_, _17765_);
  or (_17776_, _17684_, _02303_);
  and (_17777_, _17776_, _01887_);
  and (_17778_, _17777_, _17775_);
  and (_17779_, _17709_, _01860_);
  or (_17780_, _17779_, _01537_);
  or (_17781_, _17780_, _17778_);
  or (_17782_, _17677_, _01538_);
  or (_17783_, _17782_, _17682_);
  and (_17784_, _17783_, _38087_);
  and (_17785_, _17784_, _17781_);
  or (_17786_, _17785_, _17676_);
  and (_40226_, _17786_, _37580_);
  and (_17787_, _38088_, \oc8051_golden_model_1.IP [2]);
  and (_17788_, _07689_, \oc8051_golden_model_1.IP [2]);
  and (_17789_, _11020_, _03670_);
  or (_17790_, _17789_, _17788_);
  and (_17791_, _17790_, _02167_);
  nor (_17792_, _07689_, _03455_);
  or (_17794_, _17792_, _17788_);
  or (_17795_, _17794_, _05249_);
  and (_17796_, _17794_, _01999_);
  and (_17797_, _07697_, \oc8051_golden_model_1.IP [2]);
  and (_17798_, _10909_, _04324_);
  or (_17799_, _17798_, _17797_);
  or (_17800_, _17799_, _02024_);
  nor (_17801_, _10905_, _07689_);
  or (_17802_, _17801_, _17788_);
  and (_17803_, _17802_, _02001_);
  and (_17805_, _02818_, \oc8051_golden_model_1.IP [2]);
  and (_17806_, _03670_, \oc8051_golden_model_1.ACC [2]);
  or (_17807_, _17806_, _17788_);
  and (_17808_, _17807_, _02817_);
  or (_17809_, _17808_, _17805_);
  and (_17810_, _17809_, _02814_);
  or (_17811_, _17810_, _02007_);
  or (_17812_, _17811_, _17803_);
  and (_17813_, _17812_, _17800_);
  and (_17814_, _17813_, _02840_);
  or (_17816_, _17814_, _17796_);
  or (_17817_, _17816_, _02006_);
  or (_17818_, _17807_, _02021_);
  and (_17819_, _17818_, _02025_);
  and (_17820_, _17819_, _17817_);
  and (_17821_, _10894_, _04324_);
  or (_17822_, _17821_, _17797_);
  and (_17823_, _17822_, _01997_);
  or (_17824_, _17823_, _01991_);
  or (_17825_, _17824_, _17820_);
  or (_17827_, _17797_, _10924_);
  and (_17828_, _17827_, _17799_);
  or (_17829_, _17828_, _02861_);
  and (_17830_, _17829_, _02408_);
  and (_17831_, _17830_, _17825_);
  nor (_17832_, _10942_, _07697_);
  or (_17833_, _17832_, _17797_);
  and (_17834_, _17833_, _01875_);
  or (_17835_, _17834_, _05994_);
  or (_17836_, _17835_, _17831_);
  and (_17838_, _17836_, _17795_);
  or (_17839_, _17838_, _02528_);
  and (_17840_, _05043_, _03670_);
  or (_17841_, _17788_, _02888_);
  or (_17842_, _17841_, _17840_);
  and (_17843_, _17842_, _02043_);
  and (_17844_, _17843_, _17839_);
  nor (_17845_, _11000_, _07689_);
  or (_17846_, _17845_, _17788_);
  and (_17847_, _17846_, _01602_);
  or (_17849_, _17847_, _01869_);
  or (_17850_, _17849_, _17844_);
  and (_17851_, _03670_, _04724_);
  or (_17852_, _17851_, _17788_);
  or (_17853_, _17852_, _01870_);
  and (_17854_, _17853_, _17850_);
  or (_17855_, _17854_, _02079_);
  and (_17856_, _11014_, _03670_);
  or (_17857_, _17788_, _02166_);
  or (_17858_, _17857_, _17856_);
  and (_17860_, _17858_, _02912_);
  and (_17861_, _17860_, _17855_);
  or (_17862_, _17861_, _17791_);
  and (_17863_, _17862_, _02176_);
  or (_17864_, _17788_, _04156_);
  and (_17865_, _17852_, _02072_);
  and (_17866_, _17865_, _17864_);
  or (_17867_, _17866_, _17863_);
  and (_17868_, _17867_, _02907_);
  and (_17869_, _17807_, _02177_);
  and (_17871_, _17869_, _17864_);
  or (_17872_, _17871_, _02071_);
  or (_17873_, _17872_, _17868_);
  nor (_17874_, _11013_, _07689_);
  or (_17875_, _17788_, _04788_);
  or (_17876_, _17875_, _17874_);
  and (_17877_, _17876_, _04793_);
  and (_17878_, _17877_, _17873_);
  nor (_17879_, _11019_, _07689_);
  or (_17880_, _17879_, _17788_);
  and (_17881_, _17880_, _02173_);
  or (_17882_, _17881_, _02201_);
  or (_17883_, _17882_, _17878_);
  or (_17884_, _17802_, _02303_);
  and (_17885_, _17884_, _01887_);
  and (_17886_, _17885_, _17883_);
  and (_17887_, _17822_, _01860_);
  or (_17888_, _17887_, _01537_);
  or (_17889_, _17888_, _17886_);
  and (_17890_, _11072_, _03670_);
  or (_17893_, _17788_, _01538_);
  or (_17894_, _17893_, _17890_);
  and (_17895_, _17894_, _38087_);
  and (_17896_, _17895_, _17889_);
  or (_17897_, _17896_, _17787_);
  and (_40227_, _17897_, _37580_);
  and (_17898_, _38088_, \oc8051_golden_model_1.IP [3]);
  and (_17899_, _07689_, \oc8051_golden_model_1.IP [3]);
  and (_17900_, _11094_, _03670_);
  or (_17901_, _17900_, _17899_);
  and (_17903_, _17901_, _02167_);
  nor (_17904_, _07689_, _03268_);
  or (_17905_, _17904_, _17899_);
  or (_17906_, _17905_, _05249_);
  nor (_17907_, _11101_, _07689_);
  or (_17908_, _17907_, _17899_);
  or (_17909_, _17908_, _02814_);
  and (_17910_, _03670_, \oc8051_golden_model_1.ACC [3]);
  or (_17911_, _17910_, _17899_);
  and (_17912_, _17911_, _02817_);
  and (_17914_, _02818_, \oc8051_golden_model_1.IP [3]);
  or (_17915_, _17914_, _02001_);
  or (_17916_, _17915_, _17912_);
  and (_17917_, _17916_, _02024_);
  and (_17918_, _17917_, _17909_);
  and (_17919_, _07697_, \oc8051_golden_model_1.IP [3]);
  and (_17920_, _11098_, _04324_);
  or (_17921_, _17920_, _17919_);
  and (_17922_, _17921_, _02007_);
  or (_17923_, _17922_, _01999_);
  or (_17925_, _17923_, _17918_);
  or (_17926_, _17905_, _02840_);
  and (_17927_, _17926_, _17925_);
  or (_17928_, _17927_, _02006_);
  or (_17929_, _17911_, _02021_);
  and (_17930_, _17929_, _02025_);
  and (_17931_, _17930_, _17928_);
  and (_17932_, _11096_, _04324_);
  or (_17933_, _17932_, _17919_);
  and (_17934_, _17933_, _01997_);
  or (_17936_, _17934_, _01991_);
  or (_17937_, _17936_, _17931_);
  or (_17938_, _17919_, _11127_);
  and (_17939_, _17938_, _17921_);
  or (_17940_, _17939_, _02861_);
  and (_17941_, _17940_, _02408_);
  and (_17942_, _17941_, _17937_);
  nor (_17943_, _11145_, _07697_);
  or (_17944_, _17943_, _17919_);
  and (_17945_, _17944_, _01875_);
  or (_17947_, _17945_, _05994_);
  or (_17948_, _17947_, _17942_);
  and (_17949_, _17948_, _17906_);
  or (_17950_, _17949_, _02528_);
  and (_17951_, _04998_, _03670_);
  or (_17952_, _17899_, _02888_);
  or (_17953_, _17952_, _17951_);
  and (_17954_, _17953_, _02043_);
  and (_17955_, _17954_, _17950_);
  nor (_17956_, _11206_, _07689_);
  or (_17957_, _17956_, _17899_);
  and (_17958_, _17957_, _01602_);
  or (_17959_, _17958_, _01869_);
  or (_17960_, _17959_, _17955_);
  and (_17961_, _03670_, _04678_);
  or (_17962_, _17961_, _17899_);
  or (_17963_, _17962_, _01870_);
  and (_17964_, _17963_, _17960_);
  or (_17965_, _17964_, _02079_);
  and (_17966_, _11222_, _03670_);
  or (_17968_, _17899_, _02166_);
  or (_17969_, _17968_, _17966_);
  and (_17970_, _17969_, _02912_);
  and (_17971_, _17970_, _17965_);
  or (_17972_, _17971_, _17903_);
  and (_17973_, _17972_, _02176_);
  or (_17974_, _17899_, _04014_);
  and (_17975_, _17962_, _02072_);
  and (_17976_, _17975_, _17974_);
  or (_17977_, _17976_, _17973_);
  and (_17979_, _17977_, _02907_);
  and (_17980_, _17911_, _02177_);
  and (_17981_, _17980_, _17974_);
  or (_17982_, _17981_, _02071_);
  or (_17983_, _17982_, _17979_);
  nor (_17984_, _11220_, _07689_);
  or (_17985_, _17899_, _04788_);
  or (_17986_, _17985_, _17984_);
  and (_17987_, _17986_, _04793_);
  and (_17988_, _17987_, _17983_);
  nor (_17990_, _11093_, _07689_);
  or (_17991_, _17990_, _17899_);
  and (_17992_, _17991_, _02173_);
  or (_17993_, _17992_, _02201_);
  or (_17994_, _17993_, _17988_);
  or (_17995_, _17908_, _02303_);
  and (_17996_, _17995_, _01887_);
  and (_17997_, _17996_, _17994_);
  and (_17998_, _17933_, _01860_);
  or (_17999_, _17998_, _01537_);
  or (_18001_, _17999_, _17997_);
  and (_18002_, _11273_, _03670_);
  or (_18003_, _17899_, _01538_);
  or (_18004_, _18003_, _18002_);
  and (_18005_, _18004_, _38087_);
  and (_18006_, _18005_, _18001_);
  or (_18007_, _18006_, _17898_);
  and (_40228_, _18007_, _37580_);
  and (_18008_, _38088_, \oc8051_golden_model_1.IP [4]);
  and (_18009_, _07689_, \oc8051_golden_model_1.IP [4]);
  and (_18011_, _11431_, _03670_);
  or (_18012_, _18011_, _18009_);
  and (_18013_, _18012_, _02167_);
  nor (_18014_, _04211_, _07689_);
  or (_18015_, _18014_, _18009_);
  or (_18016_, _18015_, _05249_);
  and (_18017_, _07697_, \oc8051_golden_model_1.IP [4]);
  and (_18018_, _11301_, _04324_);
  or (_18019_, _18018_, _18017_);
  and (_18020_, _18019_, _01997_);
  nor (_18022_, _11317_, _07689_);
  or (_18023_, _18022_, _18009_);
  or (_18024_, _18023_, _02814_);
  and (_18025_, _03670_, \oc8051_golden_model_1.ACC [4]);
  or (_18026_, _18025_, _18009_);
  and (_18027_, _18026_, _02817_);
  and (_18028_, _02818_, \oc8051_golden_model_1.IP [4]);
  or (_18029_, _18028_, _02001_);
  or (_18030_, _18029_, _18027_);
  and (_18031_, _18030_, _02024_);
  and (_18033_, _18031_, _18024_);
  and (_18034_, _11303_, _04324_);
  or (_18035_, _18034_, _18017_);
  and (_18036_, _18035_, _02007_);
  or (_18037_, _18036_, _01999_);
  or (_18038_, _18037_, _18033_);
  or (_18039_, _18015_, _02840_);
  and (_18040_, _18039_, _18038_);
  or (_18041_, _18040_, _02006_);
  or (_18042_, _18026_, _02021_);
  and (_18044_, _18042_, _02025_);
  and (_18045_, _18044_, _18041_);
  or (_18046_, _18045_, _18020_);
  and (_18047_, _18046_, _02861_);
  and (_18048_, _11335_, _04324_);
  or (_18049_, _18048_, _18017_);
  and (_18050_, _18049_, _01991_);
  or (_18051_, _18050_, _18047_);
  and (_18052_, _18051_, _02408_);
  nor (_18053_, _11299_, _07697_);
  or (_18055_, _18053_, _18017_);
  and (_18056_, _18055_, _01875_);
  or (_18057_, _18056_, _05994_);
  or (_18058_, _18057_, _18052_);
  and (_18059_, _18058_, _18016_);
  or (_18060_, _18059_, _02528_);
  and (_18061_, _05135_, _03670_);
  or (_18062_, _18009_, _02888_);
  or (_18063_, _18062_, _18061_);
  and (_18064_, _18063_, _02043_);
  and (_18066_, _18064_, _18060_);
  nor (_18067_, _11411_, _07689_);
  or (_18068_, _18067_, _18009_);
  and (_18069_, _18068_, _01602_);
  or (_18070_, _18069_, _01869_);
  or (_18071_, _18070_, _18066_);
  and (_18072_, _04694_, _03670_);
  or (_18073_, _18072_, _18009_);
  or (_18074_, _18073_, _01870_);
  and (_18075_, _18074_, _18071_);
  or (_18077_, _18075_, _02079_);
  and (_18078_, _11425_, _03670_);
  or (_18079_, _18009_, _02166_);
  or (_18080_, _18079_, _18078_);
  and (_18081_, _18080_, _02912_);
  and (_18082_, _18081_, _18077_);
  or (_18083_, _18082_, _18013_);
  and (_18084_, _18083_, _02176_);
  or (_18085_, _18009_, _04258_);
  and (_18086_, _18073_, _02072_);
  and (_18088_, _18086_, _18085_);
  or (_18089_, _18088_, _18084_);
  and (_18090_, _18089_, _02907_);
  and (_18091_, _18026_, _02177_);
  and (_18092_, _18091_, _18085_);
  or (_18093_, _18092_, _02071_);
  or (_18094_, _18093_, _18090_);
  nor (_18095_, _11424_, _07689_);
  or (_18096_, _18009_, _04788_);
  or (_18097_, _18096_, _18095_);
  and (_18099_, _18097_, _04793_);
  and (_18100_, _18099_, _18094_);
  nor (_18101_, _11430_, _07689_);
  or (_18102_, _18101_, _18009_);
  and (_18103_, _18102_, _02173_);
  or (_18104_, _18103_, _02201_);
  or (_18105_, _18104_, _18100_);
  or (_18106_, _18023_, _02303_);
  and (_18107_, _18106_, _01887_);
  and (_18108_, _18107_, _18105_);
  and (_18110_, _18019_, _01860_);
  or (_18111_, _18110_, _01537_);
  or (_18112_, _18111_, _18108_);
  and (_18113_, _11487_, _03670_);
  or (_18114_, _18009_, _01538_);
  or (_18115_, _18114_, _18113_);
  and (_18116_, _18115_, _38087_);
  and (_18117_, _18116_, _18112_);
  or (_18118_, _18117_, _18008_);
  and (_40229_, _18118_, _37580_);
  and (_18120_, _38088_, \oc8051_golden_model_1.IP [5]);
  and (_18121_, _07689_, \oc8051_golden_model_1.IP [5]);
  and (_18122_, _11635_, _03670_);
  or (_18123_, _18122_, _18121_);
  and (_18124_, _18123_, _02167_);
  nor (_18125_, _11525_, _07689_);
  or (_18126_, _18125_, _18121_);
  or (_18127_, _18126_, _02814_);
  and (_18128_, _03670_, \oc8051_golden_model_1.ACC [5]);
  or (_18129_, _18128_, _18121_);
  and (_18130_, _18129_, _02817_);
  and (_18131_, _02818_, \oc8051_golden_model_1.IP [5]);
  or (_18132_, _18131_, _02001_);
  or (_18133_, _18132_, _18130_);
  and (_18134_, _18133_, _02024_);
  and (_18135_, _18134_, _18127_);
  and (_18136_, _07697_, \oc8051_golden_model_1.IP [5]);
  and (_18137_, _11510_, _04324_);
  or (_18138_, _18137_, _18136_);
  and (_18139_, _18138_, _02007_);
  or (_18141_, _18139_, _01999_);
  or (_18142_, _18141_, _18135_);
  nor (_18143_, _03916_, _07689_);
  or (_18144_, _18143_, _18121_);
  or (_18145_, _18144_, _02840_);
  and (_18146_, _18145_, _18142_);
  or (_18147_, _18146_, _02006_);
  or (_18148_, _18129_, _02021_);
  and (_18149_, _18148_, _02025_);
  and (_18150_, _18149_, _18147_);
  and (_18152_, _11508_, _04324_);
  or (_18153_, _18152_, _18136_);
  and (_18154_, _18153_, _01997_);
  or (_18155_, _18154_, _01991_);
  or (_18156_, _18155_, _18150_);
  or (_18157_, _18136_, _11542_);
  and (_18158_, _18157_, _18138_);
  or (_18159_, _18158_, _02861_);
  and (_18160_, _18159_, _02408_);
  and (_18161_, _18160_, _18156_);
  nor (_18163_, _11506_, _07697_);
  or (_18164_, _18163_, _18136_);
  and (_18165_, _18164_, _01875_);
  or (_18166_, _18165_, _05994_);
  or (_18167_, _18166_, _18161_);
  or (_18168_, _18144_, _05249_);
  and (_18169_, _18168_, _18167_);
  or (_18170_, _18169_, _02528_);
  and (_18171_, _05090_, _03670_);
  or (_18172_, _18121_, _02888_);
  or (_18174_, _18172_, _18171_);
  and (_18175_, _18174_, _02043_);
  and (_18176_, _18175_, _18170_);
  nor (_18177_, _11615_, _07689_);
  or (_18178_, _18177_, _18121_);
  and (_18179_, _18178_, _01602_);
  or (_18180_, _18179_, _01869_);
  or (_18181_, _18180_, _18176_);
  and (_18182_, _04672_, _03670_);
  or (_18183_, _18182_, _18121_);
  or (_18185_, _18183_, _01870_);
  and (_18186_, _18185_, _18181_);
  or (_18187_, _18186_, _02079_);
  and (_18188_, _11629_, _03670_);
  or (_18189_, _18121_, _02166_);
  or (_18190_, _18189_, _18188_);
  and (_18191_, _18190_, _02912_);
  and (_18192_, _18191_, _18187_);
  or (_18193_, _18192_, _18124_);
  and (_18194_, _18193_, _02176_);
  or (_18196_, _18121_, _03965_);
  and (_18197_, _18183_, _02072_);
  and (_18198_, _18197_, _18196_);
  or (_18199_, _18198_, _18194_);
  and (_18200_, _18199_, _02907_);
  and (_18201_, _18129_, _02177_);
  and (_18202_, _18201_, _18196_);
  or (_18203_, _18202_, _02071_);
  or (_18204_, _18203_, _18200_);
  nor (_18205_, _11628_, _07689_);
  or (_18207_, _18121_, _04788_);
  or (_18208_, _18207_, _18205_);
  and (_18209_, _18208_, _04793_);
  and (_18210_, _18209_, _18204_);
  nor (_18211_, _11634_, _07689_);
  or (_18212_, _18211_, _18121_);
  and (_18213_, _18212_, _02173_);
  or (_18214_, _18213_, _02201_);
  or (_18215_, _18214_, _18210_);
  or (_18216_, _18126_, _02303_);
  and (_18218_, _18216_, _01887_);
  and (_18219_, _18218_, _18215_);
  and (_18220_, _18153_, _01860_);
  or (_18221_, _18220_, _01537_);
  or (_18222_, _18221_, _18219_);
  and (_18223_, _11685_, _03670_);
  or (_18224_, _18121_, _01538_);
  or (_18225_, _18224_, _18223_);
  and (_18226_, _18225_, _38087_);
  and (_18227_, _18226_, _18222_);
  or (_18229_, _18227_, _18120_);
  and (_40230_, _18229_, _37580_);
  and (_18230_, _38088_, \oc8051_golden_model_1.IP [6]);
  and (_18231_, _07689_, \oc8051_golden_model_1.IP [6]);
  and (_18232_, _11709_, _03670_);
  or (_18233_, _18232_, _18231_);
  and (_18234_, _18233_, _02167_);
  nor (_18235_, _11730_, _07689_);
  or (_18236_, _18235_, _18231_);
  or (_18237_, _18236_, _02814_);
  and (_18239_, _03670_, \oc8051_golden_model_1.ACC [6]);
  or (_18240_, _18239_, _18231_);
  and (_18241_, _18240_, _02817_);
  and (_18242_, _02818_, \oc8051_golden_model_1.IP [6]);
  or (_18243_, _18242_, _02001_);
  or (_18244_, _18243_, _18241_);
  and (_18245_, _18244_, _02024_);
  and (_18246_, _18245_, _18237_);
  and (_18247_, _07697_, \oc8051_golden_model_1.IP [6]);
  and (_18248_, _11717_, _04324_);
  or (_18250_, _18248_, _18247_);
  and (_18251_, _18250_, _02007_);
  or (_18252_, _18251_, _01999_);
  or (_18253_, _18252_, _18246_);
  nor (_18254_, _03808_, _07689_);
  or (_18255_, _18254_, _18231_);
  or (_18256_, _18255_, _02840_);
  and (_18257_, _18256_, _18253_);
  or (_18258_, _18257_, _02006_);
  or (_18259_, _18240_, _02021_);
  and (_18261_, _18259_, _02025_);
  and (_18262_, _18261_, _18258_);
  and (_18263_, _11715_, _04324_);
  or (_18264_, _18263_, _18247_);
  and (_18265_, _18264_, _01997_);
  or (_18266_, _18265_, _01991_);
  or (_18267_, _18266_, _18262_);
  or (_18268_, _18247_, _11747_);
  and (_18269_, _18268_, _18250_);
  or (_18270_, _18269_, _02861_);
  and (_18272_, _18270_, _02408_);
  and (_18273_, _18272_, _18267_);
  nor (_18274_, _11713_, _07697_);
  or (_18275_, _18274_, _18247_);
  and (_18276_, _18275_, _01875_);
  or (_18277_, _18276_, _05994_);
  or (_18278_, _18277_, _18273_);
  or (_18279_, _18255_, _05249_);
  and (_18280_, _18279_, _18278_);
  or (_18281_, _18280_, _02528_);
  and (_18283_, _04861_, _03670_);
  or (_18284_, _18231_, _02888_);
  or (_18285_, _18284_, _18283_);
  and (_18286_, _18285_, _02043_);
  and (_18287_, _18286_, _18281_);
  nor (_18288_, _11820_, _07689_);
  or (_18289_, _18288_, _18231_);
  and (_18290_, _18289_, _01602_);
  or (_18291_, _18290_, _01869_);
  or (_18292_, _18291_, _18287_);
  and (_18294_, _09920_, _03670_);
  or (_18295_, _18294_, _18231_);
  or (_18296_, _18295_, _01870_);
  and (_18297_, _18296_, _18292_);
  or (_18298_, _18297_, _02079_);
  and (_18299_, _11835_, _03670_);
  or (_18300_, _18231_, _02166_);
  or (_18301_, _18300_, _18299_);
  and (_18302_, _18301_, _02912_);
  and (_18303_, _18302_, _18298_);
  or (_18304_, _18303_, _18234_);
  and (_18305_, _18304_, _02176_);
  or (_18306_, _18231_, _03863_);
  and (_18307_, _18295_, _02072_);
  and (_18308_, _18307_, _18306_);
  or (_18309_, _18308_, _18305_);
  and (_18310_, _18309_, _02907_);
  and (_18311_, _18240_, _02177_);
  and (_18312_, _18311_, _18306_);
  or (_18313_, _18312_, _02071_);
  or (_18315_, _18313_, _18310_);
  nor (_18316_, _11833_, _07689_);
  or (_18317_, _18231_, _04788_);
  or (_18318_, _18317_, _18316_);
  and (_18319_, _18318_, _04793_);
  and (_18320_, _18319_, _18315_);
  nor (_18321_, _11708_, _07689_);
  or (_18322_, _18321_, _18231_);
  and (_18323_, _18322_, _02173_);
  or (_18324_, _18323_, _02201_);
  or (_18326_, _18324_, _18320_);
  or (_18327_, _18236_, _02303_);
  and (_18328_, _18327_, _01887_);
  and (_18329_, _18328_, _18326_);
  and (_18330_, _18264_, _01860_);
  or (_18331_, _18330_, _01537_);
  or (_18332_, _18331_, _18329_);
  and (_18333_, _11887_, _03670_);
  or (_18334_, _18231_, _01538_);
  or (_18335_, _18334_, _18333_);
  and (_18336_, _18335_, _38087_);
  and (_18337_, _18336_, _18332_);
  or (_18338_, _18337_, _18230_);
  and (_40231_, _18338_, _37580_);
  and (_18339_, _07791_, \oc8051_golden_model_1.P0 [0]);
  and (_18340_, _10620_, _03832_);
  or (_18341_, _18340_, _18339_);
  and (_18342_, _18341_, _02167_);
  and (_18343_, _03832_, _03028_);
  or (_18344_, _18343_, _18339_);
  or (_18347_, _18344_, _05249_);
  nor (_18348_, _04106_, _07796_);
  or (_18349_, _18348_, _18339_);
  or (_18350_, _18349_, _02814_);
  and (_18351_, _03737_, \oc8051_golden_model_1.ACC [0]);
  or (_18352_, _18351_, _18339_);
  and (_18353_, _18352_, _02817_);
  and (_18354_, _02818_, \oc8051_golden_model_1.P0 [0]);
  or (_18355_, _18354_, _02001_);
  or (_18356_, _18355_, _18353_);
  and (_18358_, _18356_, _02024_);
  and (_18359_, _18358_, _18350_);
  and (_18360_, _07800_, \oc8051_golden_model_1.P0 [0]);
  and (_18361_, _10510_, _03656_);
  or (_18362_, _18361_, _18360_);
  and (_18363_, _18362_, _02007_);
  or (_18364_, _18363_, _18359_);
  and (_18365_, _18364_, _02840_);
  and (_18366_, _18344_, _01999_);
  or (_18367_, _18366_, _02006_);
  or (_18369_, _18367_, _18365_);
  or (_18370_, _18352_, _02021_);
  and (_18371_, _18370_, _02025_);
  and (_18372_, _18371_, _18369_);
  and (_18373_, _18339_, _01997_);
  or (_18374_, _18373_, _01991_);
  or (_18375_, _18374_, _18372_);
  or (_18376_, _18349_, _02861_);
  and (_18377_, _18376_, _02408_);
  and (_18378_, _18377_, _18375_);
  or (_18380_, _10541_, _10519_);
  and (_18381_, _18380_, _03656_);
  or (_18382_, _18381_, _18360_);
  and (_18383_, _18382_, _01875_);
  or (_18384_, _18383_, _05994_);
  or (_18385_, _18384_, _18378_);
  and (_18386_, _18385_, _18347_);
  or (_18387_, _18386_, _02528_);
  or (_18388_, _18339_, _02888_);
  and (_18389_, _04952_, _03737_);
  or (_18391_, _18389_, _18388_);
  and (_18392_, _18391_, _02043_);
  and (_18393_, _18392_, _18387_);
  and (_18394_, _04675_, \oc8051_golden_model_1.P2 [0]);
  and (_18395_, _04703_, \oc8051_golden_model_1.P0 [0]);
  or (_18396_, _18395_, _10561_);
  or (_18397_, _18396_, _18394_);
  and (_18398_, _04706_, \oc8051_golden_model_1.P1 [0]);
  and (_18399_, _04710_, \oc8051_golden_model_1.P3 [0]);
  or (_18400_, _18399_, _18398_);
  nor (_18402_, _18400_, _10562_);
  nand (_18403_, _18402_, _10570_);
  nor (_18404_, _18403_, _18397_);
  and (_18405_, _18404_, _10558_);
  nand (_18406_, _18405_, _10598_);
  or (_18407_, _18406_, _10554_);
  and (_18408_, _18407_, _03737_);
  or (_18409_, _18408_, _18339_);
  and (_18410_, _18409_, _01602_);
  or (_18411_, _18410_, _01869_);
  or (_18413_, _18411_, _18393_);
  and (_18414_, _03737_, _04562_);
  or (_18415_, _18414_, _18339_);
  or (_18416_, _18415_, _01870_);
  and (_18417_, _18416_, _18413_);
  or (_18418_, _18417_, _02079_);
  and (_18419_, _10614_, _03832_);
  or (_18420_, _18339_, _02166_);
  or (_18421_, _18420_, _18419_);
  and (_18422_, _18421_, _02912_);
  and (_18424_, _18422_, _18418_);
  or (_18425_, _18424_, _18342_);
  and (_18426_, _18425_, _02176_);
  nand (_18427_, _18415_, _02072_);
  nor (_18428_, _18427_, _18348_);
  or (_18429_, _18428_, _18426_);
  and (_18430_, _18429_, _02907_);
  or (_18431_, _18339_, _04106_);
  and (_18432_, _18352_, _02177_);
  and (_18433_, _18432_, _18431_);
  or (_18435_, _18433_, _02071_);
  or (_18436_, _18435_, _18430_);
  nor (_18437_, _10613_, _07796_);
  or (_18438_, _18339_, _04788_);
  or (_18439_, _18438_, _18437_);
  and (_18440_, _18439_, _04793_);
  and (_18441_, _18440_, _18436_);
  nor (_18442_, _10619_, _07796_);
  or (_18443_, _18442_, _18339_);
  and (_18444_, _18443_, _02173_);
  or (_18446_, _18444_, _02201_);
  or (_18447_, _18446_, _18441_);
  or (_18448_, _18349_, _02303_);
  and (_18449_, _18448_, _01887_);
  and (_18450_, _18449_, _18447_);
  and (_18451_, _18339_, _01860_);
  or (_18452_, _18451_, _01537_);
  or (_18453_, _18452_, _18450_);
  or (_18454_, _18349_, _01538_);
  and (_18455_, _18454_, _38087_);
  and (_18457_, _18455_, _18453_);
  nor (_18458_, \oc8051_golden_model_1.P0 [0], rst);
  nor (_18459_, _18458_, _03183_);
  or (_40233_, _18459_, _18457_);
  and (_18460_, _07791_, \oc8051_golden_model_1.P0 [1]);
  nor (_18461_, _07796_, _02811_);
  or (_18462_, _18461_, _18460_);
  or (_18463_, _18462_, _02840_);
  or (_18464_, _03737_, \oc8051_golden_model_1.P0 [1]);
  nand (_18465_, _10698_, _03832_);
  and (_18467_, _18465_, _18464_);
  or (_18468_, _18467_, _02814_);
  nand (_18469_, _03832_, _01613_);
  and (_18470_, _18469_, _18464_);
  and (_18471_, _18470_, _02817_);
  and (_18472_, _02818_, \oc8051_golden_model_1.P0 [1]);
  or (_18473_, _18472_, _02001_);
  or (_18474_, _18473_, _18471_);
  and (_18475_, _18474_, _02024_);
  and (_18476_, _18475_, _18468_);
  and (_18477_, _07800_, \oc8051_golden_model_1.P0 [1]);
  and (_18478_, _10710_, _03656_);
  or (_18479_, _18478_, _18477_);
  and (_18480_, _18479_, _02007_);
  or (_18481_, _18480_, _01999_);
  or (_18482_, _18481_, _18476_);
  and (_18483_, _18482_, _18463_);
  or (_18484_, _18483_, _02006_);
  or (_18485_, _18470_, _02021_);
  and (_18486_, _18485_, _02025_);
  and (_18488_, _18486_, _18484_);
  and (_18489_, _10696_, _03656_);
  or (_18490_, _18489_, _18477_);
  and (_18491_, _18490_, _01997_);
  or (_18492_, _18491_, _01991_);
  or (_18493_, _18492_, _18488_);
  and (_18494_, _18478_, _10725_);
  or (_18495_, _18477_, _02861_);
  or (_18496_, _18495_, _18494_);
  and (_18497_, _18496_, _18493_);
  and (_18499_, _18497_, _02408_);
  or (_18500_, _10741_, _10696_);
  and (_18501_, _18500_, _03656_);
  or (_18502_, _18477_, _18501_);
  and (_18503_, _18502_, _01875_);
  or (_18504_, _18503_, _05994_);
  or (_18505_, _18504_, _18499_);
  or (_18506_, _18462_, _05249_);
  and (_18507_, _18506_, _18505_);
  or (_18508_, _18507_, _02528_);
  and (_18510_, _04907_, _03737_);
  or (_18511_, _18460_, _02888_);
  or (_18512_, _18511_, _18510_);
  and (_18513_, _18512_, _02043_);
  and (_18514_, _18513_, _18508_);
  and (_18515_, _18464_, _01602_);
  and (_18516_, _04703_, \oc8051_golden_model_1.P0 [1]);
  and (_18517_, _04675_, \oc8051_golden_model_1.P2 [1]);
  or (_18518_, _18517_, _18516_);
  and (_18519_, _04706_, \oc8051_golden_model_1.P1 [1]);
  and (_18521_, _04710_, \oc8051_golden_model_1.P3 [1]);
  or (_18522_, _18521_, _18519_);
  or (_18523_, _18522_, _10784_);
  nor (_18524_, _18523_, _18518_);
  and (_18525_, _18524_, _10797_);
  and (_18526_, _18525_, _10777_);
  nand (_18527_, _18526_, _10771_);
  or (_18528_, _18527_, _10754_);
  or (_18529_, _18528_, _07796_);
  and (_18530_, _18529_, _18515_);
  or (_18532_, _18530_, _18514_);
  and (_18533_, _18532_, _01870_);
  and (_18534_, _18464_, _01869_);
  nand (_18535_, _03832_, _02687_);
  and (_18536_, _18535_, _18534_);
  or (_18537_, _18536_, _18533_);
  and (_18538_, _18537_, _02166_);
  and (_18539_, _10816_, _03737_);
  or (_18540_, _18539_, _18460_);
  and (_18541_, _18540_, _02079_);
  or (_18543_, _18541_, _18538_);
  and (_18544_, _18543_, _02912_);
  or (_18545_, _10822_, _07796_);
  and (_18546_, _18464_, _02167_);
  and (_18547_, _18546_, _18545_);
  or (_18548_, _18547_, _18544_);
  and (_18549_, _18548_, _02176_);
  and (_18550_, _10692_, _03737_);
  or (_18551_, _18550_, _18460_);
  and (_18552_, _18551_, _02072_);
  or (_18554_, _18552_, _18549_);
  and (_18555_, _18554_, _02907_);
  or (_18556_, _18460_, _04058_);
  and (_18557_, _18470_, _02177_);
  and (_18558_, _18557_, _18556_);
  or (_18559_, _18558_, _18555_);
  and (_18560_, _18559_, _02174_);
  or (_18561_, _18469_, _04058_);
  and (_18562_, _18464_, _02173_);
  and (_18563_, _18562_, _18561_);
  or (_18565_, _18563_, _02201_);
  or (_18566_, _18535_, _04058_);
  and (_18567_, _18464_, _02071_);
  and (_18568_, _18567_, _18566_);
  or (_18569_, _18568_, _18565_);
  or (_18570_, _18569_, _18560_);
  or (_18571_, _18467_, _02303_);
  and (_18572_, _18571_, _01887_);
  and (_18573_, _18572_, _18570_);
  and (_18574_, _18490_, _01860_);
  or (_18576_, _18574_, _01537_);
  or (_18577_, _18576_, _18573_);
  nor (_18578_, _18460_, _01538_);
  nand (_18579_, _18578_, _18465_);
  and (_18580_, _18579_, _38087_);
  and (_18581_, _18580_, _18577_);
  nor (_18582_, \oc8051_golden_model_1.P0 [1], rst);
  nor (_18583_, _18582_, _03183_);
  or (_40234_, _18583_, _18581_);
  and (_18584_, _07791_, \oc8051_golden_model_1.P0 [2]);
  and (_18586_, _11020_, _03832_);
  or (_18587_, _18586_, _18584_);
  and (_18588_, _18587_, _02167_);
  nor (_18589_, _07796_, _03455_);
  or (_18590_, _18589_, _18584_);
  or (_18591_, _18590_, _05249_);
  or (_18592_, _18590_, _02840_);
  nor (_18593_, _10905_, _07796_);
  or (_18594_, _18593_, _18584_);
  or (_18595_, _18594_, _02814_);
  and (_18597_, _03737_, \oc8051_golden_model_1.ACC [2]);
  or (_18598_, _18597_, _18584_);
  and (_18599_, _18598_, _02817_);
  and (_18600_, _02818_, \oc8051_golden_model_1.P0 [2]);
  or (_18601_, _18600_, _02001_);
  or (_18602_, _18601_, _18599_);
  and (_18603_, _18602_, _02024_);
  and (_18604_, _18603_, _18595_);
  and (_18605_, _07800_, \oc8051_golden_model_1.P0 [2]);
  and (_18606_, _10909_, _03656_);
  or (_18608_, _18606_, _18605_);
  and (_18609_, _18608_, _02007_);
  or (_18610_, _18609_, _01999_);
  or (_18611_, _18610_, _18604_);
  and (_18612_, _18611_, _18592_);
  or (_18613_, _18612_, _02006_);
  or (_18614_, _18598_, _02021_);
  and (_18615_, _18614_, _02025_);
  and (_18616_, _18615_, _18613_);
  and (_18617_, _10894_, _03656_);
  or (_18619_, _18617_, _18605_);
  and (_18620_, _18619_, _01997_);
  or (_18621_, _18620_, _01991_);
  or (_18622_, _18621_, _18616_);
  and (_18623_, _18606_, _10924_);
  or (_18624_, _18605_, _02861_);
  or (_18625_, _18624_, _18623_);
  and (_18626_, _18625_, _02408_);
  and (_18627_, _18626_, _18622_);
  or (_18628_, _10941_, _10894_);
  and (_18630_, _18628_, _03656_);
  or (_18631_, _18630_, _18605_);
  and (_18632_, _18631_, _01875_);
  or (_18633_, _18632_, _05994_);
  or (_18634_, _18633_, _18627_);
  and (_18635_, _18634_, _18591_);
  or (_18636_, _18635_, _02528_);
  or (_18637_, _18584_, _02888_);
  and (_18638_, _05043_, _03737_);
  or (_18639_, _18638_, _18637_);
  and (_18641_, _18639_, _02043_);
  and (_18642_, _18641_, _18636_);
  and (_18643_, _04703_, \oc8051_golden_model_1.P0 [2]);
  and (_18644_, _04675_, \oc8051_golden_model_1.P2 [2]);
  or (_18645_, _18644_, _18643_);
  and (_18646_, _04706_, \oc8051_golden_model_1.P1 [2]);
  and (_18647_, _04710_, \oc8051_golden_model_1.P3 [2]);
  or (_18648_, _18647_, _18646_);
  or (_18649_, _18648_, _10963_);
  nor (_18650_, _18649_, _18645_);
  and (_18652_, _18650_, _10981_);
  and (_18653_, _18652_, _10962_);
  nand (_18654_, _18653_, _10998_);
  or (_18655_, _18654_, _10954_);
  and (_18656_, _18655_, _03737_);
  or (_18657_, _18656_, _18584_);
  and (_18658_, _18657_, _01602_);
  or (_18659_, _18658_, _01869_);
  or (_18660_, _18659_, _18642_);
  and (_18661_, _03737_, _04724_);
  or (_18663_, _18661_, _18584_);
  or (_18664_, _18663_, _01870_);
  and (_18665_, _18664_, _18660_);
  or (_18666_, _18665_, _02079_);
  and (_18667_, _11014_, _03832_);
  or (_18668_, _18584_, _02166_);
  or (_18669_, _18668_, _18667_);
  and (_18670_, _18669_, _02912_);
  and (_18671_, _18670_, _18666_);
  or (_18672_, _18671_, _18588_);
  and (_18674_, _18672_, _02176_);
  or (_18675_, _18584_, _04156_);
  and (_18676_, _18663_, _02072_);
  and (_18677_, _18676_, _18675_);
  or (_18678_, _18677_, _18674_);
  and (_18679_, _18678_, _02907_);
  and (_18680_, _18598_, _02177_);
  and (_18681_, _18680_, _18675_);
  or (_18682_, _18681_, _02071_);
  or (_18683_, _18682_, _18679_);
  nor (_18685_, _11013_, _07796_);
  or (_18686_, _18584_, _04788_);
  or (_18687_, _18686_, _18685_);
  and (_18688_, _18687_, _04793_);
  and (_18689_, _18688_, _18683_);
  nor (_18690_, _11019_, _07796_);
  or (_18691_, _18690_, _18584_);
  and (_18692_, _18691_, _02173_);
  or (_18693_, _18692_, _02201_);
  or (_18694_, _18693_, _18689_);
  or (_18696_, _18594_, _02303_);
  and (_18697_, _18696_, _01887_);
  and (_18698_, _18697_, _18694_);
  and (_18699_, _18619_, _01860_);
  or (_18700_, _18699_, _01537_);
  or (_18701_, _18700_, _18698_);
  and (_18702_, _11072_, _03832_);
  or (_18703_, _18584_, _01538_);
  or (_18704_, _18703_, _18702_);
  and (_18705_, _18704_, _38087_);
  and (_18707_, _18705_, _18701_);
  nor (_18708_, \oc8051_golden_model_1.P0 [2], rst);
  nor (_18709_, _18708_, _03183_);
  or (_40235_, _18709_, _18707_);
  and (_18710_, _07791_, \oc8051_golden_model_1.P0 [3]);
  and (_18711_, _11094_, _03832_);
  or (_18712_, _18711_, _18710_);
  and (_18713_, _18712_, _02167_);
  nor (_18714_, _07796_, _03268_);
  or (_18715_, _18714_, _18710_);
  or (_18717_, _18715_, _05249_);
  nor (_18718_, _11101_, _07796_);
  or (_18719_, _18718_, _18710_);
  or (_18720_, _18719_, _02814_);
  and (_18721_, _03737_, \oc8051_golden_model_1.ACC [3]);
  or (_18722_, _18721_, _18710_);
  and (_18723_, _18722_, _02817_);
  and (_18724_, _02818_, \oc8051_golden_model_1.P0 [3]);
  or (_18725_, _18724_, _02001_);
  or (_18726_, _18725_, _18723_);
  and (_18728_, _18726_, _02024_);
  and (_18729_, _18728_, _18720_);
  and (_18730_, _07800_, \oc8051_golden_model_1.P0 [3]);
  and (_18731_, _11098_, _03656_);
  or (_18732_, _18731_, _18730_);
  and (_18733_, _18732_, _02007_);
  or (_18734_, _18733_, _01999_);
  or (_18735_, _18734_, _18729_);
  or (_18736_, _18715_, _02840_);
  and (_18737_, _18736_, _18735_);
  or (_18739_, _18737_, _02006_);
  or (_18740_, _18722_, _02021_);
  and (_18741_, _18740_, _02025_);
  and (_18742_, _18741_, _18739_);
  and (_18743_, _11096_, _03656_);
  or (_18744_, _18743_, _18730_);
  and (_18745_, _18744_, _01997_);
  or (_18746_, _18745_, _01991_);
  or (_18747_, _18746_, _18742_);
  or (_18748_, _18730_, _11127_);
  and (_18750_, _18748_, _18732_);
  or (_18751_, _18750_, _02861_);
  and (_18752_, _18751_, _02408_);
  and (_18753_, _18752_, _18747_);
  or (_18754_, _11096_, _11143_);
  and (_18755_, _18754_, _03656_);
  or (_18756_, _18755_, _18730_);
  and (_18757_, _18756_, _01875_);
  or (_18758_, _18757_, _05994_);
  or (_18759_, _18758_, _18753_);
  and (_18761_, _18759_, _18717_);
  or (_18762_, _18761_, _02528_);
  or (_18763_, _18710_, _02888_);
  and (_18764_, _04998_, _03737_);
  or (_18765_, _18764_, _18763_);
  and (_18766_, _18765_, _02043_);
  and (_18767_, _18766_, _18762_);
  and (_18768_, _04703_, \oc8051_golden_model_1.P0 [3]);
  and (_18769_, _04675_, \oc8051_golden_model_1.P2 [3]);
  or (_18770_, _18769_, _18768_);
  and (_18772_, _04706_, \oc8051_golden_model_1.P1 [3]);
  and (_18773_, _04710_, \oc8051_golden_model_1.P3 [3]);
  or (_18774_, _18773_, _18772_);
  or (_18775_, _18774_, _11191_);
  nor (_18776_, _18775_, _18770_);
  and (_18777_, _18776_, _11202_);
  and (_18778_, _18777_, _11183_);
  nand (_18779_, _18778_, _11176_);
  or (_18780_, _18779_, _11158_);
  and (_18781_, _18780_, _03737_);
  or (_18783_, _18781_, _18710_);
  and (_18784_, _18783_, _01602_);
  or (_18785_, _18784_, _01869_);
  or (_18786_, _18785_, _18767_);
  and (_18787_, _03737_, _04678_);
  or (_18788_, _18787_, _18710_);
  or (_18789_, _18788_, _01870_);
  and (_18790_, _18789_, _18786_);
  or (_18791_, _18790_, _02079_);
  and (_18792_, _11222_, _03832_);
  or (_18794_, _18710_, _02166_);
  or (_18795_, _18794_, _18792_);
  and (_18796_, _18795_, _02912_);
  and (_18797_, _18796_, _18791_);
  or (_18798_, _18797_, _18713_);
  and (_18799_, _18798_, _02176_);
  or (_18800_, _18710_, _04014_);
  and (_18801_, _18788_, _02072_);
  and (_18802_, _18801_, _18800_);
  or (_18803_, _18802_, _18799_);
  and (_18805_, _18803_, _02907_);
  and (_18806_, _18722_, _02177_);
  and (_18807_, _18806_, _18800_);
  or (_18808_, _18807_, _02071_);
  or (_18809_, _18808_, _18805_);
  nor (_18810_, _11220_, _07796_);
  or (_18811_, _18710_, _04788_);
  or (_18812_, _18811_, _18810_);
  and (_18813_, _18812_, _04793_);
  and (_18814_, _18813_, _18809_);
  nor (_18815_, _11093_, _07796_);
  or (_18816_, _18815_, _18710_);
  and (_18817_, _18816_, _02173_);
  or (_18818_, _18817_, _02201_);
  or (_18819_, _18818_, _18814_);
  or (_18820_, _18719_, _02303_);
  and (_18821_, _18820_, _01887_);
  and (_18822_, _18821_, _18819_);
  and (_18823_, _18744_, _01860_);
  or (_18824_, _18823_, _01537_);
  or (_18827_, _18824_, _18822_);
  and (_18828_, _11273_, _03832_);
  or (_18829_, _18710_, _01538_);
  or (_18830_, _18829_, _18828_);
  and (_18831_, _18830_, _38087_);
  and (_18832_, _18831_, _18827_);
  nor (_18833_, \oc8051_golden_model_1.P0 [3], rst);
  nor (_18834_, _18833_, _03183_);
  or (_40236_, _18834_, _18832_);
  and (_18835_, _07791_, \oc8051_golden_model_1.P0 [4]);
  and (_18837_, _11431_, _03832_);
  or (_18838_, _18837_, _18835_);
  and (_18839_, _18838_, _02167_);
  nor (_18840_, _04211_, _07796_);
  or (_18841_, _18840_, _18835_);
  or (_18842_, _18841_, _05249_);
  and (_18843_, _07800_, \oc8051_golden_model_1.P0 [4]);
  and (_18844_, _11301_, _03656_);
  or (_18845_, _18844_, _18843_);
  and (_18846_, _18845_, _01997_);
  nor (_18848_, _11317_, _07796_);
  or (_18849_, _18848_, _18835_);
  or (_18850_, _18849_, _02814_);
  and (_18851_, _03737_, \oc8051_golden_model_1.ACC [4]);
  or (_18852_, _18851_, _18835_);
  and (_18853_, _18852_, _02817_);
  and (_18854_, _02818_, \oc8051_golden_model_1.P0 [4]);
  or (_18855_, _18854_, _02001_);
  or (_18856_, _18855_, _18853_);
  and (_18857_, _18856_, _02024_);
  and (_18859_, _18857_, _18850_);
  and (_18860_, _11303_, _03656_);
  or (_18861_, _18860_, _18843_);
  and (_18862_, _18861_, _02007_);
  or (_18863_, _18862_, _01999_);
  or (_18864_, _18863_, _18859_);
  or (_18865_, _18841_, _02840_);
  and (_18866_, _18865_, _18864_);
  or (_18867_, _18866_, _02006_);
  or (_18868_, _18852_, _02021_);
  and (_18870_, _18868_, _02025_);
  and (_18871_, _18870_, _18867_);
  or (_18872_, _18871_, _18846_);
  and (_18873_, _18872_, _02861_);
  or (_18874_, _18843_, _11334_);
  and (_18875_, _18874_, _01991_);
  and (_18876_, _18875_, _18861_);
  or (_18877_, _18876_, _18873_);
  and (_18878_, _18877_, _02408_);
  or (_18879_, _11301_, _11298_);
  and (_18881_, _18879_, _03656_);
  or (_18882_, _18881_, _18843_);
  and (_18883_, _18882_, _01875_);
  or (_18884_, _18883_, _05994_);
  or (_18885_, _18884_, _18878_);
  and (_18886_, _18885_, _18842_);
  or (_18887_, _18886_, _02528_);
  or (_18888_, _18835_, _02888_);
  and (_18889_, _05135_, _03737_);
  or (_18890_, _18889_, _18888_);
  and (_18892_, _18890_, _02043_);
  and (_18893_, _18892_, _18887_);
  and (_18894_, _04675_, \oc8051_golden_model_1.P2 [4]);
  and (_18895_, _04703_, \oc8051_golden_model_1.P0 [4]);
  or (_18896_, _18895_, _11377_);
  nor (_18897_, _18896_, _18894_);
  and (_18898_, _18897_, _11374_);
  nand (_18899_, _18898_, _11365_);
  and (_18900_, _04706_, \oc8051_golden_model_1.P1 [4]);
  and (_18901_, _04710_, \oc8051_golden_model_1.P3 [4]);
  or (_18903_, _18901_, _18900_);
  or (_18904_, _18903_, _11378_);
  nor (_18905_, _18904_, _11390_);
  and (_18906_, _18905_, _11407_);
  nand (_18907_, _18906_, _11389_);
  or (_18908_, _18907_, _18899_);
  or (_18909_, _18908_, _11361_);
  and (_18910_, _18909_, _03832_);
  or (_18911_, _18910_, _18835_);
  and (_18912_, _18911_, _01602_);
  or (_18914_, _18912_, _01869_);
  or (_18915_, _18914_, _18893_);
  and (_18916_, _04694_, _03737_);
  or (_18917_, _18916_, _18835_);
  or (_18918_, _18917_, _01870_);
  and (_18919_, _18918_, _18915_);
  or (_18920_, _18919_, _02079_);
  and (_18921_, _11425_, _03832_);
  or (_18922_, _18835_, _02166_);
  or (_18923_, _18922_, _18921_);
  and (_18925_, _18923_, _02912_);
  and (_18926_, _18925_, _18920_);
  or (_18927_, _18926_, _18839_);
  and (_18928_, _18927_, _02176_);
  or (_18929_, _18835_, _04258_);
  and (_18930_, _18917_, _02072_);
  and (_18931_, _18930_, _18929_);
  or (_18932_, _18931_, _18928_);
  and (_18933_, _18932_, _02907_);
  and (_18934_, _18852_, _02177_);
  and (_18936_, _18934_, _18929_);
  or (_18937_, _18936_, _02071_);
  or (_18938_, _18937_, _18933_);
  nor (_18939_, _11424_, _07796_);
  or (_18940_, _18835_, _04788_);
  or (_18941_, _18940_, _18939_);
  and (_18942_, _18941_, _04793_);
  and (_18943_, _18942_, _18938_);
  nor (_18944_, _11430_, _07796_);
  or (_18945_, _18944_, _18835_);
  and (_18947_, _18945_, _02173_);
  or (_18948_, _18947_, _02201_);
  or (_18949_, _18948_, _18943_);
  or (_18950_, _18849_, _02303_);
  and (_18951_, _18950_, _01887_);
  and (_18952_, _18951_, _18949_);
  and (_18953_, _18845_, _01860_);
  or (_18954_, _18953_, _01537_);
  or (_18955_, _18954_, _18952_);
  and (_18956_, _11487_, _03832_);
  or (_18958_, _18835_, _01538_);
  or (_18959_, _18958_, _18956_);
  and (_18960_, _18959_, _38087_);
  and (_18961_, _18960_, _18955_);
  nor (_18962_, \oc8051_golden_model_1.P0 [4], rst);
  nor (_18963_, _18962_, _03183_);
  or (_40237_, _18963_, _18961_);
  nor (_18964_, \oc8051_golden_model_1.P0 [5], rst);
  nor (_18965_, _18964_, _03183_);
  and (_18966_, _07791_, \oc8051_golden_model_1.P0 [5]);
  and (_18968_, _11635_, _03832_);
  or (_18969_, _18968_, _18966_);
  and (_18970_, _18969_, _02167_);
  nor (_18971_, _11525_, _07796_);
  or (_18972_, _18971_, _18966_);
  or (_18973_, _18972_, _02814_);
  and (_18974_, _03737_, \oc8051_golden_model_1.ACC [5]);
  or (_18975_, _18974_, _18966_);
  and (_18976_, _18975_, _02817_);
  and (_18977_, _02818_, \oc8051_golden_model_1.P0 [5]);
  or (_18979_, _18977_, _02001_);
  or (_18980_, _18979_, _18976_);
  and (_18981_, _18980_, _02024_);
  and (_18982_, _18981_, _18973_);
  and (_18983_, _07800_, \oc8051_golden_model_1.P0 [5]);
  and (_18984_, _11510_, _03656_);
  or (_18985_, _18984_, _18983_);
  and (_18986_, _18985_, _02007_);
  or (_18987_, _18986_, _01999_);
  or (_18988_, _18987_, _18982_);
  nor (_18990_, _03916_, _07796_);
  or (_18991_, _18990_, _18966_);
  or (_18992_, _18991_, _02840_);
  and (_18993_, _18992_, _18988_);
  or (_18994_, _18993_, _02006_);
  or (_18995_, _18975_, _02021_);
  and (_18996_, _18995_, _02025_);
  and (_18997_, _18996_, _18994_);
  and (_18998_, _11508_, _03656_);
  or (_18999_, _18998_, _18983_);
  and (_19001_, _18999_, _01997_);
  or (_19002_, _19001_, _01991_);
  or (_19003_, _19002_, _18997_);
  or (_19004_, _18983_, _11542_);
  and (_19005_, _19004_, _18985_);
  or (_19006_, _19005_, _02861_);
  and (_19007_, _19006_, _02408_);
  and (_19008_, _19007_, _19003_);
  or (_19009_, _11508_, _11505_);
  and (_19010_, _19009_, _03656_);
  or (_19012_, _19010_, _18983_);
  and (_19013_, _19012_, _01875_);
  or (_19014_, _19013_, _05994_);
  or (_19015_, _19014_, _19008_);
  or (_19016_, _18991_, _05249_);
  and (_19017_, _19016_, _19015_);
  or (_19018_, _19017_, _02528_);
  and (_19019_, _05090_, _03737_);
  or (_19020_, _18966_, _02888_);
  or (_19021_, _19020_, _19019_);
  and (_19023_, _19021_, _02043_);
  and (_19024_, _19023_, _19018_);
  and (_19025_, _04703_, \oc8051_golden_model_1.P0 [5]);
  and (_19026_, _04675_, \oc8051_golden_model_1.P2 [5]);
  or (_19027_, _19026_, _19025_);
  and (_19028_, _04706_, \oc8051_golden_model_1.P1 [5]);
  and (_19029_, _04710_, \oc8051_golden_model_1.P3 [5]);
  or (_19030_, _19029_, _19028_);
  or (_19031_, _19030_, _11578_);
  nor (_19032_, _19031_, _19027_);
  and (_19034_, _19032_, _11596_);
  and (_19035_, _19034_, _11577_);
  nand (_19036_, _19035_, _11613_);
  or (_19037_, _19036_, _11569_);
  and (_19038_, _19037_, _03832_);
  or (_19039_, _19038_, _18966_);
  and (_19040_, _19039_, _01602_);
  or (_19041_, _19040_, _01869_);
  or (_19042_, _19041_, _19024_);
  and (_19043_, _04672_, _03737_);
  or (_19045_, _19043_, _18966_);
  or (_19046_, _19045_, _01870_);
  and (_19047_, _19046_, _19042_);
  or (_19048_, _19047_, _02079_);
  and (_19049_, _11629_, _03832_);
  or (_19050_, _18966_, _02166_);
  or (_19051_, _19050_, _19049_);
  and (_19052_, _19051_, _02912_);
  and (_19053_, _19052_, _19048_);
  or (_19054_, _19053_, _18970_);
  and (_19056_, _19054_, _02176_);
  or (_19057_, _18966_, _03965_);
  and (_19058_, _19045_, _02072_);
  and (_19059_, _19058_, _19057_);
  or (_19060_, _19059_, _19056_);
  and (_19061_, _19060_, _02907_);
  and (_19062_, _18975_, _02177_);
  and (_19063_, _19062_, _19057_);
  or (_19064_, _19063_, _02071_);
  or (_19065_, _19064_, _19061_);
  nor (_19067_, _11628_, _07796_);
  or (_19068_, _18966_, _04788_);
  or (_19069_, _19068_, _19067_);
  and (_19070_, _19069_, _04793_);
  and (_19071_, _19070_, _19065_);
  nor (_19072_, _11634_, _07796_);
  or (_19073_, _19072_, _18966_);
  and (_19074_, _19073_, _02173_);
  or (_19075_, _19074_, _02201_);
  or (_19076_, _19075_, _19071_);
  or (_19078_, _18972_, _02303_);
  and (_19079_, _19078_, _01887_);
  and (_19080_, _19079_, _19076_);
  and (_19081_, _18999_, _01860_);
  or (_19082_, _19081_, _01537_);
  or (_19083_, _19082_, _19080_);
  and (_19084_, _11685_, _03832_);
  or (_19085_, _18966_, _01538_);
  or (_19086_, _19085_, _19084_);
  and (_19087_, _19086_, _38087_);
  and (_19089_, _19087_, _19083_);
  or (_40238_, _19089_, _18965_);
  and (_19090_, _07791_, \oc8051_golden_model_1.P0 [6]);
  and (_19091_, _11709_, _03832_);
  or (_19092_, _19091_, _19090_);
  and (_19093_, _19092_, _02167_);
  nor (_19094_, _11730_, _07796_);
  or (_19095_, _19094_, _19090_);
  or (_19096_, _19095_, _02814_);
  and (_19097_, _03737_, \oc8051_golden_model_1.ACC [6]);
  or (_19099_, _19097_, _19090_);
  and (_19100_, _19099_, _02817_);
  and (_19101_, _02818_, \oc8051_golden_model_1.P0 [6]);
  or (_19102_, _19101_, _02001_);
  or (_19103_, _19102_, _19100_);
  and (_19104_, _19103_, _02024_);
  and (_19105_, _19104_, _19096_);
  and (_19106_, _07800_, \oc8051_golden_model_1.P0 [6]);
  and (_19107_, _11717_, _03656_);
  or (_19108_, _19107_, _19106_);
  and (_19110_, _19108_, _02007_);
  or (_19111_, _19110_, _01999_);
  or (_19112_, _19111_, _19105_);
  nor (_19113_, _03808_, _07796_);
  or (_19114_, _19113_, _19090_);
  or (_19115_, _19114_, _02840_);
  and (_19116_, _19115_, _19112_);
  or (_19117_, _19116_, _02006_);
  or (_19118_, _19099_, _02021_);
  and (_19119_, _19118_, _02025_);
  and (_19121_, _19119_, _19117_);
  and (_19122_, _11715_, _03656_);
  or (_19123_, _19122_, _19106_);
  and (_19124_, _19123_, _01997_);
  or (_19125_, _19124_, _01991_);
  or (_19126_, _19125_, _19121_);
  or (_19127_, _19106_, _11747_);
  and (_19128_, _19127_, _19108_);
  or (_19129_, _19128_, _02861_);
  and (_19130_, _19129_, _02408_);
  and (_19132_, _19130_, _19126_);
  or (_19133_, _11715_, _11712_);
  and (_19134_, _19133_, _03656_);
  or (_19135_, _19134_, _19106_);
  and (_19136_, _19135_, _01875_);
  or (_19137_, _19136_, _05994_);
  or (_19138_, _19137_, _19132_);
  or (_19139_, _19114_, _05249_);
  and (_19140_, _19139_, _19138_);
  or (_19141_, _19140_, _02528_);
  and (_19143_, _04861_, _03737_);
  or (_19144_, _19090_, _02888_);
  or (_19145_, _19144_, _19143_);
  and (_19146_, _19145_, _02043_);
  and (_19147_, _19146_, _19141_);
  and (_19148_, _04675_, \oc8051_golden_model_1.P2 [6]);
  and (_19149_, _04703_, \oc8051_golden_model_1.P0 [6]);
  or (_19150_, _19149_, _11780_);
  or (_19151_, _19150_, _19148_);
  and (_19152_, _04706_, \oc8051_golden_model_1.P1 [6]);
  and (_19154_, _04710_, \oc8051_golden_model_1.P3 [6]);
  or (_19155_, _19154_, _19152_);
  nor (_19156_, _19155_, _11781_);
  nand (_19157_, _19156_, _11789_);
  nor (_19158_, _19157_, _19151_);
  and (_19159_, _19158_, _11777_);
  nand (_19160_, _19159_, _11817_);
  or (_19161_, _19160_, _11774_);
  and (_19162_, _19161_, _03832_);
  or (_19163_, _19162_, _19090_);
  and (_19165_, _19163_, _01602_);
  or (_19166_, _19165_, _01869_);
  or (_19167_, _19166_, _19147_);
  and (_19168_, _09920_, _03737_);
  or (_19169_, _19168_, _19090_);
  or (_19170_, _19169_, _01870_);
  and (_19171_, _19170_, _19167_);
  or (_19172_, _19171_, _02079_);
  and (_19173_, _11835_, _03832_);
  or (_19174_, _19090_, _02166_);
  or (_19176_, _19174_, _19173_);
  and (_19177_, _19176_, _02912_);
  and (_19178_, _19177_, _19172_);
  or (_19179_, _19178_, _19093_);
  and (_19180_, _19179_, _02176_);
  or (_19181_, _19090_, _03863_);
  and (_19182_, _19169_, _02072_);
  and (_19183_, _19182_, _19181_);
  or (_19184_, _19183_, _19180_);
  and (_19185_, _19184_, _02907_);
  and (_19187_, _19099_, _02177_);
  and (_19188_, _19187_, _19181_);
  or (_19189_, _19188_, _02071_);
  or (_19190_, _19189_, _19185_);
  nor (_19191_, _11833_, _07796_);
  or (_19192_, _19090_, _04788_);
  or (_19193_, _19192_, _19191_);
  and (_19194_, _19193_, _04793_);
  and (_19195_, _19194_, _19190_);
  nor (_19196_, _11708_, _07796_);
  or (_19198_, _19196_, _19090_);
  and (_19199_, _19198_, _02173_);
  or (_19200_, _19199_, _02201_);
  or (_19201_, _19200_, _19195_);
  or (_19202_, _19095_, _02303_);
  and (_19203_, _19202_, _01887_);
  and (_19204_, _19203_, _19201_);
  and (_19205_, _19123_, _01860_);
  or (_19206_, _19205_, _01537_);
  or (_19207_, _19206_, _19204_);
  and (_19209_, _11887_, _03832_);
  or (_19210_, _19090_, _01538_);
  or (_19211_, _19210_, _19209_);
  and (_19212_, _19211_, _38087_);
  and (_19213_, _19212_, _19207_);
  nor (_19214_, \oc8051_golden_model_1.P0 [6], rst);
  nor (_19215_, _19214_, _03183_);
  or (_40240_, _19215_, _19213_);
  nor (_19216_, \oc8051_golden_model_1.P1 [0], rst);
  nor (_19217_, _19216_, _03183_);
  and (_19219_, _07909_, \oc8051_golden_model_1.P1 [0]);
  and (_19220_, _10620_, _03698_);
  or (_19221_, _19220_, _19219_);
  and (_19222_, _19221_, _02167_);
  and (_19223_, _03698_, _03028_);
  or (_19224_, _19223_, _19219_);
  or (_19225_, _19224_, _05249_);
  nor (_19226_, _04106_, _07909_);
  or (_19227_, _19226_, _19219_);
  or (_19228_, _19227_, _02814_);
  and (_19230_, _03698_, \oc8051_golden_model_1.ACC [0]);
  or (_19231_, _19230_, _19219_);
  and (_19232_, _19231_, _02817_);
  and (_19233_, _02818_, \oc8051_golden_model_1.P1 [0]);
  or (_19234_, _19233_, _02001_);
  or (_19235_, _19234_, _19232_);
  and (_19236_, _19235_, _02024_);
  and (_19237_, _19236_, _19228_);
  and (_19238_, _07917_, \oc8051_golden_model_1.P1 [0]);
  and (_19239_, _10510_, _04336_);
  or (_19241_, _19239_, _19238_);
  and (_19242_, _19241_, _02007_);
  or (_19243_, _19242_, _19237_);
  and (_19244_, _19243_, _02840_);
  and (_19245_, _19224_, _01999_);
  or (_19246_, _19245_, _02006_);
  or (_19247_, _19246_, _19244_);
  or (_19248_, _19231_, _02021_);
  and (_19249_, _19248_, _02025_);
  and (_19250_, _19249_, _19247_);
  and (_19252_, _19219_, _01997_);
  or (_19253_, _19252_, _01991_);
  or (_19254_, _19253_, _19250_);
  or (_19255_, _19227_, _02861_);
  and (_19256_, _19255_, _02408_);
  and (_19257_, _19256_, _19254_);
  and (_19258_, _18380_, _04336_);
  or (_19259_, _19258_, _19238_);
  and (_19260_, _19259_, _01875_);
  or (_19261_, _19260_, _05994_);
  or (_19263_, _19261_, _19257_);
  and (_19264_, _19263_, _19225_);
  or (_19265_, _19264_, _02528_);
  and (_19266_, _04952_, _03698_);
  or (_19267_, _19219_, _02888_);
  or (_19268_, _19267_, _19266_);
  and (_19269_, _19268_, _02043_);
  and (_19270_, _19269_, _19265_);
  and (_19271_, _18407_, _03698_);
  or (_19272_, _19271_, _19219_);
  and (_19274_, _19272_, _01602_);
  or (_19275_, _19274_, _01869_);
  or (_19276_, _19275_, _19270_);
  and (_19277_, _03698_, _04562_);
  or (_19278_, _19277_, _19219_);
  or (_19279_, _19278_, _01870_);
  and (_19280_, _19279_, _19276_);
  or (_19281_, _19280_, _02079_);
  and (_19282_, _10614_, _03698_);
  or (_19283_, _19219_, _02166_);
  or (_19285_, _19283_, _19282_);
  and (_19286_, _19285_, _02912_);
  and (_19287_, _19286_, _19281_);
  or (_19288_, _19287_, _19222_);
  and (_19289_, _19288_, _02176_);
  nand (_19290_, _19278_, _02072_);
  nor (_19291_, _19290_, _19226_);
  or (_19292_, _19291_, _19289_);
  and (_19293_, _19292_, _02907_);
  or (_19294_, _19219_, _04106_);
  and (_19296_, _19231_, _02177_);
  and (_19297_, _19296_, _19294_);
  or (_19298_, _19297_, _02071_);
  or (_19299_, _19298_, _19293_);
  nor (_19300_, _10613_, _07909_);
  or (_19301_, _19219_, _04788_);
  or (_19302_, _19301_, _19300_);
  and (_19303_, _19302_, _04793_);
  and (_19304_, _19303_, _19299_);
  nor (_19305_, _10619_, _07909_);
  or (_19307_, _19305_, _19219_);
  and (_19308_, _19307_, _02173_);
  or (_19309_, _19308_, _02201_);
  or (_19310_, _19309_, _19304_);
  or (_19311_, _19227_, _02303_);
  and (_19312_, _19311_, _01887_);
  and (_19313_, _19312_, _19310_);
  and (_19314_, _19219_, _01860_);
  or (_19315_, _19314_, _01537_);
  or (_19316_, _19315_, _19313_);
  or (_19318_, _19227_, _01538_);
  and (_19319_, _19318_, _38087_);
  and (_19320_, _19319_, _19316_);
  or (_40241_, _19320_, _19217_);
  and (_19321_, _07909_, \oc8051_golden_model_1.P1 [1]);
  nor (_19322_, _07909_, _02811_);
  or (_19323_, _19322_, _19321_);
  or (_19324_, _19323_, _02840_);
  or (_19325_, _03698_, \oc8051_golden_model_1.P1 [1]);
  and (_19326_, _10698_, _03698_);
  not (_19329_, _19326_);
  and (_19330_, _19329_, _19325_);
  or (_19331_, _19330_, _02814_);
  nand (_19332_, _03698_, _01613_);
  and (_19333_, _19332_, _19325_);
  and (_19334_, _19333_, _02817_);
  and (_19335_, _02818_, \oc8051_golden_model_1.P1 [1]);
  or (_19336_, _19335_, _02001_);
  or (_19337_, _19336_, _19334_);
  and (_19338_, _19337_, _02024_);
  and (_19340_, _19338_, _19331_);
  and (_19341_, _07917_, \oc8051_golden_model_1.P1 [1]);
  and (_19342_, _10710_, _04336_);
  or (_19343_, _19342_, _19341_);
  and (_19344_, _19343_, _02007_);
  or (_19345_, _19344_, _01999_);
  or (_19346_, _19345_, _19340_);
  and (_19347_, _19346_, _19324_);
  or (_19348_, _19347_, _02006_);
  or (_19349_, _19333_, _02021_);
  and (_19352_, _19349_, _02025_);
  and (_19353_, _19352_, _19348_);
  and (_19354_, _10696_, _04336_);
  or (_19355_, _19354_, _19341_);
  and (_19356_, _19355_, _01997_);
  or (_19357_, _19356_, _01991_);
  or (_19358_, _19357_, _19353_);
  and (_19359_, _19342_, _10725_);
  or (_19360_, _19341_, _02861_);
  or (_19361_, _19360_, _19359_);
  and (_19363_, _19361_, _19358_);
  and (_19364_, _19363_, _02408_);
  and (_19365_, _18500_, _04336_);
  or (_19366_, _19341_, _19365_);
  and (_19367_, _19366_, _01875_);
  or (_19368_, _19367_, _05994_);
  or (_19369_, _19368_, _19364_);
  or (_19370_, _19323_, _05249_);
  and (_19371_, _19370_, _19369_);
  or (_19372_, _19371_, _02528_);
  and (_19375_, _04907_, _03698_);
  or (_19376_, _19321_, _02888_);
  or (_19377_, _19376_, _19375_);
  and (_19378_, _19377_, _02043_);
  and (_19379_, _19378_, _19372_);
  and (_19380_, _18528_, _03698_);
  or (_19381_, _19380_, _19321_);
  and (_19382_, _19381_, _01602_);
  or (_19383_, _19382_, _19379_);
  and (_19384_, _19383_, _01870_);
  nand (_19386_, _03698_, _02687_);
  and (_19387_, _19325_, _01869_);
  and (_19388_, _19387_, _19386_);
  or (_19389_, _19388_, _19384_);
  and (_19390_, _19389_, _02166_);
  or (_19391_, _10816_, _07909_);
  and (_19392_, _19325_, _02079_);
  and (_19393_, _19392_, _19391_);
  or (_19394_, _19393_, _19390_);
  and (_19395_, _19394_, _02912_);
  or (_19398_, _10822_, _07909_);
  and (_19399_, _19325_, _02167_);
  and (_19400_, _19399_, _19398_);
  or (_19401_, _19400_, _19395_);
  and (_19402_, _19401_, _02176_);
  or (_19403_, _10692_, _07909_);
  and (_19404_, _19325_, _02072_);
  and (_19405_, _19404_, _19403_);
  or (_19406_, _19405_, _19402_);
  and (_19407_, _19406_, _02907_);
  or (_19409_, _19321_, _04058_);
  and (_19410_, _19333_, _02177_);
  and (_19411_, _19410_, _19409_);
  or (_19412_, _19411_, _19407_);
  and (_19413_, _19412_, _02174_);
  or (_19414_, _19332_, _04058_);
  and (_19415_, _19325_, _02173_);
  and (_19416_, _19415_, _19414_);
  or (_19417_, _19416_, _02201_);
  or (_19418_, _19386_, _04058_);
  and (_19420_, _19325_, _02071_);
  and (_19421_, _19420_, _19418_);
  or (_19422_, _19421_, _19417_);
  or (_19423_, _19422_, _19413_);
  or (_19424_, _19330_, _02303_);
  and (_19425_, _19424_, _01887_);
  and (_19426_, _19425_, _19423_);
  and (_19427_, _19355_, _01860_);
  or (_19428_, _19427_, _01537_);
  or (_19429_, _19428_, _19426_);
  or (_19431_, _19321_, _01538_);
  or (_19432_, _19431_, _19326_);
  and (_19433_, _19432_, _38087_);
  and (_19434_, _19433_, _19429_);
  nor (_19435_, \oc8051_golden_model_1.P1 [1], rst);
  nor (_19436_, _19435_, _03183_);
  or (_40242_, _19436_, _19434_);
  and (_19437_, _07909_, \oc8051_golden_model_1.P1 [2]);
  and (_19438_, _11020_, _03698_);
  or (_19439_, _19438_, _19437_);
  and (_19441_, _19439_, _02167_);
  nor (_19442_, _07909_, _03455_);
  or (_19443_, _19442_, _19437_);
  or (_19444_, _19443_, _05249_);
  or (_19445_, _19443_, _02840_);
  nor (_19446_, _10905_, _07909_);
  or (_19447_, _19446_, _19437_);
  or (_19448_, _19447_, _02814_);
  and (_19449_, _03698_, \oc8051_golden_model_1.ACC [2]);
  or (_19450_, _19449_, _19437_);
  and (_19452_, _19450_, _02817_);
  and (_19453_, _02818_, \oc8051_golden_model_1.P1 [2]);
  or (_19454_, _19453_, _02001_);
  or (_19455_, _19454_, _19452_);
  and (_19456_, _19455_, _02024_);
  and (_19457_, _19456_, _19448_);
  and (_19458_, _07917_, \oc8051_golden_model_1.P1 [2]);
  and (_19459_, _10909_, _04336_);
  or (_19460_, _19459_, _19458_);
  and (_19461_, _19460_, _02007_);
  or (_19463_, _19461_, _01999_);
  or (_19464_, _19463_, _19457_);
  and (_19465_, _19464_, _19445_);
  or (_19466_, _19465_, _02006_);
  or (_19467_, _19450_, _02021_);
  and (_19468_, _19467_, _02025_);
  and (_19469_, _19468_, _19466_);
  and (_19470_, _10894_, _04336_);
  or (_19471_, _19470_, _19458_);
  and (_19472_, _19471_, _01997_);
  or (_19474_, _19472_, _01991_);
  or (_19475_, _19474_, _19469_);
  and (_19476_, _19459_, _10924_);
  or (_19477_, _19458_, _02861_);
  or (_19478_, _19477_, _19476_);
  and (_19479_, _19478_, _02408_);
  and (_19480_, _19479_, _19475_);
  and (_19481_, _18628_, _04336_);
  or (_19482_, _19481_, _19458_);
  and (_19483_, _19482_, _01875_);
  or (_19485_, _19483_, _05994_);
  or (_19486_, _19485_, _19480_);
  and (_19487_, _19486_, _19444_);
  or (_19488_, _19487_, _02528_);
  and (_19489_, _05043_, _03698_);
  or (_19490_, _19437_, _02888_);
  or (_19491_, _19490_, _19489_);
  and (_19492_, _19491_, _02043_);
  and (_19493_, _19492_, _19488_);
  and (_19494_, _18655_, _03698_);
  or (_19496_, _19494_, _19437_);
  and (_19497_, _19496_, _01602_);
  or (_19498_, _19497_, _01869_);
  or (_19499_, _19498_, _19493_);
  and (_19500_, _03698_, _04724_);
  or (_19501_, _19500_, _19437_);
  or (_19502_, _19501_, _01870_);
  and (_19503_, _19502_, _19499_);
  or (_19504_, _19503_, _02079_);
  and (_19505_, _11014_, _03698_);
  or (_19507_, _19437_, _02166_);
  or (_19508_, _19507_, _19505_);
  and (_19509_, _19508_, _02912_);
  and (_19510_, _19509_, _19504_);
  or (_19511_, _19510_, _19441_);
  and (_19512_, _19511_, _02176_);
  or (_19513_, _19437_, _04156_);
  and (_19514_, _19501_, _02072_);
  and (_19515_, _19514_, _19513_);
  or (_19516_, _19515_, _19512_);
  and (_19518_, _19516_, _02907_);
  and (_19519_, _19450_, _02177_);
  and (_19520_, _19519_, _19513_);
  or (_19521_, _19520_, _02071_);
  or (_19522_, _19521_, _19518_);
  nor (_19523_, _11013_, _07909_);
  or (_19524_, _19437_, _04788_);
  or (_19525_, _19524_, _19523_);
  and (_19526_, _19525_, _04793_);
  and (_19527_, _19526_, _19522_);
  nor (_19529_, _11019_, _07909_);
  or (_19530_, _19529_, _19437_);
  and (_19531_, _19530_, _02173_);
  or (_19532_, _19531_, _02201_);
  or (_19533_, _19532_, _19527_);
  or (_19534_, _19447_, _02303_);
  and (_19535_, _19534_, _01887_);
  and (_19536_, _19535_, _19533_);
  and (_19537_, _19471_, _01860_);
  or (_19538_, _19537_, _01537_);
  or (_19540_, _19538_, _19536_);
  and (_19541_, _11072_, _03698_);
  or (_19542_, _19437_, _01538_);
  or (_19543_, _19542_, _19541_);
  and (_19544_, _19543_, _38087_);
  and (_19545_, _19544_, _19540_);
  nor (_19546_, \oc8051_golden_model_1.P1 [2], rst);
  nor (_19547_, _19546_, _03183_);
  or (_40244_, _19547_, _19545_);
  and (_19548_, _07909_, \oc8051_golden_model_1.P1 [3]);
  and (_19550_, _11094_, _03698_);
  or (_19551_, _19550_, _19548_);
  and (_19552_, _19551_, _02167_);
  nor (_19553_, _07909_, _03268_);
  or (_19554_, _19553_, _19548_);
  or (_19555_, _19554_, _05249_);
  nor (_19556_, _11101_, _07909_);
  or (_19557_, _19556_, _19548_);
  or (_19558_, _19557_, _02814_);
  and (_19559_, _03698_, \oc8051_golden_model_1.ACC [3]);
  or (_19561_, _19559_, _19548_);
  and (_19562_, _19561_, _02817_);
  and (_19563_, _02818_, \oc8051_golden_model_1.P1 [3]);
  or (_19564_, _19563_, _02001_);
  or (_19565_, _19564_, _19562_);
  and (_19566_, _19565_, _02024_);
  and (_19567_, _19566_, _19558_);
  and (_19568_, _07917_, \oc8051_golden_model_1.P1 [3]);
  and (_19569_, _11098_, _04336_);
  or (_19570_, _19569_, _19568_);
  and (_19572_, _19570_, _02007_);
  or (_19573_, _19572_, _01999_);
  or (_19574_, _19573_, _19567_);
  or (_19575_, _19554_, _02840_);
  and (_19576_, _19575_, _19574_);
  or (_19577_, _19576_, _02006_);
  or (_19578_, _19561_, _02021_);
  and (_19579_, _19578_, _02025_);
  and (_19580_, _19579_, _19577_);
  and (_19581_, _11096_, _04336_);
  or (_19583_, _19581_, _19568_);
  and (_19584_, _19583_, _01997_);
  or (_19585_, _19584_, _01991_);
  or (_19586_, _19585_, _19580_);
  or (_19587_, _19568_, _11127_);
  and (_19588_, _19587_, _19570_);
  or (_19589_, _19588_, _02861_);
  and (_19590_, _19589_, _02408_);
  and (_19591_, _19590_, _19586_);
  and (_19592_, _18754_, _04336_);
  or (_19594_, _19592_, _19568_);
  and (_19595_, _19594_, _01875_);
  or (_19596_, _19595_, _05994_);
  or (_19597_, _19596_, _19591_);
  and (_19598_, _19597_, _19555_);
  or (_19599_, _19598_, _02528_);
  and (_19600_, _04998_, _03698_);
  or (_19601_, _19548_, _02888_);
  or (_19602_, _19601_, _19600_);
  and (_19603_, _19602_, _02043_);
  and (_19605_, _19603_, _19599_);
  and (_19606_, _18780_, _03698_);
  or (_19607_, _19606_, _19548_);
  and (_19608_, _19607_, _01602_);
  or (_19609_, _19608_, _01869_);
  or (_19610_, _19609_, _19605_);
  and (_19611_, _03698_, _04678_);
  or (_19612_, _19611_, _19548_);
  or (_19613_, _19612_, _01870_);
  and (_19614_, _19613_, _19610_);
  or (_19616_, _19614_, _02079_);
  and (_19617_, _11222_, _03698_);
  or (_19618_, _19548_, _02166_);
  or (_19619_, _19618_, _19617_);
  and (_19620_, _19619_, _02912_);
  and (_19621_, _19620_, _19616_);
  or (_19622_, _19621_, _19552_);
  and (_19623_, _19622_, _02176_);
  or (_19624_, _19548_, _04014_);
  and (_19625_, _19612_, _02072_);
  and (_19627_, _19625_, _19624_);
  or (_19628_, _19627_, _19623_);
  and (_19629_, _19628_, _02907_);
  and (_19630_, _19561_, _02177_);
  and (_19631_, _19630_, _19624_);
  or (_19632_, _19631_, _02071_);
  or (_19633_, _19632_, _19629_);
  nor (_19634_, _11220_, _07909_);
  or (_19635_, _19548_, _04788_);
  or (_19636_, _19635_, _19634_);
  and (_19638_, _19636_, _04793_);
  and (_19639_, _19638_, _19633_);
  nor (_19640_, _11093_, _07909_);
  or (_19641_, _19640_, _19548_);
  and (_19642_, _19641_, _02173_);
  or (_19643_, _19642_, _02201_);
  or (_19644_, _19643_, _19639_);
  or (_19645_, _19557_, _02303_);
  and (_19646_, _19645_, _01887_);
  and (_19647_, _19646_, _19644_);
  and (_19649_, _19583_, _01860_);
  or (_19650_, _19649_, _01537_);
  or (_19651_, _19650_, _19647_);
  and (_19652_, _11273_, _03698_);
  or (_19653_, _19548_, _01538_);
  or (_19654_, _19653_, _19652_);
  and (_19655_, _19654_, _38087_);
  and (_19656_, _19655_, _19651_);
  nor (_19657_, \oc8051_golden_model_1.P1 [3], rst);
  nor (_19658_, _19657_, _03183_);
  or (_40245_, _19658_, _19656_);
  and (_19660_, _07909_, \oc8051_golden_model_1.P1 [4]);
  and (_19661_, _11431_, _03698_);
  or (_19662_, _19661_, _19660_);
  and (_19663_, _19662_, _02167_);
  nor (_19664_, _04211_, _07909_);
  or (_19665_, _19664_, _19660_);
  or (_19666_, _19665_, _05249_);
  and (_19667_, _07917_, \oc8051_golden_model_1.P1 [4]);
  and (_19668_, _11301_, _04336_);
  or (_19670_, _19668_, _19667_);
  and (_19671_, _19670_, _01997_);
  nor (_19672_, _11317_, _07909_);
  or (_19673_, _19672_, _19660_);
  or (_19674_, _19673_, _02814_);
  and (_19675_, _03698_, \oc8051_golden_model_1.ACC [4]);
  or (_19676_, _19675_, _19660_);
  and (_19677_, _19676_, _02817_);
  and (_19678_, _02818_, \oc8051_golden_model_1.P1 [4]);
  or (_19679_, _19678_, _02001_);
  or (_19681_, _19679_, _19677_);
  and (_19682_, _19681_, _02024_);
  and (_19683_, _19682_, _19674_);
  and (_19684_, _11303_, _04336_);
  or (_19685_, _19684_, _19667_);
  and (_19686_, _19685_, _02007_);
  or (_19687_, _19686_, _01999_);
  or (_19688_, _19687_, _19683_);
  or (_19689_, _19665_, _02840_);
  and (_19690_, _19689_, _19688_);
  or (_19692_, _19690_, _02006_);
  or (_19693_, _19676_, _02021_);
  and (_19694_, _19693_, _02025_);
  and (_19695_, _19694_, _19692_);
  or (_19696_, _19695_, _19671_);
  and (_19697_, _19696_, _02861_);
  or (_19698_, _19667_, _11334_);
  and (_19699_, _19698_, _01991_);
  and (_19700_, _19699_, _19685_);
  or (_19701_, _19700_, _19697_);
  and (_19703_, _19701_, _02408_);
  and (_19704_, _18879_, _04336_);
  or (_19705_, _19704_, _19667_);
  and (_19706_, _19705_, _01875_);
  or (_19707_, _19706_, _05994_);
  or (_19708_, _19707_, _19703_);
  and (_19709_, _19708_, _19666_);
  or (_19710_, _19709_, _02528_);
  and (_19711_, _05135_, _03698_);
  or (_19712_, _19660_, _02888_);
  or (_19714_, _19712_, _19711_);
  and (_19715_, _19714_, _02043_);
  and (_19716_, _19715_, _19710_);
  and (_19717_, _18909_, _03698_);
  or (_19718_, _19717_, _19660_);
  and (_19719_, _19718_, _01602_);
  or (_19720_, _19719_, _01869_);
  or (_19721_, _19720_, _19716_);
  and (_19722_, _04694_, _03698_);
  or (_19723_, _19722_, _19660_);
  or (_19725_, _19723_, _01870_);
  and (_19726_, _19725_, _19721_);
  or (_19727_, _19726_, _02079_);
  and (_19728_, _11425_, _03698_);
  or (_19729_, _19660_, _02166_);
  or (_19730_, _19729_, _19728_);
  and (_19731_, _19730_, _02912_);
  and (_19732_, _19731_, _19727_);
  or (_19733_, _19732_, _19663_);
  and (_19734_, _19733_, _02176_);
  or (_19736_, _19660_, _04258_);
  and (_19737_, _19723_, _02072_);
  and (_19738_, _19737_, _19736_);
  or (_19739_, _19738_, _19734_);
  and (_19740_, _19739_, _02907_);
  and (_19741_, _19676_, _02177_);
  and (_19742_, _19741_, _19736_);
  or (_19743_, _19742_, _02071_);
  or (_19744_, _19743_, _19740_);
  nor (_19745_, _11424_, _07909_);
  or (_19747_, _19660_, _04788_);
  or (_19748_, _19747_, _19745_);
  and (_19749_, _19748_, _04793_);
  and (_19750_, _19749_, _19744_);
  nor (_19751_, _11430_, _07909_);
  or (_19752_, _19751_, _19660_);
  and (_19753_, _19752_, _02173_);
  or (_19754_, _19753_, _02201_);
  or (_19755_, _19754_, _19750_);
  or (_19756_, _19673_, _02303_);
  and (_19758_, _19756_, _01887_);
  and (_19759_, _19758_, _19755_);
  and (_19760_, _19670_, _01860_);
  or (_19761_, _19760_, _01537_);
  or (_19762_, _19761_, _19759_);
  and (_19763_, _11487_, _03698_);
  or (_19764_, _19660_, _01538_);
  or (_19765_, _19764_, _19763_);
  and (_19766_, _19765_, _38087_);
  and (_19767_, _19766_, _19762_);
  nor (_19769_, \oc8051_golden_model_1.P1 [4], rst);
  nor (_19770_, _19769_, _03183_);
  or (_40246_, _19770_, _19767_);
  and (_19771_, _07909_, \oc8051_golden_model_1.P1 [5]);
  and (_19772_, _11635_, _03698_);
  or (_19773_, _19772_, _19771_);
  and (_19774_, _19773_, _02167_);
  nor (_19775_, _11525_, _07909_);
  or (_19776_, _19775_, _19771_);
  or (_19777_, _19776_, _02814_);
  and (_19779_, _03698_, \oc8051_golden_model_1.ACC [5]);
  or (_19780_, _19779_, _19771_);
  and (_19781_, _19780_, _02817_);
  and (_19782_, _02818_, \oc8051_golden_model_1.P1 [5]);
  or (_19783_, _19782_, _02001_);
  or (_19784_, _19783_, _19781_);
  and (_19785_, _19784_, _02024_);
  and (_19786_, _19785_, _19777_);
  and (_19787_, _07917_, \oc8051_golden_model_1.P1 [5]);
  and (_19788_, _11510_, _04336_);
  or (_19790_, _19788_, _19787_);
  and (_19791_, _19790_, _02007_);
  or (_19792_, _19791_, _01999_);
  or (_19793_, _19792_, _19786_);
  nor (_19794_, _03916_, _07909_);
  or (_19795_, _19794_, _19771_);
  or (_19796_, _19795_, _02840_);
  and (_19797_, _19796_, _19793_);
  or (_19798_, _19797_, _02006_);
  or (_19799_, _19780_, _02021_);
  and (_19801_, _19799_, _02025_);
  and (_19802_, _19801_, _19798_);
  and (_19803_, _11508_, _04336_);
  or (_19804_, _19803_, _19787_);
  and (_19805_, _19804_, _01997_);
  or (_19806_, _19805_, _01991_);
  or (_19807_, _19806_, _19802_);
  or (_19808_, _19787_, _11542_);
  and (_19809_, _19808_, _19790_);
  or (_19810_, _19809_, _02861_);
  and (_19812_, _19810_, _02408_);
  and (_19813_, _19812_, _19807_);
  and (_19814_, _19009_, _04336_);
  or (_19815_, _19814_, _19787_);
  and (_19816_, _19815_, _01875_);
  or (_19817_, _19816_, _05994_);
  or (_19818_, _19817_, _19813_);
  or (_19819_, _19795_, _05249_);
  and (_19820_, _19819_, _19818_);
  or (_19821_, _19820_, _02528_);
  and (_19823_, _05090_, _03698_);
  or (_19824_, _19771_, _02888_);
  or (_19825_, _19824_, _19823_);
  and (_19826_, _19825_, _02043_);
  and (_19827_, _19826_, _19821_);
  and (_19828_, _19037_, _03698_);
  or (_19829_, _19828_, _19771_);
  and (_19830_, _19829_, _01602_);
  or (_19831_, _19830_, _01869_);
  or (_19832_, _19831_, _19827_);
  and (_19834_, _04672_, _03698_);
  or (_19835_, _19834_, _19771_);
  or (_19836_, _19835_, _01870_);
  and (_19837_, _19836_, _19832_);
  or (_19838_, _19837_, _02079_);
  and (_19839_, _11629_, _03698_);
  or (_19840_, _19771_, _02166_);
  or (_19841_, _19840_, _19839_);
  and (_19842_, _19841_, _02912_);
  and (_19843_, _19842_, _19838_);
  or (_19845_, _19843_, _19774_);
  and (_19846_, _19845_, _02176_);
  or (_19847_, _19771_, _03965_);
  and (_19848_, _19835_, _02072_);
  and (_19849_, _19848_, _19847_);
  or (_19850_, _19849_, _19846_);
  and (_19851_, _19850_, _02907_);
  and (_19852_, _19780_, _02177_);
  and (_19853_, _19852_, _19847_);
  or (_19854_, _19853_, _02071_);
  or (_19856_, _19854_, _19851_);
  nor (_19857_, _11628_, _07909_);
  or (_19858_, _19771_, _04788_);
  or (_19859_, _19858_, _19857_);
  and (_19860_, _19859_, _04793_);
  and (_19861_, _19860_, _19856_);
  nor (_19862_, _11634_, _07909_);
  or (_19863_, _19862_, _19771_);
  and (_19864_, _19863_, _02173_);
  or (_19865_, _19864_, _02201_);
  or (_19867_, _19865_, _19861_);
  or (_19868_, _19776_, _02303_);
  and (_19869_, _19868_, _01887_);
  and (_19870_, _19869_, _19867_);
  and (_19871_, _19804_, _01860_);
  or (_19872_, _19871_, _01537_);
  or (_19873_, _19872_, _19870_);
  and (_19874_, _11685_, _03698_);
  or (_19875_, _19771_, _01538_);
  or (_19876_, _19875_, _19874_);
  and (_19878_, _19876_, _38087_);
  and (_19879_, _19878_, _19873_);
  nor (_19880_, \oc8051_golden_model_1.P1 [5], rst);
  nor (_19881_, _19880_, _03183_);
  or (_40247_, _19881_, _19879_);
  nor (_19882_, \oc8051_golden_model_1.P1 [6], rst);
  nor (_19883_, _19882_, _03183_);
  and (_19884_, _07909_, \oc8051_golden_model_1.P1 [6]);
  and (_19885_, _11709_, _03698_);
  or (_19886_, _19885_, _19884_);
  and (_19888_, _19886_, _02167_);
  nor (_19889_, _11730_, _07909_);
  or (_19890_, _19889_, _19884_);
  or (_19891_, _19890_, _02814_);
  and (_19892_, _03698_, \oc8051_golden_model_1.ACC [6]);
  or (_19893_, _19892_, _19884_);
  and (_19894_, _19893_, _02817_);
  and (_19895_, _02818_, \oc8051_golden_model_1.P1 [6]);
  or (_19896_, _19895_, _02001_);
  or (_19897_, _19896_, _19894_);
  and (_19899_, _19897_, _02024_);
  and (_19900_, _19899_, _19891_);
  and (_19901_, _07917_, \oc8051_golden_model_1.P1 [6]);
  and (_19902_, _11717_, _04336_);
  or (_19903_, _19902_, _19901_);
  and (_19904_, _19903_, _02007_);
  or (_19905_, _19904_, _01999_);
  or (_19906_, _19905_, _19900_);
  nor (_19907_, _03808_, _07909_);
  or (_19908_, _19907_, _19884_);
  or (_19910_, _19908_, _02840_);
  and (_19911_, _19910_, _19906_);
  or (_19912_, _19911_, _02006_);
  or (_19913_, _19893_, _02021_);
  and (_19914_, _19913_, _02025_);
  and (_19915_, _19914_, _19912_);
  and (_19916_, _11715_, _04336_);
  or (_19917_, _19916_, _19901_);
  and (_19918_, _19917_, _01997_);
  or (_19919_, _19918_, _01991_);
  or (_19921_, _19919_, _19915_);
  or (_19922_, _19901_, _11747_);
  and (_19923_, _19922_, _19903_);
  or (_19924_, _19923_, _02861_);
  and (_19925_, _19924_, _02408_);
  and (_19926_, _19925_, _19921_);
  and (_19927_, _19133_, _04336_);
  or (_19928_, _19927_, _19901_);
  and (_19929_, _19928_, _01875_);
  or (_19930_, _19929_, _05994_);
  or (_19932_, _19930_, _19926_);
  or (_19933_, _19908_, _05249_);
  and (_19934_, _19933_, _19932_);
  or (_19935_, _19934_, _02528_);
  and (_19936_, _04861_, _03698_);
  or (_19937_, _19884_, _02888_);
  or (_19938_, _19937_, _19936_);
  and (_19939_, _19938_, _02043_);
  and (_19940_, _19939_, _19935_);
  and (_19941_, _19161_, _03698_);
  or (_19943_, _19941_, _19884_);
  and (_19944_, _19943_, _01602_);
  or (_19945_, _19944_, _01869_);
  or (_19946_, _19945_, _19940_);
  and (_19947_, _09920_, _03698_);
  or (_19948_, _19947_, _19884_);
  or (_19949_, _19948_, _01870_);
  and (_19950_, _19949_, _19946_);
  or (_19951_, _19950_, _02079_);
  and (_19952_, _11835_, _03698_);
  or (_19954_, _19884_, _02166_);
  or (_19955_, _19954_, _19952_);
  and (_19956_, _19955_, _02912_);
  and (_19957_, _19956_, _19951_);
  or (_19958_, _19957_, _19888_);
  and (_19959_, _19958_, _02176_);
  or (_19960_, _19884_, _03863_);
  and (_19961_, _19948_, _02072_);
  and (_19962_, _19961_, _19960_);
  or (_19963_, _19962_, _19959_);
  and (_19965_, _19963_, _02907_);
  and (_19966_, _19893_, _02177_);
  and (_19967_, _19966_, _19960_);
  or (_19968_, _19967_, _02071_);
  or (_19969_, _19968_, _19965_);
  nor (_19970_, _11833_, _07909_);
  or (_19971_, _19884_, _04788_);
  or (_19972_, _19971_, _19970_);
  and (_19973_, _19972_, _04793_);
  and (_19974_, _19973_, _19969_);
  nor (_19976_, _11708_, _07909_);
  or (_19977_, _19976_, _19884_);
  and (_19978_, _19977_, _02173_);
  or (_19979_, _19978_, _02201_);
  or (_19980_, _19979_, _19974_);
  or (_19981_, _19890_, _02303_);
  and (_19982_, _19981_, _01887_);
  and (_19983_, _19982_, _19980_);
  and (_19984_, _19917_, _01860_);
  or (_19985_, _19984_, _01537_);
  or (_19987_, _19985_, _19983_);
  and (_19988_, _11887_, _03698_);
  or (_19989_, _19884_, _01538_);
  or (_19990_, _19989_, _19988_);
  and (_19991_, _19990_, _38087_);
  and (_19992_, _19991_, _19987_);
  or (_40248_, _19992_, _19883_);
  and (_19993_, _08012_, \oc8051_golden_model_1.P2 [0]);
  and (_19994_, _10620_, _03665_);
  or (_19995_, _19994_, _19993_);
  and (_19997_, _19995_, _02167_);
  and (_19998_, _03665_, _03028_);
  or (_19999_, _19998_, _19993_);
  or (_20000_, _19999_, _05249_);
  nor (_20001_, _04106_, _08012_);
  or (_20002_, _20001_, _19993_);
  or (_20003_, _20002_, _02814_);
  and (_20004_, _03665_, \oc8051_golden_model_1.ACC [0]);
  or (_20005_, _20004_, _19993_);
  and (_20006_, _20005_, _02817_);
  and (_20008_, _02818_, \oc8051_golden_model_1.P2 [0]);
  or (_20009_, _20008_, _02001_);
  or (_20010_, _20009_, _20006_);
  and (_20011_, _20010_, _02024_);
  and (_20012_, _20011_, _20003_);
  and (_20013_, _08020_, \oc8051_golden_model_1.P2 [0]);
  and (_20014_, _10510_, _04342_);
  or (_20015_, _20014_, _20013_);
  and (_20016_, _20015_, _02007_);
  or (_20017_, _20016_, _20012_);
  and (_20019_, _20017_, _02840_);
  and (_20020_, _19999_, _01999_);
  or (_20021_, _20020_, _02006_);
  or (_20022_, _20021_, _20019_);
  or (_20023_, _20005_, _02021_);
  and (_20024_, _20023_, _02025_);
  and (_20025_, _20024_, _20022_);
  and (_20026_, _19993_, _01997_);
  or (_20027_, _20026_, _01991_);
  or (_20028_, _20027_, _20025_);
  or (_20030_, _20002_, _02861_);
  and (_20031_, _20030_, _02408_);
  and (_20032_, _20031_, _20028_);
  and (_20033_, _18380_, _04342_);
  or (_20034_, _20033_, _20013_);
  and (_20035_, _20034_, _01875_);
  or (_20036_, _20035_, _05994_);
  or (_20037_, _20036_, _20032_);
  and (_20038_, _20037_, _20000_);
  or (_20039_, _20038_, _02528_);
  and (_20041_, _04952_, _03665_);
  or (_20042_, _19993_, _02888_);
  or (_20043_, _20042_, _20041_);
  and (_20044_, _20043_, _02043_);
  and (_20045_, _20044_, _20039_);
  and (_20046_, _18407_, _03665_);
  or (_20047_, _20046_, _19993_);
  and (_20048_, _20047_, _01602_);
  or (_20049_, _20048_, _01869_);
  or (_20050_, _20049_, _20045_);
  and (_20052_, _03665_, _04562_);
  or (_20053_, _20052_, _19993_);
  or (_20054_, _20053_, _01870_);
  and (_20055_, _20054_, _20050_);
  or (_20056_, _20055_, _02079_);
  and (_20057_, _10614_, _03665_);
  or (_20058_, _19993_, _02166_);
  or (_20059_, _20058_, _20057_);
  and (_20060_, _20059_, _02912_);
  and (_20061_, _20060_, _20056_);
  or (_20063_, _20061_, _19997_);
  and (_20064_, _20063_, _02176_);
  nand (_20065_, _20053_, _02072_);
  nor (_20066_, _20065_, _20001_);
  or (_20067_, _20066_, _20064_);
  and (_20068_, _20067_, _02907_);
  or (_20069_, _19993_, _04106_);
  and (_20070_, _20005_, _02177_);
  and (_20071_, _20070_, _20069_);
  or (_20072_, _20071_, _02071_);
  or (_20074_, _20072_, _20068_);
  nor (_20075_, _10613_, _08012_);
  or (_20076_, _19993_, _04788_);
  or (_20077_, _20076_, _20075_);
  and (_20078_, _20077_, _04793_);
  and (_20079_, _20078_, _20074_);
  nor (_20080_, _10619_, _08012_);
  or (_20081_, _20080_, _19993_);
  and (_20082_, _20081_, _02173_);
  or (_20083_, _20082_, _02201_);
  or (_20085_, _20083_, _20079_);
  or (_20086_, _20002_, _02303_);
  and (_20087_, _20086_, _01887_);
  and (_20088_, _20087_, _20085_);
  and (_20089_, _19993_, _01860_);
  or (_20090_, _20089_, _01537_);
  or (_20091_, _20090_, _20088_);
  or (_20092_, _20002_, _01538_);
  and (_20093_, _20092_, _38087_);
  and (_20094_, _20093_, _20091_);
  nor (_20096_, \oc8051_golden_model_1.P2 [0], rst);
  nor (_20097_, _20096_, _03183_);
  or (_40250_, _20097_, _20094_);
  nor (_20098_, \oc8051_golden_model_1.P2 [1], rst);
  nor (_20099_, _20098_, _03183_);
  and (_20100_, _08012_, \oc8051_golden_model_1.P2 [1]);
  nor (_20101_, _08012_, _02811_);
  or (_20102_, _20101_, _20100_);
  or (_20103_, _20102_, _02840_);
  or (_20104_, _03665_, \oc8051_golden_model_1.P2 [1]);
  and (_20106_, _10698_, _03665_);
  not (_20107_, _20106_);
  and (_20108_, _20107_, _20104_);
  or (_20109_, _20108_, _02814_);
  nand (_20110_, _03665_, _01613_);
  and (_20111_, _20110_, _20104_);
  and (_20112_, _20111_, _02817_);
  and (_20113_, _02818_, \oc8051_golden_model_1.P2 [1]);
  or (_20114_, _20113_, _02001_);
  or (_20115_, _20114_, _20112_);
  and (_20117_, _20115_, _02024_);
  and (_20118_, _20117_, _20109_);
  and (_20119_, _08020_, \oc8051_golden_model_1.P2 [1]);
  and (_20120_, _10710_, _04342_);
  or (_20121_, _20120_, _20119_);
  and (_20122_, _20121_, _02007_);
  or (_20123_, _20122_, _01999_);
  or (_20124_, _20123_, _20118_);
  and (_20125_, _20124_, _20103_);
  or (_20126_, _20125_, _02006_);
  or (_20128_, _20111_, _02021_);
  and (_20129_, _20128_, _02025_);
  and (_20130_, _20129_, _20126_);
  and (_20131_, _10696_, _04342_);
  or (_20132_, _20131_, _20119_);
  and (_20133_, _20132_, _01997_);
  or (_20134_, _20133_, _01991_);
  or (_20135_, _20134_, _20130_);
  and (_20136_, _20120_, _10725_);
  or (_20137_, _20119_, _02861_);
  or (_20139_, _20137_, _20136_);
  and (_20140_, _20139_, _20135_);
  and (_20141_, _20140_, _02408_);
  and (_20142_, _18500_, _04342_);
  or (_20143_, _20119_, _20142_);
  and (_20144_, _20143_, _01875_);
  or (_20145_, _20144_, _05994_);
  or (_20146_, _20145_, _20141_);
  or (_20147_, _20102_, _05249_);
  and (_20148_, _20147_, _20146_);
  or (_20150_, _20148_, _02528_);
  and (_20151_, _04907_, _03665_);
  or (_20152_, _20100_, _02888_);
  or (_20153_, _20152_, _20151_);
  and (_20154_, _20153_, _02043_);
  and (_20155_, _20154_, _20150_);
  and (_20156_, _18528_, _03665_);
  or (_20157_, _20156_, _20100_);
  and (_20158_, _20157_, _01602_);
  or (_20159_, _20158_, _20155_);
  and (_20161_, _20159_, _01870_);
  nand (_20162_, _03665_, _02687_);
  and (_20163_, _20104_, _01869_);
  and (_20164_, _20163_, _20162_);
  or (_20165_, _20164_, _20161_);
  and (_20166_, _20165_, _02166_);
  or (_20167_, _10816_, _08012_);
  and (_20168_, _20104_, _02079_);
  and (_20169_, _20168_, _20167_);
  or (_20170_, _20169_, _20166_);
  and (_20172_, _20170_, _02912_);
  or (_20173_, _10822_, _08012_);
  and (_20174_, _20104_, _02167_);
  and (_20175_, _20174_, _20173_);
  or (_20176_, _20175_, _20172_);
  and (_20177_, _20176_, _02176_);
  or (_20178_, _10692_, _08012_);
  and (_20179_, _20104_, _02072_);
  and (_20180_, _20179_, _20178_);
  or (_20181_, _20180_, _20177_);
  and (_20183_, _20181_, _02907_);
  or (_20184_, _20100_, _04058_);
  and (_20185_, _20111_, _02177_);
  and (_20186_, _20185_, _20184_);
  or (_20187_, _20186_, _20183_);
  and (_20188_, _20187_, _02174_);
  or (_20189_, _20110_, _04058_);
  and (_20190_, _20104_, _02173_);
  and (_20191_, _20190_, _20189_);
  or (_20192_, _20191_, _02201_);
  or (_20194_, _20162_, _04058_);
  and (_20195_, _20104_, _02071_);
  and (_20196_, _20195_, _20194_);
  or (_20197_, _20196_, _20192_);
  or (_20198_, _20197_, _20188_);
  or (_20199_, _20108_, _02303_);
  and (_20200_, _20199_, _01887_);
  and (_20201_, _20200_, _20198_);
  and (_20202_, _20132_, _01860_);
  or (_20203_, _20202_, _01537_);
  or (_20205_, _20203_, _20201_);
  or (_20206_, _20100_, _01538_);
  or (_20207_, _20206_, _20106_);
  and (_20208_, _20207_, _38087_);
  and (_20209_, _20208_, _20205_);
  or (_40251_, _20209_, _20099_);
  and (_20210_, _08012_, \oc8051_golden_model_1.P2 [2]);
  and (_20211_, _11020_, _03665_);
  or (_20212_, _20211_, _20210_);
  and (_20213_, _20212_, _02167_);
  nor (_20215_, _08012_, _03455_);
  or (_20216_, _20215_, _20210_);
  or (_20217_, _20216_, _05249_);
  or (_20218_, _20216_, _02840_);
  nor (_20219_, _10905_, _08012_);
  or (_20220_, _20219_, _20210_);
  or (_20221_, _20220_, _02814_);
  and (_20222_, _03665_, \oc8051_golden_model_1.ACC [2]);
  or (_20223_, _20222_, _20210_);
  and (_20224_, _20223_, _02817_);
  and (_20226_, _02818_, \oc8051_golden_model_1.P2 [2]);
  or (_20227_, _20226_, _02001_);
  or (_20228_, _20227_, _20224_);
  and (_20229_, _20228_, _02024_);
  and (_20230_, _20229_, _20221_);
  and (_20231_, _08020_, \oc8051_golden_model_1.P2 [2]);
  and (_20232_, _10909_, _04342_);
  or (_20233_, _20232_, _20231_);
  and (_20234_, _20233_, _02007_);
  or (_20235_, _20234_, _01999_);
  or (_20237_, _20235_, _20230_);
  and (_20238_, _20237_, _20218_);
  or (_20239_, _20238_, _02006_);
  or (_20240_, _20223_, _02021_);
  and (_20241_, _20240_, _02025_);
  and (_20242_, _20241_, _20239_);
  and (_20243_, _10894_, _04342_);
  or (_20244_, _20243_, _20231_);
  and (_20245_, _20244_, _01997_);
  or (_20246_, _20245_, _01991_);
  or (_20248_, _20246_, _20242_);
  and (_20249_, _20232_, _10924_);
  or (_20250_, _20231_, _02861_);
  or (_20251_, _20250_, _20249_);
  and (_20252_, _20251_, _02408_);
  and (_20253_, _20252_, _20248_);
  and (_20254_, _18628_, _04342_);
  or (_20255_, _20254_, _20231_);
  and (_20256_, _20255_, _01875_);
  or (_20257_, _20256_, _05994_);
  or (_20259_, _20257_, _20253_);
  and (_20260_, _20259_, _20217_);
  or (_20261_, _20260_, _02528_);
  and (_20262_, _05043_, _03665_);
  or (_20263_, _20210_, _02888_);
  or (_20264_, _20263_, _20262_);
  and (_20265_, _20264_, _02043_);
  and (_20266_, _20265_, _20261_);
  and (_20267_, _18655_, _03665_);
  or (_20268_, _20267_, _20210_);
  and (_20270_, _20268_, _01602_);
  or (_20271_, _20270_, _01869_);
  or (_20272_, _20271_, _20266_);
  and (_20273_, _03665_, _04724_);
  or (_20274_, _20273_, _20210_);
  or (_20275_, _20274_, _01870_);
  and (_20276_, _20275_, _20272_);
  or (_20277_, _20276_, _02079_);
  and (_20278_, _11014_, _03665_);
  or (_20279_, _20210_, _02166_);
  or (_20281_, _20279_, _20278_);
  and (_20282_, _20281_, _02912_);
  and (_20283_, _20282_, _20277_);
  or (_20284_, _20283_, _20213_);
  and (_20285_, _20284_, _02176_);
  or (_20286_, _20210_, _04156_);
  and (_20287_, _20274_, _02072_);
  and (_20288_, _20287_, _20286_);
  or (_20289_, _20288_, _20285_);
  and (_20290_, _20289_, _02907_);
  and (_20292_, _20223_, _02177_);
  and (_20293_, _20292_, _20286_);
  or (_20294_, _20293_, _02071_);
  or (_20295_, _20294_, _20290_);
  nor (_20296_, _11013_, _08012_);
  or (_20297_, _20210_, _04788_);
  or (_20298_, _20297_, _20296_);
  and (_20299_, _20298_, _04793_);
  and (_20300_, _20299_, _20295_);
  nor (_20301_, _11019_, _08012_);
  or (_20303_, _20301_, _20210_);
  and (_20304_, _20303_, _02173_);
  or (_20305_, _20304_, _02201_);
  or (_20306_, _20305_, _20300_);
  or (_20307_, _20220_, _02303_);
  and (_20308_, _20307_, _01887_);
  and (_20309_, _20308_, _20306_);
  and (_20310_, _20244_, _01860_);
  or (_20311_, _20310_, _01537_);
  or (_20312_, _20311_, _20309_);
  and (_20314_, _11072_, _03665_);
  or (_20315_, _20210_, _01538_);
  or (_20316_, _20315_, _20314_);
  and (_20317_, _20316_, _38087_);
  and (_20318_, _20317_, _20312_);
  nor (_20319_, \oc8051_golden_model_1.P2 [2], rst);
  nor (_20320_, _20319_, _03183_);
  or (_40252_, _20320_, _20318_);
  and (_20321_, _08012_, \oc8051_golden_model_1.P2 [3]);
  and (_20322_, _11094_, _03665_);
  or (_20324_, _20322_, _20321_);
  and (_20325_, _20324_, _02167_);
  nor (_20326_, _08012_, _03268_);
  or (_20327_, _20326_, _20321_);
  or (_20328_, _20327_, _05249_);
  nor (_20329_, _11101_, _08012_);
  or (_20330_, _20329_, _20321_);
  or (_20331_, _20330_, _02814_);
  and (_20332_, _03665_, \oc8051_golden_model_1.ACC [3]);
  or (_20333_, _20332_, _20321_);
  and (_20335_, _20333_, _02817_);
  and (_20336_, _02818_, \oc8051_golden_model_1.P2 [3]);
  or (_20337_, _20336_, _02001_);
  or (_20338_, _20337_, _20335_);
  and (_20339_, _20338_, _02024_);
  and (_20340_, _20339_, _20331_);
  and (_20341_, _08020_, \oc8051_golden_model_1.P2 [3]);
  and (_20342_, _11098_, _04342_);
  or (_20343_, _20342_, _20341_);
  and (_20344_, _20343_, _02007_);
  or (_20346_, _20344_, _01999_);
  or (_20347_, _20346_, _20340_);
  or (_20348_, _20327_, _02840_);
  and (_20349_, _20348_, _20347_);
  or (_20350_, _20349_, _02006_);
  or (_20351_, _20333_, _02021_);
  and (_20352_, _20351_, _02025_);
  and (_20353_, _20352_, _20350_);
  and (_20354_, _11096_, _04342_);
  or (_20355_, _20354_, _20341_);
  and (_20357_, _20355_, _01997_);
  or (_20358_, _20357_, _01991_);
  or (_20359_, _20358_, _20353_);
  or (_20360_, _20341_, _11127_);
  and (_20361_, _20360_, _20343_);
  or (_20362_, _20361_, _02861_);
  and (_20363_, _20362_, _02408_);
  and (_20364_, _20363_, _20359_);
  and (_20365_, _18754_, _04342_);
  or (_20366_, _20365_, _20341_);
  and (_20368_, _20366_, _01875_);
  or (_20369_, _20368_, _05994_);
  or (_20370_, _20369_, _20364_);
  and (_20371_, _20370_, _20328_);
  or (_20372_, _20371_, _02528_);
  and (_20373_, _04998_, _03665_);
  or (_20374_, _20321_, _02888_);
  or (_20375_, _20374_, _20373_);
  and (_20376_, _20375_, _02043_);
  and (_20377_, _20376_, _20372_);
  and (_20379_, _18780_, _03665_);
  or (_20380_, _20379_, _20321_);
  and (_20381_, _20380_, _01602_);
  or (_20382_, _20381_, _01869_);
  or (_20383_, _20382_, _20377_);
  and (_20384_, _03665_, _04678_);
  or (_20385_, _20384_, _20321_);
  or (_20386_, _20385_, _01870_);
  and (_20387_, _20386_, _20383_);
  or (_20388_, _20387_, _02079_);
  and (_20390_, _11222_, _03665_);
  or (_20391_, _20321_, _02166_);
  or (_20392_, _20391_, _20390_);
  and (_20393_, _20392_, _02912_);
  and (_20394_, _20393_, _20388_);
  or (_20395_, _20394_, _20325_);
  and (_20396_, _20395_, _02176_);
  or (_20397_, _20321_, _04014_);
  and (_20398_, _20385_, _02072_);
  and (_20399_, _20398_, _20397_);
  or (_20401_, _20399_, _20396_);
  and (_20402_, _20401_, _02907_);
  and (_20403_, _20333_, _02177_);
  and (_20404_, _20403_, _20397_);
  or (_20405_, _20404_, _02071_);
  or (_20406_, _20405_, _20402_);
  nor (_20407_, _11220_, _08012_);
  or (_20408_, _20321_, _04788_);
  or (_20409_, _20408_, _20407_);
  and (_20410_, _20409_, _04793_);
  and (_20412_, _20410_, _20406_);
  nor (_20413_, _11093_, _08012_);
  or (_20414_, _20413_, _20321_);
  and (_20415_, _20414_, _02173_);
  or (_20416_, _20415_, _02201_);
  or (_20417_, _20416_, _20412_);
  or (_20418_, _20330_, _02303_);
  and (_20419_, _20418_, _01887_);
  and (_20420_, _20419_, _20417_);
  and (_20421_, _20355_, _01860_);
  or (_20423_, _20421_, _01537_);
  or (_20424_, _20423_, _20420_);
  and (_20425_, _11273_, _03665_);
  or (_20426_, _20321_, _01538_);
  or (_20427_, _20426_, _20425_);
  and (_20428_, _20427_, _38087_);
  and (_20429_, _20428_, _20424_);
  nor (_20430_, \oc8051_golden_model_1.P2 [3], rst);
  nor (_20431_, _20430_, _03183_);
  or (_40253_, _20431_, _20429_);
  and (_20433_, _08012_, \oc8051_golden_model_1.P2 [4]);
  and (_20434_, _11431_, _03665_);
  or (_20435_, _20434_, _20433_);
  and (_20436_, _20435_, _02167_);
  nor (_20437_, _04211_, _08012_);
  or (_20438_, _20437_, _20433_);
  or (_20439_, _20438_, _05249_);
  and (_20440_, _08020_, \oc8051_golden_model_1.P2 [4]);
  and (_20441_, _11301_, _04342_);
  or (_20442_, _20441_, _20440_);
  and (_20444_, _20442_, _01997_);
  nor (_20445_, _11317_, _08012_);
  or (_20446_, _20445_, _20433_);
  or (_20447_, _20446_, _02814_);
  and (_20448_, _03665_, \oc8051_golden_model_1.ACC [4]);
  or (_20449_, _20448_, _20433_);
  and (_20450_, _20449_, _02817_);
  and (_20451_, _02818_, \oc8051_golden_model_1.P2 [4]);
  or (_20452_, _20451_, _02001_);
  or (_20453_, _20452_, _20450_);
  and (_20455_, _20453_, _02024_);
  and (_20456_, _20455_, _20447_);
  and (_20457_, _11303_, _04342_);
  or (_20458_, _20457_, _20440_);
  and (_20459_, _20458_, _02007_);
  or (_20460_, _20459_, _01999_);
  or (_20461_, _20460_, _20456_);
  or (_20462_, _20438_, _02840_);
  and (_20463_, _20462_, _20461_);
  or (_20464_, _20463_, _02006_);
  or (_20466_, _20449_, _02021_);
  and (_20467_, _20466_, _02025_);
  and (_20468_, _20467_, _20464_);
  or (_20469_, _20468_, _20444_);
  and (_20470_, _20469_, _02861_);
  or (_20471_, _20440_, _11334_);
  and (_20472_, _20471_, _01991_);
  and (_20473_, _20472_, _20458_);
  or (_20474_, _20473_, _20470_);
  and (_20475_, _20474_, _02408_);
  and (_20477_, _18879_, _04342_);
  or (_20478_, _20477_, _20440_);
  and (_20479_, _20478_, _01875_);
  or (_20480_, _20479_, _05994_);
  or (_20481_, _20480_, _20475_);
  and (_20482_, _20481_, _20439_);
  or (_20483_, _20482_, _02528_);
  and (_20484_, _05135_, _03665_);
  or (_20485_, _20433_, _02888_);
  or (_20486_, _20485_, _20484_);
  and (_20488_, _20486_, _02043_);
  and (_20489_, _20488_, _20483_);
  and (_20490_, _18909_, _03665_);
  or (_20491_, _20490_, _20433_);
  and (_20492_, _20491_, _01602_);
  or (_20493_, _20492_, _01869_);
  or (_20494_, _20493_, _20489_);
  and (_20495_, _04694_, _03665_);
  or (_20496_, _20495_, _20433_);
  or (_20497_, _20496_, _01870_);
  and (_20499_, _20497_, _20494_);
  or (_20500_, _20499_, _02079_);
  and (_20501_, _11425_, _03665_);
  or (_20502_, _20433_, _02166_);
  or (_20503_, _20502_, _20501_);
  and (_20504_, _20503_, _02912_);
  and (_20505_, _20504_, _20500_);
  or (_20506_, _20505_, _20436_);
  and (_20507_, _20506_, _02176_);
  or (_20508_, _20433_, _04258_);
  and (_20510_, _20496_, _02072_);
  and (_20511_, _20510_, _20508_);
  or (_20512_, _20511_, _20507_);
  and (_20513_, _20512_, _02907_);
  and (_20514_, _20449_, _02177_);
  and (_20515_, _20514_, _20508_);
  or (_20516_, _20515_, _02071_);
  or (_20517_, _20516_, _20513_);
  nor (_20518_, _11424_, _08012_);
  or (_20519_, _20433_, _04788_);
  or (_20521_, _20519_, _20518_);
  and (_20522_, _20521_, _04793_);
  and (_20523_, _20522_, _20517_);
  nor (_20524_, _11430_, _08012_);
  or (_20525_, _20524_, _20433_);
  and (_20526_, _20525_, _02173_);
  or (_20527_, _20526_, _02201_);
  or (_20528_, _20527_, _20523_);
  or (_20529_, _20446_, _02303_);
  and (_20530_, _20529_, _01887_);
  and (_20532_, _20530_, _20528_);
  and (_20533_, _20442_, _01860_);
  or (_20534_, _20533_, _01537_);
  or (_20535_, _20534_, _20532_);
  and (_20536_, _11487_, _03665_);
  or (_20537_, _20433_, _01538_);
  or (_20538_, _20537_, _20536_);
  and (_20539_, _20538_, _38087_);
  and (_20540_, _20539_, _20535_);
  nor (_20541_, \oc8051_golden_model_1.P2 [4], rst);
  nor (_20543_, _20541_, _03183_);
  or (_40254_, _20543_, _20540_);
  nor (_20544_, \oc8051_golden_model_1.P2 [5], rst);
  nor (_20545_, _20544_, _03183_);
  and (_20546_, _08012_, \oc8051_golden_model_1.P2 [5]);
  and (_20547_, _11635_, _03665_);
  or (_20548_, _20547_, _20546_);
  and (_20549_, _20548_, _02167_);
  nor (_20550_, _11525_, _08012_);
  or (_20551_, _20550_, _20546_);
  or (_20553_, _20551_, _02814_);
  and (_20554_, _03665_, \oc8051_golden_model_1.ACC [5]);
  or (_20555_, _20554_, _20546_);
  and (_20556_, _20555_, _02817_);
  and (_20557_, _02818_, \oc8051_golden_model_1.P2 [5]);
  or (_20558_, _20557_, _02001_);
  or (_20559_, _20558_, _20556_);
  and (_20560_, _20559_, _02024_);
  and (_20561_, _20560_, _20553_);
  and (_20562_, _08020_, \oc8051_golden_model_1.P2 [5]);
  and (_20564_, _11510_, _04342_);
  or (_20565_, _20564_, _20562_);
  and (_20566_, _20565_, _02007_);
  or (_20567_, _20566_, _01999_);
  or (_20568_, _20567_, _20561_);
  nor (_20569_, _03916_, _08012_);
  or (_20570_, _20569_, _20546_);
  or (_20571_, _20570_, _02840_);
  and (_20572_, _20571_, _20568_);
  or (_20573_, _20572_, _02006_);
  or (_20575_, _20555_, _02021_);
  and (_20576_, _20575_, _02025_);
  and (_20577_, _20576_, _20573_);
  and (_20578_, _11508_, _04342_);
  or (_20579_, _20578_, _20562_);
  and (_20580_, _20579_, _01997_);
  or (_20581_, _20580_, _01991_);
  or (_20582_, _20581_, _20577_);
  or (_20583_, _20562_, _11542_);
  and (_20584_, _20583_, _20565_);
  or (_20586_, _20584_, _02861_);
  and (_20587_, _20586_, _02408_);
  and (_20588_, _20587_, _20582_);
  and (_20589_, _19009_, _04342_);
  or (_20590_, _20589_, _20562_);
  and (_20591_, _20590_, _01875_);
  or (_20592_, _20591_, _05994_);
  or (_20593_, _20592_, _20588_);
  or (_20594_, _20570_, _05249_);
  and (_20595_, _20594_, _20593_);
  or (_20597_, _20595_, _02528_);
  and (_20598_, _05090_, _03665_);
  or (_20599_, _20546_, _02888_);
  or (_20600_, _20599_, _20598_);
  and (_20601_, _20600_, _02043_);
  and (_20602_, _20601_, _20597_);
  and (_20603_, _19037_, _03665_);
  or (_20604_, _20603_, _20546_);
  and (_20605_, _20604_, _01602_);
  or (_20606_, _20605_, _01869_);
  or (_20608_, _20606_, _20602_);
  and (_20609_, _04672_, _03665_);
  or (_20610_, _20609_, _20546_);
  or (_20611_, _20610_, _01870_);
  and (_20612_, _20611_, _20608_);
  or (_20613_, _20612_, _02079_);
  and (_20614_, _11629_, _03665_);
  or (_20615_, _20546_, _02166_);
  or (_20616_, _20615_, _20614_);
  and (_20617_, _20616_, _02912_);
  and (_20619_, _20617_, _20613_);
  or (_20620_, _20619_, _20549_);
  and (_20621_, _20620_, _02176_);
  or (_20622_, _20546_, _03965_);
  and (_20623_, _20610_, _02072_);
  and (_20624_, _20623_, _20622_);
  or (_20625_, _20624_, _20621_);
  and (_20626_, _20625_, _02907_);
  and (_20627_, _20555_, _02177_);
  and (_20628_, _20627_, _20622_);
  or (_20630_, _20628_, _02071_);
  or (_20631_, _20630_, _20626_);
  nor (_20632_, _11628_, _08012_);
  or (_20633_, _20546_, _04788_);
  or (_20634_, _20633_, _20632_);
  and (_20635_, _20634_, _04793_);
  and (_20636_, _20635_, _20631_);
  nor (_20637_, _11634_, _08012_);
  or (_20638_, _20637_, _20546_);
  and (_20639_, _20638_, _02173_);
  or (_20641_, _20639_, _02201_);
  or (_20642_, _20641_, _20636_);
  or (_20643_, _20551_, _02303_);
  and (_20644_, _20643_, _01887_);
  and (_20645_, _20644_, _20642_);
  and (_20646_, _20579_, _01860_);
  or (_20647_, _20646_, _01537_);
  or (_20648_, _20647_, _20645_);
  and (_20649_, _11685_, _03665_);
  or (_20650_, _20546_, _01538_);
  or (_20652_, _20650_, _20649_);
  and (_20653_, _20652_, _38087_);
  and (_20654_, _20653_, _20648_);
  or (_40255_, _20654_, _20545_);
  and (_20655_, _08012_, \oc8051_golden_model_1.P2 [6]);
  and (_20656_, _11709_, _03665_);
  or (_20657_, _20656_, _20655_);
  and (_20658_, _20657_, _02167_);
  nor (_20659_, _11730_, _08012_);
  or (_20660_, _20659_, _20655_);
  or (_20662_, _20660_, _02814_);
  and (_20663_, _03665_, \oc8051_golden_model_1.ACC [6]);
  or (_20664_, _20663_, _20655_);
  and (_20665_, _20664_, _02817_);
  and (_20666_, _02818_, \oc8051_golden_model_1.P2 [6]);
  or (_20667_, _20666_, _02001_);
  or (_20668_, _20667_, _20665_);
  and (_20669_, _20668_, _02024_);
  and (_20670_, _20669_, _20662_);
  and (_20671_, _08020_, \oc8051_golden_model_1.P2 [6]);
  and (_20673_, _11717_, _04342_);
  or (_20674_, _20673_, _20671_);
  and (_20675_, _20674_, _02007_);
  or (_20676_, _20675_, _01999_);
  or (_20677_, _20676_, _20670_);
  nor (_20678_, _03808_, _08012_);
  or (_20679_, _20678_, _20655_);
  or (_20680_, _20679_, _02840_);
  and (_20681_, _20680_, _20677_);
  or (_20682_, _20681_, _02006_);
  or (_20684_, _20664_, _02021_);
  and (_20685_, _20684_, _02025_);
  and (_20686_, _20685_, _20682_);
  and (_20687_, _11715_, _04342_);
  or (_20688_, _20687_, _20671_);
  and (_20689_, _20688_, _01997_);
  or (_20690_, _20689_, _01991_);
  or (_20691_, _20690_, _20686_);
  or (_20692_, _20671_, _11747_);
  and (_20693_, _20692_, _20674_);
  or (_20695_, _20693_, _02861_);
  and (_20696_, _20695_, _02408_);
  and (_20697_, _20696_, _20691_);
  and (_20698_, _19133_, _04342_);
  or (_20699_, _20698_, _20671_);
  and (_20700_, _20699_, _01875_);
  or (_20701_, _20700_, _05994_);
  or (_20702_, _20701_, _20697_);
  or (_20703_, _20679_, _05249_);
  and (_20704_, _20703_, _20702_);
  or (_20706_, _20704_, _02528_);
  and (_20707_, _04861_, _03665_);
  or (_20708_, _20655_, _02888_);
  or (_20709_, _20708_, _20707_);
  and (_20710_, _20709_, _02043_);
  and (_20711_, _20710_, _20706_);
  and (_20712_, _19161_, _03665_);
  or (_20713_, _20712_, _20655_);
  and (_20714_, _20713_, _01602_);
  or (_20715_, _20714_, _01869_);
  or (_20717_, _20715_, _20711_);
  and (_20718_, _09920_, _03665_);
  or (_20719_, _20718_, _20655_);
  or (_20720_, _20719_, _01870_);
  and (_20721_, _20720_, _20717_);
  or (_20722_, _20721_, _02079_);
  and (_20723_, _11835_, _03665_);
  or (_20724_, _20655_, _02166_);
  or (_20725_, _20724_, _20723_);
  and (_20726_, _20725_, _02912_);
  and (_20728_, _20726_, _20722_);
  or (_20729_, _20728_, _20658_);
  and (_20730_, _20729_, _02176_);
  or (_20731_, _20655_, _03863_);
  and (_20732_, _20719_, _02072_);
  and (_20733_, _20732_, _20731_);
  or (_20734_, _20733_, _20730_);
  and (_20735_, _20734_, _02907_);
  and (_20736_, _20664_, _02177_);
  and (_20737_, _20736_, _20731_);
  or (_20739_, _20737_, _02071_);
  or (_20740_, _20739_, _20735_);
  nor (_20741_, _11833_, _08012_);
  or (_20742_, _20655_, _04788_);
  or (_20743_, _20742_, _20741_);
  and (_20744_, _20743_, _04793_);
  and (_20745_, _20744_, _20740_);
  nor (_20746_, _11708_, _08012_);
  or (_20747_, _20746_, _20655_);
  and (_20748_, _20747_, _02173_);
  or (_20750_, _20748_, _02201_);
  or (_20751_, _20750_, _20745_);
  or (_20752_, _20660_, _02303_);
  and (_20753_, _20752_, _01887_);
  and (_20754_, _20753_, _20751_);
  and (_20755_, _20688_, _01860_);
  or (_20756_, _20755_, _01537_);
  or (_20757_, _20756_, _20754_);
  and (_20758_, _11887_, _03665_);
  or (_20759_, _20655_, _01538_);
  or (_20761_, _20759_, _20758_);
  and (_20762_, _20761_, _38087_);
  and (_20763_, _20762_, _20757_);
  nor (_20764_, \oc8051_golden_model_1.P2 [6], rst);
  nor (_20765_, _20764_, _03183_);
  or (_40256_, _20765_, _20763_);
  and (_20766_, _08115_, \oc8051_golden_model_1.P3 [0]);
  and (_20767_, _10620_, _03646_);
  or (_20768_, _20767_, _20766_);
  and (_20769_, _20768_, _02167_);
  and (_20771_, _03646_, _03028_);
  or (_20772_, _20771_, _20766_);
  or (_20773_, _20772_, _05249_);
  nor (_20774_, _04106_, _08115_);
  or (_20775_, _20774_, _20766_);
  or (_20776_, _20775_, _02814_);
  and (_20777_, _03646_, \oc8051_golden_model_1.ACC [0]);
  or (_20778_, _20777_, _20766_);
  and (_20779_, _20778_, _02817_);
  and (_20780_, _02818_, \oc8051_golden_model_1.P3 [0]);
  or (_20782_, _20780_, _02001_);
  or (_20783_, _20782_, _20779_);
  and (_20784_, _20783_, _02024_);
  and (_20785_, _20784_, _20776_);
  and (_20786_, _08123_, \oc8051_golden_model_1.P3 [0]);
  and (_20787_, _10510_, _04338_);
  or (_20788_, _20787_, _20786_);
  and (_20789_, _20788_, _02007_);
  or (_20790_, _20789_, _20785_);
  and (_20791_, _20790_, _02840_);
  and (_20793_, _20772_, _01999_);
  or (_20794_, _20793_, _02006_);
  or (_20795_, _20794_, _20791_);
  or (_20796_, _20778_, _02021_);
  and (_20797_, _20796_, _02025_);
  and (_20798_, _20797_, _20795_);
  and (_20799_, _20766_, _01997_);
  or (_20800_, _20799_, _01991_);
  or (_20801_, _20800_, _20798_);
  or (_20802_, _20775_, _02861_);
  and (_20804_, _20802_, _02408_);
  and (_20805_, _20804_, _20801_);
  and (_20806_, _18380_, _04338_);
  or (_20807_, _20806_, _20786_);
  and (_20808_, _20807_, _01875_);
  or (_20809_, _20808_, _05994_);
  or (_20810_, _20809_, _20805_);
  and (_20811_, _20810_, _20773_);
  or (_20812_, _20811_, _02528_);
  and (_20813_, _04952_, _03646_);
  or (_20815_, _20766_, _02888_);
  or (_20816_, _20815_, _20813_);
  and (_20817_, _20816_, _02043_);
  and (_20818_, _20817_, _20812_);
  and (_20819_, _18407_, _03646_);
  or (_20820_, _20819_, _20766_);
  and (_20821_, _20820_, _01602_);
  or (_20822_, _20821_, _01869_);
  or (_20823_, _20822_, _20818_);
  and (_20824_, _03646_, _04562_);
  or (_20826_, _20824_, _20766_);
  or (_20827_, _20826_, _01870_);
  and (_20828_, _20827_, _20823_);
  or (_20829_, _20828_, _02079_);
  and (_20830_, _10614_, _03646_);
  or (_20831_, _20766_, _02166_);
  or (_20832_, _20831_, _20830_);
  and (_20833_, _20832_, _02912_);
  and (_20834_, _20833_, _20829_);
  or (_20835_, _20834_, _20769_);
  and (_20837_, _20835_, _02176_);
  nand (_20838_, _20826_, _02072_);
  nor (_20839_, _20838_, _20774_);
  or (_20840_, _20839_, _20837_);
  and (_20841_, _20840_, _02907_);
  or (_20842_, _20766_, _04106_);
  and (_20843_, _20778_, _02177_);
  and (_20844_, _20843_, _20842_);
  or (_20845_, _20844_, _02071_);
  or (_20846_, _20845_, _20841_);
  nor (_20848_, _10613_, _08115_);
  or (_20849_, _20766_, _04788_);
  or (_20850_, _20849_, _20848_);
  and (_20851_, _20850_, _04793_);
  and (_20852_, _20851_, _20846_);
  nor (_20853_, _10619_, _08115_);
  or (_20854_, _20853_, _20766_);
  and (_20855_, _20854_, _02173_);
  or (_20856_, _20855_, _02201_);
  or (_20857_, _20856_, _20852_);
  or (_20859_, _20775_, _02303_);
  and (_20860_, _20859_, _01887_);
  and (_20861_, _20860_, _20857_);
  and (_20862_, _20766_, _01860_);
  or (_20863_, _20862_, _01537_);
  or (_20864_, _20863_, _20861_);
  or (_20865_, _20775_, _01538_);
  and (_20866_, _20865_, _38087_);
  and (_20867_, _20866_, _20864_);
  nor (_20868_, \oc8051_golden_model_1.P3 [0], rst);
  nor (_20870_, _20868_, _03183_);
  or (_40258_, _20870_, _20867_);
  and (_20871_, _08115_, \oc8051_golden_model_1.P3 [1]);
  nor (_20872_, _08115_, _02811_);
  or (_20873_, _20872_, _20871_);
  or (_20874_, _20873_, _02840_);
  or (_20875_, _03646_, \oc8051_golden_model_1.P3 [1]);
  and (_20876_, _10698_, _03646_);
  not (_20877_, _20876_);
  and (_20878_, _20877_, _20875_);
  or (_20880_, _20878_, _02814_);
  nand (_20881_, _03646_, _01613_);
  and (_20882_, _20881_, _20875_);
  and (_20883_, _20882_, _02817_);
  and (_20884_, _02818_, \oc8051_golden_model_1.P3 [1]);
  or (_20885_, _20884_, _02001_);
  or (_20886_, _20885_, _20883_);
  and (_20887_, _20886_, _02024_);
  and (_20888_, _20887_, _20880_);
  and (_20889_, _08123_, \oc8051_golden_model_1.P3 [1]);
  and (_20891_, _10710_, _04338_);
  or (_20892_, _20891_, _20889_);
  and (_20893_, _20892_, _02007_);
  or (_20894_, _20893_, _01999_);
  or (_20895_, _20894_, _20888_);
  and (_20896_, _20895_, _20874_);
  or (_20897_, _20896_, _02006_);
  or (_20898_, _20882_, _02021_);
  and (_20899_, _20898_, _02025_);
  and (_20900_, _20899_, _20897_);
  and (_20902_, _10696_, _04338_);
  or (_20903_, _20902_, _20889_);
  and (_20904_, _20903_, _01997_);
  or (_20905_, _20904_, _01991_);
  or (_20906_, _20905_, _20900_);
  and (_20907_, _20891_, _10725_);
  or (_20908_, _20889_, _02861_);
  or (_20909_, _20908_, _20907_);
  and (_20910_, _20909_, _20906_);
  and (_20911_, _20910_, _02408_);
  and (_20913_, _18500_, _04338_);
  or (_20914_, _20889_, _20913_);
  and (_20915_, _20914_, _01875_);
  or (_20916_, _20915_, _05994_);
  or (_20917_, _20916_, _20911_);
  or (_20918_, _20873_, _05249_);
  and (_20919_, _20918_, _20917_);
  or (_20920_, _20919_, _02528_);
  and (_20921_, _04907_, _03646_);
  or (_20922_, _20871_, _02888_);
  or (_20924_, _20922_, _20921_);
  and (_20925_, _20924_, _02043_);
  and (_20926_, _20925_, _20920_);
  and (_20927_, _18528_, _03646_);
  or (_20928_, _20927_, _20871_);
  and (_20929_, _20928_, _01602_);
  or (_20930_, _20929_, _20926_);
  and (_20931_, _20930_, _01870_);
  nand (_20932_, _03646_, _02687_);
  and (_20933_, _20875_, _01869_);
  and (_20935_, _20933_, _20932_);
  or (_20936_, _20935_, _20931_);
  and (_20937_, _20936_, _02166_);
  or (_20938_, _10816_, _08115_);
  and (_20939_, _20875_, _02079_);
  and (_20940_, _20939_, _20938_);
  or (_20941_, _20940_, _20937_);
  and (_20942_, _20941_, _02912_);
  or (_20943_, _10822_, _08115_);
  and (_20944_, _20875_, _02167_);
  and (_20946_, _20944_, _20943_);
  or (_20947_, _20946_, _20942_);
  and (_20948_, _20947_, _02176_);
  or (_20949_, _10692_, _08115_);
  and (_20950_, _20875_, _02072_);
  and (_20951_, _20950_, _20949_);
  or (_20952_, _20951_, _20948_);
  and (_20953_, _20952_, _02907_);
  or (_20954_, _20871_, _04058_);
  and (_20955_, _20882_, _02177_);
  and (_20957_, _20955_, _20954_);
  or (_20958_, _20957_, _20953_);
  and (_20959_, _20958_, _02174_);
  or (_20960_, _20881_, _04058_);
  and (_20961_, _20875_, _02173_);
  and (_20962_, _20961_, _20960_);
  or (_20963_, _20962_, _02201_);
  or (_20964_, _20932_, _04058_);
  and (_20965_, _20875_, _02071_);
  and (_20966_, _20965_, _20964_);
  or (_20968_, _20966_, _20963_);
  or (_20969_, _20968_, _20959_);
  or (_20970_, _20878_, _02303_);
  and (_20971_, _20970_, _01887_);
  and (_20972_, _20971_, _20969_);
  and (_20973_, _20903_, _01860_);
  or (_20974_, _20973_, _01537_);
  or (_20975_, _20974_, _20972_);
  or (_20976_, _20871_, _01538_);
  or (_20977_, _20976_, _20876_);
  and (_20979_, _20977_, _38087_);
  and (_20980_, _20979_, _20975_);
  nor (_20981_, \oc8051_golden_model_1.P3 [1], rst);
  nor (_20982_, _20981_, _03183_);
  or (_40259_, _20982_, _20980_);
  and (_20983_, _08115_, \oc8051_golden_model_1.P3 [2]);
  and (_20984_, _11020_, _03646_);
  or (_20985_, _20984_, _20983_);
  and (_20986_, _20985_, _02167_);
  nor (_20987_, _08115_, _03455_);
  or (_20989_, _20987_, _20983_);
  or (_20990_, _20989_, _05249_);
  and (_20991_, _20989_, _01999_);
  and (_20992_, _08123_, \oc8051_golden_model_1.P3 [2]);
  and (_20993_, _10909_, _04338_);
  or (_20994_, _20993_, _20992_);
  or (_20995_, _20994_, _02024_);
  nor (_20996_, _10905_, _08115_);
  or (_20997_, _20996_, _20983_);
  and (_20998_, _20997_, _02001_);
  and (_21000_, _02818_, \oc8051_golden_model_1.P3 [2]);
  and (_21001_, _03646_, \oc8051_golden_model_1.ACC [2]);
  or (_21002_, _21001_, _20983_);
  and (_21003_, _21002_, _02817_);
  or (_21004_, _21003_, _21000_);
  and (_21005_, _21004_, _02814_);
  or (_21006_, _21005_, _02007_);
  or (_21007_, _21006_, _20998_);
  and (_21008_, _21007_, _20995_);
  and (_21009_, _21008_, _02840_);
  or (_21011_, _21009_, _20991_);
  or (_21012_, _21011_, _02006_);
  or (_21013_, _21002_, _02021_);
  and (_21014_, _21013_, _02025_);
  and (_21015_, _21014_, _21012_);
  and (_21016_, _10894_, _04338_);
  or (_21017_, _21016_, _20992_);
  and (_21018_, _21017_, _01997_);
  or (_21019_, _21018_, _01991_);
  or (_21020_, _21019_, _21015_);
  or (_21022_, _20992_, _10924_);
  and (_21023_, _21022_, _20994_);
  or (_21024_, _21023_, _02861_);
  and (_21025_, _21024_, _02408_);
  and (_21026_, _21025_, _21020_);
  and (_21027_, _18628_, _04338_);
  or (_21028_, _21027_, _20992_);
  and (_21029_, _21028_, _01875_);
  or (_21030_, _21029_, _05994_);
  or (_21031_, _21030_, _21026_);
  and (_21033_, _21031_, _20990_);
  or (_21034_, _21033_, _02528_);
  and (_21035_, _05043_, _03646_);
  or (_21036_, _20983_, _02888_);
  or (_21037_, _21036_, _21035_);
  and (_21038_, _21037_, _02043_);
  and (_21039_, _21038_, _21034_);
  and (_21040_, _18655_, _03646_);
  or (_21041_, _21040_, _20983_);
  and (_21042_, _21041_, _01602_);
  or (_21044_, _21042_, _01869_);
  or (_21045_, _21044_, _21039_);
  and (_21046_, _03646_, _04724_);
  or (_21047_, _21046_, _20983_);
  or (_21048_, _21047_, _01870_);
  and (_21049_, _21048_, _21045_);
  or (_21050_, _21049_, _02079_);
  and (_21051_, _11014_, _03646_);
  or (_21052_, _20983_, _02166_);
  or (_21053_, _21052_, _21051_);
  and (_21055_, _21053_, _02912_);
  and (_21056_, _21055_, _21050_);
  or (_21057_, _21056_, _20986_);
  and (_21058_, _21057_, _02176_);
  or (_21059_, _20983_, _04156_);
  and (_21060_, _21047_, _02072_);
  and (_21061_, _21060_, _21059_);
  or (_21062_, _21061_, _21058_);
  and (_21063_, _21062_, _02907_);
  and (_21064_, _21002_, _02177_);
  and (_21066_, _21064_, _21059_);
  or (_21067_, _21066_, _02071_);
  or (_21068_, _21067_, _21063_);
  nor (_21069_, _11013_, _08115_);
  or (_21070_, _20983_, _04788_);
  or (_21071_, _21070_, _21069_);
  and (_21072_, _21071_, _04793_);
  and (_21073_, _21072_, _21068_);
  nor (_21074_, _11019_, _08115_);
  or (_21075_, _21074_, _20983_);
  and (_21077_, _21075_, _02173_);
  or (_21078_, _21077_, _02201_);
  or (_21079_, _21078_, _21073_);
  or (_21080_, _20997_, _02303_);
  and (_21081_, _21080_, _01887_);
  and (_21082_, _21081_, _21079_);
  and (_21083_, _21017_, _01860_);
  or (_21084_, _21083_, _01537_);
  or (_21085_, _21084_, _21082_);
  and (_21086_, _11072_, _03646_);
  or (_21088_, _20983_, _01538_);
  or (_21089_, _21088_, _21086_);
  and (_21090_, _21089_, _38087_);
  and (_21091_, _21090_, _21085_);
  nor (_21092_, \oc8051_golden_model_1.P3 [2], rst);
  nor (_21093_, _21092_, _03183_);
  or (_40260_, _21093_, _21091_);
  and (_21094_, _08115_, \oc8051_golden_model_1.P3 [3]);
  and (_21095_, _11094_, _03646_);
  or (_21096_, _21095_, _21094_);
  and (_21098_, _21096_, _02167_);
  nor (_21099_, _08115_, _03268_);
  or (_21100_, _21099_, _21094_);
  or (_21101_, _21100_, _05249_);
  nor (_21102_, _11101_, _08115_);
  or (_21103_, _21102_, _21094_);
  or (_21104_, _21103_, _02814_);
  and (_21105_, _03646_, \oc8051_golden_model_1.ACC [3]);
  or (_21106_, _21105_, _21094_);
  and (_21107_, _21106_, _02817_);
  and (_21109_, _02818_, \oc8051_golden_model_1.P3 [3]);
  or (_21110_, _21109_, _02001_);
  or (_21111_, _21110_, _21107_);
  and (_21112_, _21111_, _02024_);
  and (_21113_, _21112_, _21104_);
  and (_21114_, _08123_, \oc8051_golden_model_1.P3 [3]);
  and (_21115_, _11098_, _04338_);
  or (_21116_, _21115_, _21114_);
  and (_21117_, _21116_, _02007_);
  or (_21118_, _21117_, _01999_);
  or (_21120_, _21118_, _21113_);
  or (_21121_, _21100_, _02840_);
  and (_21122_, _21121_, _21120_);
  or (_21123_, _21122_, _02006_);
  or (_21124_, _21106_, _02021_);
  and (_21125_, _21124_, _02025_);
  and (_21126_, _21125_, _21123_);
  and (_21127_, _11096_, _04338_);
  or (_21128_, _21127_, _21114_);
  and (_21129_, _21128_, _01997_);
  or (_21131_, _21129_, _01991_);
  or (_21132_, _21131_, _21126_);
  or (_21133_, _21114_, _11127_);
  and (_21134_, _21133_, _21116_);
  or (_21135_, _21134_, _02861_);
  and (_21136_, _21135_, _02408_);
  and (_21137_, _21136_, _21132_);
  and (_21138_, _18754_, _04338_);
  or (_21139_, _21138_, _21114_);
  and (_21140_, _21139_, _01875_);
  or (_21142_, _21140_, _05994_);
  or (_21143_, _21142_, _21137_);
  and (_21144_, _21143_, _21101_);
  or (_21145_, _21144_, _02528_);
  and (_21146_, _04998_, _03646_);
  or (_21147_, _21094_, _02888_);
  or (_21148_, _21147_, _21146_);
  and (_21149_, _21148_, _02043_);
  and (_21150_, _21149_, _21145_);
  and (_21151_, _18780_, _03646_);
  or (_21153_, _21151_, _21094_);
  and (_21154_, _21153_, _01602_);
  or (_21155_, _21154_, _01869_);
  or (_21156_, _21155_, _21150_);
  and (_21157_, _03646_, _04678_);
  or (_21158_, _21157_, _21094_);
  or (_21159_, _21158_, _01870_);
  and (_21160_, _21159_, _21156_);
  or (_21161_, _21160_, _02079_);
  and (_21162_, _11222_, _03646_);
  or (_21164_, _21094_, _02166_);
  or (_21165_, _21164_, _21162_);
  and (_21166_, _21165_, _02912_);
  and (_21167_, _21166_, _21161_);
  or (_21168_, _21167_, _21098_);
  and (_21169_, _21168_, _02176_);
  or (_21170_, _21094_, _04014_);
  and (_21171_, _21158_, _02072_);
  and (_21172_, _21171_, _21170_);
  or (_21173_, _21172_, _21169_);
  and (_21175_, _21173_, _02907_);
  and (_21176_, _21106_, _02177_);
  and (_21177_, _21176_, _21170_);
  or (_21178_, _21177_, _02071_);
  or (_21179_, _21178_, _21175_);
  nor (_21180_, _11220_, _08115_);
  or (_21181_, _21094_, _04788_);
  or (_21182_, _21181_, _21180_);
  and (_21183_, _21182_, _04793_);
  and (_21184_, _21183_, _21179_);
  nor (_21186_, _11093_, _08115_);
  or (_21187_, _21186_, _21094_);
  and (_21188_, _21187_, _02173_);
  or (_21189_, _21188_, _02201_);
  or (_21190_, _21189_, _21184_);
  or (_21191_, _21103_, _02303_);
  and (_21192_, _21191_, _01887_);
  and (_21193_, _21192_, _21190_);
  and (_21194_, _21128_, _01860_);
  or (_21195_, _21194_, _01537_);
  or (_21197_, _21195_, _21193_);
  and (_21198_, _11273_, _03646_);
  or (_21199_, _21094_, _01538_);
  or (_21200_, _21199_, _21198_);
  and (_21201_, _21200_, _38087_);
  and (_21202_, _21201_, _21197_);
  nor (_21203_, \oc8051_golden_model_1.P3 [3], rst);
  nor (_21204_, _21203_, _03183_);
  or (_40261_, _21204_, _21202_);
  nor (_21205_, \oc8051_golden_model_1.P3 [4], rst);
  nor (_21207_, _21205_, _03183_);
  and (_21208_, _08115_, \oc8051_golden_model_1.P3 [4]);
  and (_21209_, _11431_, _03646_);
  or (_21210_, _21209_, _21208_);
  and (_21211_, _21210_, _02167_);
  nor (_21212_, _04211_, _08115_);
  or (_21213_, _21212_, _21208_);
  or (_21214_, _21213_, _05249_);
  and (_21215_, _08123_, \oc8051_golden_model_1.P3 [4]);
  and (_21216_, _11301_, _04338_);
  or (_21218_, _21216_, _21215_);
  and (_21219_, _21218_, _01997_);
  nor (_21220_, _11317_, _08115_);
  or (_21221_, _21220_, _21208_);
  or (_21222_, _21221_, _02814_);
  and (_21223_, _03646_, \oc8051_golden_model_1.ACC [4]);
  or (_21224_, _21223_, _21208_);
  and (_21225_, _21224_, _02817_);
  and (_21226_, _02818_, \oc8051_golden_model_1.P3 [4]);
  or (_21227_, _21226_, _02001_);
  or (_21229_, _21227_, _21225_);
  and (_21230_, _21229_, _02024_);
  and (_21231_, _21230_, _21222_);
  and (_21232_, _11303_, _04338_);
  or (_21233_, _21232_, _21215_);
  and (_21234_, _21233_, _02007_);
  or (_21235_, _21234_, _01999_);
  or (_21236_, _21235_, _21231_);
  or (_21237_, _21213_, _02840_);
  and (_21238_, _21237_, _21236_);
  or (_21240_, _21238_, _02006_);
  or (_21241_, _21224_, _02021_);
  and (_21242_, _21241_, _02025_);
  and (_21243_, _21242_, _21240_);
  or (_21244_, _21243_, _21219_);
  and (_21245_, _21244_, _02861_);
  and (_21246_, _11335_, _04338_);
  or (_21247_, _21246_, _21215_);
  and (_21248_, _21247_, _01991_);
  or (_21249_, _21248_, _21245_);
  and (_21251_, _21249_, _02408_);
  and (_21252_, _18879_, _04338_);
  or (_21253_, _21252_, _21215_);
  and (_21254_, _21253_, _01875_);
  or (_21255_, _21254_, _05994_);
  or (_21256_, _21255_, _21251_);
  and (_21257_, _21256_, _21214_);
  or (_21258_, _21257_, _02528_);
  and (_21259_, _05135_, _03646_);
  or (_21260_, _21208_, _02888_);
  or (_21262_, _21260_, _21259_);
  and (_21263_, _21262_, _02043_);
  and (_21264_, _21263_, _21258_);
  and (_21265_, _18909_, _03646_);
  or (_21266_, _21265_, _21208_);
  and (_21267_, _21266_, _01602_);
  or (_21268_, _21267_, _01869_);
  or (_21269_, _21268_, _21264_);
  and (_21270_, _04694_, _03646_);
  or (_21271_, _21270_, _21208_);
  or (_21273_, _21271_, _01870_);
  and (_21274_, _21273_, _21269_);
  or (_21275_, _21274_, _02079_);
  and (_21276_, _11425_, _03646_);
  or (_21277_, _21208_, _02166_);
  or (_21278_, _21277_, _21276_);
  and (_21279_, _21278_, _02912_);
  and (_21280_, _21279_, _21275_);
  or (_21281_, _21280_, _21211_);
  and (_21282_, _21281_, _02176_);
  or (_21284_, _21208_, _04258_);
  and (_21285_, _21271_, _02072_);
  and (_21286_, _21285_, _21284_);
  or (_21287_, _21286_, _21282_);
  and (_21288_, _21287_, _02907_);
  and (_21289_, _21224_, _02177_);
  and (_21290_, _21289_, _21284_);
  or (_21291_, _21290_, _02071_);
  or (_21292_, _21291_, _21288_);
  nor (_21293_, _11424_, _08115_);
  or (_21295_, _21208_, _04788_);
  or (_21296_, _21295_, _21293_);
  and (_21297_, _21296_, _04793_);
  and (_21298_, _21297_, _21292_);
  nor (_21299_, _11430_, _08115_);
  or (_21300_, _21299_, _21208_);
  and (_21301_, _21300_, _02173_);
  or (_21302_, _21301_, _02201_);
  or (_21303_, _21302_, _21298_);
  or (_21304_, _21221_, _02303_);
  and (_21306_, _21304_, _01887_);
  and (_21307_, _21306_, _21303_);
  and (_21308_, _21218_, _01860_);
  or (_21309_, _21308_, _01537_);
  or (_21310_, _21309_, _21307_);
  and (_21311_, _11487_, _03646_);
  or (_21312_, _21208_, _01538_);
  or (_21313_, _21312_, _21311_);
  and (_21314_, _21313_, _38087_);
  and (_21315_, _21314_, _21310_);
  or (_40263_, _21315_, _21207_);
  and (_21317_, _08115_, \oc8051_golden_model_1.P3 [5]);
  and (_21318_, _11635_, _03646_);
  or (_21319_, _21318_, _21317_);
  and (_21320_, _21319_, _02167_);
  nor (_21321_, _11525_, _08115_);
  or (_21322_, _21321_, _21317_);
  or (_21323_, _21322_, _02814_);
  and (_21324_, _03646_, \oc8051_golden_model_1.ACC [5]);
  or (_21325_, _21324_, _21317_);
  and (_21327_, _21325_, _02817_);
  and (_21328_, _02818_, \oc8051_golden_model_1.P3 [5]);
  or (_21329_, _21328_, _02001_);
  or (_21330_, _21329_, _21327_);
  and (_21331_, _21330_, _02024_);
  and (_21332_, _21331_, _21323_);
  and (_21333_, _08123_, \oc8051_golden_model_1.P3 [5]);
  and (_21334_, _11510_, _04338_);
  or (_21335_, _21334_, _21333_);
  and (_21336_, _21335_, _02007_);
  or (_21338_, _21336_, _01999_);
  or (_21339_, _21338_, _21332_);
  nor (_21340_, _03916_, _08115_);
  or (_21341_, _21340_, _21317_);
  or (_21342_, _21341_, _02840_);
  and (_21343_, _21342_, _21339_);
  or (_21344_, _21343_, _02006_);
  or (_21345_, _21325_, _02021_);
  and (_21346_, _21345_, _02025_);
  and (_21347_, _21346_, _21344_);
  and (_21349_, _11508_, _04338_);
  or (_21350_, _21349_, _21333_);
  and (_21351_, _21350_, _01997_);
  or (_21352_, _21351_, _01991_);
  or (_21353_, _21352_, _21347_);
  or (_21354_, _21333_, _11542_);
  and (_21355_, _21354_, _21335_);
  or (_21356_, _21355_, _02861_);
  and (_21357_, _21356_, _02408_);
  and (_21358_, _21357_, _21353_);
  and (_21360_, _19009_, _04338_);
  or (_21361_, _21360_, _21333_);
  and (_21362_, _21361_, _01875_);
  or (_21363_, _21362_, _05994_);
  or (_21364_, _21363_, _21358_);
  or (_21365_, _21341_, _05249_);
  and (_21366_, _21365_, _21364_);
  or (_21367_, _21366_, _02528_);
  and (_21368_, _05090_, _03646_);
  or (_21369_, _21317_, _02888_);
  or (_21371_, _21369_, _21368_);
  and (_21372_, _21371_, _02043_);
  and (_21373_, _21372_, _21367_);
  and (_21374_, _19037_, _03646_);
  or (_21375_, _21374_, _21317_);
  and (_21376_, _21375_, _01602_);
  or (_21377_, _21376_, _01869_);
  or (_21378_, _21377_, _21373_);
  and (_21379_, _04672_, _03646_);
  or (_21380_, _21379_, _21317_);
  or (_21382_, _21380_, _01870_);
  and (_21383_, _21382_, _21378_);
  or (_21384_, _21383_, _02079_);
  and (_21385_, _11629_, _03646_);
  or (_21386_, _21317_, _02166_);
  or (_21387_, _21386_, _21385_);
  and (_21388_, _21387_, _02912_);
  and (_21389_, _21388_, _21384_);
  or (_21390_, _21389_, _21320_);
  and (_21391_, _21390_, _02176_);
  or (_21393_, _21317_, _03965_);
  and (_21394_, _21380_, _02072_);
  and (_21395_, _21394_, _21393_);
  or (_21396_, _21395_, _21391_);
  and (_21397_, _21396_, _02907_);
  and (_21398_, _21325_, _02177_);
  and (_21399_, _21398_, _21393_);
  or (_21400_, _21399_, _02071_);
  or (_21401_, _21400_, _21397_);
  nor (_21402_, _11628_, _08115_);
  or (_21404_, _21317_, _04788_);
  or (_21405_, _21404_, _21402_);
  and (_21406_, _21405_, _04793_);
  and (_21407_, _21406_, _21401_);
  nor (_21408_, _11634_, _08115_);
  or (_21409_, _21408_, _21317_);
  and (_21410_, _21409_, _02173_);
  or (_21411_, _21410_, _02201_);
  or (_21412_, _21411_, _21407_);
  or (_21413_, _21322_, _02303_);
  and (_21415_, _21413_, _01887_);
  and (_21416_, _21415_, _21412_);
  and (_21417_, _21350_, _01860_);
  or (_21418_, _21417_, _01537_);
  or (_21419_, _21418_, _21416_);
  and (_21420_, _11685_, _03646_);
  or (_21421_, _21317_, _01538_);
  or (_21422_, _21421_, _21420_);
  and (_21423_, _21422_, _38087_);
  and (_21424_, _21423_, _21419_);
  nor (_21426_, \oc8051_golden_model_1.P3 [5], rst);
  nor (_21427_, _21426_, _03183_);
  or (_40264_, _21427_, _21424_);
  and (_21428_, _08115_, \oc8051_golden_model_1.P3 [6]);
  and (_21429_, _11709_, _03646_);
  or (_21430_, _21429_, _21428_);
  and (_21431_, _21430_, _02167_);
  nor (_21432_, _11730_, _08115_);
  or (_21433_, _21432_, _21428_);
  or (_21434_, _21433_, _02814_);
  and (_21436_, _03646_, \oc8051_golden_model_1.ACC [6]);
  or (_21437_, _21436_, _21428_);
  and (_21438_, _21437_, _02817_);
  and (_21439_, _02818_, \oc8051_golden_model_1.P3 [6]);
  or (_21440_, _21439_, _02001_);
  or (_21441_, _21440_, _21438_);
  and (_21442_, _21441_, _02024_);
  and (_21443_, _21442_, _21434_);
  and (_21444_, _08123_, \oc8051_golden_model_1.P3 [6]);
  and (_21445_, _11717_, _04338_);
  or (_21447_, _21445_, _21444_);
  and (_21448_, _21447_, _02007_);
  or (_21449_, _21448_, _01999_);
  or (_21450_, _21449_, _21443_);
  nor (_21451_, _03808_, _08115_);
  or (_21452_, _21451_, _21428_);
  or (_21453_, _21452_, _02840_);
  and (_21454_, _21453_, _21450_);
  or (_21455_, _21454_, _02006_);
  or (_21456_, _21437_, _02021_);
  and (_21458_, _21456_, _02025_);
  and (_21459_, _21458_, _21455_);
  and (_21460_, _11715_, _04338_);
  or (_21461_, _21460_, _21444_);
  and (_21462_, _21461_, _01997_);
  or (_21463_, _21462_, _01991_);
  or (_21464_, _21463_, _21459_);
  or (_21465_, _21444_, _11747_);
  and (_21466_, _21465_, _21447_);
  or (_21467_, _21466_, _02861_);
  and (_21469_, _21467_, _02408_);
  and (_21470_, _21469_, _21464_);
  and (_21471_, _19133_, _04338_);
  or (_21472_, _21471_, _21444_);
  and (_21473_, _21472_, _01875_);
  or (_21474_, _21473_, _05994_);
  or (_21475_, _21474_, _21470_);
  or (_21476_, _21452_, _05249_);
  and (_21477_, _21476_, _21475_);
  or (_21478_, _21477_, _02528_);
  and (_21480_, _04861_, _03646_);
  or (_21481_, _21428_, _02888_);
  or (_21482_, _21481_, _21480_);
  and (_21483_, _21482_, _02043_);
  and (_21484_, _21483_, _21478_);
  and (_21485_, _19161_, _03646_);
  or (_21486_, _21485_, _21428_);
  and (_21487_, _21486_, _01602_);
  or (_21488_, _21487_, _01869_);
  or (_21489_, _21488_, _21484_);
  and (_21491_, _09920_, _03646_);
  or (_21492_, _21491_, _21428_);
  or (_21493_, _21492_, _01870_);
  and (_21494_, _21493_, _21489_);
  or (_21495_, _21494_, _02079_);
  and (_21496_, _11835_, _03646_);
  or (_21497_, _21428_, _02166_);
  or (_21498_, _21497_, _21496_);
  and (_21499_, _21498_, _02912_);
  and (_21500_, _21499_, _21495_);
  or (_21502_, _21500_, _21431_);
  and (_21503_, _21502_, _02176_);
  or (_21504_, _21428_, _03863_);
  and (_21505_, _21492_, _02072_);
  and (_21506_, _21505_, _21504_);
  or (_21507_, _21506_, _21503_);
  and (_21508_, _21507_, _02907_);
  and (_21509_, _21437_, _02177_);
  and (_21510_, _21509_, _21504_);
  or (_21511_, _21510_, _02071_);
  or (_21513_, _21511_, _21508_);
  nor (_21514_, _11833_, _08115_);
  or (_21515_, _21428_, _04788_);
  or (_21516_, _21515_, _21514_);
  and (_21517_, _21516_, _04793_);
  and (_21518_, _21517_, _21513_);
  nor (_21519_, _11708_, _08115_);
  or (_21520_, _21519_, _21428_);
  and (_21521_, _21520_, _02173_);
  or (_21522_, _21521_, _02201_);
  or (_21524_, _21522_, _21518_);
  or (_21525_, _21433_, _02303_);
  and (_21526_, _21525_, _01887_);
  and (_21527_, _21526_, _21524_);
  and (_21528_, _21461_, _01860_);
  or (_21529_, _21528_, _01537_);
  or (_21530_, _21529_, _21527_);
  and (_21531_, _11887_, _03646_);
  or (_21532_, _21428_, _01538_);
  or (_21533_, _21532_, _21531_);
  and (_21535_, _21533_, _38087_);
  and (_21536_, _21535_, _21530_);
  nor (_21537_, \oc8051_golden_model_1.P3 [6], rst);
  nor (_21538_, _21537_, _03183_);
  or (_40265_, _21538_, _21536_);
  not (_21539_, \oc8051_golden_model_1.PSW [0]);
  nor (_21540_, _38087_, _21539_);
  nor (_21541_, _06126_, _06125_);
  nor (_21542_, _21541_, _06026_);
  and (_21543_, _21541_, _06026_);
  nor (_21545_, _21543_, _21542_);
  nor (_21546_, _06044_, _06043_);
  nor (_21547_, _21546_, _13937_);
  and (_21548_, _21546_, _13937_);
  nor (_21549_, _21548_, _21547_);
  and (_21550_, _21549_, _21545_);
  nor (_21551_, _21549_, _21545_);
  nor (_21552_, _21551_, _21550_);
  or (_21553_, _21552_, _04776_);
  nand (_21554_, _21552_, _04776_);
  and (_21556_, _21554_, _21553_);
  or (_21557_, _21556_, _05172_);
  nand (_21558_, _13793_, _13523_);
  or (_21559_, _13793_, _13523_);
  and (_21560_, _21559_, _21558_);
  and (_21561_, _21560_, _14097_);
  nor (_21562_, _21560_, _14097_);
  or (_21563_, _21562_, _21561_);
  nor (_21564_, _21563_, _14408_);
  and (_21565_, _21563_, _14408_);
  nor (_21567_, _21565_, _21564_);
  or (_21568_, _21567_, _14612_);
  nand (_21569_, _21567_, _14612_);
  and (_21570_, _21569_, _21568_);
  nor (_21571_, _21570_, _14917_);
  and (_21572_, _21570_, _14917_);
  or (_21573_, _21572_, _21571_);
  and (_21574_, _21573_, _15332_);
  nor (_21575_, _21573_, _15332_);
  nor (_21576_, _21575_, _21574_);
  and (_21578_, _21576_, _06540_);
  nor (_21579_, _21576_, _06540_);
  or (_21580_, _21579_, _21578_);
  or (_21581_, _21580_, _06777_);
  not (_21582_, _14038_);
  nor (_21583_, _13756_, _13452_);
  and (_21584_, _13756_, _13452_);
  nor (_21585_, _21584_, _21583_);
  nor (_21586_, _21585_, _21582_);
  and (_21587_, _21585_, _21582_);
  or (_21589_, _21587_, _21586_);
  and (_21590_, _21589_, _14357_);
  nor (_21591_, _21589_, _14357_);
  or (_21592_, _21591_, _21590_);
  and (_21593_, _21592_, _14659_);
  nor (_21594_, _21592_, _14659_);
  or (_21595_, _21594_, _21593_);
  and (_21596_, _21595_, _14981_);
  nor (_21597_, _21595_, _14981_);
  or (_21598_, _21597_, _21596_);
  and (_21600_, _21598_, _15304_);
  nor (_21601_, _21598_, _15304_);
  or (_21602_, _21601_, _21600_);
  and (_21603_, _21602_, _06687_);
  nor (_21604_, _21602_, _06687_);
  or (_21605_, _21604_, _21603_);
  and (_21606_, _21605_, _01997_);
  and (_21607_, \oc8051_golden_model_1.ACC [2], \oc8051_golden_model_1.ACC [0]);
  nor (_21608_, \oc8051_golden_model_1.ACC [2], \oc8051_golden_model_1.ACC [0]);
  or (_21609_, _21608_, _21607_);
  and (_21611_, _21609_, _13731_);
  nor (_21612_, _21609_, _13731_);
  nor (_21613_, _21612_, _21611_);
  and (_21614_, _14635_, _14334_);
  nor (_21615_, _14635_, _14334_);
  nor (_21616_, _21615_, _21614_);
  nor (_21617_, _21616_, _21613_);
  and (_21618_, _21616_, _21613_);
  or (_21619_, _21618_, _21617_);
  nor (_21620_, _21619_, _14959_);
  and (_21622_, _21619_, _14959_);
  or (_21623_, _21622_, _21620_);
  nor (_21624_, _15280_, _06661_);
  and (_21625_, _15280_, _06661_);
  nor (_21626_, _21625_, _21624_);
  nand (_21627_, _21626_, _21623_);
  or (_21628_, _21626_, _21623_);
  and (_21629_, _21628_, _21627_);
  or (_21630_, _21629_, _06642_);
  and (_21631_, _06884_, _06867_);
  nor (_21633_, _21631_, _06885_);
  and (_21634_, _21633_, _06804_);
  nor (_21635_, _21633_, _06804_);
  nor (_21636_, _21635_, _21634_);
  and (_21637_, _06839_, _06816_);
  and (_21638_, _06838_, _06817_);
  nor (_21639_, _21638_, _21637_);
  and (_21640_, _06850_, _06791_);
  nor (_21641_, _06850_, _06791_);
  or (_21642_, _21641_, _21640_);
  and (_21644_, _21642_, _21639_);
  nor (_21645_, _21642_, _21639_);
  or (_21646_, _21645_, _21644_);
  nor (_21647_, _21646_, _21636_);
  and (_21648_, _21646_, _21636_);
  nor (_21649_, _21648_, _21647_);
  and (_21650_, _21649_, _04528_);
  nor (_21651_, _21649_, _04528_);
  or (_21652_, _21651_, _21650_);
  and (_21653_, _21652_, _02003_);
  nor (_21655_, _05180_, _05044_);
  not (_21656_, _21655_);
  nand (_21657_, _21656_, _10690_);
  or (_21658_, _21656_, _10690_);
  and (_21659_, _21658_, _21657_);
  not (_21660_, _21659_);
  nor (_21661_, _05182_, _05136_);
  nand (_21662_, _21661_, _04861_);
  or (_21663_, _21661_, _04861_);
  and (_21664_, _21663_, _21662_);
  nand (_21666_, _21664_, _21660_);
  or (_21667_, _21664_, _21660_);
  nand (_21668_, _21667_, _21666_);
  nor (_21669_, _21668_, _04483_);
  and (_21670_, _21668_, _04483_);
  or (_21671_, _21670_, _21669_);
  or (_21672_, _21671_, _06621_);
  nor (_21673_, _10700_, _05160_);
  and (_21674_, _10700_, _05160_);
  nor (_21675_, _21674_, _21673_);
  nor (_21677_, _08779_, _10103_);
  nor (_21678_, _05162_, _04373_);
  and (_21679_, _21678_, _03916_);
  nor (_21680_, _21678_, _03916_);
  or (_21681_, _21680_, _21679_);
  nand (_21682_, _21681_, _21677_);
  or (_21683_, _21681_, _21677_);
  and (_21684_, _21683_, _21682_);
  or (_21685_, _21684_, _21675_);
  nand (_21686_, _21684_, _21675_);
  and (_21688_, _21686_, _21685_);
  and (_21689_, _21688_, _06623_);
  nor (_21690_, _10112_, _06625_);
  and (_21691_, _21690_, _09224_);
  or (_21692_, _21691_, _21556_);
  nand (_21693_, _21691_, _21539_);
  and (_21694_, _21693_, _21692_);
  or (_21695_, _21694_, _06620_);
  and (_21696_, _21695_, _13461_);
  or (_21697_, _21696_, _21689_);
  and (_21699_, _21697_, _06618_);
  and (_21700_, _21699_, _21672_);
  or (_21701_, _21700_, _21653_);
  nor (_21702_, _04380_, _10140_);
  and (_21703_, _21702_, _10136_);
  and (_21704_, _21703_, _21701_);
  not (_21705_, _21702_);
  and (_21706_, _21705_, _21556_);
  or (_21707_, _21706_, _01883_);
  or (_21708_, _21707_, _21704_);
  nor (_21710_, _21546_, \oc8051_golden_model_1.ACC [6]);
  and (_21711_, _21546_, \oc8051_golden_model_1.ACC [6]);
  nor (_21712_, _21711_, _21710_);
  nor (_21713_, _21712_, \oc8051_golden_model_1.ACC [7]);
  and (_21714_, _21712_, \oc8051_golden_model_1.ACC [7]);
  nor (_21715_, _21714_, _21713_);
  and (_21716_, _21715_, _21659_);
  nor (_21717_, _21715_, _21659_);
  or (_21718_, _21717_, _21716_);
  or (_21719_, _21718_, _04394_);
  and (_21721_, _21719_, _02814_);
  and (_21722_, _21721_, _21708_);
  nor (_21723_, _14629_, _14312_);
  and (_21724_, _14629_, _14312_);
  nor (_21725_, _21724_, _21723_);
  and (_21726_, _21725_, _15273_);
  nor (_21727_, _21725_, _15273_);
  nor (_21728_, _21727_, _21726_);
  not (_21729_, _13475_);
  nor (_21730_, _13725_, _21729_);
  and (_21732_, _13725_, _21729_);
  nor (_21733_, _21732_, _21730_);
  and (_21734_, _21733_, _14006_);
  nor (_21735_, _21733_, _14006_);
  nor (_21736_, _21735_, _21734_);
  and (_21737_, _21736_, _14953_);
  nor (_21738_, _21736_, _14953_);
  or (_21739_, _21738_, _21737_);
  and (_21740_, _21739_, _06638_);
  nor (_21741_, _21739_, _06638_);
  or (_21743_, _21741_, _21740_);
  nand (_21744_, _21743_, _21728_);
  or (_21745_, _21743_, _21728_);
  and (_21746_, _21745_, _21744_);
  and (_21747_, _21746_, _02001_);
  or (_21748_, _21747_, _06636_);
  or (_21749_, _21748_, _21722_);
  and (_21750_, _21749_, _21630_);
  or (_21751_, _21750_, _08516_);
  or (_21752_, _21556_, _08517_);
  and (_21754_, _21752_, _02024_);
  and (_21755_, _21754_, _21751_);
  nor (_21756_, _14338_, _14020_);
  and (_21757_, _14338_, _14020_);
  nor (_21758_, _21757_, _21756_);
  and (_21759_, _21758_, _14963_);
  nor (_21760_, _21758_, _14963_);
  nor (_21761_, _21760_, _21759_);
  and (_21762_, _13738_, _13481_);
  nor (_21763_, _13738_, _13481_);
  or (_21765_, _21763_, _21762_);
  not (_21766_, _21765_);
  and (_21767_, _15286_, _14641_);
  nor (_21768_, _15286_, _14641_);
  or (_21769_, _21768_, _21767_);
  and (_21770_, _21769_, _21766_);
  nor (_21771_, _21769_, _21766_);
  nor (_21772_, _21771_, _21770_);
  nor (_21773_, _21772_, _21761_);
  and (_21774_, _21772_, _21761_);
  nor (_21776_, _21774_, _21773_);
  and (_21777_, _21776_, _06667_);
  nor (_21778_, _21776_, _06667_);
  or (_21779_, _21778_, _21777_);
  and (_21780_, _21779_, _02007_);
  or (_21781_, _21780_, _21755_);
  and (_21782_, _21781_, _01558_);
  and (_21783_, _21556_, _03279_);
  or (_21784_, _21783_, _21782_);
  or (_21785_, _21784_, _01999_);
  and (_21787_, _13696_, _13454_);
  nor (_21788_, _13696_, _13454_);
  nor (_21789_, _21788_, _21787_);
  and (_21790_, _21789_, _13971_);
  nor (_21791_, _21789_, _13971_);
  or (_21792_, _21791_, _21790_);
  and (_21793_, _21792_, _14291_);
  nor (_21794_, _21792_, _14291_);
  or (_21795_, _21794_, _21793_);
  not (_21796_, _15217_);
  nor (_21798_, _14903_, _14599_);
  and (_21799_, _14903_, _14599_);
  nor (_21800_, _21799_, _21798_);
  nor (_21801_, _21800_, _21796_);
  and (_21802_, _21800_, _21796_);
  nor (_21803_, _21802_, _21801_);
  nor (_21804_, _21803_, _21795_);
  and (_21805_, _21803_, _21795_);
  or (_21806_, _21805_, _21804_);
  nand (_21807_, _21806_, _06474_);
  or (_21809_, _21806_, _06474_);
  and (_21810_, _21809_, _21807_);
  or (_21811_, _21810_, _02840_);
  and (_21812_, _21811_, _06613_);
  and (_21813_, _21812_, _21785_);
  or (_21814_, _21688_, _02850_);
  and (_21815_, _21814_, _10157_);
  or (_21816_, _21815_, _21813_);
  or (_21817_, _21671_, _06675_);
  and (_21818_, _21817_, _02021_);
  and (_21820_, _21818_, _21816_);
  and (_21821_, _21652_, _02006_);
  or (_21822_, _21821_, _10165_);
  or (_21823_, _21822_, _21820_);
  or (_21824_, _21556_, _10163_);
  and (_21825_, _21824_, _02025_);
  and (_21826_, _21825_, _21823_);
  or (_21827_, _21826_, _21606_);
  and (_21828_, _10168_, _08537_);
  and (_21829_, _21828_, _21827_);
  not (_21831_, _21828_);
  nand (_21832_, _21831_, _21556_);
  nor (_21833_, _08493_, _02050_);
  and (_21834_, _08441_, _21833_);
  and (_21835_, _21834_, _09867_);
  nand (_21836_, _21835_, _21832_);
  or (_21837_, _21836_, _21829_);
  or (_21838_, _21835_, _21556_);
  and (_21839_, _21838_, _02861_);
  and (_21840_, _21839_, _21837_);
  not (_21842_, _14043_);
  and (_21843_, _21842_, _13761_);
  nor (_21844_, _21842_, _13761_);
  nor (_21845_, _21844_, _21843_);
  not (_21846_, _21845_);
  nor (_21847_, _14308_, _21729_);
  and (_21848_, _14308_, _21729_);
  nor (_21849_, _21848_, _21847_);
  not (_21850_, _21849_);
  not (_21851_, _14936_);
  and (_21853_, _21851_, _14664_);
  nor (_21854_, _21851_, _14664_);
  nor (_21855_, _21854_, _21853_);
  and (_21856_, _21855_, _21850_);
  nor (_21857_, _21855_, _21850_);
  nor (_21858_, _21857_, _21856_);
  nor (_21859_, _21858_, _21846_);
  and (_21860_, _21858_, _21846_);
  nor (_21861_, _21860_, _21859_);
  not (_21862_, _15309_);
  and (_21864_, _21862_, _06692_);
  nor (_21865_, _21862_, _06692_);
  nor (_21866_, _21865_, _21864_);
  nand (_21867_, _21866_, _21861_);
  or (_21868_, _21866_, _21861_);
  and (_21869_, _21868_, _01991_);
  nand (_21870_, _21869_, _21867_);
  nor (_21871_, _01992_, _03131_);
  and (_21872_, _21871_, _01988_);
  nand (_21873_, _21872_, _21870_);
  or (_21875_, _21873_, _21840_);
  or (_21876_, _21872_, _21556_);
  nand (_21877_, _21876_, _21875_);
  nor (_21878_, _10204_, _02871_);
  and (_21879_, _21878_, _01974_);
  nand (_21880_, _21879_, _21877_);
  or (_21881_, _21879_, _21556_);
  and (_21882_, _21881_, _05285_);
  and (_21883_, _21882_, _21880_);
  nor (_21884_, _01967_, _10213_);
  and (_21886_, _21884_, _07417_);
  nor (_21887_, _13767_, _13505_);
  and (_21888_, _13767_, _13505_);
  or (_21889_, _21888_, _21887_);
  nor (_21890_, _21889_, _14048_);
  and (_21891_, _21889_, _14048_);
  nor (_21892_, _21891_, _21890_);
  nor (_21893_, _21892_, _14364_);
  and (_21894_, _21892_, _14364_);
  or (_21895_, _21894_, _21893_);
  nor (_21897_, _21895_, _14669_);
  and (_21898_, _21895_, _14669_);
  or (_21899_, _21898_, _21897_);
  nor (_21900_, _21899_, _14988_);
  and (_21901_, _21899_, _14988_);
  or (_21902_, _21901_, _21900_);
  nor (_21903_, _21902_, _15314_);
  and (_21904_, _21902_, _15314_);
  or (_21905_, _21904_, _21903_);
  or (_21906_, _21905_, _06697_);
  nand (_21908_, _21905_, _06697_);
  and (_21909_, _21908_, _05279_);
  nand (_21910_, _21909_, _21906_);
  nand (_21911_, _21910_, _21886_);
  or (_21912_, _21911_, _21883_);
  or (_21913_, _21886_, _21556_);
  and (_21914_, _21913_, _08248_);
  and (_21915_, _21914_, _21912_);
  nand (_21916_, _21556_, _01966_);
  nand (_21917_, _21916_, _08771_);
  or (_21919_, _21917_, _21915_);
  not (_21920_, _06769_);
  nor (_21921_, _13776_, _13510_);
  and (_21922_, _13776_, _13510_);
  nor (_21923_, _21922_, _21921_);
  or (_21924_, _21923_, _14378_);
  nand (_21925_, _21923_, _14378_);
  and (_21926_, _21925_, _21924_);
  or (_21927_, _21926_, _14066_);
  nand (_21928_, _21926_, _14066_);
  and (_21930_, _21928_, _21927_);
  or (_21931_, _21930_, _14686_);
  nand (_21932_, _21930_, _14686_);
  and (_21933_, _21932_, _21931_);
  nor (_21934_, _21933_, _15004_);
  and (_21935_, _21933_, _15004_);
  or (_21936_, _21935_, _21934_);
  nor (_21937_, _21936_, _15256_);
  and (_21938_, _21936_, _15256_);
  or (_21939_, _21938_, _21937_);
  nor (_21941_, _21939_, _21920_);
  and (_21942_, _21939_, _21920_);
  or (_21943_, _21942_, _21941_);
  or (_21944_, _21943_, _08771_);
  and (_21945_, _21944_, _08778_);
  and (_21946_, _21945_, _21919_);
  and (_21947_, _21943_, _08777_);
  or (_21948_, _21947_, _06609_);
  or (_21949_, _21948_, _21946_);
  not (_21950_, _06608_);
  or (_21952_, _13784_, _13438_);
  nand (_21953_, _13784_, _13438_);
  and (_21954_, _21953_, _21952_);
  nor (_21955_, _21954_, _13987_);
  and (_21956_, _21954_, _13987_);
  or (_21957_, _21956_, _21955_);
  nor (_21958_, _21957_, _14303_);
  and (_21959_, _21957_, _14303_);
  or (_21960_, _21959_, _21958_);
  and (_21961_, _14931_, _14703_);
  nor (_21963_, _14931_, _14703_);
  or (_21964_, _21963_, _21961_);
  and (_21965_, _21964_, _21960_);
  nor (_21966_, _21964_, _21960_);
  nor (_21967_, _21966_, _21965_);
  nor (_21968_, _21967_, _15243_);
  and (_21969_, _21967_, _15243_);
  nor (_21970_, _21969_, _21968_);
  and (_21971_, _21970_, _21950_);
  nor (_21972_, _21970_, _21950_);
  or (_21974_, _21972_, _21971_);
  or (_21975_, _21974_, _08245_);
  and (_21976_, _21975_, _02036_);
  and (_21977_, _21976_, _21949_);
  not (_21978_, _06949_);
  nand (_21979_, _13704_, _13518_);
  or (_21980_, _13704_, _13518_);
  and (_21981_, _21980_, _21979_);
  and (_21982_, _21981_, _14081_);
  nor (_21983_, _21981_, _14081_);
  nor (_21985_, _21983_, _21982_);
  nor (_21986_, _21985_, _14394_);
  and (_21987_, _21985_, _14394_);
  or (_21988_, _21987_, _21986_);
  and (_21989_, _21988_, _14714_);
  nor (_21990_, _21988_, _14714_);
  nor (_21991_, _21990_, _21989_);
  nor (_21992_, _21991_, _15023_);
  and (_21993_, _21991_, _15023_);
  or (_21994_, _21993_, _21992_);
  and (_21996_, _21994_, _15229_);
  nor (_21997_, _21994_, _15229_);
  nor (_21998_, _21997_, _21996_);
  nand (_21999_, _21998_, _21978_);
  or (_22000_, _21998_, _21978_);
  and (_22001_, _22000_, _21999_);
  and (_22002_, _22001_, _01963_);
  or (_22003_, _22002_, _21977_);
  or (_22004_, _22003_, _06476_);
  and (_22005_, _22004_, _21581_);
  or (_22007_, _22005_, _01549_);
  nor (_22008_, _03621_, _01923_);
  nor (_22009_, _03631_, _03623_);
  nor (_22010_, _03642_, _03689_);
  nor (_22011_, _03627_, _03658_);
  nor (_22012_, _22011_, _22010_);
  and (_22013_, _22011_, _22010_);
  nor (_22014_, _22013_, _22012_);
  nor (_22015_, _22014_, _22009_);
  and (_22016_, _22014_, _22009_);
  nor (_22018_, _22016_, _22015_);
  not (_22019_, _22018_);
  nor (_22020_, _22019_, _22008_);
  and (_22021_, _22019_, _22008_);
  or (_22022_, _22021_, _22020_);
  or (_22023_, _22022_, _01550_);
  and (_22024_, _22023_, _02408_);
  and (_22025_, _22024_, _22007_);
  not (_22026_, _14416_);
  and (_22027_, _22026_, _14105_);
  nor (_22029_, _22026_, _14105_);
  nor (_22030_, _22029_, _22027_);
  nor (_22031_, _15033_, _14724_);
  and (_22032_, _15033_, _14724_);
  nor (_22033_, _22032_, _22031_);
  nor (_22034_, _22033_, _22030_);
  and (_22035_, _22033_, _22030_);
  nor (_22036_, _22035_, _22034_);
  and (_22037_, _13801_, _13531_);
  nor (_22038_, _13801_, _13531_);
  nor (_22040_, _22038_, _22037_);
  and (_22041_, _15340_, _06960_);
  nor (_22042_, _15340_, _06960_);
  nor (_22043_, _22042_, _22041_);
  not (_22044_, _22043_);
  and (_22045_, _22044_, _22040_);
  nor (_22046_, _22044_, _22040_);
  nor (_22047_, _22046_, _22045_);
  nand (_22048_, _22047_, _22036_);
  or (_22049_, _22047_, _22036_);
  and (_22051_, _22049_, _01875_);
  nand (_22052_, _22051_, _22048_);
  nor (_22053_, _02080_, _01604_);
  nand (_22054_, _22053_, _22052_);
  or (_22055_, _22054_, _22025_);
  or (_22056_, _22053_, _21556_);
  and (_22057_, _22056_, _05249_);
  and (_22058_, _22057_, _22055_);
  and (_22059_, _21810_, _05994_);
  or (_22060_, _22059_, _02528_);
  or (_22062_, _22060_, _22058_);
  not (_22063_, _15040_);
  and (_22064_, _22063_, _14731_);
  nor (_22065_, _22063_, _14731_);
  nor (_22066_, _22065_, _22064_);
  and (_22067_, _13808_, _13538_);
  nor (_22068_, _13808_, _13538_);
  nor (_22069_, _22068_, _22067_);
  and (_22070_, _22069_, _14112_);
  nor (_22071_, _22069_, _14112_);
  or (_22073_, _22071_, _22070_);
  and (_22074_, _22073_, _14423_);
  nor (_22075_, _22073_, _14423_);
  or (_22076_, _22075_, _22074_);
  nor (_22077_, _22076_, _22066_);
  and (_22078_, _22076_, _22066_);
  nor (_22079_, _22078_, _22077_);
  and (_22080_, _22079_, _15347_);
  nor (_22081_, _22079_, _15347_);
  or (_22082_, _22081_, _22080_);
  nor (_22084_, _22082_, _06967_);
  and (_22085_, _22082_, _06967_);
  or (_22086_, _22085_, _02888_);
  or (_22087_, _22086_, _22084_);
  and (_22088_, _22087_, _02043_);
  and (_22089_, _22088_, _22062_);
  and (_22090_, _13813_, _13543_);
  nor (_22091_, _13813_, _13543_);
  nor (_22092_, _22091_, _22090_);
  and (_22093_, _22092_, _14117_);
  nor (_22095_, _22092_, _14117_);
  or (_22096_, _22095_, _22093_);
  nand (_22097_, _22096_, _14428_);
  or (_22098_, _22096_, _14428_);
  and (_22099_, _22098_, _22097_);
  nor (_22100_, _15352_, _15045_);
  and (_22101_, _15352_, _15045_);
  nor (_22102_, _22101_, _22100_);
  not (_22103_, _14736_);
  and (_22104_, _22103_, _06972_);
  nor (_22106_, _22103_, _06972_);
  nor (_22107_, _22106_, _22104_);
  nor (_22108_, _22107_, _22102_);
  and (_22109_, _22107_, _22102_);
  nor (_22110_, _22109_, _22108_);
  nand (_22111_, _22110_, _22099_);
  or (_22112_, _22110_, _22099_);
  and (_22113_, _22112_, _01602_);
  and (_22114_, _22113_, _22111_);
  or (_22115_, _22114_, _06008_);
  or (_22117_, _22115_, _22089_);
  and (_22118_, _06059_, _15357_);
  nor (_22119_, _06059_, _15357_);
  nor (_22120_, _22119_, _22118_);
  not (_22121_, _22120_);
  nor (_22122_, _06146_, _06097_);
  and (_22123_, _06146_, _06097_);
  nor (_22124_, _22123_, _22122_);
  not (_22125_, _22124_);
  and (_22126_, _22125_, _06198_);
  nor (_22128_, _22125_, _06198_);
  nor (_22129_, _22128_, _22126_);
  and (_22130_, _22129_, _22121_);
  nor (_22131_, _22129_, _22121_);
  nor (_22132_, _22131_, _22130_);
  nor (_22133_, _06274_, _06977_);
  and (_22134_, _06274_, _06977_);
  nor (_22135_, _22134_, _22133_);
  and (_22136_, _22135_, _22132_);
  nor (_22137_, _22135_, _22132_);
  nor (_22139_, _22137_, _22136_);
  not (_22140_, _22139_);
  nor (_22141_, _22140_, _06353_);
  and (_22142_, _22140_, _06353_);
  or (_22143_, _22142_, _06355_);
  or (_22144_, _22143_, _22141_);
  and (_22145_, _22144_, _01609_);
  and (_22146_, _22145_, _22117_);
  nand (_22147_, _22022_, _01608_);
  and (_22148_, _01977_, _01637_);
  and (_22150_, _02065_, _01637_);
  nor (_22151_, _22150_, _22148_);
  and (_22152_, _10254_, _10247_);
  and (_22153_, _22152_, _22151_);
  nand (_22154_, _22153_, _22147_);
  or (_22155_, _22154_, _22146_);
  or (_22156_, _22153_, _21556_);
  nand (_22157_, _22156_, _22155_);
  nor (_22158_, _02899_, _02895_);
  nand (_22159_, _22158_, _22157_);
  or (_22161_, _22158_, _21556_);
  and (_22162_, _22161_, _01870_);
  and (_22163_, _22162_, _22159_);
  nor (_22164_, _14439_, _14128_);
  and (_22165_, _14439_, _14128_);
  nor (_22166_, _22165_, _22164_);
  nor (_22167_, _13824_, _13554_);
  and (_22168_, _13824_, _13554_);
  or (_22169_, _22168_, _22167_);
  nor (_22170_, _22169_, _22166_);
  and (_22172_, _22169_, _22166_);
  nor (_22173_, _22172_, _22170_);
  not (_22174_, _15365_);
  nor (_22175_, _15056_, _14747_);
  and (_22176_, _15056_, _14747_);
  nor (_22177_, _22176_, _22175_);
  nor (_22178_, _22177_, _22174_);
  and (_22179_, _22177_, _22174_);
  nor (_22180_, _22179_, _22178_);
  nor (_22181_, _22180_, _22173_);
  and (_22183_, _22180_, _22173_);
  or (_22184_, _22183_, _22181_);
  or (_22185_, _22184_, _06466_);
  nand (_22186_, _22184_, _06466_);
  and (_22187_, _22186_, _01869_);
  and (_22188_, _22187_, _22185_);
  or (_22189_, _22188_, _22163_);
  and (_22190_, _22189_, _06985_);
  nand (_22191_, _22022_, _06984_);
  and (_22192_, _10306_, _10268_);
  and (_22194_, _22192_, _10311_);
  nand (_22195_, _22194_, _22191_);
  or (_22196_, _22195_, _22190_);
  and (_22197_, _14276_, _06427_);
  nor (_22198_, _14276_, _06427_);
  nor (_22199_, _22198_, _22197_);
  and (_22200_, _13561_, _06432_);
  nor (_22201_, _22200_, _14059_);
  nor (_22202_, _22201_, _22199_);
  and (_22203_, _22201_, _22199_);
  nor (_22205_, _22203_, _22202_);
  and (_22206_, _06419_, _06415_);
  nor (_22207_, _06419_, _06415_);
  nor (_22208_, _22207_, _22206_);
  nor (_22209_, _22208_, _22205_);
  and (_22210_, _22208_, _22205_);
  nor (_22211_, _22210_, _22209_);
  nand (_22212_, _22211_, _15214_);
  or (_22213_, _22211_, _15214_);
  and (_22214_, _22213_, _22212_);
  nor (_22216_, _22214_, _06408_);
  and (_22217_, _22214_, _06408_);
  or (_22218_, _22217_, _22216_);
  or (_22219_, _22218_, _10325_);
  or (_22220_, _22194_, _21556_);
  and (_22221_, _22220_, _10323_);
  and (_22222_, _22221_, _22219_);
  and (_22223_, _22222_, _22196_);
  and (_22224_, _22218_, _13828_);
  or (_22225_, _22224_, _02579_);
  or (_22227_, _22225_, _22223_);
  nor (_22228_, _14288_, _07229_);
  and (_22229_, _14288_, _07229_);
  nor (_22230_, _22229_, _22228_);
  and (_22231_, _13573_, _07233_);
  nor (_22232_, _22231_, _13980_);
  nor (_22233_, _22232_, _22230_);
  and (_22234_, _22232_, _22230_);
  nor (_22235_, _22234_, _22233_);
  nor (_22236_, _07218_, _07222_);
  and (_22238_, _07218_, _07222_);
  nor (_22239_, _22238_, _22236_);
  nor (_22240_, _22239_, _22235_);
  and (_22241_, _22239_, _22235_);
  nor (_22242_, _22241_, _22240_);
  nor (_22243_, _22242_, _07215_);
  and (_22244_, _22242_, _07215_);
  or (_22245_, _22244_, _22243_);
  nor (_22246_, _22245_, _07008_);
  and (_22247_, _22245_, _07008_);
  or (_22249_, _22247_, _22246_);
  or (_22250_, _22249_, _07006_);
  and (_22251_, _22250_, _07014_);
  and (_22252_, _22251_, _22227_);
  and (_22253_, _10822_, _10620_);
  nor (_22254_, _10822_, _10620_);
  or (_22255_, _22254_, _22253_);
  nor (_22256_, _11094_, _11020_);
  and (_22257_, _11094_, _11020_);
  nor (_22258_, _22257_, _22256_);
  nor (_22260_, _22258_, _22255_);
  and (_22261_, _22258_, _22255_);
  nor (_22262_, _22261_, _22260_);
  not (_22263_, _22262_);
  nor (_22264_, _11635_, _11431_);
  and (_22265_, _11635_, _11431_);
  nor (_22266_, _22265_, _22264_);
  nor (_22267_, _11709_, _04779_);
  and (_22268_, _11709_, _04779_);
  nor (_22269_, _22268_, _22267_);
  not (_22271_, _22269_);
  and (_22272_, _22271_, _22266_);
  nor (_22273_, _22271_, _22266_);
  nor (_22274_, _22273_, _22272_);
  nor (_22275_, _22274_, _22263_);
  and (_22276_, _22274_, _22263_);
  or (_22277_, _22276_, _07012_);
  or (_22278_, _22277_, _22275_);
  and (_22279_, _22278_, _10330_);
  or (_22280_, _22279_, _22252_);
  and (_22282_, _15165_, _07308_);
  nor (_22283_, _15165_, _07308_);
  nor (_22284_, _22283_, _22282_);
  and (_22285_, _08661_, _07322_);
  nor (_22286_, _22285_, _08662_);
  nor (_22287_, _22286_, _07318_);
  and (_22288_, _22286_, _07318_);
  nor (_22289_, _22288_, _22287_);
  and (_22290_, _07313_, _08629_);
  nor (_22291_, _07313_, _08629_);
  nor (_22293_, _22291_, _22290_);
  nor (_22294_, _22293_, _22289_);
  and (_22295_, _22293_, _22289_);
  nor (_22296_, _22295_, _22294_);
  nor (_22297_, _22296_, _22284_);
  and (_22298_, _22296_, _22284_);
  or (_22299_, _22298_, _22297_);
  or (_22300_, _22299_, _07020_);
  nand (_22301_, _22299_, _07020_);
  and (_22302_, _22301_, _22300_);
  or (_22304_, _22302_, _07013_);
  and (_22305_, _22304_, _02166_);
  and (_22306_, _22305_, _22280_);
  nor (_22307_, _13693_, _13584_);
  and (_22308_, _13693_, _13584_);
  nor (_22309_, _22308_, _22307_);
  and (_22310_, _22309_, _13968_);
  nor (_22311_, _22309_, _13968_);
  or (_22312_, _22311_, _22310_);
  nand (_22313_, _22312_, _14286_);
  or (_22315_, _22312_, _14286_);
  and (_22316_, _22315_, _22313_);
  nor (_22317_, _15210_, _14894_);
  and (_22318_, _15210_, _14894_);
  nor (_22319_, _22318_, _22317_);
  not (_22320_, _14596_);
  and (_22321_, _22320_, _06470_);
  nor (_22322_, _22320_, _06470_);
  nor (_22323_, _22322_, _22321_);
  nor (_22324_, _22323_, _22319_);
  and (_22326_, _22323_, _22319_);
  nor (_22327_, _22326_, _22324_);
  nand (_22328_, _22327_, _22316_);
  or (_22329_, _22327_, _22316_);
  and (_22330_, _22329_, _02079_);
  and (_22331_, _22330_, _22328_);
  or (_22332_, _22331_, _22306_);
  and (_22333_, _22332_, _02912_);
  nand (_22334_, _21556_, _02167_);
  or (_22335_, _22334_, _03680_);
  nor (_22337_, _10343_, _01645_);
  nand (_22338_, _22337_, _22335_);
  or (_22339_, _22338_, _22333_);
  or (_22340_, _22337_, _21556_);
  and (_22341_, _22340_, _07027_);
  and (_22342_, _22341_, _22339_);
  not (_22343_, _06407_);
  or (_22344_, _06433_, _06429_);
  nand (_22345_, _06433_, _06429_);
  and (_22346_, _22345_, _22344_);
  nor (_22348_, _06425_, _06424_);
  and (_22349_, _06425_, _06424_);
  nor (_22350_, _22349_, _22348_);
  not (_22351_, _22350_);
  and (_22352_, _22351_, _22346_);
  nor (_22353_, _22351_, _22346_);
  nor (_22354_, _22353_, _22352_);
  nor (_22355_, _06417_, _06413_);
  and (_22356_, _06417_, _06413_);
  nor (_22357_, _22356_, _22355_);
  nor (_22359_, _22357_, _06410_);
  and (_22360_, _22357_, _06410_);
  nor (_22361_, _22360_, _22359_);
  not (_22362_, _22361_);
  and (_22363_, _22362_, _22354_);
  nor (_22364_, _22362_, _22354_);
  or (_22365_, _22364_, _22363_);
  nor (_22366_, _22365_, _22343_);
  and (_22367_, _22365_, _22343_);
  or (_22368_, _22367_, _22366_);
  and (_22370_, _22368_, _07026_);
  or (_22371_, _22370_, _07031_);
  or (_22372_, _22371_, _22342_);
  not (_22373_, _07007_);
  or (_22374_, _07234_, _07231_);
  nand (_22375_, _07234_, _07231_);
  and (_22376_, _22375_, _22374_);
  and (_22377_, _07226_, _07227_);
  nor (_22378_, _07226_, _07227_);
  nor (_22379_, _22378_, _22377_);
  and (_22381_, _22379_, _22376_);
  nor (_22382_, _22379_, _22376_);
  nor (_22383_, _22382_, _22381_);
  nor (_22384_, _07216_, _07220_);
  and (_22385_, _07216_, _07220_);
  nor (_22386_, _22385_, _22384_);
  nor (_22387_, _22386_, _07213_);
  and (_22388_, _22386_, _07213_);
  nor (_22389_, _22388_, _22387_);
  nor (_22390_, _22389_, _22383_);
  and (_22392_, _22389_, _22383_);
  or (_22393_, _22392_, _22390_);
  nor (_22394_, _22393_, _22373_);
  and (_22395_, _22393_, _22373_);
  or (_22396_, _22395_, _22394_);
  or (_22397_, _22396_, _07036_);
  and (_22398_, _22397_, _07035_);
  and (_22399_, _22398_, _22372_);
  nor (_22400_, _10820_, _10618_);
  and (_22401_, _10820_, _10618_);
  nor (_22403_, _22401_, _22400_);
  not (_22404_, _11092_);
  and (_22405_, _22404_, _11018_);
  nor (_22406_, _22404_, _11018_);
  nor (_22407_, _22406_, _22405_);
  and (_22408_, _22407_, _22403_);
  nor (_22409_, _22407_, _22403_);
  nor (_22410_, _22409_, _22408_);
  not (_22411_, _11707_);
  nor (_22412_, _11633_, _11429_);
  and (_22414_, _11633_, _11429_);
  nor (_22415_, _22414_, _22412_);
  nor (_22416_, _22415_, _22411_);
  and (_22417_, _22415_, _22411_);
  nor (_22418_, _22417_, _22416_);
  and (_22419_, _22418_, _22410_);
  nor (_22420_, _22418_, _22410_);
  or (_22421_, _22420_, _22419_);
  nor (_22422_, _22421_, _04777_);
  and (_22423_, _22421_, _04777_);
  or (_22425_, _22423_, _07040_);
  or (_22426_, _22425_, _22422_);
  and (_22427_, _22426_, _07042_);
  or (_22428_, _22427_, _22399_);
  not (_22429_, _07311_);
  or (_22430_, _07323_, _07320_);
  nand (_22431_, _07323_, _07320_);
  and (_22432_, _22431_, _22430_);
  not (_22433_, _07314_);
  and (_22434_, _22433_, _07316_);
  nor (_22436_, _22433_, _07316_);
  nor (_22437_, _22436_, _22434_);
  not (_22438_, _22437_);
  and (_22439_, _22438_, _22432_);
  nor (_22440_, _22438_, _22432_);
  nor (_22441_, _22440_, _22439_);
  nand (_22442_, _22441_, _22429_);
  or (_22443_, _22441_, _22429_);
  and (_22444_, _22443_, _22442_);
  or (_22445_, _22444_, _07309_);
  nand (_22447_, _22444_, _07309_);
  and (_22448_, _22447_, _22445_);
  or (_22449_, _22448_, _07306_);
  nand (_22450_, _22448_, _07306_);
  and (_22451_, _22450_, _22449_);
  and (_22452_, _22451_, _07018_);
  nor (_22453_, _22451_, _07018_);
  or (_22454_, _22453_, _22452_);
  or (_22455_, _22454_, _07046_);
  and (_22456_, _22455_, _02176_);
  and (_22458_, _22456_, _22428_);
  and (_22459_, _10364_, _09292_);
  nor (_22460_, _14176_, _13605_);
  and (_22461_, _14176_, _13605_);
  nor (_22462_, _22461_, _22460_);
  nor (_22463_, _15406_, _14795_);
  and (_22464_, _15406_, _14795_);
  nor (_22465_, _22464_, _22463_);
  and (_22466_, _22465_, _22462_);
  nor (_22467_, _22465_, _22462_);
  nor (_22469_, _22467_, _22466_);
  or (_22470_, _14489_, _13689_);
  nand (_22471_, _14489_, _13689_);
  and (_22472_, _22471_, _22470_);
  or (_22473_, _22472_, _15105_);
  nand (_22474_, _22472_, _15105_);
  and (_22475_, _22474_, _22473_);
  and (_22476_, _22475_, _06467_);
  nor (_22477_, _22475_, _06467_);
  or (_22478_, _22477_, _22476_);
  nand (_22480_, _22478_, _22469_);
  or (_22481_, _22478_, _22469_);
  and (_22482_, _22481_, _02072_);
  nand (_22483_, _22482_, _22480_);
  nand (_22484_, _22483_, _22459_);
  or (_22485_, _22484_, _22458_);
  nor (_22486_, _21556_, _22459_);
  nor (_22487_, _22486_, _14591_);
  and (_22488_, _22487_, _22485_);
  nor (_22489_, _13440_, _06430_);
  and (_22491_, _13440_, _06430_);
  nor (_22492_, _22491_, _22489_);
  and (_22493_, _14180_, _06421_);
  and (_22494_, _06426_, _06422_);
  nor (_22495_, _22494_, _22493_);
  and (_22496_, _22495_, _22492_);
  nor (_22497_, _22495_, _22492_);
  nor (_22498_, _22497_, _22496_);
  not (_22499_, _06414_);
  nor (_22500_, _06418_, _06411_);
  and (_22502_, _06418_, _06411_);
  nor (_22503_, _22502_, _22500_);
  nor (_22504_, _22503_, _22499_);
  and (_22505_, _22503_, _22499_);
  nor (_22506_, _22505_, _22504_);
  and (_22507_, _22506_, _22498_);
  nor (_22508_, _22506_, _22498_);
  or (_22509_, _22508_, _22507_);
  and (_22510_, _22509_, _06406_);
  nor (_22511_, _22509_, _06406_);
  or (_22513_, _22511_, _22510_);
  and (_22514_, _22513_, _14591_);
  or (_22515_, _22514_, _06462_);
  or (_22516_, _22515_, _22488_);
  nor (_22517_, _13572_, _07232_);
  and (_22518_, _13572_, _07232_);
  nor (_22519_, _22518_, _22517_);
  not (_22520_, _22519_);
  and (_22521_, _07224_, _07228_);
  nor (_22522_, _07224_, _07228_);
  nor (_22524_, _22522_, _22521_);
  nor (_22525_, _22524_, _22520_);
  and (_22526_, _22524_, _22520_);
  nor (_22527_, _22526_, _22525_);
  not (_22528_, _07217_);
  nor (_22529_, _07221_, _07214_);
  and (_22530_, _07221_, _07214_);
  nor (_22531_, _22530_, _22529_);
  nor (_22532_, _22531_, _22528_);
  and (_22533_, _22531_, _22528_);
  nor (_22535_, _22533_, _22532_);
  nor (_22536_, _22535_, _22527_);
  and (_22537_, _22535_, _22527_);
  nor (_22538_, _22537_, _22536_);
  and (_22539_, _22538_, _06461_);
  nor (_22540_, _22538_, _06461_);
  or (_22541_, _22540_, _22539_);
  or (_22542_, _22541_, _09855_);
  and (_22543_, _22542_, _02172_);
  and (_22544_, _22543_, _22516_);
  nor (_22546_, _10821_, _10619_);
  and (_22547_, _10821_, _10619_);
  nor (_22548_, _22547_, _22546_);
  and (_22549_, _22548_, _11019_);
  nor (_22550_, _22548_, _11019_);
  or (_22551_, _22550_, _22549_);
  nand (_22552_, _22551_, _11093_);
  or (_22553_, _22551_, _11093_);
  and (_22554_, _22553_, _22552_);
  nor (_22555_, _11634_, _11430_);
  and (_22557_, _11634_, _11430_);
  nor (_22558_, _22557_, _22555_);
  nor (_22559_, _22558_, _11708_);
  and (_22560_, _22558_, _11708_);
  nor (_22561_, _22560_, _22559_);
  not (_22562_, _22561_);
  nor (_22563_, _22562_, _22554_);
  and (_22564_, _22562_, _22554_);
  nor (_22565_, _22564_, _22563_);
  or (_22566_, _22565_, _04778_);
  nand (_22568_, _22565_, _04778_);
  and (_22569_, _22568_, _02171_);
  and (_22570_, _22569_, _22566_);
  or (_22571_, _22570_, _07069_);
  or (_22572_, _22571_, _22544_);
  nor (_22573_, _08660_, _07321_);
  and (_22574_, _08660_, _07321_);
  nor (_22575_, _22574_, _22573_);
  not (_22576_, _07315_);
  and (_22577_, _22576_, _07317_);
  nor (_22579_, _22576_, _07317_);
  nor (_22580_, _22579_, _22577_);
  and (_22581_, _22580_, _22575_);
  nor (_22582_, _22580_, _22575_);
  nor (_22583_, _22582_, _22581_);
  not (_22584_, _07312_);
  nor (_22585_, _07310_, _07307_);
  and (_22586_, _07310_, _07307_);
  nor (_22587_, _22586_, _22585_);
  nor (_22588_, _22587_, _22584_);
  and (_22590_, _22587_, _22584_);
  nor (_22591_, _22590_, _22588_);
  and (_22592_, _22591_, _22583_);
  nor (_22593_, _22591_, _22583_);
  or (_22594_, _22593_, _22592_);
  nor (_22595_, _22594_, _07019_);
  and (_22596_, _22594_, _07019_);
  or (_22597_, _22596_, _22595_);
  or (_22598_, _22597_, _07070_);
  and (_22599_, _22598_, _04788_);
  and (_22601_, _22599_, _22572_);
  and (_22602_, _09850_, _09849_);
  not (_22603_, _15427_);
  and (_22604_, _22603_, _07078_);
  nor (_22605_, _22603_, _07078_);
  nor (_22606_, _22605_, _22604_);
  not (_22607_, _14890_);
  and (_22608_, _22607_, _14810_);
  nor (_22609_, _22607_, _14810_);
  nor (_22610_, _22609_, _22608_);
  not (_22612_, _22610_);
  nor (_22613_, _13885_, _13627_);
  and (_22614_, _13885_, _13627_);
  or (_22615_, _22614_, _22613_);
  and (_22616_, _22615_, _14199_);
  nor (_22617_, _22615_, _14199_);
  or (_22618_, _22617_, _22616_);
  nand (_22619_, _22618_, _14283_);
  or (_22620_, _22618_, _14283_);
  and (_22621_, _22620_, _22619_);
  nor (_22623_, _22621_, _22612_);
  and (_22624_, _22621_, _22612_);
  nor (_22625_, _22624_, _22623_);
  and (_22626_, _22625_, _22606_);
  nor (_22627_, _22625_, _22606_);
  or (_22628_, _22627_, _04788_);
  or (_22629_, _22628_, _22626_);
  nand (_22630_, _22629_, _22602_);
  or (_22631_, _22630_, _22601_);
  or (_22632_, _21556_, _22602_);
  and (_22634_, _22632_, _07084_);
  and (_22635_, _22634_, _22631_);
  nor (_22636_, _13890_, _13510_);
  and (_22637_, _13890_, _13510_);
  or (_22638_, _22637_, _22636_);
  nor (_22639_, _22638_, _14204_);
  and (_22640_, _22638_, _14204_);
  nor (_22641_, _22640_, _22639_);
  nor (_22642_, _22641_, _14512_);
  and (_22643_, _22641_, _14512_);
  or (_22645_, _22643_, _22642_);
  nor (_22646_, _22645_, _14815_);
  and (_22647_, _22645_, _14815_);
  or (_22648_, _22647_, _22646_);
  and (_22649_, _22648_, _15124_);
  nor (_22650_, _22648_, _15124_);
  or (_22651_, _22650_, _22649_);
  nor (_22652_, _22651_, _15432_);
  and (_22653_, _22651_, _15432_);
  or (_22654_, _22653_, _22652_);
  not (_22656_, _22654_);
  nor (_22657_, _22656_, _07111_);
  and (_22658_, _22656_, _07111_);
  or (_22659_, _22658_, _22657_);
  and (_22660_, _22659_, _07085_);
  or (_22661_, _22660_, _07114_);
  or (_22662_, _22661_, _22635_);
  nor (_22663_, _13895_, _13438_);
  and (_22664_, _13895_, _13438_);
  or (_22665_, _22664_, _22663_);
  nor (_22667_, _22665_, _13961_);
  and (_22668_, _22665_, _13961_);
  nor (_22669_, _22668_, _22667_);
  nor (_22670_, _22669_, _14517_);
  and (_22671_, _22669_, _14517_);
  or (_22672_, _22671_, _22670_);
  nor (_22673_, _22672_, _14820_);
  and (_22674_, _22672_, _14820_);
  or (_22675_, _22674_, _22673_);
  and (_22676_, _22675_, _15129_);
  nor (_22677_, _22675_, _15129_);
  nor (_22678_, _22677_, _22676_);
  and (_22679_, _22678_, _15437_);
  nor (_22680_, _22678_, _15437_);
  or (_22681_, _22680_, _22679_);
  and (_22682_, _22681_, _07140_);
  nor (_22683_, _22681_, _07140_);
  or (_22684_, _22683_, _22682_);
  or (_22685_, _22684_, _07116_);
  and (_22686_, _22685_, _02165_);
  and (_22688_, _22686_, _22662_);
  and (_22689_, _13900_, _13518_);
  nor (_22690_, _13900_, _13518_);
  nor (_22691_, _22690_, _22689_);
  nor (_22692_, _22691_, _14211_);
  and (_22693_, _22691_, _14211_);
  nor (_22694_, _22693_, _22692_);
  and (_22695_, _22694_, _14522_);
  nor (_22696_, _22694_, _14522_);
  nor (_22697_, _22696_, _22695_);
  nor (_22699_, _22697_, _14825_);
  and (_22700_, _22697_, _14825_);
  or (_22701_, _22700_, _22699_);
  nor (_22702_, _22701_, _15134_);
  and (_22703_, _22701_, _15134_);
  or (_22704_, _22703_, _22702_);
  and (_22705_, _22704_, _15442_);
  nor (_22706_, _22704_, _15442_);
  or (_22707_, _22706_, _22705_);
  nand (_22708_, _22707_, _07171_);
  or (_22710_, _22707_, _07171_);
  and (_22711_, _22710_, _02164_);
  and (_22712_, _22711_, _22708_);
  or (_22713_, _22712_, _07144_);
  or (_22714_, _22713_, _22688_);
  nor (_22715_, _13905_, _13523_);
  and (_22716_, _13905_, _13523_);
  or (_22717_, _22716_, _22715_);
  nor (_22718_, _22717_, _14216_);
  and (_22719_, _22717_, _14216_);
  nor (_22721_, _22719_, _22718_);
  and (_22722_, _22721_, _14527_);
  nor (_22723_, _22721_, _14527_);
  nor (_22724_, _22723_, _22722_);
  nor (_22725_, _22724_, _14588_);
  and (_22726_, _22724_, _14588_);
  or (_22727_, _22726_, _22725_);
  nor (_22728_, _22727_, _15139_);
  and (_22729_, _22727_, _15139_);
  or (_22730_, _22729_, _22728_);
  nor (_22732_, _22730_, _15447_);
  and (_22733_, _22730_, _15447_);
  or (_22734_, _22733_, _22732_);
  nor (_22735_, _22734_, _07202_);
  and (_22736_, _22734_, _07202_);
  or (_22737_, _22736_, _07177_);
  or (_22738_, _22737_, _22735_);
  and (_22739_, _22738_, _07176_);
  and (_22740_, _22739_, _22714_);
  nor (_22741_, _13699_, _13698_);
  nor (_22743_, _14012_, \oc8051_golden_model_1.ACC [3]);
  and (_22744_, _14012_, \oc8051_golden_model_1.ACC [3]);
  nor (_22745_, _22744_, _22743_);
  and (_22746_, _22745_, _21712_);
  nor (_22747_, _22745_, _21712_);
  nor (_22748_, _22747_, _22746_);
  not (_22749_, _22748_);
  nand (_22750_, _22749_, _22741_);
  or (_22751_, _22749_, _22741_);
  and (_22752_, _22751_, _22750_);
  nand (_22754_, _22752_, _07175_);
  nor (_22755_, _02185_, _01636_);
  and (_22756_, _22755_, _10403_);
  nand (_22757_, _22756_, _22754_);
  or (_22758_, _22757_, _22740_);
  or (_22759_, _22756_, _21556_);
  and (_22760_, _22759_, _06458_);
  and (_22761_, _22760_, _22758_);
  not (_22762_, _13440_);
  and (_22763_, _22762_, _06432_);
  nor (_22765_, _22762_, _06432_);
  nor (_22766_, _22765_, _22763_);
  and (_22767_, _22766_, _14224_);
  nor (_22768_, _22766_, _14224_);
  nor (_22769_, _22768_, _22767_);
  and (_22770_, _22769_, _14279_);
  nor (_22771_, _22769_, _14279_);
  nor (_22772_, _22771_, _22770_);
  and (_22773_, _22772_, _14835_);
  nor (_22774_, _22772_, _14835_);
  nor (_22776_, _22774_, _22773_);
  and (_22777_, _22776_, _15148_);
  nor (_22778_, _22776_, _15148_);
  nor (_22779_, _22778_, _22777_);
  nor (_22780_, _22779_, _15455_);
  and (_22781_, _22779_, _15455_);
  or (_22782_, _22781_, _22780_);
  and (_22783_, _22782_, _06449_);
  nor (_22784_, _22782_, _06449_);
  or (_22785_, _22784_, _22783_);
  and (_22787_, _22785_, _06459_);
  or (_22788_, _22787_, _07210_);
  or (_22789_, _22788_, _22761_);
  not (_22790_, _13572_);
  and (_22791_, _22790_, _07233_);
  nor (_22792_, _22790_, _07233_);
  nor (_22793_, _22792_, _22791_);
  and (_22794_, _22793_, _14229_);
  nor (_22795_, _22793_, _14229_);
  nor (_22796_, _22795_, _22794_);
  and (_22798_, _22796_, _14538_);
  nor (_22799_, _22796_, _14538_);
  nor (_22800_, _22799_, _22798_);
  and (_22801_, _22800_, _14840_);
  nor (_22802_, _22800_, _14840_);
  nor (_22803_, _22802_, _22801_);
  nor (_22804_, _22803_, _15156_);
  and (_22805_, _22803_, _15156_);
  or (_22806_, _22805_, _22804_);
  and (_22807_, _22806_, _15460_);
  nor (_22809_, _22806_, _15460_);
  or (_22810_, _22809_, _22807_);
  nor (_22811_, _22810_, _07249_);
  and (_22812_, _22810_, _07249_);
  or (_22813_, _22812_, _07212_);
  or (_22814_, _22813_, _22811_);
  and (_22815_, _22814_, _07254_);
  and (_22816_, _22815_, _22789_);
  nor (_22817_, _13923_, _08622_);
  and (_22818_, _13923_, _08622_);
  or (_22820_, _22818_, _22817_);
  and (_22821_, _22820_, _14234_);
  nor (_22822_, _22820_, _14234_);
  nor (_22823_, _22822_, _22821_);
  and (_22824_, _22823_, _14544_);
  nor (_22825_, _22823_, _14544_);
  or (_22826_, _22825_, _22824_);
  nor (_22827_, _22826_, _14845_);
  and (_22828_, _22826_, _14845_);
  or (_22829_, _22828_, _22827_);
  nor (_22831_, _22829_, _15161_);
  and (_22832_, _22829_, _15161_);
  or (_22833_, _22832_, _22831_);
  nor (_22834_, _22833_, _15465_);
  and (_22835_, _22833_, _15465_);
  or (_22836_, _22835_, _22834_);
  and (_22837_, _22836_, _07300_);
  nor (_22838_, _22836_, _07300_);
  or (_22839_, _22838_, _22837_);
  and (_22840_, _22839_, _01890_);
  nor (_22842_, _08660_, _07322_);
  and (_22843_, _08660_, _07322_);
  nor (_22844_, _22843_, _22842_);
  nor (_22845_, _22844_, _14239_);
  and (_22846_, _22844_, _14239_);
  or (_22847_, _22846_, _22845_);
  and (_22848_, _22847_, _14550_);
  nor (_22849_, _22847_, _14550_);
  nor (_22850_, _22849_, _22848_);
  nor (_22851_, _22850_, _14850_);
  and (_22853_, _22850_, _14850_);
  or (_22854_, _22853_, _22851_);
  and (_22855_, _22854_, _15168_);
  nor (_22856_, _22854_, _15168_);
  nor (_22857_, _22856_, _22855_);
  nor (_22858_, _22857_, _15470_);
  and (_22859_, _22857_, _15470_);
  nor (_22860_, _22859_, _22858_);
  nand (_22861_, _22860_, _07338_);
  or (_22862_, _22860_, _07338_);
  and (_22864_, _22862_, _22861_);
  nand (_22865_, _22864_, _07253_);
  nor (_22866_, _02082_, _01653_);
  nor (_22867_, _07304_, _01888_);
  and (_22868_, _22867_, _22866_);
  nand (_22869_, _22868_, _22865_);
  or (_22870_, _22869_, _22840_);
  or (_22871_, _22870_, _22816_);
  or (_22872_, _22868_, _21556_);
  and (_22873_, _22872_, _10438_);
  and (_22875_, _22873_, _22871_);
  and (_22876_, _21556_, _10435_);
  or (_22877_, _22876_, _02201_);
  or (_22878_, _22877_, _22875_);
  or (_22879_, _21746_, _02303_);
  and (_22880_, _22879_, _07346_);
  and (_22881_, _22880_, _22878_);
  not (_22882_, _07351_);
  and (_22883_, _14012_, _22882_);
  and (_22884_, _22883_, \oc8051_golden_model_1.ACC [3]);
  nor (_22886_, _22883_, \oc8051_golden_model_1.ACC [3]);
  nor (_22887_, _22886_, _22884_);
  and (_22888_, _22887_, _14862_);
  nor (_22889_, _22887_, _14862_);
  nor (_22890_, _22889_, _22888_);
  and (_22891_, _15178_, _06026_);
  nor (_22892_, _15178_, _06026_);
  nor (_22893_, _22892_, _22891_);
  nor (_22894_, _22893_, _22890_);
  and (_22895_, _22893_, _22890_);
  or (_22897_, _22895_, _22894_);
  nor (_22898_, _22897_, _07357_);
  and (_22899_, _22897_, _07357_);
  or (_22900_, _22899_, _22898_);
  and (_22901_, _22900_, _07345_);
  or (_22902_, _22901_, _22881_);
  and (_22903_, _22902_, _08922_);
  and (_22904_, \oc8051_golden_model_1.PSW [7], \oc8051_golden_model_1.ACC [7]);
  nor (_22905_, _22904_, _06658_);
  or (_22906_, _22905_, _22748_);
  nand (_22908_, _22905_, _22748_);
  and (_22909_, _22908_, _22906_);
  nand (_22910_, _22909_, _07350_);
  nand (_22911_, _22910_, _02942_);
  or (_22912_, _22911_, _22903_);
  or (_22913_, _21556_, _02942_);
  and (_22914_, _22913_, _01887_);
  and (_22915_, _22914_, _22912_);
  and (_22916_, _21605_, _01860_);
  or (_22917_, _22916_, _05171_);
  or (_22919_, _22917_, _22915_);
  and (_22920_, _22919_, _21557_);
  or (_22921_, _22920_, _02952_);
  or (_22922_, _21556_, _05178_);
  and (_22923_, _22922_, _01538_);
  and (_22924_, _22923_, _22921_);
  not (_22925_, _14572_);
  nor (_22926_, _14873_, _22925_);
  and (_22927_, _14873_, _22925_);
  nor (_22928_, _22927_, _22926_);
  nor (_22930_, _22928_, _15491_);
  and (_22931_, _22928_, _15491_);
  nor (_22932_, _22931_, _22930_);
  not (_22933_, _22932_);
  nor (_22934_, _13947_, _13475_);
  and (_22935_, _13947_, _13475_);
  nor (_22936_, _22935_, _22934_);
  nor (_22937_, _22936_, _14261_);
  and (_22938_, _22936_, _14261_);
  nor (_22939_, _22938_, _22937_);
  and (_22941_, _22939_, _15190_);
  nor (_22942_, _22939_, _15190_);
  or (_22943_, _22942_, _22941_);
  and (_22944_, _22943_, _07370_);
  nor (_22945_, _22943_, _07370_);
  or (_22946_, _22945_, _22944_);
  nand (_22947_, _22946_, _22933_);
  or (_22948_, _22946_, _22933_);
  and (_22949_, _22948_, _01537_);
  and (_22950_, _22949_, _22947_);
  or (_22952_, _22950_, _22924_);
  and (_22953_, _22952_, _07368_);
  nor (_22954_, _09829_, _01651_);
  nor (_22955_, _07374_, _02057_);
  and (_22956_, _22955_, _22954_);
  not (_22957_, _07375_);
  and (_22958_, _14012_, _22957_);
  and (_22959_, _22958_, _01689_);
  nor (_22960_, _22958_, _01689_);
  nor (_22961_, _22960_, _22959_);
  nor (_22963_, _22961_, _14878_);
  and (_22964_, _22961_, _14878_);
  or (_22965_, _22964_, _22963_);
  and (_22966_, _22965_, _15496_);
  nor (_22967_, _22965_, _15496_);
  nor (_22968_, _22967_, _22966_);
  not (_22969_, _22968_);
  nor (_22970_, _15195_, _07382_);
  and (_22971_, _15195_, _07382_);
  nor (_22972_, _22971_, _22970_);
  nand (_22974_, _22972_, _22969_);
  or (_22975_, _22972_, _22969_);
  and (_22976_, _22975_, _07367_);
  nand (_22977_, _22976_, _22974_);
  nand (_22978_, _22977_, _22956_);
  or (_22979_, _22978_, _22953_);
  or (_22980_, _22956_, _21556_);
  and (_22981_, _22980_, _38087_);
  and (_22982_, _22981_, _22979_);
  or (_22983_, _22982_, _21540_);
  and (_40267_, _22983_, _37580_);
  and (_22985_, _38088_, \oc8051_golden_model_1.PSW [1]);
  and (_22986_, _08232_, \oc8051_golden_model_1.PSW [1]);
  nor (_22987_, _08232_, _02811_);
  or (_22988_, _22987_, _22986_);
  or (_22989_, _22988_, _02840_);
  or (_22990_, _03676_, \oc8051_golden_model_1.PSW [1]);
  and (_22991_, _10698_, _03676_);
  not (_22992_, _22991_);
  and (_22993_, _22992_, _22990_);
  or (_22995_, _22993_, _02814_);
  nand (_22996_, _03676_, _01613_);
  and (_22997_, _22996_, _22990_);
  and (_22998_, _22997_, _02817_);
  and (_22999_, _02818_, \oc8051_golden_model_1.PSW [1]);
  or (_23000_, _22999_, _02001_);
  or (_23001_, _23000_, _22998_);
  and (_23002_, _23001_, _02024_);
  and (_23003_, _23002_, _22995_);
  not (_23004_, _04321_);
  and (_23006_, _23004_, \oc8051_golden_model_1.PSW [1]);
  and (_23007_, _10710_, _04321_);
  or (_23008_, _23007_, _23006_);
  and (_23009_, _23008_, _02007_);
  or (_23010_, _23009_, _01999_);
  or (_23011_, _23010_, _23003_);
  and (_23012_, _23011_, _22989_);
  or (_23013_, _23012_, _02006_);
  or (_23014_, _22997_, _02021_);
  and (_23015_, _23014_, _02025_);
  and (_23017_, _23015_, _23013_);
  and (_23018_, _10696_, _04321_);
  or (_23019_, _23018_, _23006_);
  and (_23020_, _23019_, _01997_);
  or (_23021_, _23020_, _01991_);
  or (_23022_, _23021_, _23017_);
  and (_23023_, _23007_, _10725_);
  or (_23024_, _23006_, _02861_);
  or (_23025_, _23024_, _23023_);
  and (_23026_, _23025_, _23022_);
  and (_23028_, _23026_, _02408_);
  nor (_23029_, _10742_, _23004_);
  or (_23030_, _23006_, _23029_);
  and (_23031_, _23030_, _01875_);
  or (_23032_, _23031_, _05994_);
  or (_23033_, _23032_, _23028_);
  or (_23034_, _22988_, _05249_);
  and (_23035_, _23034_, _23033_);
  or (_23036_, _23035_, _02528_);
  and (_23037_, _04907_, _03676_);
  or (_23039_, _22986_, _02888_);
  or (_23040_, _23039_, _23037_);
  and (_23041_, _23040_, _02043_);
  and (_23042_, _23041_, _23036_);
  nor (_23043_, _10802_, _08232_);
  or (_23044_, _23043_, _22986_);
  and (_23045_, _23044_, _01602_);
  or (_23046_, _23045_, _23042_);
  and (_23047_, _23046_, _01870_);
  nand (_23048_, _03676_, _02687_);
  and (_23050_, _22990_, _01869_);
  and (_23051_, _23050_, _23048_);
  or (_23052_, _23051_, _23047_);
  and (_23053_, _23052_, _02166_);
  or (_23054_, _10816_, _08232_);
  and (_23055_, _22990_, _02079_);
  and (_23056_, _23055_, _23054_);
  or (_23057_, _23056_, _23053_);
  and (_23058_, _23057_, _02912_);
  or (_23059_, _10822_, _08232_);
  and (_23061_, _22990_, _02167_);
  and (_23062_, _23061_, _23059_);
  or (_23063_, _23062_, _23058_);
  and (_23064_, _23063_, _02176_);
  or (_23065_, _10692_, _08232_);
  and (_23066_, _22990_, _02072_);
  and (_23067_, _23066_, _23065_);
  or (_23068_, _23067_, _23064_);
  and (_23069_, _23068_, _02907_);
  or (_23070_, _22986_, _04058_);
  and (_23072_, _22997_, _02177_);
  and (_23073_, _23072_, _23070_);
  or (_23074_, _23073_, _23069_);
  and (_23075_, _23074_, _02174_);
  or (_23076_, _22996_, _04058_);
  and (_23077_, _22990_, _02173_);
  and (_23078_, _23077_, _23076_);
  or (_23079_, _23078_, _02201_);
  or (_23080_, _23048_, _04058_);
  and (_23081_, _22990_, _02071_);
  and (_23083_, _23081_, _23080_);
  or (_23084_, _23083_, _23079_);
  or (_23085_, _23084_, _23075_);
  or (_23086_, _22993_, _02303_);
  and (_23087_, _23086_, _01887_);
  and (_23088_, _23087_, _23085_);
  and (_23089_, _23019_, _01860_);
  or (_23090_, _23089_, _01537_);
  or (_23091_, _23090_, _23088_);
  or (_23092_, _22986_, _01538_);
  or (_23094_, _23092_, _22991_);
  and (_23095_, _23094_, _38087_);
  and (_23096_, _23095_, _23091_);
  or (_23097_, _23096_, _22985_);
  and (_40268_, _23097_, _37580_);
  and (_23098_, _38088_, \oc8051_golden_model_1.PSW [2]);
  nor (_23099_, _06704_, _22343_);
  nor (_23100_, _06705_, \oc8051_golden_model_1.ACC [7]);
  nor (_23101_, _23100_, _08866_);
  nor (_23102_, _23101_, _23099_);
  and (_23104_, _23102_, _07111_);
  and (_23105_, _23099_, _07108_);
  or (_23106_, _23105_, _07084_);
  or (_23107_, _23106_, _23104_);
  and (_23108_, _08232_, \oc8051_golden_model_1.PSW [2]);
  and (_23109_, _11020_, _03676_);
  or (_23110_, _23109_, _23108_);
  and (_23111_, _23110_, _02167_);
  nor (_23112_, _08232_, _03455_);
  or (_23113_, _23112_, _23108_);
  or (_23115_, _23113_, _05249_);
  nor (_23116_, _06542_, _22373_);
  nor (_23117_, _06544_, \oc8051_golden_model_1.ACC [7]);
  or (_23118_, _23117_, _23116_);
  and (_23119_, _23118_, _08243_);
  nor (_23120_, _23118_, _08243_);
  nor (_23121_, _23120_, _23119_);
  nor (_23122_, _23121_, _21950_);
  and (_23123_, _23121_, _21950_);
  or (_23124_, _23123_, _08245_);
  or (_23126_, _23124_, _23122_);
  and (_23127_, _08785_, _06706_);
  nor (_23128_, _08785_, _06706_);
  or (_23129_, _23128_, _23127_);
  or (_23130_, _23129_, _06766_);
  nand (_23131_, _23129_, _06766_);
  and (_23132_, _23131_, _23130_);
  and (_23133_, _23132_, _06699_);
  and (_23134_, _23004_, \oc8051_golden_model_1.PSW [2]);
  and (_23135_, _10894_, _04321_);
  or (_23137_, _23135_, _23134_);
  and (_23138_, _23137_, _01997_);
  or (_23139_, _23113_, _02840_);
  nor (_23140_, _10905_, _08232_);
  or (_23141_, _23140_, _23108_);
  or (_23142_, _23141_, _02814_);
  and (_23143_, _03676_, \oc8051_golden_model_1.ACC [2]);
  or (_23144_, _23143_, _23108_);
  and (_23145_, _23144_, _02817_);
  and (_23146_, _02818_, \oc8051_golden_model_1.PSW [2]);
  or (_23148_, _23146_, _02001_);
  or (_23149_, _23148_, _23145_);
  and (_23150_, _23149_, _02024_);
  and (_23151_, _23150_, _23142_);
  and (_23152_, _10909_, _04321_);
  or (_23153_, _23152_, _23134_);
  and (_23154_, _23153_, _02007_);
  or (_23155_, _23154_, _01999_);
  or (_23156_, _23155_, _23151_);
  and (_23157_, _23156_, _23139_);
  or (_23159_, _23157_, _02006_);
  or (_23160_, _23144_, _02021_);
  and (_23161_, _23160_, _02025_);
  and (_23162_, _23161_, _23159_);
  or (_23163_, _23162_, _23138_);
  and (_23164_, _23163_, _02861_);
  and (_23165_, _23152_, _10924_);
  or (_23166_, _23165_, _23134_);
  and (_23167_, _23166_, _01991_);
  or (_23168_, _23167_, _05279_);
  or (_23170_, _23168_, _23164_);
  or (_23171_, _12772_, _12667_);
  or (_23172_, _23171_, _12892_);
  or (_23173_, _23172_, _13011_);
  or (_23174_, _23173_, _13129_);
  or (_23175_, _23174_, _13249_);
  or (_23176_, _23175_, _13366_);
  or (_23177_, _23176_, _05988_);
  and (_23178_, _23177_, _06700_);
  and (_23179_, _23178_, _23170_);
  or (_23181_, _23179_, _06609_);
  or (_23182_, _23181_, _23133_);
  and (_23183_, _23182_, _02036_);
  and (_23184_, _23183_, _23126_);
  nor (_23185_, _06888_, \oc8051_golden_model_1.ACC [7]);
  nor (_23186_, _06887_, _08914_);
  or (_23187_, _23186_, _23185_);
  nor (_23188_, _23187_, _08799_);
  and (_23189_, _23187_, _08799_);
  nor (_23190_, _23189_, _23188_);
  and (_23192_, _23190_, _21978_);
  nor (_23193_, _23190_, _21978_);
  or (_23194_, _23193_, _23192_);
  or (_23195_, _23194_, _06476_);
  and (_23196_, _23195_, _06776_);
  or (_23197_, _23196_, _23184_);
  nor (_23198_, _06480_, _08224_);
  nor (_23199_, _06481_, \oc8051_golden_model_1.ACC [7]);
  nor (_23200_, _23199_, _23198_);
  not (_23201_, _23200_);
  nor (_23203_, _23201_, _08811_);
  and (_23204_, _23201_, _08811_);
  or (_23205_, _23204_, _23203_);
  nor (_23206_, _23205_, _06540_);
  and (_23207_, _23205_, _06540_);
  or (_23208_, _23207_, _23206_);
  or (_23209_, _23208_, _06777_);
  and (_23210_, _23209_, _02408_);
  and (_23211_, _23210_, _23197_);
  nor (_23212_, _10942_, _23004_);
  or (_23213_, _23212_, _23134_);
  and (_23214_, _23213_, _01875_);
  or (_23215_, _23214_, _05994_);
  or (_23216_, _23215_, _23211_);
  and (_23217_, _23216_, _23115_);
  or (_23218_, _23217_, _02528_);
  and (_23219_, _05043_, _03676_);
  or (_23220_, _23108_, _02888_);
  or (_23221_, _23220_, _23219_);
  and (_23222_, _23221_, _02043_);
  and (_23224_, _23222_, _23218_);
  nor (_23225_, _11000_, _08232_);
  or (_23226_, _23225_, _23108_);
  and (_23227_, _23226_, _01602_);
  or (_23228_, _23227_, _06008_);
  or (_23229_, _23228_, _23224_);
  nand (_23230_, _06024_, _06020_);
  nand (_23231_, _23230_, _06008_);
  and (_23232_, _23231_, _23229_);
  and (_23233_, _23232_, _01870_);
  and (_23235_, _03676_, _04724_);
  or (_23236_, _23235_, _23108_);
  and (_23237_, _23236_, _01869_);
  or (_23238_, _23237_, _02079_);
  or (_23239_, _23238_, _23233_);
  and (_23240_, _11014_, _03676_);
  or (_23241_, _23108_, _02166_);
  or (_23242_, _23241_, _23240_);
  and (_23243_, _23242_, _02912_);
  and (_23244_, _23243_, _23239_);
  or (_23246_, _23244_, _23111_);
  and (_23247_, _23246_, _02176_);
  or (_23248_, _23108_, _04156_);
  and (_23249_, _23236_, _02072_);
  and (_23250_, _23249_, _23248_);
  or (_23251_, _23250_, _23247_);
  and (_23252_, _23251_, _02907_);
  and (_23253_, _23144_, _02177_);
  and (_23254_, _23253_, _23248_);
  or (_23255_, _23254_, _02071_);
  or (_23257_, _23255_, _23252_);
  nor (_23258_, _11013_, _08232_);
  or (_23259_, _23108_, _04788_);
  or (_23260_, _23259_, _23258_);
  and (_23261_, _23260_, _04793_);
  and (_23262_, _23261_, _23257_);
  nor (_23263_, _11019_, _08232_);
  or (_23264_, _23263_, _23108_);
  and (_23265_, _23264_, _02173_);
  or (_23266_, _23265_, _07085_);
  or (_23268_, _23266_, _23262_);
  and (_23269_, _23268_, _23107_);
  or (_23270_, _23269_, _07114_);
  nor (_23271_, _23118_, _08873_);
  nor (_23272_, _23271_, _23116_);
  and (_23273_, _23272_, _07140_);
  and (_23274_, _23116_, _07137_);
  or (_23275_, _23274_, _07116_);
  or (_23276_, _23275_, _23273_);
  and (_23277_, _23276_, _02165_);
  and (_23279_, _23277_, _23270_);
  and (_23280_, _23186_, _07168_);
  nor (_23281_, _23187_, _08879_);
  nor (_23282_, _23281_, _23186_);
  and (_23283_, _23282_, _07171_);
  or (_23284_, _23283_, _23280_);
  and (_23285_, _23284_, _02164_);
  or (_23286_, _23285_, _07144_);
  or (_23287_, _23286_, _23279_);
  nor (_23288_, _23201_, _08886_);
  or (_23290_, _23288_, _23198_);
  nand (_23291_, _23290_, _07202_);
  or (_23292_, _23290_, _07202_);
  and (_23293_, _23292_, _23291_);
  or (_23294_, _23293_, _07177_);
  nand (_23295_, _23294_, _23287_);
  nand (_23296_, _23295_, _06457_);
  or (_23297_, _08897_, _06445_);
  or (_23298_, _06446_, _06406_);
  and (_23299_, _23298_, _23297_);
  or (_23301_, _23299_, _06457_);
  and (_23302_, _23301_, _23296_);
  or (_23303_, _23302_, _06450_);
  or (_23304_, _23299_, _06451_);
  and (_23305_, _23304_, _07212_);
  and (_23306_, _23305_, _23303_);
  or (_23307_, _07246_, _06461_);
  or (_23308_, _08906_, _07245_);
  and (_23309_, _23308_, _07210_);
  and (_23310_, _23309_, _23307_);
  or (_23311_, _23310_, _23306_);
  and (_23312_, _23311_, _07254_);
  or (_23313_, _07297_, _07257_);
  and (_23314_, _23313_, _08916_);
  nand (_23315_, _07335_, _08224_);
  and (_23316_, _23315_, _08226_);
  or (_23317_, _23316_, _02201_);
  or (_23318_, _23317_, _23314_);
  or (_23319_, _23318_, _23312_);
  or (_23320_, _23141_, _02303_);
  and (_23322_, _23320_, _01887_);
  and (_23323_, _23322_, _23319_);
  and (_23324_, _23137_, _01860_);
  or (_23325_, _23324_, _01537_);
  or (_23326_, _23325_, _23323_);
  and (_23327_, _11072_, _03676_);
  or (_23328_, _23108_, _01538_);
  or (_23329_, _23328_, _23327_);
  and (_23330_, _23329_, _38087_);
  and (_23331_, _23330_, _23326_);
  or (_23333_, _23331_, _23098_);
  and (_40269_, _23333_, _37580_);
  not (_23334_, \oc8051_golden_model_1.PSW [3]);
  nor (_23335_, _38087_, _23334_);
  nor (_23336_, _03676_, _23334_);
  and (_23337_, _11094_, _03676_);
  or (_23338_, _23337_, _23336_);
  and (_23339_, _23338_, _02167_);
  nor (_23340_, _08232_, _03268_);
  or (_23341_, _23340_, _23336_);
  or (_23343_, _23341_, _05249_);
  nor (_23344_, _11101_, _08232_);
  or (_23345_, _23344_, _23336_);
  or (_23346_, _23345_, _02814_);
  and (_23347_, _03676_, \oc8051_golden_model_1.ACC [3]);
  or (_23348_, _23347_, _23336_);
  and (_23349_, _23348_, _02817_);
  nor (_23350_, _02817_, _23334_);
  or (_23351_, _23350_, _02001_);
  or (_23352_, _23351_, _23349_);
  and (_23354_, _23352_, _02024_);
  and (_23355_, _23354_, _23346_);
  nor (_23356_, _04321_, _23334_);
  and (_23357_, _11098_, _04321_);
  or (_23358_, _23357_, _23356_);
  and (_23359_, _23358_, _02007_);
  or (_23360_, _23359_, _01999_);
  or (_23361_, _23360_, _23355_);
  or (_23362_, _23341_, _02840_);
  and (_23363_, _23362_, _23361_);
  or (_23365_, _23363_, _02006_);
  or (_23366_, _23348_, _02021_);
  and (_23367_, _23366_, _02025_);
  and (_23368_, _23367_, _23365_);
  and (_23369_, _11096_, _04321_);
  or (_23370_, _23369_, _23356_);
  and (_23371_, _23370_, _01997_);
  or (_23372_, _23371_, _01991_);
  or (_23373_, _23372_, _23368_);
  or (_23374_, _23356_, _11127_);
  and (_23376_, _23374_, _23358_);
  or (_23377_, _23376_, _02861_);
  and (_23378_, _23377_, _02408_);
  and (_23379_, _23378_, _23373_);
  nor (_23380_, _11145_, _23004_);
  or (_23381_, _23380_, _23356_);
  and (_23382_, _23381_, _01875_);
  or (_23383_, _23382_, _05994_);
  or (_23384_, _23383_, _23379_);
  and (_23385_, _23384_, _23343_);
  or (_23386_, _23385_, _02528_);
  and (_23387_, _04998_, _03676_);
  or (_23388_, _23336_, _02888_);
  or (_23389_, _23388_, _23387_);
  and (_23390_, _23389_, _02043_);
  and (_23391_, _23390_, _23386_);
  nor (_23392_, _11206_, _08232_);
  or (_23393_, _23392_, _23336_);
  and (_23394_, _23393_, _01602_);
  or (_23395_, _23394_, _01869_);
  or (_23397_, _23395_, _23391_);
  and (_23398_, _03676_, _04678_);
  or (_23399_, _23398_, _23336_);
  or (_23400_, _23399_, _01870_);
  and (_23401_, _23400_, _23397_);
  or (_23402_, _23401_, _02079_);
  and (_23403_, _11222_, _03676_);
  or (_23404_, _23336_, _02166_);
  or (_23405_, _23404_, _23403_);
  and (_23406_, _23405_, _02912_);
  and (_23408_, _23406_, _23402_);
  or (_23409_, _23408_, _23339_);
  and (_23410_, _23409_, _02176_);
  or (_23411_, _23336_, _04014_);
  and (_23412_, _23399_, _02072_);
  and (_23413_, _23412_, _23411_);
  or (_23414_, _23413_, _23410_);
  and (_23415_, _23414_, _02907_);
  and (_23416_, _23348_, _02177_);
  and (_23417_, _23416_, _23411_);
  or (_23419_, _23417_, _02071_);
  or (_23420_, _23419_, _23415_);
  nor (_23421_, _11220_, _08232_);
  or (_23422_, _23336_, _04788_);
  or (_23423_, _23422_, _23421_);
  and (_23424_, _23423_, _04793_);
  and (_23425_, _23424_, _23420_);
  nor (_23426_, _11093_, _08232_);
  or (_23427_, _23426_, _23336_);
  and (_23428_, _23427_, _02173_);
  or (_23430_, _23428_, _02201_);
  or (_23431_, _23430_, _23425_);
  or (_23432_, _23345_, _02303_);
  and (_23433_, _23432_, _01887_);
  and (_23434_, _23433_, _23431_);
  and (_23435_, _23370_, _01860_);
  or (_23436_, _23435_, _01537_);
  or (_23437_, _23436_, _23434_);
  and (_23438_, _11273_, _03676_);
  or (_23439_, _23336_, _01538_);
  or (_23441_, _23439_, _23438_);
  and (_23442_, _23441_, _38087_);
  and (_23443_, _23442_, _23437_);
  or (_23444_, _23443_, _23335_);
  and (_40270_, _23444_, _37580_);
  and (_23445_, _38088_, \oc8051_golden_model_1.PSW [4]);
  and (_23446_, _08232_, \oc8051_golden_model_1.PSW [4]);
  and (_23447_, _11431_, _03676_);
  or (_23448_, _23447_, _23446_);
  and (_23449_, _23448_, _02167_);
  nor (_23451_, _04211_, _08232_);
  or (_23452_, _23451_, _23446_);
  or (_23453_, _23452_, _05249_);
  and (_23454_, _23004_, \oc8051_golden_model_1.PSW [4]);
  and (_23455_, _11301_, _04321_);
  or (_23456_, _23455_, _23454_);
  and (_23457_, _23456_, _01997_);
  nor (_23458_, _11317_, _08232_);
  or (_23459_, _23458_, _23446_);
  or (_23460_, _23459_, _02814_);
  and (_23461_, _03676_, \oc8051_golden_model_1.ACC [4]);
  or (_23462_, _23461_, _23446_);
  and (_23463_, _23462_, _02817_);
  and (_23464_, _02818_, \oc8051_golden_model_1.PSW [4]);
  or (_23465_, _23464_, _02001_);
  or (_23466_, _23465_, _23463_);
  and (_23467_, _23466_, _02024_);
  and (_23468_, _23467_, _23460_);
  and (_23469_, _11303_, _04321_);
  or (_23470_, _23469_, _23454_);
  and (_23472_, _23470_, _02007_);
  or (_23473_, _23472_, _01999_);
  or (_23474_, _23473_, _23468_);
  or (_23475_, _23452_, _02840_);
  and (_23476_, _23475_, _23474_);
  or (_23477_, _23476_, _02006_);
  or (_23478_, _23462_, _02021_);
  and (_23479_, _23478_, _02025_);
  and (_23480_, _23479_, _23477_);
  or (_23481_, _23480_, _23457_);
  and (_23483_, _23481_, _02861_);
  and (_23484_, _11335_, _04321_);
  or (_23485_, _23484_, _23454_);
  and (_23486_, _23485_, _01991_);
  or (_23487_, _23486_, _23483_);
  and (_23488_, _23487_, _02408_);
  nor (_23489_, _11299_, _23004_);
  or (_23490_, _23489_, _23454_);
  and (_23491_, _23490_, _01875_);
  or (_23492_, _23491_, _05994_);
  or (_23494_, _23492_, _23488_);
  and (_23495_, _23494_, _23453_);
  or (_23496_, _23495_, _02528_);
  and (_23497_, _05135_, _03676_);
  or (_23498_, _23446_, _02888_);
  or (_23499_, _23498_, _23497_);
  and (_23500_, _23499_, _02043_);
  and (_23501_, _23500_, _23496_);
  nor (_23502_, _11411_, _08232_);
  or (_23503_, _23502_, _23446_);
  and (_23505_, _23503_, _01602_);
  or (_23506_, _23505_, _01869_);
  or (_23507_, _23506_, _23501_);
  and (_23508_, _04694_, _03676_);
  or (_23509_, _23508_, _23446_);
  or (_23510_, _23509_, _01870_);
  and (_23511_, _23510_, _23507_);
  or (_23512_, _23511_, _02079_);
  and (_23513_, _11425_, _03676_);
  or (_23514_, _23446_, _02166_);
  or (_23516_, _23514_, _23513_);
  and (_23517_, _23516_, _02912_);
  and (_23518_, _23517_, _23512_);
  or (_23519_, _23518_, _23449_);
  and (_23520_, _23519_, _02176_);
  or (_23521_, _23446_, _04258_);
  and (_23522_, _23509_, _02072_);
  and (_23523_, _23522_, _23521_);
  or (_23524_, _23523_, _23520_);
  and (_23525_, _23524_, _02907_);
  and (_23527_, _23462_, _02177_);
  and (_23528_, _23527_, _23521_);
  or (_23529_, _23528_, _02071_);
  or (_23530_, _23529_, _23525_);
  nor (_23531_, _11424_, _08232_);
  or (_23532_, _23446_, _04788_);
  or (_23533_, _23532_, _23531_);
  and (_23534_, _23533_, _04793_);
  and (_23535_, _23534_, _23530_);
  nor (_23536_, _11430_, _08232_);
  or (_23537_, _23536_, _23446_);
  and (_23538_, _23537_, _02173_);
  or (_23539_, _23538_, _02201_);
  or (_23540_, _23539_, _23535_);
  or (_23541_, _23459_, _02303_);
  and (_23542_, _23541_, _01887_);
  and (_23543_, _23542_, _23540_);
  and (_23544_, _23456_, _01860_);
  or (_23545_, _23544_, _01537_);
  or (_23546_, _23545_, _23543_);
  and (_23548_, _11487_, _03676_);
  or (_23549_, _23446_, _01538_);
  or (_23550_, _23549_, _23548_);
  and (_23551_, _23550_, _38087_);
  and (_23552_, _23551_, _23546_);
  or (_23553_, _23552_, _23445_);
  and (_40271_, _23553_, _37580_);
  and (_23554_, _38088_, \oc8051_golden_model_1.PSW [5]);
  and (_23555_, _08232_, \oc8051_golden_model_1.PSW [5]);
  and (_23556_, _11635_, _03676_);
  or (_23558_, _23556_, _23555_);
  and (_23559_, _23558_, _02167_);
  nor (_23560_, _11525_, _08232_);
  or (_23561_, _23560_, _23555_);
  or (_23562_, _23561_, _02814_);
  and (_23563_, _03676_, \oc8051_golden_model_1.ACC [5]);
  or (_23564_, _23563_, _23555_);
  and (_23565_, _23564_, _02817_);
  and (_23566_, _02818_, \oc8051_golden_model_1.PSW [5]);
  or (_23567_, _23566_, _02001_);
  or (_23569_, _23567_, _23565_);
  and (_23570_, _23569_, _02024_);
  and (_23571_, _23570_, _23562_);
  and (_23572_, _23004_, \oc8051_golden_model_1.PSW [5]);
  and (_23573_, _11510_, _04321_);
  or (_23574_, _23573_, _23572_);
  and (_23575_, _23574_, _02007_);
  or (_23576_, _23575_, _01999_);
  or (_23577_, _23576_, _23571_);
  nor (_23578_, _03916_, _08232_);
  or (_23580_, _23578_, _23555_);
  or (_23581_, _23580_, _02840_);
  and (_23582_, _23581_, _23577_);
  or (_23583_, _23582_, _02006_);
  or (_23584_, _23564_, _02021_);
  and (_23585_, _23584_, _02025_);
  and (_23586_, _23585_, _23583_);
  and (_23587_, _11508_, _04321_);
  or (_23588_, _23587_, _23572_);
  and (_23589_, _23588_, _01997_);
  or (_23591_, _23589_, _01991_);
  or (_23592_, _23591_, _23586_);
  or (_23593_, _23572_, _11542_);
  and (_23594_, _23593_, _23574_);
  or (_23595_, _23594_, _02861_);
  and (_23596_, _23595_, _02408_);
  and (_23597_, _23596_, _23592_);
  nor (_23598_, _11506_, _23004_);
  or (_23599_, _23598_, _23572_);
  and (_23600_, _23599_, _01875_);
  or (_23602_, _23600_, _05994_);
  or (_23603_, _23602_, _23597_);
  or (_23604_, _23580_, _05249_);
  and (_23605_, _23604_, _23603_);
  or (_23606_, _23605_, _02528_);
  and (_23607_, _05090_, _03676_);
  or (_23608_, _23555_, _02888_);
  or (_23609_, _23608_, _23607_);
  and (_23610_, _23609_, _02043_);
  and (_23611_, _23610_, _23606_);
  nor (_23612_, _11615_, _08232_);
  or (_23613_, _23612_, _23555_);
  and (_23614_, _23613_, _01602_);
  or (_23615_, _23614_, _01869_);
  or (_23616_, _23615_, _23611_);
  and (_23617_, _04672_, _03676_);
  or (_23618_, _23617_, _23555_);
  or (_23619_, _23618_, _01870_);
  and (_23620_, _23619_, _23616_);
  or (_23621_, _23620_, _02079_);
  and (_23623_, _11629_, _03676_);
  or (_23624_, _23555_, _02166_);
  or (_23625_, _23624_, _23623_);
  and (_23626_, _23625_, _02912_);
  and (_23627_, _23626_, _23621_);
  or (_23628_, _23627_, _23559_);
  and (_23629_, _23628_, _02176_);
  or (_23630_, _23555_, _03965_);
  and (_23631_, _23618_, _02072_);
  and (_23632_, _23631_, _23630_);
  or (_23634_, _23632_, _23629_);
  and (_23635_, _23634_, _02907_);
  and (_23636_, _23564_, _02177_);
  and (_23637_, _23636_, _23630_);
  or (_23638_, _23637_, _02071_);
  or (_23639_, _23638_, _23635_);
  nor (_23640_, _11628_, _08232_);
  or (_23641_, _23555_, _04788_);
  or (_23642_, _23641_, _23640_);
  and (_23643_, _23642_, _04793_);
  and (_23645_, _23643_, _23639_);
  nor (_23646_, _11634_, _08232_);
  or (_23647_, _23646_, _23555_);
  and (_23648_, _23647_, _02173_);
  or (_23649_, _23648_, _02201_);
  or (_23650_, _23649_, _23645_);
  or (_23651_, _23561_, _02303_);
  and (_23652_, _23651_, _01887_);
  and (_23653_, _23652_, _23650_);
  and (_23654_, _23588_, _01860_);
  or (_23656_, _23654_, _01537_);
  or (_23657_, _23656_, _23653_);
  and (_23658_, _11685_, _03676_);
  or (_23659_, _23555_, _01538_);
  or (_23660_, _23659_, _23658_);
  and (_23661_, _23660_, _38087_);
  and (_23662_, _23661_, _23657_);
  or (_23663_, _23662_, _23554_);
  and (_40272_, _23663_, _37580_);
  nor (_23664_, _38087_, _14331_);
  or (_23666_, _07329_, _07256_);
  or (_23667_, _07161_, _06854_);
  and (_23668_, _23667_, _02164_);
  or (_23669_, _07102_, _06721_);
  and (_23670_, _23669_, _07083_);
  or (_23671_, _23670_, _07084_);
  nor (_23672_, _03676_, _14331_);
  and (_23673_, _11709_, _03676_);
  or (_23674_, _23673_, _23672_);
  and (_23675_, _23674_, _02167_);
  nor (_23677_, _03808_, _08232_);
  or (_23678_, _23677_, _23672_);
  or (_23679_, _23678_, _05249_);
  or (_23680_, _06533_, _06478_);
  and (_23681_, _23680_, _06476_);
  or (_23682_, _06721_, _06700_);
  or (_23683_, _23682_, _06759_);
  nor (_23684_, _04321_, _14331_);
  and (_23685_, _11715_, _04321_);
  or (_23686_, _23685_, _23684_);
  and (_23687_, _23686_, _01997_);
  nor (_23688_, _11730_, _08232_);
  or (_23689_, _23688_, _23672_);
  or (_23690_, _23689_, _02814_);
  and (_23691_, _03676_, \oc8051_golden_model_1.ACC [6]);
  or (_23692_, _23691_, _23672_);
  and (_23693_, _23692_, _02817_);
  nor (_23694_, _02817_, _14331_);
  or (_23695_, _23694_, _02001_);
  or (_23696_, _23695_, _23693_);
  and (_23698_, _23696_, _02024_);
  and (_23699_, _23698_, _23690_);
  and (_23700_, _11717_, _04321_);
  or (_23701_, _23700_, _23684_);
  and (_23702_, _23701_, _02007_);
  or (_23703_, _23702_, _01999_);
  or (_23704_, _23703_, _23699_);
  or (_23705_, _23678_, _02840_);
  and (_23706_, _23705_, _23704_);
  or (_23707_, _23706_, _02006_);
  or (_23709_, _23692_, _02021_);
  and (_23710_, _23709_, _02025_);
  and (_23711_, _23710_, _23707_);
  or (_23712_, _23711_, _23687_);
  and (_23713_, _23712_, _02861_);
  or (_23714_, _23684_, _11747_);
  and (_23715_, _23714_, _01991_);
  and (_23716_, _23715_, _23701_);
  or (_23717_, _23716_, _06699_);
  or (_23718_, _23717_, _23713_);
  and (_23720_, _23718_, _23683_);
  or (_23721_, _23720_, _06609_);
  or (_23722_, _08245_, _06561_);
  or (_23723_, _23722_, _06598_);
  and (_23724_, _23723_, _23721_);
  or (_23725_, _23724_, _01963_);
  or (_23726_, _06854_, _02036_);
  or (_23727_, _23726_, _06936_);
  and (_23728_, _23727_, _06777_);
  and (_23729_, _23728_, _23725_);
  or (_23731_, _23729_, _23681_);
  and (_23732_, _23731_, _02408_);
  nor (_23733_, _11713_, _23004_);
  or (_23734_, _23733_, _23684_);
  and (_23735_, _23734_, _01875_);
  or (_23736_, _23735_, _05994_);
  or (_23737_, _23736_, _23732_);
  and (_23738_, _23737_, _23679_);
  or (_23739_, _23738_, _02528_);
  and (_23740_, _04861_, _03676_);
  or (_23742_, _23672_, _02888_);
  or (_23743_, _23742_, _23740_);
  and (_23744_, _23743_, _02043_);
  and (_23745_, _23744_, _23739_);
  nor (_23746_, _11820_, _08232_);
  or (_23747_, _23746_, _23672_);
  and (_23748_, _23747_, _01602_);
  or (_23749_, _23748_, _01869_);
  or (_23750_, _23749_, _23745_);
  and (_23751_, _09920_, _03676_);
  or (_23753_, _23751_, _23672_);
  or (_23754_, _23753_, _01870_);
  and (_23755_, _23754_, _23750_);
  or (_23756_, _23755_, _02079_);
  and (_23757_, _11835_, _03676_);
  or (_23758_, _23672_, _02166_);
  or (_23759_, _23758_, _23757_);
  and (_23760_, _23759_, _02912_);
  and (_23761_, _23760_, _23756_);
  or (_23762_, _23761_, _23675_);
  and (_23763_, _23762_, _02176_);
  or (_23764_, _23672_, _03863_);
  and (_23765_, _23753_, _02072_);
  and (_23766_, _23765_, _23764_);
  or (_23767_, _23766_, _23763_);
  and (_23768_, _23767_, _02907_);
  and (_23769_, _23692_, _02177_);
  and (_23770_, _23769_, _23764_);
  or (_23771_, _23770_, _02071_);
  or (_23772_, _23771_, _23768_);
  nor (_23774_, _11833_, _08232_);
  or (_23775_, _23672_, _04788_);
  or (_23776_, _23775_, _23774_);
  and (_23777_, _23776_, _04793_);
  and (_23778_, _23777_, _23772_);
  nor (_23779_, _11708_, _08232_);
  or (_23780_, _23779_, _23672_);
  nand (_23781_, _23780_, _02173_);
  nand (_23782_, _23781_, _07081_);
  or (_23783_, _23782_, _23778_);
  and (_23785_, _23783_, _23671_);
  and (_23786_, _23669_, _07082_);
  or (_23787_, _23786_, _07114_);
  or (_23788_, _23787_, _23785_);
  or (_23789_, _07116_, _06561_);
  or (_23790_, _23789_, _07131_);
  and (_23791_, _23790_, _02165_);
  and (_23792_, _23791_, _23788_);
  or (_23793_, _23792_, _23668_);
  and (_23794_, _23793_, _07177_);
  or (_23796_, _07193_, _06478_);
  and (_23797_, _23796_, _07144_);
  or (_23798_, _23797_, _06459_);
  or (_23799_, _23798_, _23794_);
  or (_23800_, _06458_, _06439_);
  and (_23801_, _23800_, _23799_);
  or (_23802_, _23801_, _07210_);
  or (_23803_, _07240_, _07212_);
  and (_23804_, _23803_, _01891_);
  and (_23805_, _23804_, _23802_);
  or (_23807_, _07291_, _07253_);
  and (_23808_, _23807_, _07255_);
  or (_23809_, _23808_, _23805_);
  and (_23810_, _23809_, _23666_);
  or (_23811_, _23810_, _02201_);
  or (_23812_, _23689_, _02303_);
  and (_23813_, _23812_, _01887_);
  and (_23814_, _23813_, _23811_);
  and (_23815_, _23686_, _01860_);
  or (_23816_, _23815_, _01537_);
  or (_23818_, _23816_, _23814_);
  and (_23819_, _11887_, _03676_);
  or (_23820_, _23672_, _01538_);
  or (_23821_, _23820_, _23819_);
  and (_23822_, _23821_, _38087_);
  and (_23823_, _23822_, _23818_);
  or (_23824_, _23823_, _23664_);
  and (_40273_, _23824_, _37580_);
  not (_23825_, \oc8051_golden_model_1.PCON [0]);
  nor (_23826_, _38087_, _23825_);
  nor (_23828_, _04106_, _08941_);
  nor (_23829_, _03662_, _23825_);
  and (_23830_, _03662_, _04562_);
  or (_23831_, _23830_, _23829_);
  nand (_23832_, _23831_, _02072_);
  nor (_23833_, _23832_, _23828_);
  and (_23834_, _03662_, \oc8051_golden_model_1.ACC [0]);
  or (_23835_, _23834_, _23829_);
  and (_23836_, _23835_, _02006_);
  or (_23837_, _23836_, _05994_);
  or (_23839_, _23829_, _23828_);
  and (_23840_, _23839_, _02001_);
  nor (_23841_, _02817_, _23825_);
  and (_23842_, _23835_, _02817_);
  or (_23843_, _23842_, _23841_);
  and (_23844_, _23843_, _02814_);
  or (_23845_, _23844_, _01999_);
  or (_23846_, _23845_, _23840_);
  and (_23847_, _23846_, _02021_);
  or (_23848_, _23847_, _23837_);
  and (_23850_, _03662_, _03028_);
  and (_23851_, _05249_, _02840_);
  or (_23852_, _23851_, _23829_);
  or (_23853_, _23852_, _23850_);
  and (_23854_, _23853_, _23848_);
  or (_23855_, _23854_, _02528_);
  and (_23856_, _04952_, _03662_);
  or (_23857_, _23829_, _02888_);
  or (_23858_, _23857_, _23856_);
  and (_23859_, _23858_, _23855_);
  or (_23861_, _23859_, _01602_);
  nor (_23862_, _10600_, _08941_);
  or (_23863_, _23862_, _23829_);
  or (_23864_, _23863_, _02043_);
  and (_23865_, _23864_, _01870_);
  and (_23866_, _23865_, _23861_);
  and (_23867_, _23831_, _01869_);
  or (_23868_, _23867_, _02079_);
  or (_23869_, _23868_, _23866_);
  and (_23870_, _10614_, _03662_);
  or (_23872_, _23870_, _23829_);
  or (_23873_, _23872_, _02166_);
  and (_23874_, _23873_, _23869_);
  or (_23875_, _23874_, _02167_);
  and (_23876_, _10620_, _03662_);
  or (_23877_, _23829_, _02912_);
  or (_23878_, _23877_, _23876_);
  and (_23879_, _23878_, _02176_);
  and (_23880_, _23879_, _23875_);
  or (_23881_, _23880_, _23833_);
  and (_23883_, _23881_, _02907_);
  or (_23884_, _23829_, _04106_);
  and (_23885_, _23835_, _02177_);
  and (_23886_, _23885_, _23884_);
  or (_23887_, _23886_, _02071_);
  or (_23888_, _23887_, _23883_);
  nor (_23889_, _10613_, _08941_);
  or (_23890_, _23829_, _04788_);
  or (_23891_, _23890_, _23889_);
  and (_23892_, _23891_, _04793_);
  and (_23894_, _23892_, _23888_);
  nor (_23895_, _10619_, _08941_);
  or (_23896_, _23895_, _23829_);
  and (_23897_, _23896_, _02173_);
  or (_23898_, _23897_, _15577_);
  or (_23899_, _23898_, _23894_);
  or (_23900_, _23839_, _02743_);
  and (_23901_, _23900_, _38087_);
  and (_23902_, _23901_, _23899_);
  or (_23903_, _23902_, _23826_);
  and (_40274_, _23903_, _37580_);
  not (_23904_, \oc8051_golden_model_1.PCON [1]);
  nor (_23905_, _38087_, _23904_);
  or (_23906_, _03662_, \oc8051_golden_model_1.PCON [1]);
  and (_23907_, _10698_, _03662_);
  not (_23908_, _23907_);
  and (_23909_, _23908_, _23906_);
  or (_23910_, _23909_, _02814_);
  nand (_23911_, _03662_, _01613_);
  and (_23912_, _23911_, _23906_);
  and (_23914_, _23912_, _02817_);
  nor (_23915_, _02817_, _23904_);
  or (_23916_, _23915_, _02001_);
  or (_23917_, _23916_, _23914_);
  and (_23918_, _23917_, _02840_);
  and (_23919_, _23918_, _23910_);
  nand (_23920_, _03662_, _02811_);
  and (_23921_, _23920_, _23906_);
  and (_23922_, _23921_, _01999_);
  or (_23923_, _23922_, _23919_);
  and (_23925_, _23923_, _02021_);
  and (_23926_, _23912_, _02006_);
  or (_23927_, _23926_, _05994_);
  or (_23928_, _23927_, _23925_);
  or (_23929_, _23921_, _05249_);
  and (_23930_, _23929_, _02888_);
  and (_23931_, _23930_, _23928_);
  or (_23932_, _04907_, _08941_);
  and (_23933_, _23906_, _02528_);
  and (_23934_, _23933_, _23932_);
  or (_23936_, _23934_, _23931_);
  and (_23937_, _23936_, _02043_);
  nand (_23938_, _10802_, _03662_);
  and (_23939_, _23906_, _01602_);
  and (_23940_, _23939_, _23938_);
  or (_23941_, _23940_, _23937_);
  and (_23942_, _23941_, _01870_);
  nand (_23943_, _03662_, _02687_);
  and (_23944_, _23906_, _01869_);
  and (_23945_, _23944_, _23943_);
  or (_23947_, _23945_, _23942_);
  and (_23948_, _23947_, _02166_);
  or (_23949_, _10816_, _08941_);
  and (_23950_, _23906_, _02079_);
  and (_23951_, _23950_, _23949_);
  or (_23952_, _23951_, _23948_);
  and (_23953_, _23952_, _02912_);
  or (_23954_, _10822_, _08941_);
  and (_23955_, _23906_, _02167_);
  and (_23956_, _23955_, _23954_);
  or (_23958_, _23956_, _23953_);
  and (_23959_, _23958_, _02176_);
  or (_23960_, _10692_, _08941_);
  and (_23961_, _23906_, _02072_);
  and (_23962_, _23961_, _23960_);
  or (_23963_, _23962_, _23959_);
  and (_23964_, _23963_, _02907_);
  nor (_23965_, _03662_, _23904_);
  or (_23966_, _23965_, _04058_);
  and (_23967_, _23912_, _02177_);
  and (_23969_, _23967_, _23966_);
  or (_23970_, _23969_, _23964_);
  and (_23971_, _23970_, _02174_);
  or (_23972_, _23911_, _04058_);
  and (_23973_, _23906_, _02173_);
  and (_23974_, _23973_, _23972_);
  or (_23975_, _23974_, _02201_);
  or (_23976_, _23943_, _04058_);
  and (_23977_, _23906_, _02071_);
  and (_23978_, _23977_, _23976_);
  or (_23979_, _23978_, _23975_);
  or (_23980_, _23979_, _23971_);
  or (_23981_, _23909_, _02303_);
  and (_23982_, _23981_, _23980_);
  or (_23983_, _23982_, _01537_);
  or (_23984_, _23965_, _01538_);
  or (_23985_, _23984_, _23907_);
  and (_23986_, _23985_, _38087_);
  and (_23987_, _23986_, _23983_);
  or (_23988_, _23987_, _23905_);
  and (_40275_, _23988_, _37580_);
  not (_23990_, \oc8051_golden_model_1.PCON [2]);
  nor (_23991_, _38087_, _23990_);
  nor (_23992_, _03662_, _23990_);
  nor (_23993_, _11019_, _08941_);
  or (_23994_, _23993_, _23992_);
  and (_23995_, _23994_, _02173_);
  or (_23996_, _23992_, _04156_);
  and (_23997_, _03662_, _04724_);
  or (_23998_, _23997_, _23992_);
  and (_24000_, _23998_, _02072_);
  and (_24001_, _24000_, _23996_);
  and (_24002_, _11020_, _03662_);
  or (_24003_, _24002_, _23992_);
  and (_24004_, _24003_, _02167_);
  nor (_24005_, _08941_, _03455_);
  or (_24006_, _24005_, _23992_);
  or (_24007_, _24006_, _05249_);
  nor (_24008_, _10905_, _08941_);
  or (_24009_, _24008_, _23992_);
  or (_24011_, _24009_, _02814_);
  and (_24012_, _03662_, \oc8051_golden_model_1.ACC [2]);
  or (_24013_, _24012_, _23992_);
  and (_24014_, _24013_, _02817_);
  nor (_24015_, _02817_, _23990_);
  or (_24016_, _24015_, _02001_);
  or (_24017_, _24016_, _24014_);
  and (_24018_, _24017_, _02840_);
  and (_24019_, _24018_, _24011_);
  and (_24020_, _24006_, _01999_);
  or (_24022_, _24020_, _24019_);
  and (_24023_, _24022_, _02021_);
  and (_24024_, _24013_, _02006_);
  or (_24025_, _24024_, _05994_);
  or (_24026_, _24025_, _24023_);
  and (_24027_, _24026_, _24007_);
  or (_24028_, _24027_, _02528_);
  and (_24029_, _05043_, _03662_);
  or (_24030_, _23992_, _02888_);
  or (_24031_, _24030_, _24029_);
  and (_24033_, _24031_, _24028_);
  or (_24034_, _24033_, _01602_);
  nor (_24035_, _11000_, _08941_);
  or (_24036_, _23992_, _02043_);
  or (_24037_, _24036_, _24035_);
  and (_24038_, _24037_, _01870_);
  and (_24039_, _24038_, _24034_);
  and (_24040_, _23998_, _01869_);
  or (_24041_, _24040_, _02079_);
  or (_24042_, _24041_, _24039_);
  and (_24044_, _11014_, _03662_);
  or (_24045_, _23992_, _02166_);
  or (_24046_, _24045_, _24044_);
  and (_24047_, _24046_, _02912_);
  and (_24048_, _24047_, _24042_);
  or (_24049_, _24048_, _24004_);
  and (_24050_, _24049_, _02176_);
  or (_24051_, _24050_, _24001_);
  and (_24052_, _24051_, _02907_);
  and (_24053_, _24013_, _02177_);
  and (_24055_, _24053_, _23996_);
  or (_24056_, _24055_, _02071_);
  or (_24057_, _24056_, _24052_);
  nor (_24058_, _11013_, _08941_);
  or (_24059_, _23992_, _04788_);
  or (_24060_, _24059_, _24058_);
  and (_24061_, _24060_, _04793_);
  and (_24062_, _24061_, _24057_);
  or (_24063_, _24062_, _23995_);
  and (_24064_, _24063_, _02303_);
  and (_24066_, _24009_, _02201_);
  or (_24067_, _24066_, _01537_);
  or (_24068_, _24067_, _24064_);
  and (_24069_, _11072_, _03662_);
  or (_24070_, _23992_, _01538_);
  or (_24071_, _24070_, _24069_);
  and (_24072_, _24071_, _38087_);
  and (_24073_, _24072_, _24068_);
  or (_24074_, _24073_, _23991_);
  and (_40276_, _24074_, _37580_);
  or (_24075_, _38087_, \oc8051_golden_model_1.PCON [3]);
  and (_24076_, _24075_, _37580_);
  and (_24077_, _08941_, \oc8051_golden_model_1.PCON [3]);
  or (_24078_, _24077_, _04014_);
  and (_24079_, _03662_, _04678_);
  or (_24080_, _24079_, _24077_);
  and (_24081_, _24080_, _02072_);
  and (_24082_, _24081_, _24078_);
  and (_24083_, _11094_, _03662_);
  or (_24084_, _24083_, _24077_);
  and (_24086_, _24084_, _02167_);
  nor (_24087_, _11101_, _08941_);
  or (_24088_, _24087_, _24077_);
  or (_24089_, _24088_, _02814_);
  and (_24090_, _03662_, \oc8051_golden_model_1.ACC [3]);
  or (_24091_, _24090_, _24077_);
  and (_24092_, _24091_, _02817_);
  and (_24093_, _02818_, \oc8051_golden_model_1.PCON [3]);
  or (_24094_, _24093_, _02001_);
  or (_24095_, _24094_, _24092_);
  and (_24097_, _24095_, _02840_);
  and (_24098_, _24097_, _24089_);
  nor (_24099_, _08941_, _03268_);
  or (_24100_, _24099_, _24077_);
  and (_24101_, _24100_, _01999_);
  or (_24102_, _24101_, _24098_);
  and (_24103_, _24102_, _02021_);
  and (_24104_, _24091_, _02006_);
  or (_24105_, _24104_, _05994_);
  or (_24106_, _24105_, _24103_);
  or (_24108_, _24100_, _05249_);
  and (_24109_, _24108_, _24106_);
  or (_24110_, _24109_, _02528_);
  and (_24111_, _04998_, _03662_);
  or (_24112_, _24077_, _02888_);
  or (_24113_, _24112_, _24111_);
  and (_24114_, _24113_, _02043_);
  and (_24115_, _24114_, _24110_);
  nor (_24116_, _11206_, _08941_);
  or (_24117_, _24116_, _24077_);
  and (_24119_, _24117_, _01602_);
  or (_24120_, _24119_, _01869_);
  or (_24121_, _24120_, _24115_);
  or (_24122_, _24080_, _01870_);
  and (_24123_, _24122_, _24121_);
  or (_24124_, _24123_, _02079_);
  and (_24125_, _11222_, _03662_);
  or (_24126_, _24077_, _02166_);
  or (_24127_, _24126_, _24125_);
  and (_24128_, _24127_, _02912_);
  and (_24130_, _24128_, _24124_);
  or (_24131_, _24130_, _24086_);
  and (_24132_, _24131_, _02176_);
  or (_24133_, _24132_, _24082_);
  and (_24134_, _24133_, _02907_);
  and (_24135_, _24091_, _02177_);
  and (_24136_, _24135_, _24078_);
  or (_24137_, _24136_, _02071_);
  or (_24138_, _24137_, _24134_);
  nor (_24139_, _11220_, _08941_);
  or (_24141_, _24077_, _04788_);
  or (_24142_, _24141_, _24139_);
  and (_24143_, _24142_, _04793_);
  and (_24144_, _24143_, _24138_);
  nor (_24145_, _11093_, _08941_);
  or (_24146_, _24145_, _24077_);
  and (_24147_, _24146_, _02173_);
  or (_24148_, _24147_, _02201_);
  or (_24149_, _24148_, _24144_);
  or (_24150_, _24088_, _02303_);
  and (_24152_, _24150_, _01538_);
  and (_24153_, _24152_, _24149_);
  and (_24154_, _11273_, _03662_);
  or (_24155_, _24154_, _24077_);
  and (_24156_, _24155_, _01537_);
  or (_24157_, _24156_, _38088_);
  or (_24158_, _24157_, _24153_);
  and (_40277_, _24158_, _24076_);
  or (_24159_, _38087_, \oc8051_golden_model_1.PCON [4]);
  and (_24160_, _24159_, _37580_);
  and (_24161_, _08941_, \oc8051_golden_model_1.PCON [4]);
  and (_24162_, _11431_, _03662_);
  or (_24163_, _24162_, _24161_);
  and (_24164_, _24163_, _02167_);
  nor (_24165_, _11317_, _08941_);
  or (_24166_, _24165_, _24161_);
  or (_24167_, _24166_, _02814_);
  and (_24168_, _03662_, \oc8051_golden_model_1.ACC [4]);
  or (_24169_, _24168_, _24161_);
  and (_24170_, _24169_, _02817_);
  and (_24172_, _02818_, \oc8051_golden_model_1.PCON [4]);
  or (_24173_, _24172_, _02001_);
  or (_24174_, _24173_, _24170_);
  and (_24175_, _24174_, _02840_);
  and (_24176_, _24175_, _24167_);
  nor (_24177_, _04211_, _08941_);
  or (_24178_, _24177_, _24161_);
  and (_24179_, _24178_, _01999_);
  or (_24180_, _24179_, _24176_);
  and (_24181_, _24180_, _02021_);
  and (_24183_, _24169_, _02006_);
  or (_24184_, _24183_, _05994_);
  or (_24185_, _24184_, _24181_);
  or (_24186_, _24178_, _05249_);
  and (_24187_, _24186_, _24185_);
  or (_24188_, _24187_, _02528_);
  and (_24189_, _05135_, _03662_);
  or (_24190_, _24161_, _02888_);
  or (_24191_, _24190_, _24189_);
  and (_24192_, _24191_, _02043_);
  and (_24194_, _24192_, _24188_);
  nor (_24195_, _11411_, _08941_);
  or (_24196_, _24195_, _24161_);
  and (_24197_, _24196_, _01602_);
  or (_24198_, _24197_, _01869_);
  or (_24199_, _24198_, _24194_);
  and (_24200_, _04694_, _03662_);
  or (_24201_, _24200_, _24161_);
  or (_24202_, _24201_, _01870_);
  and (_24203_, _24202_, _24199_);
  or (_24205_, _24203_, _02079_);
  and (_24206_, _11425_, _03662_);
  or (_24207_, _24161_, _02166_);
  or (_24208_, _24207_, _24206_);
  and (_24209_, _24208_, _02912_);
  and (_24210_, _24209_, _24205_);
  or (_24211_, _24210_, _24164_);
  and (_24212_, _24211_, _02176_);
  or (_24213_, _24161_, _04258_);
  and (_24214_, _24201_, _02072_);
  and (_24216_, _24214_, _24213_);
  or (_24217_, _24216_, _24212_);
  and (_24218_, _24217_, _02907_);
  and (_24219_, _24169_, _02177_);
  and (_24220_, _24219_, _24213_);
  or (_24221_, _24220_, _02071_);
  or (_24222_, _24221_, _24218_);
  nor (_24223_, _11424_, _08941_);
  or (_24224_, _24161_, _04788_);
  or (_24225_, _24224_, _24223_);
  and (_24227_, _24225_, _04793_);
  and (_24228_, _24227_, _24222_);
  nor (_24229_, _11430_, _08941_);
  or (_24230_, _24229_, _24161_);
  and (_24231_, _24230_, _02173_);
  or (_24232_, _24231_, _02201_);
  or (_24233_, _24232_, _24228_);
  or (_24234_, _24166_, _02303_);
  and (_24235_, _24234_, _01538_);
  and (_24236_, _24235_, _24233_);
  and (_24238_, _11487_, _03662_);
  or (_24239_, _24238_, _24161_);
  and (_24240_, _24239_, _01537_);
  or (_24241_, _24240_, _38088_);
  or (_24242_, _24241_, _24236_);
  and (_40278_, _24242_, _24160_);
  or (_24243_, _38087_, \oc8051_golden_model_1.PCON [5]);
  and (_24244_, _24243_, _37580_);
  and (_24245_, _08941_, \oc8051_golden_model_1.PCON [5]);
  and (_24246_, _11635_, _03662_);
  or (_24247_, _24246_, _24245_);
  and (_24248_, _24247_, _02167_);
  nor (_24249_, _11525_, _08941_);
  or (_24250_, _24249_, _24245_);
  or (_24251_, _24250_, _02814_);
  and (_24252_, _03662_, \oc8051_golden_model_1.ACC [5]);
  or (_24253_, _24252_, _24245_);
  and (_24254_, _24253_, _02817_);
  and (_24255_, _02818_, \oc8051_golden_model_1.PCON [5]);
  or (_24256_, _24255_, _02001_);
  or (_24258_, _24256_, _24254_);
  and (_24259_, _24258_, _02840_);
  and (_24260_, _24259_, _24251_);
  nor (_24261_, _03916_, _08941_);
  or (_24262_, _24261_, _24245_);
  and (_24263_, _24262_, _01999_);
  or (_24264_, _24263_, _24260_);
  and (_24265_, _24264_, _02021_);
  and (_24266_, _24253_, _02006_);
  or (_24267_, _24266_, _05994_);
  or (_24269_, _24267_, _24265_);
  or (_24270_, _24262_, _05249_);
  and (_24271_, _24270_, _24269_);
  or (_24272_, _24271_, _02528_);
  and (_24273_, _05090_, _03662_);
  or (_24274_, _24245_, _02888_);
  or (_24275_, _24274_, _24273_);
  and (_24276_, _24275_, _02043_);
  and (_24277_, _24276_, _24272_);
  nor (_24278_, _11615_, _08941_);
  or (_24280_, _24278_, _24245_);
  and (_24281_, _24280_, _01602_);
  or (_24282_, _24281_, _01869_);
  or (_24283_, _24282_, _24277_);
  and (_24284_, _04672_, _03662_);
  or (_24285_, _24284_, _24245_);
  or (_24286_, _24285_, _01870_);
  and (_24287_, _24286_, _24283_);
  or (_24288_, _24287_, _02079_);
  and (_24289_, _11629_, _03662_);
  or (_24291_, _24245_, _02166_);
  or (_24292_, _24291_, _24289_);
  and (_24293_, _24292_, _02912_);
  and (_24294_, _24293_, _24288_);
  or (_24295_, _24294_, _24248_);
  and (_24296_, _24295_, _02176_);
  or (_24297_, _24245_, _03965_);
  and (_24298_, _24285_, _02072_);
  and (_24299_, _24298_, _24297_);
  or (_24300_, _24299_, _24296_);
  and (_24302_, _24300_, _02907_);
  and (_24303_, _24253_, _02177_);
  and (_24304_, _24303_, _24297_);
  or (_24305_, _24304_, _02071_);
  or (_24306_, _24305_, _24302_);
  nor (_24307_, _11628_, _08941_);
  or (_24308_, _24245_, _04788_);
  or (_24309_, _24308_, _24307_);
  and (_24310_, _24309_, _04793_);
  and (_24311_, _24310_, _24306_);
  nor (_24313_, _11634_, _08941_);
  or (_24314_, _24313_, _24245_);
  and (_24315_, _24314_, _02173_);
  or (_24316_, _24315_, _02201_);
  or (_24317_, _24316_, _24311_);
  or (_24318_, _24250_, _02303_);
  and (_24319_, _24318_, _01538_);
  and (_24320_, _24319_, _24317_);
  and (_24321_, _11685_, _03662_);
  or (_24322_, _24321_, _24245_);
  and (_24324_, _24322_, _01537_);
  or (_24325_, _24324_, _38088_);
  or (_24326_, _24325_, _24320_);
  and (_40279_, _24326_, _24244_);
  or (_24327_, _38087_, \oc8051_golden_model_1.PCON [6]);
  and (_24328_, _24327_, _37580_);
  and (_24329_, _08941_, \oc8051_golden_model_1.PCON [6]);
  and (_24330_, _11709_, _03662_);
  or (_24331_, _24330_, _24329_);
  and (_24332_, _24331_, _02167_);
  nor (_24333_, _11730_, _08941_);
  or (_24334_, _24333_, _24329_);
  or (_24335_, _24334_, _02814_);
  and (_24336_, _03662_, \oc8051_golden_model_1.ACC [6]);
  or (_24337_, _24336_, _24329_);
  and (_24338_, _24337_, _02817_);
  and (_24339_, _02818_, \oc8051_golden_model_1.PCON [6]);
  or (_24340_, _24339_, _02001_);
  or (_24341_, _24340_, _24338_);
  and (_24342_, _24341_, _02840_);
  and (_24344_, _24342_, _24335_);
  nor (_24345_, _03808_, _08941_);
  or (_24346_, _24345_, _24329_);
  and (_24347_, _24346_, _01999_);
  or (_24348_, _24347_, _24344_);
  and (_24349_, _24348_, _02021_);
  and (_24350_, _24337_, _02006_);
  or (_24351_, _24350_, _05994_);
  or (_24352_, _24351_, _24349_);
  or (_24353_, _24346_, _05249_);
  and (_24355_, _24353_, _24352_);
  or (_24356_, _24355_, _02528_);
  and (_24357_, _04861_, _03662_);
  or (_24358_, _24329_, _02888_);
  or (_24359_, _24358_, _24357_);
  and (_24360_, _24359_, _02043_);
  and (_24361_, _24360_, _24356_);
  nor (_24362_, _11820_, _08941_);
  or (_24363_, _24362_, _24329_);
  and (_24364_, _24363_, _01602_);
  or (_24366_, _24364_, _01869_);
  or (_24367_, _24366_, _24361_);
  and (_24368_, _09920_, _03662_);
  or (_24369_, _24368_, _24329_);
  or (_24370_, _24369_, _01870_);
  and (_24371_, _24370_, _24367_);
  or (_24372_, _24371_, _02079_);
  and (_24373_, _11835_, _03662_);
  or (_24374_, _24329_, _02166_);
  or (_24375_, _24374_, _24373_);
  and (_24377_, _24375_, _02912_);
  and (_24378_, _24377_, _24372_);
  or (_24379_, _24378_, _24332_);
  and (_24380_, _24379_, _02176_);
  or (_24381_, _24329_, _03863_);
  and (_24382_, _24369_, _02072_);
  and (_24383_, _24382_, _24381_);
  or (_24384_, _24383_, _24380_);
  and (_24385_, _24384_, _02907_);
  and (_24386_, _24337_, _02177_);
  and (_24388_, _24386_, _24381_);
  or (_24389_, _24388_, _02071_);
  or (_24390_, _24389_, _24385_);
  nor (_24391_, _11833_, _08941_);
  or (_24392_, _24329_, _04788_);
  or (_24393_, _24392_, _24391_);
  and (_24394_, _24393_, _04793_);
  and (_24395_, _24394_, _24390_);
  nor (_24396_, _11708_, _08941_);
  or (_24397_, _24396_, _24329_);
  and (_24399_, _24397_, _02173_);
  or (_24400_, _24399_, _02201_);
  or (_24401_, _24400_, _24395_);
  or (_24402_, _24334_, _02303_);
  and (_24403_, _24402_, _01538_);
  and (_24404_, _24403_, _24401_);
  and (_24405_, _11887_, _03662_);
  or (_24406_, _24405_, _24329_);
  and (_24407_, _24406_, _01537_);
  or (_24408_, _24407_, _38088_);
  or (_24410_, _24408_, _24404_);
  and (_40281_, _24410_, _24328_);
  and (_24411_, _38088_, \oc8051_golden_model_1.SBUF [0]);
  and (_24412_, _09019_, \oc8051_golden_model_1.SBUF [0]);
  and (_24413_, _03625_, \oc8051_golden_model_1.ACC [0]);
  or (_24414_, _24413_, _24412_);
  and (_24415_, _24414_, _02006_);
  or (_24416_, _24415_, _05994_);
  nor (_24417_, _04106_, _09019_);
  or (_24418_, _24417_, _24412_);
  and (_24419_, _24418_, _02001_);
  and (_24420_, _02818_, \oc8051_golden_model_1.SBUF [0]);
  and (_24421_, _24414_, _02817_);
  or (_24422_, _24421_, _24420_);
  and (_24423_, _24422_, _02814_);
  or (_24424_, _24423_, _01999_);
  or (_24425_, _24424_, _24419_);
  and (_24426_, _24425_, _02021_);
  or (_24427_, _24426_, _24416_);
  and (_24428_, _03625_, _03028_);
  or (_24430_, _24412_, _23851_);
  or (_24431_, _24430_, _24428_);
  and (_24432_, _24431_, _24427_);
  or (_24433_, _24432_, _02528_);
  and (_24434_, _04952_, _03625_);
  or (_24435_, _24412_, _02888_);
  or (_24436_, _24435_, _24434_);
  and (_24437_, _24436_, _24433_);
  or (_24438_, _24437_, _01602_);
  nor (_24439_, _10600_, _09019_);
  or (_24441_, _24439_, _24412_);
  or (_24442_, _24441_, _02043_);
  and (_24443_, _24442_, _01870_);
  and (_24444_, _24443_, _24438_);
  and (_24445_, _03625_, _04562_);
  or (_24446_, _24445_, _24412_);
  and (_24447_, _24446_, _01869_);
  or (_24448_, _24447_, _02079_);
  or (_24449_, _24448_, _24444_);
  and (_24450_, _10614_, _03625_);
  or (_24452_, _24450_, _24412_);
  or (_24453_, _24452_, _02166_);
  and (_24454_, _24453_, _24449_);
  or (_24455_, _24454_, _02167_);
  and (_24456_, _10620_, _03625_);
  or (_24457_, _24412_, _02912_);
  or (_24458_, _24457_, _24456_);
  and (_24459_, _24458_, _02176_);
  and (_24460_, _24459_, _24455_);
  nand (_24461_, _24446_, _02072_);
  nor (_24463_, _24461_, _24417_);
  or (_24464_, _24463_, _24460_);
  and (_24465_, _24464_, _02907_);
  or (_24466_, _24412_, _04106_);
  and (_24467_, _24414_, _02177_);
  and (_24468_, _24467_, _24466_);
  or (_24469_, _24468_, _02071_);
  or (_24470_, _24469_, _24465_);
  nor (_24471_, _10613_, _09019_);
  or (_24472_, _24412_, _04788_);
  or (_24474_, _24472_, _24471_);
  and (_24475_, _24474_, _04793_);
  and (_24476_, _24475_, _24470_);
  nor (_24477_, _10619_, _09019_);
  or (_24478_, _24477_, _24412_);
  and (_24479_, _24478_, _02173_);
  or (_24480_, _24479_, _15577_);
  or (_24481_, _24480_, _24476_);
  or (_24482_, _24418_, _02743_);
  and (_24483_, _24482_, _38087_);
  and (_24485_, _24483_, _24481_);
  or (_24486_, _24485_, _24411_);
  and (_40282_, _24486_, _37580_);
  and (_24487_, _38088_, \oc8051_golden_model_1.SBUF [1]);
  or (_24488_, _03625_, \oc8051_golden_model_1.SBUF [1]);
  and (_24489_, _10698_, _03625_);
  not (_24490_, _24489_);
  and (_24491_, _24490_, _24488_);
  or (_24492_, _24491_, _02814_);
  nand (_24493_, _03625_, _01613_);
  and (_24495_, _24493_, _24488_);
  and (_24496_, _24495_, _02817_);
  and (_24497_, _02818_, \oc8051_golden_model_1.SBUF [1]);
  or (_24498_, _24497_, _02001_);
  or (_24499_, _24498_, _24496_);
  and (_24500_, _24499_, _02840_);
  and (_24501_, _24500_, _24492_);
  nand (_24502_, _03625_, _02811_);
  and (_24503_, _24502_, _24488_);
  and (_24504_, _24503_, _01999_);
  or (_24505_, _24504_, _24501_);
  and (_24506_, _24505_, _02021_);
  and (_24507_, _24495_, _02006_);
  or (_24508_, _24507_, _05994_);
  or (_24509_, _24508_, _24506_);
  or (_24510_, _24503_, _05249_);
  and (_24511_, _24510_, _02888_);
  and (_24512_, _24511_, _24509_);
  or (_24513_, _04907_, _09019_);
  and (_24514_, _24488_, _02528_);
  and (_24516_, _24514_, _24513_);
  or (_24517_, _24516_, _24512_);
  and (_24518_, _24517_, _02043_);
  nand (_24519_, _10802_, _03625_);
  and (_24520_, _24488_, _01602_);
  and (_24521_, _24520_, _24519_);
  or (_24522_, _24521_, _24518_);
  and (_24523_, _24522_, _01870_);
  nand (_24524_, _03625_, _02687_);
  and (_24525_, _24488_, _01869_);
  and (_24527_, _24525_, _24524_);
  or (_24528_, _24527_, _24523_);
  and (_24529_, _24528_, _02166_);
  or (_24530_, _10816_, _09019_);
  and (_24531_, _24488_, _02079_);
  and (_24532_, _24531_, _24530_);
  or (_24533_, _24532_, _24529_);
  and (_24534_, _24533_, _02912_);
  or (_24535_, _10822_, _09019_);
  and (_24536_, _24488_, _02167_);
  and (_24538_, _24536_, _24535_);
  or (_24539_, _24538_, _24534_);
  and (_24540_, _24539_, _02176_);
  or (_24541_, _10692_, _09019_);
  and (_24542_, _24488_, _02072_);
  and (_24543_, _24542_, _24541_);
  or (_24544_, _24543_, _24540_);
  and (_24545_, _24544_, _02907_);
  and (_24546_, _09019_, \oc8051_golden_model_1.SBUF [1]);
  or (_24547_, _24546_, _04058_);
  and (_24549_, _24495_, _02177_);
  and (_24550_, _24549_, _24547_);
  or (_24551_, _24550_, _24545_);
  and (_24552_, _24551_, _02174_);
  or (_24553_, _24493_, _04058_);
  and (_24554_, _24488_, _02173_);
  and (_24555_, _24554_, _24553_);
  or (_24556_, _24555_, _02201_);
  or (_24557_, _24524_, _04058_);
  and (_24558_, _24488_, _02071_);
  and (_24560_, _24558_, _24557_);
  or (_24561_, _24560_, _24556_);
  or (_24562_, _24561_, _24552_);
  or (_24563_, _24491_, _02303_);
  and (_24564_, _24563_, _24562_);
  or (_24565_, _24564_, _01537_);
  or (_24566_, _24546_, _01538_);
  or (_24567_, _24566_, _24489_);
  and (_24568_, _24567_, _38087_);
  and (_24569_, _24568_, _24565_);
  or (_24571_, _24569_, _24487_);
  and (_40283_, _24571_, _37580_);
  and (_24572_, _38088_, \oc8051_golden_model_1.SBUF [2]);
  and (_24573_, _09019_, \oc8051_golden_model_1.SBUF [2]);
  nor (_24574_, _11019_, _09019_);
  or (_24575_, _24574_, _24573_);
  and (_24576_, _24575_, _02173_);
  and (_24577_, _11020_, _03625_);
  or (_24578_, _24577_, _24573_);
  and (_24579_, _24578_, _02167_);
  nor (_24581_, _10905_, _09019_);
  or (_24582_, _24581_, _24573_);
  or (_24583_, _24582_, _02814_);
  and (_24584_, _03625_, \oc8051_golden_model_1.ACC [2]);
  or (_24585_, _24584_, _24573_);
  and (_24586_, _24585_, _02817_);
  and (_24587_, _02818_, \oc8051_golden_model_1.SBUF [2]);
  or (_24588_, _24587_, _02001_);
  or (_24589_, _24588_, _24586_);
  and (_24590_, _24589_, _02840_);
  and (_24591_, _24590_, _24583_);
  nor (_24592_, _09019_, _03455_);
  or (_24593_, _24592_, _24573_);
  and (_24594_, _24593_, _01999_);
  or (_24595_, _24594_, _24591_);
  and (_24596_, _24595_, _02021_);
  and (_24597_, _24585_, _02006_);
  or (_24598_, _24597_, _05994_);
  or (_24599_, _24598_, _24596_);
  or (_24600_, _24593_, _05249_);
  and (_24602_, _24600_, _24599_);
  or (_24603_, _24602_, _02528_);
  and (_24604_, _05043_, _03625_);
  or (_24605_, _24573_, _02888_);
  or (_24606_, _24605_, _24604_);
  and (_24607_, _24606_, _24603_);
  or (_24608_, _24607_, _01602_);
  nor (_24609_, _11000_, _09019_);
  or (_24610_, _24573_, _02043_);
  or (_24611_, _24610_, _24609_);
  and (_24613_, _24611_, _01870_);
  and (_24614_, _24613_, _24608_);
  and (_24615_, _03625_, _04724_);
  or (_24616_, _24615_, _24573_);
  and (_24617_, _24616_, _01869_);
  or (_24618_, _24617_, _02079_);
  or (_24619_, _24618_, _24614_);
  and (_24620_, _11014_, _03625_);
  or (_24621_, _24573_, _02166_);
  or (_24622_, _24621_, _24620_);
  and (_24624_, _24622_, _02912_);
  and (_24625_, _24624_, _24619_);
  or (_24626_, _24625_, _24579_);
  and (_24627_, _24626_, _02176_);
  or (_24628_, _24573_, _04156_);
  and (_24629_, _24616_, _02072_);
  and (_24630_, _24629_, _24628_);
  or (_24631_, _24630_, _24627_);
  and (_24632_, _24631_, _02907_);
  and (_24633_, _24585_, _02177_);
  and (_24634_, _24633_, _24628_);
  or (_24635_, _24634_, _02071_);
  or (_24636_, _24635_, _24632_);
  nor (_24637_, _11013_, _09019_);
  or (_24638_, _24573_, _04788_);
  or (_24639_, _24638_, _24637_);
  and (_24640_, _24639_, _04793_);
  and (_24641_, _24640_, _24636_);
  or (_24642_, _24641_, _24576_);
  and (_24643_, _24642_, _02303_);
  and (_24645_, _24582_, _02201_);
  or (_24646_, _24645_, _01537_);
  or (_24647_, _24646_, _24643_);
  and (_24648_, _11072_, _03625_);
  or (_24649_, _24573_, _01538_);
  or (_24650_, _24649_, _24648_);
  and (_24651_, _24650_, _38087_);
  and (_24652_, _24651_, _24647_);
  or (_24653_, _24652_, _24572_);
  and (_40285_, _24653_, _37580_);
  or (_24655_, _38087_, \oc8051_golden_model_1.SBUF [3]);
  and (_24656_, _24655_, _37580_);
  and (_24657_, _09019_, \oc8051_golden_model_1.SBUF [3]);
  or (_24658_, _24657_, _04014_);
  and (_24659_, _03625_, _04678_);
  or (_24660_, _24659_, _24657_);
  and (_24661_, _24660_, _02072_);
  and (_24662_, _24661_, _24658_);
  and (_24663_, _11094_, _03625_);
  or (_24664_, _24663_, _24657_);
  and (_24666_, _24664_, _02167_);
  nor (_24667_, _11101_, _09019_);
  or (_24668_, _24667_, _24657_);
  or (_24669_, _24668_, _02814_);
  and (_24670_, _03625_, \oc8051_golden_model_1.ACC [3]);
  or (_24671_, _24670_, _24657_);
  and (_24672_, _24671_, _02817_);
  and (_24673_, _02818_, \oc8051_golden_model_1.SBUF [3]);
  or (_24674_, _24673_, _02001_);
  or (_24675_, _24674_, _24672_);
  and (_24676_, _24675_, _02840_);
  and (_24677_, _24676_, _24669_);
  nor (_24678_, _09019_, _03268_);
  or (_24679_, _24678_, _24657_);
  and (_24680_, _24679_, _01999_);
  or (_24681_, _24680_, _24677_);
  and (_24682_, _24681_, _02021_);
  and (_24683_, _24671_, _02006_);
  or (_24684_, _24683_, _05994_);
  or (_24685_, _24684_, _24682_);
  or (_24687_, _24679_, _05249_);
  and (_24688_, _24687_, _24685_);
  or (_24689_, _24688_, _02528_);
  and (_24690_, _04998_, _03625_);
  or (_24691_, _24657_, _02888_);
  or (_24692_, _24691_, _24690_);
  and (_24693_, _24692_, _02043_);
  and (_24694_, _24693_, _24689_);
  nor (_24695_, _11206_, _09019_);
  or (_24696_, _24695_, _24657_);
  and (_24698_, _24696_, _01602_);
  or (_24699_, _24698_, _01869_);
  or (_24700_, _24699_, _24694_);
  or (_24701_, _24660_, _01870_);
  and (_24702_, _24701_, _24700_);
  or (_24703_, _24702_, _02079_);
  and (_24704_, _11222_, _03625_);
  or (_24705_, _24657_, _02166_);
  or (_24706_, _24705_, _24704_);
  and (_24707_, _24706_, _02912_);
  and (_24709_, _24707_, _24703_);
  or (_24710_, _24709_, _24666_);
  and (_24711_, _24710_, _02176_);
  or (_24712_, _24711_, _24662_);
  and (_24713_, _24712_, _02907_);
  and (_24714_, _24671_, _02177_);
  and (_24715_, _24714_, _24658_);
  or (_24716_, _24715_, _02071_);
  or (_24717_, _24716_, _24713_);
  nor (_24718_, _11220_, _09019_);
  or (_24719_, _24657_, _04788_);
  or (_24720_, _24719_, _24718_);
  and (_24721_, _24720_, _04793_);
  and (_24722_, _24721_, _24717_);
  nor (_24723_, _11093_, _09019_);
  or (_24724_, _24723_, _24657_);
  and (_24725_, _24724_, _02173_);
  or (_24726_, _24725_, _02201_);
  or (_24727_, _24726_, _24722_);
  or (_24728_, _24668_, _02303_);
  and (_24730_, _24728_, _01538_);
  and (_24731_, _24730_, _24727_);
  and (_24732_, _11273_, _03625_);
  or (_24733_, _24732_, _24657_);
  and (_24734_, _24733_, _01537_);
  or (_24735_, _24734_, _38088_);
  or (_24736_, _24735_, _24731_);
  and (_40286_, _24736_, _24656_);
  or (_24737_, _38087_, \oc8051_golden_model_1.SBUF [4]);
  and (_24738_, _24737_, _37580_);
  and (_24740_, _09019_, \oc8051_golden_model_1.SBUF [4]);
  and (_24741_, _11431_, _03625_);
  or (_24742_, _24741_, _24740_);
  and (_24743_, _24742_, _02167_);
  nor (_24744_, _11317_, _09019_);
  or (_24745_, _24744_, _24740_);
  or (_24746_, _24745_, _02814_);
  and (_24747_, _03625_, \oc8051_golden_model_1.ACC [4]);
  or (_24748_, _24747_, _24740_);
  and (_24749_, _24748_, _02817_);
  and (_24751_, _02818_, \oc8051_golden_model_1.SBUF [4]);
  or (_24752_, _24751_, _02001_);
  or (_24753_, _24752_, _24749_);
  and (_24754_, _24753_, _02840_);
  and (_24755_, _24754_, _24746_);
  nor (_24756_, _04211_, _09019_);
  or (_24757_, _24756_, _24740_);
  and (_24758_, _24757_, _01999_);
  or (_24759_, _24758_, _24755_);
  and (_24760_, _24759_, _02021_);
  and (_24761_, _24748_, _02006_);
  or (_24762_, _24761_, _05994_);
  or (_24763_, _24762_, _24760_);
  or (_24764_, _24757_, _05249_);
  and (_24765_, _24764_, _24763_);
  or (_24766_, _24765_, _02528_);
  and (_24767_, _05135_, _03625_);
  or (_24768_, _24740_, _02888_);
  or (_24769_, _24768_, _24767_);
  and (_24770_, _24769_, _02043_);
  and (_24772_, _24770_, _24766_);
  nor (_24773_, _11411_, _09019_);
  or (_24774_, _24773_, _24740_);
  and (_24775_, _24774_, _01602_);
  or (_24776_, _24775_, _01869_);
  or (_24777_, _24776_, _24772_);
  and (_24778_, _04694_, _03625_);
  or (_24779_, _24778_, _24740_);
  or (_24780_, _24779_, _01870_);
  and (_24781_, _24780_, _24777_);
  or (_24783_, _24781_, _02079_);
  and (_24784_, _11425_, _03625_);
  or (_24785_, _24740_, _02166_);
  or (_24786_, _24785_, _24784_);
  and (_24787_, _24786_, _02912_);
  and (_24788_, _24787_, _24783_);
  or (_24789_, _24788_, _24743_);
  and (_24790_, _24789_, _02176_);
  or (_24791_, _24740_, _04258_);
  and (_24792_, _24779_, _02072_);
  and (_24794_, _24792_, _24791_);
  or (_24795_, _24794_, _24790_);
  and (_24796_, _24795_, _02907_);
  and (_24797_, _24748_, _02177_);
  and (_24798_, _24797_, _24791_);
  or (_24799_, _24798_, _02071_);
  or (_24800_, _24799_, _24796_);
  nor (_24801_, _11424_, _09019_);
  or (_24802_, _24740_, _04788_);
  or (_24803_, _24802_, _24801_);
  and (_24804_, _24803_, _04793_);
  and (_24805_, _24804_, _24800_);
  nor (_24806_, _11430_, _09019_);
  or (_24807_, _24806_, _24740_);
  and (_24808_, _24807_, _02173_);
  or (_24809_, _24808_, _02201_);
  or (_24810_, _24809_, _24805_);
  or (_24811_, _24745_, _02303_);
  and (_24812_, _24811_, _01538_);
  and (_24813_, _24812_, _24810_);
  and (_24815_, _11487_, _03625_);
  or (_24816_, _24815_, _24740_);
  and (_24817_, _24816_, _01537_);
  or (_24818_, _24817_, _38088_);
  or (_24819_, _24818_, _24813_);
  and (_40287_, _24819_, _24738_);
  or (_24820_, _38087_, \oc8051_golden_model_1.SBUF [5]);
  and (_24821_, _24820_, _37580_);
  and (_24822_, _09019_, \oc8051_golden_model_1.SBUF [5]);
  and (_24823_, _11635_, _03625_);
  or (_24825_, _24823_, _24822_);
  and (_24826_, _24825_, _02167_);
  nor (_24827_, _11525_, _09019_);
  or (_24828_, _24827_, _24822_);
  or (_24829_, _24828_, _02814_);
  and (_24830_, _03625_, \oc8051_golden_model_1.ACC [5]);
  or (_24831_, _24830_, _24822_);
  and (_24832_, _24831_, _02817_);
  and (_24833_, _02818_, \oc8051_golden_model_1.SBUF [5]);
  or (_24834_, _24833_, _02001_);
  or (_24836_, _24834_, _24832_);
  and (_24837_, _24836_, _02840_);
  and (_24838_, _24837_, _24829_);
  nor (_24839_, _03916_, _09019_);
  or (_24840_, _24839_, _24822_);
  and (_24841_, _24840_, _01999_);
  or (_24842_, _24841_, _24838_);
  and (_24843_, _24842_, _02021_);
  and (_24844_, _24831_, _02006_);
  or (_24845_, _24844_, _05994_);
  or (_24846_, _24845_, _24843_);
  or (_24847_, _24840_, _05249_);
  and (_24848_, _24847_, _24846_);
  or (_24849_, _24848_, _02528_);
  and (_24850_, _05090_, _03625_);
  or (_24851_, _24822_, _02888_);
  or (_24852_, _24851_, _24850_);
  and (_24853_, _24852_, _02043_);
  and (_24854_, _24853_, _24849_);
  nor (_24855_, _11615_, _09019_);
  or (_24857_, _24855_, _24822_);
  and (_24858_, _24857_, _01602_);
  or (_24859_, _24858_, _01869_);
  or (_24860_, _24859_, _24854_);
  and (_24861_, _04672_, _03625_);
  or (_24862_, _24861_, _24822_);
  or (_24863_, _24862_, _01870_);
  and (_24864_, _24863_, _24860_);
  or (_24865_, _24864_, _02079_);
  and (_24866_, _11629_, _03625_);
  or (_24868_, _24822_, _02166_);
  or (_24869_, _24868_, _24866_);
  and (_24870_, _24869_, _02912_);
  and (_24871_, _24870_, _24865_);
  or (_24872_, _24871_, _24826_);
  and (_24873_, _24872_, _02176_);
  or (_24874_, _24822_, _03965_);
  and (_24875_, _24862_, _02072_);
  and (_24876_, _24875_, _24874_);
  or (_24877_, _24876_, _24873_);
  and (_24879_, _24877_, _02907_);
  and (_24880_, _24831_, _02177_);
  and (_24881_, _24880_, _24874_);
  or (_24882_, _24881_, _02071_);
  or (_24883_, _24882_, _24879_);
  nor (_24884_, _11628_, _09019_);
  or (_24885_, _24822_, _04788_);
  or (_24886_, _24885_, _24884_);
  and (_24887_, _24886_, _04793_);
  and (_24888_, _24887_, _24883_);
  nor (_24889_, _11634_, _09019_);
  or (_24890_, _24889_, _24822_);
  and (_24891_, _24890_, _02173_);
  or (_24892_, _24891_, _02201_);
  or (_24893_, _24892_, _24888_);
  or (_24894_, _24828_, _02303_);
  and (_24895_, _24894_, _01538_);
  and (_24896_, _24895_, _24893_);
  and (_24897_, _11685_, _03625_);
  or (_24898_, _24897_, _24822_);
  and (_24900_, _24898_, _01537_);
  or (_24901_, _24900_, _38088_);
  or (_24902_, _24901_, _24896_);
  and (_40288_, _24902_, _24821_);
  or (_24903_, _38087_, \oc8051_golden_model_1.SBUF [6]);
  and (_24904_, _24903_, _37580_);
  and (_24905_, _09019_, \oc8051_golden_model_1.SBUF [6]);
  and (_24906_, _11709_, _03625_);
  or (_24907_, _24906_, _24905_);
  and (_24908_, _24907_, _02167_);
  nor (_24910_, _03808_, _09019_);
  or (_24911_, _24910_, _24905_);
  or (_24912_, _24911_, _05249_);
  nor (_24913_, _11730_, _09019_);
  or (_24914_, _24913_, _24905_);
  or (_24915_, _24914_, _02814_);
  and (_24916_, _03625_, \oc8051_golden_model_1.ACC [6]);
  or (_24917_, _24916_, _24905_);
  and (_24918_, _24917_, _02817_);
  and (_24919_, _02818_, \oc8051_golden_model_1.SBUF [6]);
  or (_24921_, _24919_, _02001_);
  or (_24922_, _24921_, _24918_);
  and (_24923_, _24922_, _02840_);
  and (_24924_, _24923_, _24915_);
  and (_24925_, _24911_, _01999_);
  or (_24926_, _24925_, _24924_);
  and (_24927_, _24926_, _02021_);
  and (_24928_, _24917_, _02006_);
  or (_24929_, _24928_, _05994_);
  or (_24930_, _24929_, _24927_);
  and (_24932_, _24930_, _24912_);
  or (_24933_, _24932_, _02528_);
  and (_24934_, _04861_, _03625_);
  or (_24935_, _24905_, _02888_);
  or (_24936_, _24935_, _24934_);
  and (_24937_, _24936_, _02043_);
  and (_24938_, _24937_, _24933_);
  nor (_24939_, _11820_, _09019_);
  or (_24940_, _24939_, _24905_);
  and (_24941_, _24940_, _01602_);
  or (_24943_, _24941_, _01869_);
  or (_24944_, _24943_, _24938_);
  and (_24945_, _09920_, _03625_);
  or (_24946_, _24945_, _24905_);
  or (_24947_, _24946_, _01870_);
  and (_24948_, _24947_, _24944_);
  or (_24949_, _24948_, _02079_);
  and (_24950_, _11835_, _03625_);
  or (_24951_, _24905_, _02166_);
  or (_24952_, _24951_, _24950_);
  and (_24954_, _24952_, _02912_);
  and (_24955_, _24954_, _24949_);
  or (_24956_, _24955_, _24908_);
  and (_24957_, _24956_, _02176_);
  or (_24958_, _24905_, _03863_);
  and (_24959_, _24946_, _02072_);
  and (_24960_, _24959_, _24958_);
  or (_24961_, _24960_, _24957_);
  and (_24962_, _24961_, _02907_);
  and (_24963_, _24917_, _02177_);
  and (_24965_, _24963_, _24958_);
  or (_24966_, _24965_, _02071_);
  or (_24967_, _24966_, _24962_);
  nor (_24968_, _11833_, _09019_);
  or (_24969_, _24905_, _04788_);
  or (_24970_, _24969_, _24968_);
  and (_24971_, _24970_, _04793_);
  and (_24972_, _24971_, _24967_);
  nor (_24973_, _11708_, _09019_);
  or (_24974_, _24973_, _24905_);
  and (_24976_, _24974_, _02173_);
  or (_24977_, _24976_, _02201_);
  or (_24978_, _24977_, _24972_);
  or (_24979_, _24914_, _02303_);
  and (_24980_, _24979_, _01538_);
  and (_24981_, _24980_, _24978_);
  and (_24982_, _11887_, _03625_);
  or (_24983_, _24982_, _24905_);
  and (_24984_, _24983_, _01537_);
  or (_24985_, _24984_, _38088_);
  or (_24987_, _24985_, _24981_);
  and (_40289_, _24987_, _24904_);
  and (_24988_, _38088_, \oc8051_golden_model_1.SCON [0]);
  and (_24989_, _09096_, \oc8051_golden_model_1.SCON [0]);
  and (_24990_, _10620_, _03716_);
  or (_24991_, _24990_, _24989_);
  and (_24992_, _24991_, _02167_);
  and (_24993_, _03716_, _03028_);
  or (_24994_, _24993_, _24989_);
  or (_24995_, _24994_, _05249_);
  nor (_24997_, _04106_, _09096_);
  or (_24998_, _24997_, _24989_);
  or (_24999_, _24998_, _02814_);
  and (_25000_, _03716_, \oc8051_golden_model_1.ACC [0]);
  or (_25001_, _25000_, _24989_);
  and (_25002_, _25001_, _02817_);
  and (_25003_, _02818_, \oc8051_golden_model_1.SCON [0]);
  or (_25004_, _25003_, _02001_);
  or (_25005_, _25004_, _25002_);
  and (_25006_, _25005_, _02024_);
  and (_25008_, _25006_, _24999_);
  and (_25009_, _09104_, \oc8051_golden_model_1.SCON [0]);
  and (_25010_, _10510_, _04331_);
  or (_25011_, _25010_, _25009_);
  and (_25012_, _25011_, _02007_);
  or (_25013_, _25012_, _25008_);
  and (_25014_, _25013_, _02840_);
  and (_25015_, _24994_, _01999_);
  or (_25016_, _25015_, _02006_);
  or (_25017_, _25016_, _25014_);
  or (_25019_, _25001_, _02021_);
  and (_25020_, _25019_, _02025_);
  and (_25021_, _25020_, _25017_);
  and (_25022_, _24989_, _01997_);
  or (_25023_, _25022_, _01991_);
  or (_25024_, _25023_, _25021_);
  or (_25025_, _24998_, _02861_);
  and (_25026_, _25025_, _02408_);
  and (_25027_, _25026_, _25024_);
  nor (_25028_, _10542_, _09104_);
  or (_25030_, _25028_, _25009_);
  and (_25031_, _25030_, _01875_);
  or (_25032_, _25031_, _05994_);
  or (_25033_, _25032_, _25027_);
  and (_25034_, _25033_, _24995_);
  or (_25035_, _25034_, _02528_);
  and (_25036_, _04952_, _03716_);
  or (_25037_, _24989_, _02888_);
  or (_25038_, _25037_, _25036_);
  and (_25039_, _25038_, _02043_);
  and (_25041_, _25039_, _25035_);
  nor (_25042_, _10600_, _09096_);
  or (_25043_, _25042_, _24989_);
  and (_25044_, _25043_, _01602_);
  or (_25045_, _25044_, _01869_);
  or (_25046_, _25045_, _25041_);
  and (_25047_, _03716_, _04562_);
  or (_25048_, _25047_, _24989_);
  or (_25049_, _25048_, _01870_);
  and (_25050_, _25049_, _25046_);
  or (_25052_, _25050_, _02079_);
  and (_25053_, _10614_, _03716_);
  or (_25054_, _24989_, _02166_);
  or (_25055_, _25054_, _25053_);
  and (_25056_, _25055_, _02912_);
  and (_25057_, _25056_, _25052_);
  or (_25058_, _25057_, _24992_);
  and (_25059_, _25058_, _02176_);
  nand (_25060_, _25048_, _02072_);
  nor (_25061_, _25060_, _24997_);
  or (_25063_, _25061_, _25059_);
  and (_25064_, _25063_, _02907_);
  or (_25065_, _24989_, _04106_);
  and (_25066_, _25001_, _02177_);
  and (_25067_, _25066_, _25065_);
  or (_25068_, _25067_, _02071_);
  or (_25069_, _25068_, _25064_);
  nor (_25070_, _10613_, _09096_);
  or (_25071_, _24989_, _04788_);
  or (_25072_, _25071_, _25070_);
  and (_25074_, _25072_, _04793_);
  and (_25075_, _25074_, _25069_);
  nor (_25076_, _10619_, _09096_);
  or (_25077_, _25076_, _24989_);
  and (_25078_, _25077_, _02173_);
  or (_25079_, _25078_, _02201_);
  or (_25080_, _25079_, _25075_);
  or (_25081_, _24998_, _02303_);
  and (_25082_, _25081_, _01887_);
  and (_25083_, _25082_, _25080_);
  and (_25085_, _24989_, _01860_);
  or (_25086_, _25085_, _01537_);
  or (_25087_, _25086_, _25083_);
  or (_25088_, _24998_, _01538_);
  and (_25089_, _25088_, _38087_);
  and (_25090_, _25089_, _25087_);
  or (_25091_, _25090_, _24988_);
  and (_40291_, _25091_, _37580_);
  and (_25092_, _38088_, \oc8051_golden_model_1.SCON [1]);
  and (_25093_, _09096_, \oc8051_golden_model_1.SCON [1]);
  nor (_25095_, _09096_, _02811_);
  or (_25096_, _25095_, _25093_);
  and (_25097_, _25096_, _01999_);
  and (_25098_, _09104_, \oc8051_golden_model_1.SCON [1]);
  and (_25099_, _10710_, _04331_);
  or (_25100_, _25099_, _25098_);
  or (_25101_, _25100_, _02024_);
  or (_25102_, _03716_, \oc8051_golden_model_1.SCON [1]);
  and (_25103_, _10698_, _03716_);
  not (_25104_, _25103_);
  and (_25106_, _25104_, _25102_);
  and (_25107_, _25106_, _02001_);
  nand (_25108_, _03716_, _01613_);
  and (_25109_, _25108_, _25102_);
  and (_25110_, _25109_, _02817_);
  and (_25111_, _02818_, \oc8051_golden_model_1.SCON [1]);
  or (_25112_, _25111_, _25110_);
  and (_25113_, _25112_, _02814_);
  or (_25114_, _25113_, _02007_);
  or (_25115_, _25114_, _25107_);
  and (_25117_, _25115_, _25101_);
  and (_25118_, _25117_, _02840_);
  or (_25119_, _25118_, _25097_);
  or (_25120_, _25119_, _02006_);
  or (_25121_, _25109_, _02021_);
  and (_25122_, _25121_, _02025_);
  and (_25123_, _25122_, _25120_);
  and (_25124_, _10696_, _04331_);
  or (_25125_, _25124_, _25098_);
  and (_25126_, _25125_, _01997_);
  or (_25128_, _25126_, _01991_);
  or (_25129_, _25128_, _25123_);
  or (_25130_, _25098_, _10725_);
  and (_25131_, _25130_, _25100_);
  or (_25132_, _25131_, _02861_);
  and (_25133_, _25132_, _02408_);
  and (_25134_, _25133_, _25129_);
  nor (_25135_, _10742_, _09104_);
  or (_25136_, _25135_, _25098_);
  and (_25137_, _25136_, _01875_);
  or (_25139_, _25137_, _05994_);
  or (_25140_, _25139_, _25134_);
  or (_25141_, _25096_, _05249_);
  and (_25142_, _25141_, _25140_);
  or (_25143_, _25142_, _02528_);
  and (_25144_, _04907_, _03716_);
  or (_25145_, _25093_, _02888_);
  or (_25146_, _25145_, _25144_);
  and (_25147_, _25146_, _02043_);
  and (_25148_, _25147_, _25143_);
  nor (_25149_, _10802_, _09096_);
  or (_25150_, _25149_, _25093_);
  and (_25151_, _25150_, _01602_);
  or (_25152_, _25151_, _25148_);
  and (_25153_, _25152_, _01870_);
  nand (_25154_, _03716_, _02687_);
  and (_25155_, _25102_, _01869_);
  and (_25156_, _25155_, _25154_);
  or (_25157_, _25156_, _25153_);
  and (_25158_, _25157_, _02166_);
  or (_25160_, _10816_, _09096_);
  and (_25161_, _25102_, _02079_);
  and (_25162_, _25161_, _25160_);
  or (_25163_, _25162_, _25158_);
  and (_25164_, _25163_, _02912_);
  or (_25165_, _10822_, _09096_);
  and (_25166_, _25102_, _02167_);
  and (_25167_, _25166_, _25165_);
  or (_25168_, _25167_, _25164_);
  and (_25169_, _25168_, _02176_);
  or (_25171_, _10692_, _09096_);
  and (_25172_, _25102_, _02072_);
  and (_25173_, _25172_, _25171_);
  or (_25174_, _25173_, _25169_);
  and (_25175_, _25174_, _02907_);
  or (_25176_, _25093_, _04058_);
  and (_25177_, _25109_, _02177_);
  and (_25178_, _25177_, _25176_);
  or (_25179_, _25178_, _25175_);
  and (_25180_, _25179_, _02174_);
  or (_25182_, _25108_, _04058_);
  and (_25183_, _25102_, _02173_);
  and (_25184_, _25183_, _25182_);
  or (_25185_, _25184_, _02201_);
  or (_25186_, _25154_, _04058_);
  and (_25187_, _25102_, _02071_);
  and (_25188_, _25187_, _25186_);
  or (_25189_, _25188_, _25185_);
  or (_25190_, _25189_, _25180_);
  or (_25191_, _25106_, _02303_);
  and (_25193_, _25191_, _01887_);
  and (_25194_, _25193_, _25190_);
  and (_25195_, _25125_, _01860_);
  or (_25196_, _25195_, _01537_);
  or (_25197_, _25196_, _25194_);
  or (_25198_, _25093_, _01538_);
  or (_25199_, _25198_, _25103_);
  and (_25200_, _25199_, _38087_);
  and (_25201_, _25200_, _25197_);
  or (_25202_, _25201_, _25092_);
  and (_40292_, _25202_, _37580_);
  and (_25204_, _38088_, \oc8051_golden_model_1.SCON [2]);
  and (_25205_, _09096_, \oc8051_golden_model_1.SCON [2]);
  and (_25206_, _11020_, _03716_);
  or (_25207_, _25206_, _25205_);
  and (_25208_, _25207_, _02167_);
  nor (_25209_, _09096_, _03455_);
  or (_25210_, _25209_, _25205_);
  or (_25211_, _25210_, _05249_);
  or (_25212_, _25210_, _02840_);
  nor (_25214_, _10905_, _09096_);
  or (_25215_, _25214_, _25205_);
  or (_25216_, _25215_, _02814_);
  and (_25217_, _03716_, \oc8051_golden_model_1.ACC [2]);
  or (_25218_, _25217_, _25205_);
  and (_25219_, _25218_, _02817_);
  and (_25220_, _02818_, \oc8051_golden_model_1.SCON [2]);
  or (_25221_, _25220_, _02001_);
  or (_25222_, _25221_, _25219_);
  and (_25223_, _25222_, _02024_);
  and (_25225_, _25223_, _25216_);
  and (_25226_, _09104_, \oc8051_golden_model_1.SCON [2]);
  and (_25227_, _10909_, _04331_);
  or (_25228_, _25227_, _25226_);
  and (_25229_, _25228_, _02007_);
  or (_25230_, _25229_, _01999_);
  or (_25231_, _25230_, _25225_);
  and (_25232_, _25231_, _25212_);
  or (_25233_, _25232_, _02006_);
  or (_25234_, _25218_, _02021_);
  and (_25236_, _25234_, _02025_);
  and (_25237_, _25236_, _25233_);
  and (_25238_, _10894_, _04331_);
  or (_25239_, _25238_, _25226_);
  and (_25240_, _25239_, _01997_);
  or (_25241_, _25240_, _01991_);
  or (_25242_, _25241_, _25237_);
  and (_25243_, _25227_, _10924_);
  or (_25244_, _25226_, _02861_);
  or (_25245_, _25244_, _25243_);
  and (_25247_, _25245_, _02408_);
  and (_25248_, _25247_, _25242_);
  nor (_25249_, _10942_, _09104_);
  or (_25250_, _25249_, _25226_);
  and (_25251_, _25250_, _01875_);
  or (_25252_, _25251_, _05994_);
  or (_25253_, _25252_, _25248_);
  and (_25254_, _25253_, _25211_);
  or (_25255_, _25254_, _02528_);
  and (_25256_, _05043_, _03716_);
  or (_25258_, _25205_, _02888_);
  or (_25259_, _25258_, _25256_);
  and (_25260_, _25259_, _02043_);
  and (_25261_, _25260_, _25255_);
  nor (_25262_, _11000_, _09096_);
  or (_25263_, _25262_, _25205_);
  and (_25264_, _25263_, _01602_);
  or (_25265_, _25264_, _01869_);
  or (_25266_, _25265_, _25261_);
  and (_25267_, _03716_, _04724_);
  or (_25269_, _25267_, _25205_);
  or (_25270_, _25269_, _01870_);
  and (_25271_, _25270_, _25266_);
  or (_25272_, _25271_, _02079_);
  and (_25273_, _11014_, _03716_);
  or (_25274_, _25205_, _02166_);
  or (_25275_, _25274_, _25273_);
  and (_25276_, _25275_, _02912_);
  and (_25277_, _25276_, _25272_);
  or (_25278_, _25277_, _25208_);
  and (_25279_, _25278_, _02176_);
  or (_25280_, _25205_, _04156_);
  and (_25281_, _25269_, _02072_);
  and (_25282_, _25281_, _25280_);
  or (_25283_, _25282_, _25279_);
  and (_25284_, _25283_, _02907_);
  and (_25285_, _25218_, _02177_);
  and (_25286_, _25285_, _25280_);
  or (_25287_, _25286_, _02071_);
  or (_25288_, _25287_, _25284_);
  nor (_25290_, _11013_, _09096_);
  or (_25291_, _25205_, _04788_);
  or (_25292_, _25291_, _25290_);
  and (_25293_, _25292_, _04793_);
  and (_25294_, _25293_, _25288_);
  nor (_25295_, _11019_, _09096_);
  or (_25296_, _25295_, _25205_);
  and (_25297_, _25296_, _02173_);
  or (_25298_, _25297_, _02201_);
  or (_25299_, _25298_, _25294_);
  or (_25301_, _25215_, _02303_);
  and (_25302_, _25301_, _01887_);
  and (_25303_, _25302_, _25299_);
  and (_25304_, _25239_, _01860_);
  or (_25305_, _25304_, _01537_);
  or (_25306_, _25305_, _25303_);
  and (_25307_, _11072_, _03716_);
  or (_25308_, _25205_, _01538_);
  or (_25309_, _25308_, _25307_);
  and (_25310_, _25309_, _38087_);
  and (_25312_, _25310_, _25306_);
  or (_25313_, _25312_, _25204_);
  and (_40293_, _25313_, _37580_);
  and (_25314_, _38088_, \oc8051_golden_model_1.SCON [3]);
  and (_25315_, _09096_, \oc8051_golden_model_1.SCON [3]);
  and (_25316_, _11094_, _03716_);
  or (_25317_, _25316_, _25315_);
  and (_25318_, _25317_, _02167_);
  nor (_25319_, _09096_, _03268_);
  or (_25320_, _25319_, _25315_);
  or (_25322_, _25320_, _05249_);
  nor (_25323_, _11101_, _09096_);
  or (_25324_, _25323_, _25315_);
  or (_25325_, _25324_, _02814_);
  and (_25326_, _03716_, \oc8051_golden_model_1.ACC [3]);
  or (_25327_, _25326_, _25315_);
  and (_25328_, _25327_, _02817_);
  and (_25329_, _02818_, \oc8051_golden_model_1.SCON [3]);
  or (_25330_, _25329_, _02001_);
  or (_25331_, _25330_, _25328_);
  and (_25333_, _25331_, _02024_);
  and (_25334_, _25333_, _25325_);
  and (_25335_, _09104_, \oc8051_golden_model_1.SCON [3]);
  and (_25336_, _11098_, _04331_);
  or (_25337_, _25336_, _25335_);
  and (_25338_, _25337_, _02007_);
  or (_25339_, _25338_, _01999_);
  or (_25340_, _25339_, _25334_);
  or (_25341_, _25320_, _02840_);
  and (_25342_, _25341_, _25340_);
  or (_25344_, _25342_, _02006_);
  or (_25345_, _25327_, _02021_);
  and (_25346_, _25345_, _02025_);
  and (_25347_, _25346_, _25344_);
  and (_25348_, _11096_, _04331_);
  or (_25349_, _25348_, _25335_);
  and (_25350_, _25349_, _01997_);
  or (_25351_, _25350_, _01991_);
  or (_25352_, _25351_, _25347_);
  or (_25353_, _25335_, _11127_);
  and (_25355_, _25353_, _25337_);
  or (_25356_, _25355_, _02861_);
  and (_25357_, _25356_, _02408_);
  and (_25358_, _25357_, _25352_);
  nor (_25359_, _11145_, _09104_);
  or (_25360_, _25359_, _25335_);
  and (_25361_, _25360_, _01875_);
  or (_25362_, _25361_, _05994_);
  or (_25363_, _25362_, _25358_);
  and (_25364_, _25363_, _25322_);
  or (_25366_, _25364_, _02528_);
  and (_25367_, _04998_, _03716_);
  or (_25368_, _25315_, _02888_);
  or (_25369_, _25368_, _25367_);
  and (_25370_, _25369_, _02043_);
  and (_25371_, _25370_, _25366_);
  nor (_25372_, _11206_, _09096_);
  or (_25373_, _25372_, _25315_);
  and (_25374_, _25373_, _01602_);
  or (_25375_, _25374_, _01869_);
  or (_25377_, _25375_, _25371_);
  and (_25378_, _03716_, _04678_);
  or (_25379_, _25378_, _25315_);
  or (_25380_, _25379_, _01870_);
  and (_25381_, _25380_, _25377_);
  or (_25382_, _25381_, _02079_);
  and (_25383_, _11222_, _03716_);
  or (_25384_, _25315_, _02166_);
  or (_25385_, _25384_, _25383_);
  and (_25386_, _25385_, _02912_);
  and (_25388_, _25386_, _25382_);
  or (_25389_, _25388_, _25318_);
  and (_25390_, _25389_, _02176_);
  or (_25391_, _25315_, _04014_);
  and (_25392_, _25379_, _02072_);
  and (_25393_, _25392_, _25391_);
  or (_25394_, _25393_, _25390_);
  and (_25395_, _25394_, _02907_);
  and (_25396_, _25327_, _02177_);
  and (_25397_, _25396_, _25391_);
  or (_25399_, _25397_, _02071_);
  or (_25400_, _25399_, _25395_);
  nor (_25401_, _11220_, _09096_);
  or (_25402_, _25315_, _04788_);
  or (_25403_, _25402_, _25401_);
  and (_25404_, _25403_, _04793_);
  and (_25405_, _25404_, _25400_);
  nor (_25406_, _11093_, _09096_);
  or (_25407_, _25406_, _25315_);
  and (_25408_, _25407_, _02173_);
  or (_25410_, _25408_, _02201_);
  or (_25411_, _25410_, _25405_);
  or (_25412_, _25324_, _02303_);
  and (_25413_, _25412_, _01887_);
  and (_25414_, _25413_, _25411_);
  and (_25415_, _25349_, _01860_);
  or (_25416_, _25415_, _01537_);
  or (_25417_, _25416_, _25414_);
  and (_25418_, _11273_, _03716_);
  or (_25419_, _25315_, _01538_);
  or (_25421_, _25419_, _25418_);
  and (_25422_, _25421_, _38087_);
  and (_25423_, _25422_, _25417_);
  or (_25424_, _25423_, _25314_);
  and (_40294_, _25424_, _37580_);
  and (_25425_, _38088_, \oc8051_golden_model_1.SCON [4]);
  and (_25426_, _09096_, \oc8051_golden_model_1.SCON [4]);
  and (_25427_, _11431_, _03716_);
  or (_25428_, _25427_, _25426_);
  and (_25429_, _25428_, _02167_);
  nor (_25430_, _04211_, _09096_);
  or (_25431_, _25430_, _25426_);
  or (_25432_, _25431_, _05249_);
  and (_25433_, _09104_, \oc8051_golden_model_1.SCON [4]);
  and (_25434_, _11301_, _04331_);
  or (_25435_, _25434_, _25433_);
  and (_25436_, _25435_, _01997_);
  nor (_25437_, _11317_, _09096_);
  or (_25438_, _25437_, _25426_);
  or (_25439_, _25438_, _02814_);
  and (_25441_, _03716_, \oc8051_golden_model_1.ACC [4]);
  or (_25442_, _25441_, _25426_);
  and (_25443_, _25442_, _02817_);
  and (_25444_, _02818_, \oc8051_golden_model_1.SCON [4]);
  or (_25445_, _25444_, _02001_);
  or (_25446_, _25445_, _25443_);
  and (_25447_, _25446_, _02024_);
  and (_25448_, _25447_, _25439_);
  and (_25449_, _11303_, _04331_);
  or (_25450_, _25449_, _25433_);
  and (_25452_, _25450_, _02007_);
  or (_25453_, _25452_, _01999_);
  or (_25454_, _25453_, _25448_);
  or (_25455_, _25431_, _02840_);
  and (_25456_, _25455_, _25454_);
  or (_25457_, _25456_, _02006_);
  or (_25458_, _25442_, _02021_);
  and (_25459_, _25458_, _02025_);
  and (_25460_, _25459_, _25457_);
  or (_25461_, _25460_, _25436_);
  and (_25463_, _25461_, _02861_);
  or (_25464_, _25433_, _11334_);
  and (_25465_, _25464_, _01991_);
  and (_25466_, _25465_, _25450_);
  or (_25467_, _25466_, _25463_);
  and (_25468_, _25467_, _02408_);
  nor (_25469_, _11299_, _09104_);
  or (_25470_, _25469_, _25433_);
  and (_25471_, _25470_, _01875_);
  or (_25472_, _25471_, _05994_);
  or (_25474_, _25472_, _25468_);
  and (_25475_, _25474_, _25432_);
  or (_25476_, _25475_, _02528_);
  and (_25477_, _05135_, _03716_);
  or (_25478_, _25426_, _02888_);
  or (_25479_, _25478_, _25477_);
  and (_25480_, _25479_, _02043_);
  and (_25481_, _25480_, _25476_);
  nor (_25482_, _11411_, _09096_);
  or (_25483_, _25482_, _25426_);
  and (_25485_, _25483_, _01602_);
  or (_25486_, _25485_, _01869_);
  or (_25487_, _25486_, _25481_);
  and (_25488_, _04694_, _03716_);
  or (_25489_, _25488_, _25426_);
  or (_25490_, _25489_, _01870_);
  and (_25491_, _25490_, _25487_);
  or (_25492_, _25491_, _02079_);
  and (_25493_, _11425_, _03716_);
  or (_25494_, _25426_, _02166_);
  or (_25496_, _25494_, _25493_);
  and (_25497_, _25496_, _02912_);
  and (_25498_, _25497_, _25492_);
  or (_25499_, _25498_, _25429_);
  and (_25500_, _25499_, _02176_);
  or (_25501_, _25426_, _04258_);
  and (_25502_, _25489_, _02072_);
  and (_25503_, _25502_, _25501_);
  or (_25504_, _25503_, _25500_);
  and (_25505_, _25504_, _02907_);
  and (_25507_, _25442_, _02177_);
  and (_25508_, _25507_, _25501_);
  or (_25509_, _25508_, _02071_);
  or (_25510_, _25509_, _25505_);
  nor (_25511_, _11424_, _09096_);
  or (_25512_, _25426_, _04788_);
  or (_25513_, _25512_, _25511_);
  and (_25514_, _25513_, _04793_);
  and (_25515_, _25514_, _25510_);
  nor (_25516_, _11430_, _09096_);
  or (_25518_, _25516_, _25426_);
  and (_25519_, _25518_, _02173_);
  or (_25520_, _25519_, _02201_);
  or (_25521_, _25520_, _25515_);
  or (_25522_, _25438_, _02303_);
  and (_25523_, _25522_, _01887_);
  and (_25524_, _25523_, _25521_);
  and (_25525_, _25435_, _01860_);
  or (_25526_, _25525_, _01537_);
  or (_25527_, _25526_, _25524_);
  and (_25529_, _11487_, _03716_);
  or (_25530_, _25426_, _01538_);
  or (_25531_, _25530_, _25529_);
  and (_25532_, _25531_, _38087_);
  and (_25533_, _25532_, _25527_);
  or (_25534_, _25533_, _25425_);
  and (_40295_, _25534_, _37580_);
  and (_25535_, _38088_, \oc8051_golden_model_1.SCON [5]);
  and (_25536_, _09096_, \oc8051_golden_model_1.SCON [5]);
  and (_25537_, _11635_, _03716_);
  or (_25539_, _25537_, _25536_);
  and (_25540_, _25539_, _02167_);
  nor (_25541_, _11525_, _09096_);
  or (_25542_, _25541_, _25536_);
  or (_25543_, _25542_, _02814_);
  and (_25544_, _03716_, \oc8051_golden_model_1.ACC [5]);
  or (_25545_, _25544_, _25536_);
  and (_25546_, _25545_, _02817_);
  and (_25547_, _02818_, \oc8051_golden_model_1.SCON [5]);
  or (_25548_, _25547_, _02001_);
  or (_25550_, _25548_, _25546_);
  and (_25551_, _25550_, _02024_);
  and (_25552_, _25551_, _25543_);
  and (_25553_, _09104_, \oc8051_golden_model_1.SCON [5]);
  and (_25554_, _11510_, _04331_);
  or (_25555_, _25554_, _25553_);
  and (_25556_, _25555_, _02007_);
  or (_25557_, _25556_, _01999_);
  or (_25558_, _25557_, _25552_);
  nor (_25559_, _03916_, _09096_);
  or (_25561_, _25559_, _25536_);
  or (_25562_, _25561_, _02840_);
  and (_25563_, _25562_, _25558_);
  or (_25564_, _25563_, _02006_);
  or (_25565_, _25545_, _02021_);
  and (_25566_, _25565_, _02025_);
  and (_25567_, _25566_, _25564_);
  and (_25568_, _11508_, _04331_);
  or (_25569_, _25568_, _25553_);
  and (_25570_, _25569_, _01997_);
  or (_25572_, _25570_, _01991_);
  or (_25573_, _25572_, _25567_);
  or (_25574_, _25553_, _11542_);
  and (_25575_, _25574_, _25555_);
  or (_25576_, _25575_, _02861_);
  and (_25577_, _25576_, _02408_);
  and (_25578_, _25577_, _25573_);
  nor (_25579_, _11506_, _09104_);
  or (_25580_, _25579_, _25553_);
  and (_25581_, _25580_, _01875_);
  or (_25583_, _25581_, _05994_);
  or (_25584_, _25583_, _25578_);
  or (_25585_, _25561_, _05249_);
  and (_25586_, _25585_, _25584_);
  or (_25587_, _25586_, _02528_);
  and (_25588_, _05090_, _03716_);
  or (_25589_, _25536_, _02888_);
  or (_25590_, _25589_, _25588_);
  and (_25591_, _25590_, _02043_);
  and (_25592_, _25591_, _25587_);
  nor (_25594_, _11615_, _09096_);
  or (_25595_, _25594_, _25536_);
  and (_25596_, _25595_, _01602_);
  or (_25597_, _25596_, _01869_);
  or (_25598_, _25597_, _25592_);
  and (_25599_, _04672_, _03716_);
  or (_25600_, _25599_, _25536_);
  or (_25601_, _25600_, _01870_);
  and (_25602_, _25601_, _25598_);
  or (_25603_, _25602_, _02079_);
  and (_25604_, _11629_, _03716_);
  or (_25605_, _25536_, _02166_);
  or (_25606_, _25605_, _25604_);
  and (_25607_, _25606_, _02912_);
  and (_25608_, _25607_, _25603_);
  or (_25609_, _25608_, _25540_);
  and (_25610_, _25609_, _02176_);
  or (_25611_, _25536_, _03965_);
  and (_25612_, _25600_, _02072_);
  and (_25613_, _25612_, _25611_);
  or (_25615_, _25613_, _25610_);
  and (_25616_, _25615_, _02907_);
  and (_25617_, _25545_, _02177_);
  and (_25618_, _25617_, _25611_);
  or (_25619_, _25618_, _02071_);
  or (_25620_, _25619_, _25616_);
  nor (_25621_, _11628_, _09096_);
  or (_25622_, _25536_, _04788_);
  or (_25623_, _25622_, _25621_);
  and (_25624_, _25623_, _04793_);
  and (_25626_, _25624_, _25620_);
  nor (_25627_, _11634_, _09096_);
  or (_25628_, _25627_, _25536_);
  and (_25629_, _25628_, _02173_);
  or (_25630_, _25629_, _02201_);
  or (_25631_, _25630_, _25626_);
  or (_25632_, _25542_, _02303_);
  and (_25633_, _25632_, _01887_);
  and (_25634_, _25633_, _25631_);
  and (_25635_, _25569_, _01860_);
  or (_25637_, _25635_, _01537_);
  or (_25638_, _25637_, _25634_);
  and (_25639_, _11685_, _03716_);
  or (_25640_, _25536_, _01538_);
  or (_25641_, _25640_, _25639_);
  and (_25642_, _25641_, _38087_);
  and (_25643_, _25642_, _25638_);
  or (_25644_, _25643_, _25535_);
  and (_40296_, _25644_, _37580_);
  and (_25645_, _38088_, \oc8051_golden_model_1.SCON [6]);
  and (_25647_, _09096_, \oc8051_golden_model_1.SCON [6]);
  and (_25648_, _11709_, _03716_);
  or (_25649_, _25648_, _25647_);
  and (_25650_, _25649_, _02167_);
  nor (_25651_, _11730_, _09096_);
  or (_25652_, _25651_, _25647_);
  or (_25653_, _25652_, _02814_);
  and (_25654_, _03716_, \oc8051_golden_model_1.ACC [6]);
  or (_25655_, _25654_, _25647_);
  and (_25656_, _25655_, _02817_);
  and (_25658_, _02818_, \oc8051_golden_model_1.SCON [6]);
  or (_25659_, _25658_, _02001_);
  or (_25660_, _25659_, _25656_);
  and (_25661_, _25660_, _02024_);
  and (_25662_, _25661_, _25653_);
  and (_25663_, _09104_, \oc8051_golden_model_1.SCON [6]);
  and (_25664_, _11717_, _04331_);
  or (_25665_, _25664_, _25663_);
  and (_25666_, _25665_, _02007_);
  or (_25667_, _25666_, _01999_);
  or (_25669_, _25667_, _25662_);
  nor (_25670_, _03808_, _09096_);
  or (_25671_, _25670_, _25647_);
  or (_25672_, _25671_, _02840_);
  and (_25673_, _25672_, _25669_);
  or (_25674_, _25673_, _02006_);
  or (_25675_, _25655_, _02021_);
  and (_25676_, _25675_, _02025_);
  and (_25677_, _25676_, _25674_);
  and (_25678_, _11715_, _04331_);
  or (_25680_, _25678_, _25663_);
  and (_25681_, _25680_, _01997_);
  or (_25682_, _25681_, _01991_);
  or (_25683_, _25682_, _25677_);
  or (_25684_, _25663_, _11747_);
  and (_25685_, _25684_, _25665_);
  or (_25686_, _25685_, _02861_);
  and (_25687_, _25686_, _02408_);
  and (_25688_, _25687_, _25683_);
  nor (_25689_, _11713_, _09104_);
  or (_25690_, _25689_, _25663_);
  and (_25691_, _25690_, _01875_);
  or (_25692_, _25691_, _05994_);
  or (_25693_, _25692_, _25688_);
  or (_25694_, _25671_, _05249_);
  and (_25695_, _25694_, _25693_);
  or (_25696_, _25695_, _02528_);
  and (_25697_, _04861_, _03716_);
  or (_25698_, _25647_, _02888_);
  or (_25699_, _25698_, _25697_);
  and (_25701_, _25699_, _02043_);
  and (_25702_, _25701_, _25696_);
  nor (_25703_, _11820_, _09096_);
  or (_25704_, _25703_, _25647_);
  and (_25705_, _25704_, _01602_);
  or (_25706_, _25705_, _01869_);
  or (_25707_, _25706_, _25702_);
  and (_25708_, _09920_, _03716_);
  or (_25709_, _25708_, _25647_);
  or (_25710_, _25709_, _01870_);
  and (_25712_, _25710_, _25707_);
  or (_25713_, _25712_, _02079_);
  and (_25714_, _11835_, _03716_);
  or (_25715_, _25647_, _02166_);
  or (_25716_, _25715_, _25714_);
  and (_25717_, _25716_, _02912_);
  and (_25718_, _25717_, _25713_);
  or (_25719_, _25718_, _25650_);
  and (_25720_, _25719_, _02176_);
  or (_25721_, _25647_, _03863_);
  and (_25723_, _25709_, _02072_);
  and (_25724_, _25723_, _25721_);
  or (_25725_, _25724_, _25720_);
  and (_25726_, _25725_, _02907_);
  and (_25727_, _25655_, _02177_);
  and (_25728_, _25727_, _25721_);
  or (_25729_, _25728_, _02071_);
  or (_25730_, _25729_, _25726_);
  nor (_25731_, _11833_, _09096_);
  or (_25732_, _25647_, _04788_);
  or (_25734_, _25732_, _25731_);
  and (_25735_, _25734_, _04793_);
  and (_25736_, _25735_, _25730_);
  nor (_25737_, _11708_, _09096_);
  or (_25738_, _25737_, _25647_);
  and (_25739_, _25738_, _02173_);
  or (_25740_, _25739_, _02201_);
  or (_25741_, _25740_, _25736_);
  or (_25742_, _25652_, _02303_);
  and (_25743_, _25742_, _01887_);
  and (_25745_, _25743_, _25741_);
  and (_25746_, _25680_, _01860_);
  or (_25747_, _25746_, _01537_);
  or (_25748_, _25747_, _25745_);
  and (_25749_, _11887_, _03716_);
  or (_25750_, _25647_, _01538_);
  or (_25751_, _25750_, _25749_);
  and (_25752_, _25751_, _38087_);
  and (_25753_, _25752_, _25748_);
  or (_25754_, _25753_, _25645_);
  and (_40297_, _25754_, _37580_);
  nor (_25756_, _03745_, _01864_);
  nor (_25757_, _04106_, _09213_);
  or (_25758_, _25757_, _25756_);
  or (_25759_, _25758_, _02814_);
  and (_25760_, _03745_, \oc8051_golden_model_1.ACC [0]);
  or (_25761_, _25760_, _25756_);
  and (_25762_, _25761_, _02817_);
  nor (_25763_, _02817_, _01864_);
  or (_25764_, _25763_, _02001_);
  or (_25766_, _25764_, _25762_);
  and (_25767_, _25766_, _02840_);
  and (_25768_, _25767_, _25759_);
  or (_25769_, _25768_, _02481_);
  or (_25770_, _25761_, _02021_);
  and (_25771_, _25770_, _01880_);
  and (_25772_, _25771_, _25769_);
  nand (_25773_, _05249_, _03051_);
  or (_25774_, _25773_, _25772_);
  and (_25775_, _03853_, _03028_);
  or (_25777_, _25756_, _05249_);
  or (_25778_, _25777_, _25775_);
  and (_25779_, _25778_, _25774_);
  or (_25780_, _25779_, _02528_);
  or (_25781_, _25756_, _02888_);
  and (_25782_, _04952_, _03745_);
  or (_25783_, _25782_, _25781_);
  and (_25784_, _25783_, _25780_);
  or (_25785_, _25784_, _01602_);
  nor (_25786_, _10600_, _09213_);
  or (_25787_, _25756_, _02043_);
  or (_25788_, _25787_, _25786_);
  and (_25789_, _25788_, _01870_);
  and (_25790_, _25789_, _25785_);
  and (_25791_, _03745_, _04562_);
  or (_25792_, _25791_, _25756_);
  and (_25793_, _25792_, _01869_);
  or (_25794_, _25793_, _02079_);
  or (_25795_, _25794_, _25790_);
  and (_25796_, _10614_, _03745_);
  or (_25798_, _25796_, _25756_);
  or (_25799_, _25798_, _02166_);
  and (_25800_, _25799_, _25795_);
  or (_25801_, _25800_, _02167_);
  and (_25802_, _10620_, _03853_);
  or (_25803_, _25756_, _02912_);
  or (_25804_, _25803_, _25802_);
  and (_25805_, _25804_, _02176_);
  and (_25806_, _25805_, _25801_);
  nand (_25807_, _25792_, _02072_);
  nor (_25809_, _25807_, _25757_);
  or (_25810_, _25809_, _25806_);
  and (_25811_, _25810_, _02907_);
  or (_25812_, _25756_, _04106_);
  and (_25813_, _25761_, _02177_);
  and (_25814_, _25813_, _25812_);
  or (_25815_, _25814_, _02071_);
  or (_25816_, _25815_, _25811_);
  nor (_25817_, _10613_, _09213_);
  or (_25818_, _25756_, _04788_);
  or (_25820_, _25818_, _25817_);
  and (_25821_, _25820_, _04793_);
  and (_25822_, _25821_, _25816_);
  nor (_25823_, _10619_, _09213_);
  or (_25824_, _25823_, _25756_);
  and (_25825_, _25824_, _02173_);
  or (_25826_, _25825_, _15577_);
  or (_25827_, _25826_, _25822_);
  or (_25828_, _25758_, _02743_);
  and (_25829_, _25828_, _38087_);
  and (_25831_, _25829_, _25827_);
  nor (_25832_, _38087_, _01864_);
  or (_25833_, _25832_, rst);
  or (_40299_, _25833_, _25831_);
  nor (_25834_, _03745_, _01862_);
  and (_25835_, _10698_, _03853_);
  or (_25836_, _25835_, _25834_);
  and (_25837_, _25836_, _01537_);
  or (_25838_, _22755_, _01862_);
  not (_25839_, _25835_);
  or (_25841_, _03745_, \oc8051_golden_model_1.SP [1]);
  and (_25842_, _25841_, _25839_);
  or (_25843_, _25842_, _02814_);
  and (_25844_, _03745_, \oc8051_golden_model_1.ACC [1]);
  or (_25845_, _25844_, _25834_);
  or (_25846_, _25845_, _02818_);
  nor (_25847_, _09224_, \oc8051_golden_model_1.SP [1]);
  and (_25848_, _01562_, \oc8051_golden_model_1.SP [1]);
  or (_25849_, _25848_, _25847_);
  and (_25850_, _25849_, _25846_);
  or (_25852_, _25850_, _02001_);
  and (_25853_, _25852_, _01558_);
  and (_25854_, _25853_, _25843_);
  nor (_25855_, _01558_, \oc8051_golden_model_1.SP [1]);
  or (_25856_, _25855_, _01999_);
  or (_25857_, _25856_, _25854_);
  nand (_25858_, _01999_, _01867_);
  and (_25859_, _25858_, _25857_);
  or (_25860_, _25859_, _02006_);
  or (_25861_, _25845_, _02021_);
  and (_25863_, _25861_, _01880_);
  and (_25864_, _25863_, _25860_);
  or (_25865_, _03132_, _01879_);
  or (_25866_, _25865_, _25864_);
  nand (_25867_, _03132_, \oc8051_golden_model_1.SP [1]);
  and (_25868_, _25867_, _05249_);
  and (_25869_, _25868_, _25866_);
  nand (_25870_, _03853_, _02811_);
  and (_25871_, _25841_, _05994_);
  and (_25872_, _25871_, _25870_);
  or (_25874_, _25872_, _02528_);
  or (_25875_, _25874_, _25869_);
  or (_25876_, _25834_, _02888_);
  and (_25877_, _04907_, _03745_);
  or (_25878_, _25877_, _25876_);
  and (_25879_, _25878_, _02043_);
  and (_25880_, _25879_, _25875_);
  and (_25881_, _25841_, _01602_);
  nand (_25882_, _10802_, _03853_);
  and (_25883_, _25882_, _25881_);
  or (_25885_, _25883_, _25880_);
  and (_25886_, _25885_, _01870_);
  and (_25887_, _25841_, _01869_);
  nand (_25888_, _03853_, _02687_);
  and (_25889_, _25888_, _25887_);
  or (_25890_, _25889_, _01638_);
  or (_25891_, _25890_, _25886_);
  nand (_25892_, _01638_, \oc8051_golden_model_1.SP [1]);
  and (_25893_, _25892_, _02166_);
  and (_25894_, _25893_, _25891_);
  or (_25896_, _10816_, _09213_);
  and (_25897_, _25841_, _02079_);
  and (_25898_, _25897_, _25896_);
  or (_25899_, _25898_, _25894_);
  and (_25900_, _25899_, _02912_);
  or (_25901_, _10822_, _09213_);
  and (_25902_, _25841_, _02167_);
  and (_25903_, _25902_, _25901_);
  or (_25904_, _25903_, _25900_);
  and (_25905_, _25904_, _02176_);
  or (_25907_, _10692_, _09213_);
  and (_25908_, _25841_, _02072_);
  and (_25909_, _25908_, _25907_);
  or (_25910_, _25909_, _25905_);
  and (_25911_, _25910_, _09292_);
  and (_25912_, _01632_, _01862_);
  or (_25913_, _25834_, _04058_);
  and (_25914_, _25845_, _02177_);
  and (_25915_, _25914_, _25913_);
  or (_25916_, _25915_, _25912_);
  or (_25918_, _25916_, _25911_);
  and (_25919_, _25918_, _02174_);
  nand (_25920_, _10821_, _03853_);
  and (_25921_, _25841_, _02173_);
  and (_25922_, _25921_, _25920_);
  or (_25923_, _25888_, _04058_);
  and (_25924_, _25841_, _02071_);
  nand (_25925_, _25924_, _25923_);
  nand (_25926_, _25925_, _22755_);
  or (_25927_, _25926_, _25922_);
  or (_25929_, _25927_, _25919_);
  and (_25930_, _25929_, _25838_);
  or (_25931_, _25930_, _01888_);
  nor (_25932_, _02703_, _02201_);
  and (_25933_, _25932_, _25931_);
  and (_25934_, _25842_, _02201_);
  or (_25935_, _25934_, _03370_);
  or (_25936_, _25935_, _25933_);
  or (_25937_, _02942_, _01862_);
  and (_25938_, _25937_, _01538_);
  and (_25939_, _25938_, _25936_);
  or (_25940_, _25939_, _25837_);
  and (_25941_, _25940_, _38087_);
  nor (_25942_, _38087_, _01862_);
  or (_25943_, _25942_, rst);
  or (_40300_, _25943_, _25941_);
  nor (_25944_, _38087_, _02346_);
  or (_25945_, _25944_, rst);
  nor (_25946_, _03745_, _02346_);
  and (_25947_, _11020_, _03853_);
  or (_25949_, _25947_, _25946_);
  and (_25950_, _25949_, _02167_);
  nand (_25951_, _10678_, _01638_);
  nor (_25952_, _09213_, _03455_);
  or (_25953_, _25946_, _05249_);
  or (_25954_, _25953_, _25952_);
  nor (_25955_, _10905_, _09213_);
  or (_25956_, _25955_, _25946_);
  or (_25957_, _25956_, _02814_);
  and (_25958_, _03745_, \oc8051_golden_model_1.ACC [2]);
  or (_25960_, _25958_, _25946_);
  and (_25961_, _25960_, _02817_);
  and (_25962_, _09224_, \oc8051_golden_model_1.SP [2]);
  nor (_25963_, _10678_, _01562_);
  or (_25964_, _25963_, _02001_);
  or (_25965_, _25964_, _25962_);
  or (_25966_, _25965_, _25961_);
  and (_25967_, _25966_, _01558_);
  and (_25968_, _25967_, _25957_);
  nor (_25969_, _10678_, _01558_);
  or (_25971_, _25969_, _01999_);
  or (_25972_, _25971_, _25968_);
  nand (_25973_, _04412_, _01999_);
  and (_25974_, _25973_, _25972_);
  or (_25975_, _25974_, _02006_);
  or (_25976_, _25960_, _02021_);
  and (_25977_, _25976_, _01880_);
  and (_25978_, _25977_, _25975_);
  or (_25979_, _03395_, _03131_);
  or (_25980_, _25979_, _25978_);
  nor (_25982_, _03548_, _01565_);
  nor (_25983_, _25982_, _01604_);
  and (_25984_, _25983_, _25980_);
  nand (_25985_, _03548_, _01604_);
  nand (_25986_, _25985_, _05249_);
  or (_25987_, _25986_, _25984_);
  and (_25988_, _25987_, _25954_);
  or (_25989_, _25988_, _02528_);
  or (_25990_, _25946_, _02888_);
  and (_25991_, _05043_, _03745_);
  or (_25993_, _25991_, _25990_);
  and (_25994_, _25993_, _02043_);
  and (_25995_, _25994_, _25989_);
  not (_25996_, _03745_);
  nor (_25997_, _11000_, _25996_);
  or (_25998_, _25997_, _25946_);
  and (_25999_, _25998_, _01602_);
  or (_26000_, _25999_, _01869_);
  or (_26001_, _26000_, _25995_);
  and (_26002_, _03745_, _04724_);
  or (_26004_, _26002_, _25946_);
  or (_26005_, _26004_, _01870_);
  and (_26006_, _26005_, _26001_);
  or (_26007_, _26006_, _01638_);
  and (_26008_, _26007_, _25951_);
  or (_26009_, _26008_, _02079_);
  and (_26010_, _11014_, _03853_);
  or (_26011_, _25946_, _02166_);
  or (_26012_, _26011_, _26010_);
  and (_26013_, _26012_, _02912_);
  and (_26015_, _26013_, _26009_);
  or (_26016_, _26015_, _25950_);
  and (_26017_, _26016_, _02176_);
  or (_26018_, _25946_, _04156_);
  and (_26019_, _26004_, _02072_);
  and (_26020_, _26019_, _26018_);
  or (_26021_, _26020_, _26017_);
  and (_26022_, _26021_, _09292_);
  and (_26023_, _25960_, _02177_);
  and (_26024_, _26023_, _26018_);
  and (_26026_, _03548_, _01632_);
  or (_26027_, _26026_, _02071_);
  or (_26028_, _26027_, _26024_);
  or (_26029_, _26028_, _26022_);
  nor (_26030_, _11013_, _25996_);
  or (_26031_, _26030_, _25946_);
  or (_26032_, _26031_, _04788_);
  and (_26033_, _26032_, _26029_);
  or (_26034_, _26033_, _02173_);
  nor (_26035_, _11019_, _09213_);
  or (_26037_, _25946_, _04793_);
  or (_26038_, _26037_, _26035_);
  and (_26039_, _26038_, _09305_);
  and (_26040_, _26039_, _26034_);
  and (_26041_, _10678_, _02185_);
  or (_26042_, _26041_, _01636_);
  or (_26043_, _26042_, _26040_);
  nand (_26044_, _10678_, _01636_);
  and (_26045_, _26044_, _01889_);
  and (_26046_, _26045_, _26043_);
  and (_26048_, _10678_, _01888_);
  or (_26049_, _26048_, _02201_);
  or (_26050_, _26049_, _26046_);
  or (_26051_, _25956_, _02303_);
  and (_26052_, _26051_, _02942_);
  and (_26053_, _26052_, _26050_);
  nor (_26054_, _10678_, _02942_);
  or (_26055_, _26054_, _01537_);
  or (_26056_, _26055_, _26053_);
  and (_26057_, _11072_, _03853_);
  or (_26059_, _25946_, _01538_);
  or (_26060_, _26059_, _26057_);
  and (_26061_, _26060_, _38087_);
  and (_26062_, _26061_, _26056_);
  or (_40301_, _26062_, _25945_);
  nor (_26063_, _38087_, _01998_);
  or (_26064_, _03552_, _02942_);
  nor (_26065_, _03745_, _01998_);
  and (_26066_, _11094_, _03853_);
  or (_26067_, _26066_, _26065_);
  and (_26069_, _26067_, _02167_);
  nand (_26070_, _12061_, _01638_);
  nor (_26071_, _09213_, _03268_);
  or (_26072_, _26065_, _02528_);
  or (_26073_, _26072_, _26071_);
  and (_26074_, _26073_, _09212_);
  nor (_26075_, _11101_, _09213_);
  or (_26076_, _26075_, _26065_);
  or (_26077_, _26076_, _02814_);
  and (_26078_, _03745_, \oc8051_golden_model_1.ACC [3]);
  or (_26080_, _26078_, _26065_);
  and (_26081_, _26080_, _02817_);
  and (_26082_, _09224_, \oc8051_golden_model_1.SP [3]);
  nor (_26083_, _12061_, _01562_);
  or (_26084_, _26083_, _02001_);
  or (_26085_, _26084_, _26082_);
  or (_26086_, _26085_, _26081_);
  and (_26087_, _26086_, _01558_);
  and (_26088_, _26087_, _26077_);
  nor (_26089_, _12061_, _01558_);
  or (_26091_, _26089_, _01999_);
  or (_26092_, _26091_, _26088_);
  nand (_26093_, _04401_, _01999_);
  and (_26094_, _26093_, _26092_);
  or (_26095_, _26094_, _02006_);
  or (_26096_, _26080_, _02021_);
  and (_26097_, _26096_, _01880_);
  and (_26098_, _26097_, _26095_);
  or (_26099_, _03319_, _03132_);
  or (_26100_, _26099_, _26098_);
  nand (_26102_, _12061_, _03132_);
  and (_26103_, _26102_, _05249_);
  and (_26104_, _26103_, _26100_);
  or (_26105_, _26104_, _26074_);
  or (_26106_, _26065_, _02888_);
  and (_26107_, _04998_, _03745_);
  or (_26108_, _26107_, _26106_);
  and (_26109_, _26108_, _02043_);
  and (_26110_, _26109_, _26105_);
  nor (_26111_, _11206_, _25996_);
  or (_26113_, _26111_, _26065_);
  and (_26114_, _26113_, _01602_);
  or (_26115_, _26114_, _01869_);
  or (_26116_, _26115_, _26110_);
  and (_26117_, _03745_, _04678_);
  or (_26118_, _26117_, _26065_);
  or (_26119_, _26118_, _01870_);
  and (_26120_, _26119_, _26116_);
  or (_26121_, _26120_, _01638_);
  and (_26122_, _26121_, _26070_);
  or (_26124_, _26122_, _02079_);
  and (_26125_, _11222_, _03853_);
  or (_26126_, _26065_, _02166_);
  or (_26127_, _26126_, _26125_);
  and (_26128_, _26127_, _02912_);
  and (_26129_, _26128_, _26124_);
  or (_26130_, _26129_, _26069_);
  and (_26131_, _26130_, _02176_);
  or (_26132_, _26065_, _04014_);
  and (_26133_, _26118_, _02072_);
  and (_26135_, _26133_, _26132_);
  or (_26136_, _26135_, _26131_);
  and (_26137_, _26136_, _09292_);
  and (_26138_, _26080_, _02177_);
  and (_26139_, _26138_, _26132_);
  and (_26140_, _03552_, _01632_);
  or (_26141_, _26140_, _02071_);
  or (_26142_, _26141_, _26139_);
  or (_26143_, _26142_, _26137_);
  nor (_26144_, _11220_, _25996_);
  or (_26146_, _26144_, _26065_);
  or (_26147_, _26146_, _04788_);
  and (_26148_, _26147_, _26143_);
  or (_26149_, _26148_, _02173_);
  nor (_26150_, _11093_, _09213_);
  or (_26151_, _26065_, _04793_);
  or (_26152_, _26151_, _26150_);
  and (_26153_, _26152_, _09305_);
  and (_26154_, _26153_, _26149_);
  nor (_26155_, _04398_, _01998_);
  or (_26157_, _26155_, _04399_);
  and (_26158_, _26157_, _02185_);
  or (_26159_, _26158_, _01636_);
  or (_26160_, _26159_, _26154_);
  nand (_26161_, _12061_, _01636_);
  and (_26162_, _26161_, _26160_);
  or (_26163_, _26162_, _01888_);
  or (_26164_, _26157_, _01889_);
  and (_26165_, _26164_, _02303_);
  and (_26166_, _26165_, _26163_);
  and (_26168_, _26076_, _02201_);
  or (_26169_, _26168_, _03370_);
  or (_26170_, _26169_, _26166_);
  and (_26171_, _26170_, _26064_);
  or (_26172_, _26171_, _01537_);
  and (_26173_, _11273_, _03853_);
  or (_26174_, _26065_, _01538_);
  or (_26175_, _26174_, _26173_);
  and (_26176_, _26175_, _38087_);
  and (_26177_, _26176_, _26172_);
  or (_26179_, _26177_, _26063_);
  and (_40302_, _26179_, _37580_);
  nor (_26180_, _38087_, _09237_);
  nor (_26181_, _03549_, \oc8051_golden_model_1.SP [4]);
  nor (_26182_, _26181_, _09200_);
  or (_26183_, _26182_, _02942_);
  nor (_26184_, _03745_, _09237_);
  and (_26185_, _11431_, _03853_);
  or (_26186_, _26185_, _26184_);
  and (_26187_, _26186_, _02167_);
  nor (_26189_, _04211_, _09213_);
  or (_26190_, _26184_, _02528_);
  or (_26191_, _26190_, _26189_);
  and (_26192_, _26191_, _09212_);
  nor (_26193_, _11317_, _09213_);
  or (_26194_, _26193_, _26184_);
  or (_26195_, _26194_, _02814_);
  and (_26196_, _03745_, \oc8051_golden_model_1.ACC [4]);
  or (_26197_, _26196_, _26184_);
  and (_26198_, _26197_, _02817_);
  and (_26200_, _09224_, \oc8051_golden_model_1.SP [4]);
  and (_26201_, _26182_, _02823_);
  or (_26202_, _26201_, _02001_);
  or (_26203_, _26202_, _26200_);
  or (_26204_, _26203_, _26198_);
  and (_26205_, _26204_, _01558_);
  and (_26206_, _26205_, _26195_);
  and (_26207_, _26182_, _03279_);
  or (_26208_, _26207_, _01999_);
  or (_26209_, _26208_, _26206_);
  and (_26211_, _09238_, _01864_);
  nor (_26212_, _04400_, _09237_);
  nor (_26213_, _26212_, _26211_);
  nand (_26214_, _26213_, _01999_);
  and (_26215_, _26214_, _26209_);
  or (_26216_, _26215_, _02006_);
  or (_26217_, _26197_, _02021_);
  and (_26218_, _26217_, _01880_);
  and (_26219_, _26218_, _26216_);
  and (_26220_, _03275_, \oc8051_golden_model_1.SP [4]);
  nor (_26222_, _03275_, \oc8051_golden_model_1.SP [4]);
  nor (_26223_, _26222_, _26220_);
  and (_26224_, _26223_, _01878_);
  or (_26225_, _26224_, _03132_);
  or (_26226_, _26225_, _26219_);
  or (_26227_, _26182_, _03133_);
  and (_26228_, _26227_, _05249_);
  and (_26229_, _26228_, _26226_);
  or (_26230_, _26229_, _26192_);
  or (_26231_, _26184_, _02888_);
  and (_26232_, _05135_, _03745_);
  or (_26233_, _26232_, _26231_);
  and (_26234_, _26233_, _02043_);
  and (_26235_, _26234_, _26230_);
  nor (_26236_, _11411_, _25996_);
  or (_26237_, _26236_, _26184_);
  and (_26238_, _26237_, _01602_);
  or (_26239_, _26238_, _01869_);
  or (_26240_, _26239_, _26235_);
  and (_26241_, _04694_, _03745_);
  or (_26243_, _26241_, _26184_);
  or (_26244_, _26243_, _01870_);
  and (_26245_, _26244_, _26240_);
  or (_26246_, _26245_, _01638_);
  or (_26247_, _26182_, _09277_);
  and (_26248_, _26247_, _26246_);
  or (_26249_, _26248_, _02079_);
  and (_26250_, _11425_, _03853_);
  or (_26251_, _26184_, _02166_);
  or (_26252_, _26251_, _26250_);
  and (_26254_, _26252_, _02912_);
  and (_26255_, _26254_, _26249_);
  or (_26256_, _26255_, _26187_);
  and (_26257_, _26256_, _02176_);
  or (_26258_, _26184_, _04258_);
  and (_26259_, _26243_, _02072_);
  and (_26260_, _26259_, _26258_);
  or (_26261_, _26260_, _26257_);
  and (_26262_, _26261_, _09292_);
  and (_26263_, _26197_, _02177_);
  and (_26265_, _26263_, _26258_);
  and (_26266_, _26182_, _01632_);
  or (_26267_, _26266_, _02071_);
  or (_26268_, _26267_, _26265_);
  or (_26269_, _26268_, _26262_);
  nor (_26270_, _11424_, _25996_);
  or (_26271_, _26270_, _26184_);
  or (_26272_, _26271_, _04788_);
  and (_26273_, _26272_, _26269_);
  or (_26274_, _26273_, _02173_);
  nor (_26276_, _11430_, _09213_);
  or (_26277_, _26184_, _04793_);
  or (_26278_, _26277_, _26276_);
  and (_26279_, _26278_, _09305_);
  and (_26280_, _26279_, _26274_);
  nor (_26281_, _04399_, _09237_);
  or (_26282_, _26281_, _09238_);
  and (_26283_, _26282_, _02185_);
  or (_26284_, _26283_, _01636_);
  or (_26285_, _26284_, _26280_);
  or (_26287_, _26182_, _04799_);
  and (_26288_, _26287_, _26285_);
  or (_26289_, _26288_, _01888_);
  or (_26290_, _26282_, _01889_);
  and (_26291_, _26290_, _02303_);
  and (_26292_, _26291_, _26289_);
  and (_26293_, _26194_, _02201_);
  or (_26294_, _26293_, _03370_);
  or (_26295_, _26294_, _26292_);
  and (_26296_, _26295_, _26183_);
  or (_26298_, _26296_, _01537_);
  and (_26299_, _11487_, _03853_);
  or (_26300_, _26184_, _01538_);
  or (_26301_, _26300_, _26299_);
  and (_26302_, _26301_, _38087_);
  and (_26303_, _26302_, _26298_);
  or (_26304_, _26303_, _26180_);
  and (_40304_, _26304_, _37580_);
  nor (_26305_, _38087_, _09236_);
  nor (_26306_, _09200_, \oc8051_golden_model_1.SP [5]);
  nor (_26308_, _26306_, _09201_);
  or (_26309_, _26308_, _02942_);
  nor (_26310_, _03745_, _09236_);
  and (_26311_, _11635_, _03853_);
  or (_26312_, _26311_, _26310_);
  and (_26313_, _26312_, _02167_);
  nor (_26314_, _03916_, _09213_);
  or (_26315_, _26310_, _02528_);
  or (_26316_, _26315_, _26314_);
  and (_26317_, _26316_, _09212_);
  nor (_26319_, _11525_, _09213_);
  or (_26320_, _26319_, _26310_);
  or (_26321_, _26320_, _02814_);
  and (_26322_, _03745_, \oc8051_golden_model_1.ACC [5]);
  or (_26323_, _26322_, _26310_);
  and (_26324_, _26323_, _02817_);
  and (_26325_, _09224_, \oc8051_golden_model_1.SP [5]);
  and (_26326_, _26308_, _02823_);
  or (_26327_, _26326_, _02001_);
  or (_26328_, _26327_, _26325_);
  or (_26330_, _26328_, _26324_);
  and (_26331_, _26330_, _01558_);
  and (_26332_, _26331_, _26321_);
  and (_26333_, _26308_, _03279_);
  or (_26334_, _26333_, _01999_);
  or (_26335_, _26334_, _26332_);
  and (_26336_, _09239_, _01864_);
  nor (_26337_, _26211_, _09236_);
  nor (_26338_, _26337_, _26336_);
  nand (_26339_, _26338_, _01999_);
  and (_26341_, _26339_, _26335_);
  or (_26342_, _26341_, _02006_);
  or (_26343_, _26323_, _02021_);
  and (_26344_, _26343_, _01880_);
  and (_26345_, _26344_, _26342_);
  and (_26346_, _09201_, \oc8051_golden_model_1.SP [0]);
  nor (_26347_, _26220_, \oc8051_golden_model_1.SP [5]);
  nor (_26348_, _26347_, _26346_);
  and (_26349_, _26348_, _01878_);
  or (_26350_, _26349_, _03132_);
  or (_26352_, _26350_, _26345_);
  or (_26353_, _26308_, _03133_);
  and (_26354_, _26353_, _05249_);
  and (_26355_, _26354_, _26352_);
  or (_26356_, _26355_, _26317_);
  or (_26357_, _26310_, _02888_);
  and (_26358_, _05090_, _03745_);
  or (_26359_, _26358_, _26357_);
  and (_26360_, _26359_, _02043_);
  and (_26361_, _26360_, _26356_);
  nor (_26363_, _11615_, _25996_);
  or (_26364_, _26363_, _26310_);
  and (_26365_, _26364_, _01602_);
  or (_26366_, _26365_, _01869_);
  or (_26367_, _26366_, _26361_);
  and (_26368_, _04672_, _03745_);
  or (_26369_, _26368_, _26310_);
  or (_26370_, _26369_, _01870_);
  and (_26371_, _26370_, _26367_);
  or (_26372_, _26371_, _01638_);
  or (_26374_, _26308_, _09277_);
  and (_26375_, _26374_, _26372_);
  or (_26376_, _26375_, _02079_);
  and (_26377_, _11629_, _03853_);
  or (_26378_, _26310_, _02166_);
  or (_26379_, _26378_, _26377_);
  and (_26380_, _26379_, _02912_);
  and (_26381_, _26380_, _26376_);
  or (_26382_, _26381_, _26313_);
  and (_26383_, _26382_, _02176_);
  or (_26384_, _26310_, _03965_);
  and (_26385_, _26369_, _02072_);
  and (_26386_, _26385_, _26384_);
  or (_26387_, _26386_, _26383_);
  and (_26388_, _26387_, _09292_);
  and (_26389_, _26323_, _02177_);
  and (_26390_, _26389_, _26384_);
  and (_26391_, _26308_, _01632_);
  or (_26392_, _26391_, _02071_);
  or (_26393_, _26392_, _26390_);
  or (_26395_, _26393_, _26388_);
  nor (_26396_, _11628_, _25996_);
  or (_26397_, _26396_, _26310_);
  or (_26398_, _26397_, _04788_);
  and (_26399_, _26398_, _26395_);
  or (_26400_, _26399_, _02173_);
  nor (_26401_, _11634_, _09213_);
  or (_26402_, _26310_, _04793_);
  or (_26403_, _26402_, _26401_);
  and (_26404_, _26403_, _09305_);
  and (_26406_, _26404_, _26400_);
  nor (_26407_, _09238_, _09236_);
  or (_26408_, _26407_, _09239_);
  and (_26409_, _26408_, _02185_);
  or (_26410_, _26409_, _01636_);
  or (_26411_, _26410_, _26406_);
  or (_26412_, _26308_, _04799_);
  and (_26413_, _26412_, _26411_);
  or (_26414_, _26413_, _01888_);
  or (_26415_, _26408_, _01889_);
  and (_26417_, _26415_, _02303_);
  and (_26418_, _26417_, _26414_);
  and (_26419_, _26320_, _02201_);
  or (_26420_, _26419_, _03370_);
  or (_26421_, _26420_, _26418_);
  and (_26422_, _26421_, _26309_);
  or (_26423_, _26422_, _01537_);
  and (_26424_, _11685_, _03853_);
  or (_26425_, _26310_, _01538_);
  or (_26426_, _26425_, _26424_);
  and (_26428_, _26426_, _38087_);
  and (_26429_, _26428_, _26423_);
  or (_26430_, _26429_, _26305_);
  and (_40305_, _26430_, _37580_);
  nor (_26431_, _38087_, _09235_);
  nor (_26432_, _03745_, _09235_);
  and (_26433_, _11709_, _03853_);
  or (_26434_, _26433_, _26432_);
  and (_26435_, _26434_, _02167_);
  nor (_26436_, _11730_, _09213_);
  or (_26438_, _26436_, _26432_);
  or (_26439_, _26438_, _02814_);
  and (_26440_, _03745_, \oc8051_golden_model_1.ACC [6]);
  or (_26441_, _26440_, _26432_);
  and (_26442_, _26441_, _02817_);
  and (_26443_, _09224_, \oc8051_golden_model_1.SP [6]);
  nor (_26444_, _09201_, \oc8051_golden_model_1.SP [6]);
  nor (_26445_, _26444_, _09202_);
  and (_26446_, _26445_, _02823_);
  or (_26447_, _26446_, _02001_);
  or (_26449_, _26447_, _26443_);
  or (_26450_, _26449_, _26442_);
  and (_26451_, _26450_, _01558_);
  and (_26452_, _26451_, _26439_);
  and (_26453_, _26445_, _03279_);
  or (_26454_, _26453_, _01999_);
  or (_26455_, _26454_, _26452_);
  nor (_26456_, _26336_, _09235_);
  nor (_26457_, _26456_, _09241_);
  nand (_26458_, _26457_, _01999_);
  and (_26460_, _26458_, _26455_);
  or (_26461_, _26460_, _02006_);
  or (_26462_, _26441_, _02021_);
  and (_26463_, _26462_, _01880_);
  and (_26464_, _26463_, _26461_);
  nor (_26465_, _26346_, \oc8051_golden_model_1.SP [6]);
  nor (_26466_, _26465_, _09251_);
  and (_26467_, _26466_, _01878_);
  or (_26468_, _26467_, _26464_);
  and (_26469_, _26468_, _03133_);
  nand (_26471_, _26445_, _03132_);
  nand (_26472_, _26471_, _05249_);
  or (_26473_, _26472_, _26469_);
  nor (_26474_, _03808_, _09213_);
  or (_26475_, _26432_, _05249_);
  or (_26476_, _26475_, _26474_);
  and (_26477_, _26476_, _26473_);
  or (_26478_, _26477_, _02528_);
  and (_26479_, _04861_, _03745_);
  or (_26480_, _26432_, _02888_);
  or (_26482_, _26480_, _26479_);
  and (_26483_, _26482_, _02043_);
  and (_26484_, _26483_, _26478_);
  nor (_26485_, _11820_, _09213_);
  or (_26486_, _26485_, _26432_);
  and (_26487_, _26486_, _01602_);
  or (_26488_, _26487_, _01869_);
  or (_26489_, _26488_, _26484_);
  and (_26490_, _09920_, _03745_);
  or (_26491_, _26490_, _26432_);
  or (_26493_, _26491_, _01870_);
  and (_26494_, _26493_, _26489_);
  or (_26495_, _26494_, _01638_);
  or (_26496_, _26445_, _09277_);
  and (_26497_, _26496_, _26495_);
  or (_26498_, _26497_, _02079_);
  and (_26499_, _11835_, _03853_);
  or (_26500_, _26432_, _02166_);
  or (_26501_, _26500_, _26499_);
  and (_26502_, _26501_, _02912_);
  and (_26504_, _26502_, _26498_);
  or (_26505_, _26504_, _26435_);
  and (_26506_, _26505_, _02176_);
  or (_26507_, _26432_, _03863_);
  and (_26508_, _26491_, _02072_);
  and (_26509_, _26508_, _26507_);
  or (_26510_, _26509_, _26506_);
  and (_26511_, _26510_, _09292_);
  and (_26512_, _26441_, _02177_);
  and (_26513_, _26512_, _26507_);
  and (_26515_, _26445_, _01632_);
  or (_26516_, _26515_, _02071_);
  or (_26517_, _26516_, _26513_);
  or (_26518_, _26517_, _26511_);
  nor (_26519_, _11833_, _25996_);
  or (_26520_, _26519_, _26432_);
  or (_26521_, _26520_, _04788_);
  and (_26522_, _26521_, _26518_);
  or (_26523_, _26522_, _02173_);
  nor (_26524_, _11708_, _09213_);
  or (_26525_, _26432_, _04793_);
  or (_26526_, _26525_, _26524_);
  and (_26527_, _26526_, _09305_);
  and (_26528_, _26527_, _26523_);
  nor (_26529_, _09239_, _09235_);
  or (_26530_, _26529_, _09240_);
  and (_26531_, _26530_, _02185_);
  or (_26532_, _26531_, _01636_);
  or (_26533_, _26532_, _26528_);
  or (_26534_, _26445_, _04799_);
  and (_26536_, _26534_, _01889_);
  and (_26537_, _26536_, _26533_);
  and (_26538_, _26530_, _01888_);
  or (_26539_, _26538_, _02201_);
  or (_26540_, _26539_, _26537_);
  or (_26541_, _26438_, _02303_);
  and (_26542_, _26541_, _02942_);
  and (_26543_, _26542_, _26540_);
  and (_26544_, _26445_, _03370_);
  or (_26545_, _26544_, _01537_);
  or (_26547_, _26545_, _26543_);
  and (_26548_, _11887_, _03853_);
  or (_26549_, _26432_, _01538_);
  or (_26550_, _26549_, _26548_);
  and (_26551_, _26550_, _38087_);
  and (_26552_, _26551_, _26547_);
  or (_26553_, _26552_, _26431_);
  and (_40306_, _26553_, _37580_);
  and (_26554_, _38088_, \oc8051_golden_model_1.TCON [0]);
  and (_26555_, _09335_, \oc8051_golden_model_1.TCON [0]);
  and (_26557_, _10620_, _03693_);
  or (_26558_, _26557_, _26555_);
  and (_26559_, _26558_, _02167_);
  and (_26560_, _03693_, _03028_);
  or (_26561_, _26560_, _26555_);
  or (_26562_, _26561_, _05249_);
  nor (_26563_, _04106_, _09335_);
  or (_26564_, _26563_, _26555_);
  or (_26565_, _26564_, _02814_);
  and (_26566_, _03693_, \oc8051_golden_model_1.ACC [0]);
  or (_26568_, _26566_, _26555_);
  and (_26569_, _26568_, _02817_);
  and (_26570_, _02818_, \oc8051_golden_model_1.TCON [0]);
  or (_26571_, _26570_, _02001_);
  or (_26572_, _26571_, _26569_);
  and (_26573_, _26572_, _02024_);
  and (_26574_, _26573_, _26565_);
  and (_26575_, _09343_, \oc8051_golden_model_1.TCON [0]);
  and (_26576_, _10510_, _04315_);
  or (_26577_, _26576_, _26575_);
  and (_26579_, _26577_, _02007_);
  or (_26580_, _26579_, _26574_);
  and (_26581_, _26580_, _02840_);
  and (_26582_, _26561_, _01999_);
  or (_26583_, _26582_, _02006_);
  or (_26584_, _26583_, _26581_);
  or (_26585_, _26568_, _02021_);
  and (_26586_, _26585_, _02025_);
  and (_26587_, _26586_, _26584_);
  and (_26588_, _26555_, _01997_);
  or (_26590_, _26588_, _01991_);
  or (_26591_, _26590_, _26587_);
  or (_26592_, _26564_, _02861_);
  and (_26593_, _26592_, _02408_);
  and (_26594_, _26593_, _26591_);
  nor (_26595_, _10542_, _09343_);
  or (_26596_, _26595_, _26575_);
  and (_26597_, _26596_, _01875_);
  or (_26598_, _26597_, _05994_);
  or (_26599_, _26598_, _26594_);
  and (_26601_, _26599_, _26562_);
  or (_26602_, _26601_, _02528_);
  and (_26603_, _04952_, _03693_);
  or (_26604_, _26555_, _02888_);
  or (_26605_, _26604_, _26603_);
  and (_26606_, _26605_, _02043_);
  and (_26607_, _26606_, _26602_);
  nor (_26608_, _10600_, _09335_);
  or (_26609_, _26608_, _26555_);
  and (_26610_, _26609_, _01602_);
  or (_26612_, _26610_, _01869_);
  or (_26613_, _26612_, _26607_);
  and (_26614_, _03693_, _04562_);
  or (_26615_, _26614_, _26555_);
  or (_26616_, _26615_, _01870_);
  and (_26617_, _26616_, _26613_);
  or (_26618_, _26617_, _02079_);
  and (_26619_, _10614_, _03693_);
  or (_26620_, _26555_, _02166_);
  or (_26621_, _26620_, _26619_);
  and (_26623_, _26621_, _02912_);
  and (_26624_, _26623_, _26618_);
  or (_26625_, _26624_, _26559_);
  and (_26626_, _26625_, _02176_);
  nand (_26627_, _26615_, _02072_);
  nor (_26628_, _26627_, _26563_);
  or (_26629_, _26628_, _26626_);
  and (_26630_, _26629_, _02907_);
  or (_26631_, _26555_, _04106_);
  and (_26632_, _26568_, _02177_);
  and (_26634_, _26632_, _26631_);
  or (_26635_, _26634_, _02071_);
  or (_26636_, _26635_, _26630_);
  nor (_26637_, _10613_, _09335_);
  or (_26638_, _26555_, _04788_);
  or (_26639_, _26638_, _26637_);
  and (_26640_, _26639_, _04793_);
  and (_26641_, _26640_, _26636_);
  nor (_26642_, _10619_, _09335_);
  or (_26643_, _26642_, _26555_);
  and (_26645_, _26643_, _02173_);
  or (_26646_, _26645_, _02201_);
  or (_26647_, _26646_, _26641_);
  or (_26648_, _26564_, _02303_);
  and (_26649_, _26648_, _01887_);
  and (_26650_, _26649_, _26647_);
  and (_26651_, _26555_, _01860_);
  or (_26652_, _26651_, _01537_);
  or (_26653_, _26652_, _26650_);
  or (_26654_, _26564_, _01538_);
  and (_26656_, _26654_, _38087_);
  and (_26657_, _26656_, _26653_);
  or (_26658_, _26657_, _26554_);
  and (_40308_, _26658_, _37580_);
  and (_26659_, _09335_, \oc8051_golden_model_1.TCON [1]);
  nor (_26660_, _09335_, _02811_);
  or (_26661_, _26660_, _26659_);
  or (_26662_, _26661_, _02840_);
  or (_26663_, _03693_, \oc8051_golden_model_1.TCON [1]);
  and (_26664_, _10698_, _03693_);
  not (_26666_, _26664_);
  and (_26667_, _26666_, _26663_);
  or (_26668_, _26667_, _02814_);
  nand (_26669_, _03693_, _01613_);
  and (_26670_, _26669_, _26663_);
  and (_26671_, _26670_, _02817_);
  and (_26672_, _02818_, \oc8051_golden_model_1.TCON [1]);
  or (_26673_, _26672_, _02001_);
  or (_26674_, _26673_, _26671_);
  and (_26675_, _26674_, _02024_);
  and (_26676_, _26675_, _26668_);
  and (_26677_, _09343_, \oc8051_golden_model_1.TCON [1]);
  and (_26678_, _10710_, _04315_);
  or (_26679_, _26678_, _26677_);
  and (_26680_, _26679_, _02007_);
  or (_26681_, _26680_, _01999_);
  or (_26682_, _26681_, _26676_);
  and (_26683_, _26682_, _26662_);
  or (_26684_, _26683_, _02006_);
  or (_26685_, _26670_, _02021_);
  and (_26687_, _26685_, _02025_);
  and (_26688_, _26687_, _26684_);
  and (_26689_, _10696_, _04315_);
  or (_26690_, _26689_, _26677_);
  and (_26691_, _26690_, _01997_);
  or (_26692_, _26691_, _01991_);
  or (_26693_, _26692_, _26688_);
  and (_26694_, _26678_, _10725_);
  or (_26695_, _26677_, _02861_);
  or (_26696_, _26695_, _26694_);
  and (_26698_, _26696_, _26693_);
  and (_26699_, _26698_, _02408_);
  nor (_26700_, _10742_, _09343_);
  or (_26701_, _26677_, _26700_);
  and (_26702_, _26701_, _01875_);
  or (_26703_, _26702_, _05994_);
  or (_26704_, _26703_, _26699_);
  or (_26705_, _26661_, _05249_);
  and (_26706_, _26705_, _26704_);
  or (_26707_, _26706_, _02528_);
  and (_26709_, _04907_, _03693_);
  or (_26710_, _26659_, _02888_);
  or (_26711_, _26710_, _26709_);
  and (_26712_, _26711_, _02043_);
  and (_26713_, _26712_, _26707_);
  nor (_26714_, _10802_, _09335_);
  or (_26715_, _26714_, _26659_);
  and (_26716_, _26715_, _01602_);
  or (_26717_, _26716_, _26713_);
  and (_26718_, _26717_, _01870_);
  nand (_26720_, _03693_, _02687_);
  and (_26721_, _26663_, _01869_);
  and (_26722_, _26721_, _26720_);
  or (_26723_, _26722_, _26718_);
  and (_26724_, _26723_, _02166_);
  or (_26725_, _10816_, _09335_);
  and (_26726_, _26663_, _02079_);
  and (_26727_, _26726_, _26725_);
  or (_26728_, _26727_, _26724_);
  and (_26729_, _26728_, _02912_);
  or (_26731_, _10822_, _09335_);
  and (_26732_, _26663_, _02167_);
  and (_26733_, _26732_, _26731_);
  or (_26734_, _26733_, _26729_);
  and (_26735_, _26734_, _02176_);
  or (_26736_, _10692_, _09335_);
  and (_26737_, _26663_, _02072_);
  and (_26738_, _26737_, _26736_);
  or (_26739_, _26738_, _26735_);
  and (_26740_, _26739_, _02907_);
  or (_26742_, _26659_, _04058_);
  and (_26743_, _26670_, _02177_);
  and (_26744_, _26743_, _26742_);
  or (_26745_, _26744_, _26740_);
  and (_26746_, _26745_, _02174_);
  or (_26747_, _26669_, _04058_);
  and (_26748_, _26663_, _02173_);
  and (_26749_, _26748_, _26747_);
  or (_26750_, _26749_, _02201_);
  or (_26751_, _26720_, _04058_);
  and (_26753_, _26663_, _02071_);
  and (_26754_, _26753_, _26751_);
  or (_26755_, _26754_, _26750_);
  or (_26756_, _26755_, _26746_);
  or (_26757_, _26667_, _02303_);
  and (_26758_, _26757_, _01887_);
  and (_26759_, _26758_, _26756_);
  and (_26760_, _26690_, _01860_);
  or (_26761_, _26760_, _01537_);
  or (_26762_, _26761_, _26759_);
  or (_26764_, _26659_, _01538_);
  or (_26765_, _26764_, _26664_);
  and (_26766_, _26765_, _38087_);
  and (_26767_, _26766_, _26762_);
  nor (_26768_, \oc8051_golden_model_1.TCON [1], rst);
  nor (_26769_, _26768_, _03183_);
  or (_40309_, _26769_, _26767_);
  and (_26770_, _38088_, \oc8051_golden_model_1.TCON [2]);
  and (_26771_, _09335_, \oc8051_golden_model_1.TCON [2]);
  and (_26772_, _11020_, _03693_);
  or (_26774_, _26772_, _26771_);
  and (_26775_, _26774_, _02167_);
  nor (_26776_, _09335_, _03455_);
  or (_26777_, _26776_, _26771_);
  or (_26778_, _26777_, _05249_);
  or (_26779_, _26777_, _02840_);
  nor (_26780_, _10905_, _09335_);
  or (_26781_, _26780_, _26771_);
  or (_26782_, _26781_, _02814_);
  and (_26783_, _03693_, \oc8051_golden_model_1.ACC [2]);
  or (_26785_, _26783_, _26771_);
  and (_26786_, _26785_, _02817_);
  and (_26787_, _02818_, \oc8051_golden_model_1.TCON [2]);
  or (_26788_, _26787_, _02001_);
  or (_26789_, _26788_, _26786_);
  and (_26790_, _26789_, _02024_);
  and (_26791_, _26790_, _26782_);
  and (_26792_, _09343_, \oc8051_golden_model_1.TCON [2]);
  and (_26793_, _10909_, _04315_);
  or (_26794_, _26793_, _26792_);
  and (_26796_, _26794_, _02007_);
  or (_26797_, _26796_, _01999_);
  or (_26798_, _26797_, _26791_);
  and (_26799_, _26798_, _26779_);
  or (_26800_, _26799_, _02006_);
  or (_26801_, _26785_, _02021_);
  and (_26802_, _26801_, _02025_);
  and (_26803_, _26802_, _26800_);
  and (_26804_, _10894_, _04315_);
  or (_26805_, _26804_, _26792_);
  and (_26807_, _26805_, _01997_);
  or (_26808_, _26807_, _01991_);
  or (_26809_, _26808_, _26803_);
  and (_26810_, _26793_, _10924_);
  or (_26811_, _26792_, _02861_);
  or (_26812_, _26811_, _26810_);
  and (_26813_, _26812_, _02408_);
  and (_26814_, _26813_, _26809_);
  nor (_26815_, _10942_, _09343_);
  or (_26816_, _26815_, _26792_);
  and (_26818_, _26816_, _01875_);
  or (_26819_, _26818_, _05994_);
  or (_26820_, _26819_, _26814_);
  and (_26821_, _26820_, _26778_);
  or (_26822_, _26821_, _02528_);
  and (_26823_, _05043_, _03693_);
  or (_26824_, _26771_, _02888_);
  or (_26825_, _26824_, _26823_);
  and (_26826_, _26825_, _02043_);
  and (_26827_, _26826_, _26822_);
  nor (_26828_, _11000_, _09335_);
  or (_26829_, _26828_, _26771_);
  and (_26830_, _26829_, _01602_);
  or (_26831_, _26830_, _01869_);
  or (_26832_, _26831_, _26827_);
  and (_26833_, _03693_, _04724_);
  or (_26834_, _26833_, _26771_);
  or (_26835_, _26834_, _01870_);
  and (_26836_, _26835_, _26832_);
  or (_26837_, _26836_, _02079_);
  and (_26839_, _11014_, _03693_);
  or (_26840_, _26771_, _02166_);
  or (_26841_, _26840_, _26839_);
  and (_26842_, _26841_, _02912_);
  and (_26843_, _26842_, _26837_);
  or (_26844_, _26843_, _26775_);
  and (_26845_, _26844_, _02176_);
  or (_26846_, _26771_, _04156_);
  and (_26847_, _26834_, _02072_);
  and (_26848_, _26847_, _26846_);
  or (_26850_, _26848_, _26845_);
  and (_26851_, _26850_, _02907_);
  and (_26852_, _26785_, _02177_);
  and (_26853_, _26852_, _26846_);
  or (_26854_, _26853_, _02071_);
  or (_26855_, _26854_, _26851_);
  nor (_26856_, _11013_, _09335_);
  or (_26857_, _26771_, _04788_);
  or (_26858_, _26857_, _26856_);
  and (_26859_, _26858_, _04793_);
  and (_26861_, _26859_, _26855_);
  nor (_26862_, _11019_, _09335_);
  or (_26863_, _26862_, _26771_);
  and (_26864_, _26863_, _02173_);
  or (_26865_, _26864_, _02201_);
  or (_26866_, _26865_, _26861_);
  or (_26867_, _26781_, _02303_);
  and (_26868_, _26867_, _01887_);
  and (_26869_, _26868_, _26866_);
  and (_26870_, _26805_, _01860_);
  or (_26872_, _26870_, _01537_);
  or (_26873_, _26872_, _26869_);
  and (_26874_, _11072_, _03693_);
  or (_26875_, _26771_, _01538_);
  or (_26876_, _26875_, _26874_);
  and (_26877_, _26876_, _38087_);
  and (_26878_, _26877_, _26873_);
  or (_26879_, _26878_, _26770_);
  and (_40310_, _26879_, _37580_);
  and (_26880_, _38088_, \oc8051_golden_model_1.TCON [3]);
  and (_26882_, _09335_, \oc8051_golden_model_1.TCON [3]);
  and (_26883_, _11094_, _03693_);
  or (_26884_, _26883_, _26882_);
  and (_26885_, _26884_, _02167_);
  nor (_26886_, _09335_, _03268_);
  or (_26887_, _26886_, _26882_);
  or (_26888_, _26887_, _05249_);
  nor (_26889_, _11101_, _09335_);
  or (_26890_, _26889_, _26882_);
  or (_26891_, _26890_, _02814_);
  and (_26893_, _03693_, \oc8051_golden_model_1.ACC [3]);
  or (_26894_, _26893_, _26882_);
  and (_26895_, _26894_, _02817_);
  and (_26896_, _02818_, \oc8051_golden_model_1.TCON [3]);
  or (_26897_, _26896_, _02001_);
  or (_26898_, _26897_, _26895_);
  and (_26899_, _26898_, _02024_);
  and (_26900_, _26899_, _26891_);
  and (_26901_, _09343_, \oc8051_golden_model_1.TCON [3]);
  and (_26902_, _11098_, _04315_);
  or (_26904_, _26902_, _26901_);
  and (_26905_, _26904_, _02007_);
  or (_26906_, _26905_, _01999_);
  or (_26907_, _26906_, _26900_);
  or (_26908_, _26887_, _02840_);
  and (_26909_, _26908_, _26907_);
  or (_26910_, _26909_, _02006_);
  or (_26911_, _26894_, _02021_);
  and (_26912_, _26911_, _02025_);
  and (_26913_, _26912_, _26910_);
  and (_26915_, _11096_, _04315_);
  or (_26916_, _26915_, _26901_);
  and (_26917_, _26916_, _01997_);
  or (_26918_, _26917_, _01991_);
  or (_26919_, _26918_, _26913_);
  or (_26920_, _26901_, _11127_);
  and (_26921_, _26920_, _26904_);
  or (_26922_, _26921_, _02861_);
  and (_26923_, _26922_, _02408_);
  and (_26924_, _26923_, _26919_);
  nor (_26926_, _11145_, _09343_);
  or (_26927_, _26926_, _26901_);
  and (_26928_, _26927_, _01875_);
  or (_26929_, _26928_, _05994_);
  or (_26930_, _26929_, _26924_);
  and (_26931_, _26930_, _26888_);
  or (_26932_, _26931_, _02528_);
  and (_26933_, _04998_, _03693_);
  or (_26934_, _26882_, _02888_);
  or (_26935_, _26934_, _26933_);
  and (_26937_, _26935_, _02043_);
  and (_26938_, _26937_, _26932_);
  nor (_26939_, _11206_, _09335_);
  or (_26940_, _26939_, _26882_);
  and (_26941_, _26940_, _01602_);
  or (_26942_, _26941_, _01869_);
  or (_26943_, _26942_, _26938_);
  and (_26944_, _03693_, _04678_);
  or (_26945_, _26944_, _26882_);
  or (_26946_, _26945_, _01870_);
  and (_26948_, _26946_, _26943_);
  or (_26949_, _26948_, _02079_);
  and (_26950_, _11222_, _03693_);
  or (_26951_, _26882_, _02166_);
  or (_26952_, _26951_, _26950_);
  and (_26953_, _26952_, _02912_);
  and (_26954_, _26953_, _26949_);
  or (_26955_, _26954_, _26885_);
  and (_26956_, _26955_, _02176_);
  or (_26957_, _26882_, _04014_);
  and (_26959_, _26945_, _02072_);
  and (_26960_, _26959_, _26957_);
  or (_26961_, _26960_, _26956_);
  and (_26962_, _26961_, _02907_);
  and (_26963_, _26894_, _02177_);
  and (_26964_, _26963_, _26957_);
  or (_26965_, _26964_, _02071_);
  or (_26966_, _26965_, _26962_);
  nor (_26967_, _11220_, _09335_);
  or (_26968_, _26882_, _04788_);
  or (_26970_, _26968_, _26967_);
  and (_26971_, _26970_, _04793_);
  and (_26972_, _26971_, _26966_);
  nor (_26973_, _11093_, _09335_);
  or (_26974_, _26973_, _26882_);
  and (_26975_, _26974_, _02173_);
  or (_26976_, _26975_, _02201_);
  or (_26977_, _26976_, _26972_);
  or (_26978_, _26890_, _02303_);
  and (_26979_, _26978_, _01887_);
  and (_26980_, _26979_, _26977_);
  and (_26981_, _26916_, _01860_);
  or (_26982_, _26981_, _01537_);
  or (_26983_, _26982_, _26980_);
  and (_26984_, _11273_, _03693_);
  or (_26985_, _26882_, _01538_);
  or (_26986_, _26985_, _26984_);
  and (_26987_, _26986_, _38087_);
  and (_26988_, _26987_, _26983_);
  or (_26989_, _26988_, _26880_);
  and (_40311_, _26989_, _37580_);
  and (_26991_, _38088_, \oc8051_golden_model_1.TCON [4]);
  and (_26992_, _09335_, \oc8051_golden_model_1.TCON [4]);
  and (_26993_, _11431_, _03693_);
  or (_26994_, _26993_, _26992_);
  and (_26995_, _26994_, _02167_);
  nor (_26996_, _04211_, _09335_);
  or (_26997_, _26996_, _26992_);
  or (_26998_, _26997_, _05249_);
  and (_26999_, _09343_, \oc8051_golden_model_1.TCON [4]);
  and (_27001_, _11301_, _04315_);
  or (_27002_, _27001_, _26999_);
  and (_27003_, _27002_, _01997_);
  nor (_27004_, _11317_, _09335_);
  or (_27005_, _27004_, _26992_);
  or (_27006_, _27005_, _02814_);
  and (_27007_, _03693_, \oc8051_golden_model_1.ACC [4]);
  or (_27008_, _27007_, _26992_);
  and (_27009_, _27008_, _02817_);
  and (_27010_, _02818_, \oc8051_golden_model_1.TCON [4]);
  or (_27012_, _27010_, _02001_);
  or (_27013_, _27012_, _27009_);
  and (_27014_, _27013_, _02024_);
  and (_27015_, _27014_, _27006_);
  and (_27016_, _11303_, _04315_);
  or (_27017_, _27016_, _26999_);
  and (_27018_, _27017_, _02007_);
  or (_27019_, _27018_, _01999_);
  or (_27020_, _27019_, _27015_);
  or (_27021_, _26997_, _02840_);
  and (_27023_, _27021_, _27020_);
  or (_27024_, _27023_, _02006_);
  or (_27025_, _27008_, _02021_);
  and (_27026_, _27025_, _02025_);
  and (_27027_, _27026_, _27024_);
  or (_27028_, _27027_, _27003_);
  and (_27029_, _27028_, _02861_);
  or (_27030_, _26999_, _11334_);
  and (_27031_, _27030_, _01991_);
  and (_27032_, _27031_, _27017_);
  or (_27034_, _27032_, _27029_);
  and (_27035_, _27034_, _02408_);
  nor (_27036_, _11299_, _09343_);
  or (_27037_, _27036_, _26999_);
  and (_27038_, _27037_, _01875_);
  or (_27039_, _27038_, _05994_);
  or (_27040_, _27039_, _27035_);
  and (_27041_, _27040_, _26998_);
  or (_27042_, _27041_, _02528_);
  and (_27043_, _05135_, _03693_);
  or (_27045_, _26992_, _02888_);
  or (_27046_, _27045_, _27043_);
  and (_27047_, _27046_, _02043_);
  and (_27048_, _27047_, _27042_);
  nor (_27049_, _11411_, _09335_);
  or (_27050_, _27049_, _26992_);
  and (_27051_, _27050_, _01602_);
  or (_27052_, _27051_, _01869_);
  or (_27053_, _27052_, _27048_);
  and (_27054_, _04694_, _03693_);
  or (_27056_, _27054_, _26992_);
  or (_27057_, _27056_, _01870_);
  and (_27058_, _27057_, _27053_);
  or (_27059_, _27058_, _02079_);
  and (_27060_, _11425_, _03693_);
  or (_27061_, _26992_, _02166_);
  or (_27062_, _27061_, _27060_);
  and (_27063_, _27062_, _02912_);
  and (_27064_, _27063_, _27059_);
  or (_27065_, _27064_, _26995_);
  and (_27067_, _27065_, _02176_);
  or (_27068_, _26992_, _04258_);
  and (_27069_, _27056_, _02072_);
  and (_27070_, _27069_, _27068_);
  or (_27071_, _27070_, _27067_);
  and (_27072_, _27071_, _02907_);
  and (_27073_, _27008_, _02177_);
  and (_27074_, _27073_, _27068_);
  or (_27075_, _27074_, _02071_);
  or (_27076_, _27075_, _27072_);
  nor (_27078_, _11424_, _09335_);
  or (_27079_, _26992_, _04788_);
  or (_27080_, _27079_, _27078_);
  and (_27081_, _27080_, _04793_);
  and (_27082_, _27081_, _27076_);
  nor (_27083_, _11430_, _09335_);
  or (_27084_, _27083_, _26992_);
  and (_27085_, _27084_, _02173_);
  or (_27086_, _27085_, _02201_);
  or (_27087_, _27086_, _27082_);
  or (_27089_, _27005_, _02303_);
  and (_27090_, _27089_, _01887_);
  and (_27091_, _27090_, _27087_);
  and (_27092_, _27002_, _01860_);
  or (_27093_, _27092_, _01537_);
  or (_27094_, _27093_, _27091_);
  and (_27095_, _11487_, _03693_);
  or (_27096_, _26992_, _01538_);
  or (_27097_, _27096_, _27095_);
  and (_27098_, _27097_, _38087_);
  and (_27100_, _27098_, _27094_);
  or (_27101_, _27100_, _26991_);
  and (_40312_, _27101_, _37580_);
  and (_27102_, _38088_, \oc8051_golden_model_1.TCON [5]);
  and (_27103_, _09335_, \oc8051_golden_model_1.TCON [5]);
  and (_27104_, _11635_, _03693_);
  or (_27105_, _27104_, _27103_);
  and (_27106_, _27105_, _02167_);
  nor (_27107_, _11525_, _09335_);
  or (_27108_, _27107_, _27103_);
  or (_27110_, _27108_, _02814_);
  and (_27111_, _03693_, \oc8051_golden_model_1.ACC [5]);
  or (_27112_, _27111_, _27103_);
  and (_27113_, _27112_, _02817_);
  and (_27114_, _02818_, \oc8051_golden_model_1.TCON [5]);
  or (_27115_, _27114_, _02001_);
  or (_27116_, _27115_, _27113_);
  and (_27117_, _27116_, _02024_);
  and (_27118_, _27117_, _27110_);
  and (_27119_, _09343_, \oc8051_golden_model_1.TCON [5]);
  and (_27121_, _11510_, _04315_);
  or (_27122_, _27121_, _27119_);
  and (_27123_, _27122_, _02007_);
  or (_27124_, _27123_, _01999_);
  or (_27125_, _27124_, _27118_);
  nor (_27126_, _03916_, _09335_);
  or (_27127_, _27126_, _27103_);
  or (_27128_, _27127_, _02840_);
  and (_27129_, _27128_, _27125_);
  or (_27130_, _27129_, _02006_);
  or (_27131_, _27112_, _02021_);
  and (_27132_, _27131_, _02025_);
  and (_27133_, _27132_, _27130_);
  and (_27134_, _11508_, _04315_);
  or (_27135_, _27134_, _27119_);
  and (_27136_, _27135_, _01997_);
  or (_27137_, _27136_, _01991_);
  or (_27138_, _27137_, _27133_);
  or (_27139_, _27119_, _11542_);
  and (_27140_, _27139_, _27122_);
  or (_27142_, _27140_, _02861_);
  and (_27143_, _27142_, _02408_);
  and (_27144_, _27143_, _27138_);
  nor (_27145_, _11506_, _09343_);
  or (_27146_, _27145_, _27119_);
  and (_27147_, _27146_, _01875_);
  or (_27148_, _27147_, _05994_);
  or (_27149_, _27148_, _27144_);
  or (_27150_, _27127_, _05249_);
  and (_27151_, _27150_, _27149_);
  or (_27153_, _27151_, _02528_);
  and (_27154_, _05090_, _03693_);
  or (_27155_, _27103_, _02888_);
  or (_27156_, _27155_, _27154_);
  and (_27157_, _27156_, _02043_);
  and (_27158_, _27157_, _27153_);
  nor (_27159_, _11615_, _09335_);
  or (_27160_, _27159_, _27103_);
  and (_27161_, _27160_, _01602_);
  or (_27162_, _27161_, _01869_);
  or (_27164_, _27162_, _27158_);
  and (_27165_, _04672_, _03693_);
  or (_27166_, _27165_, _27103_);
  or (_27167_, _27166_, _01870_);
  and (_27168_, _27167_, _27164_);
  or (_27169_, _27168_, _02079_);
  and (_27170_, _11629_, _03693_);
  or (_27171_, _27103_, _02166_);
  or (_27172_, _27171_, _27170_);
  and (_27173_, _27172_, _02912_);
  and (_27175_, _27173_, _27169_);
  or (_27176_, _27175_, _27106_);
  and (_27177_, _27176_, _02176_);
  or (_27178_, _27103_, _03965_);
  and (_27179_, _27166_, _02072_);
  and (_27180_, _27179_, _27178_);
  or (_27181_, _27180_, _27177_);
  and (_27182_, _27181_, _02907_);
  and (_27183_, _27112_, _02177_);
  and (_27184_, _27183_, _27178_);
  or (_27186_, _27184_, _02071_);
  or (_27187_, _27186_, _27182_);
  nor (_27188_, _11628_, _09335_);
  or (_27189_, _27103_, _04788_);
  or (_27190_, _27189_, _27188_);
  and (_27191_, _27190_, _04793_);
  and (_27192_, _27191_, _27187_);
  nor (_27193_, _11634_, _09335_);
  or (_27194_, _27193_, _27103_);
  and (_27195_, _27194_, _02173_);
  or (_27197_, _27195_, _02201_);
  or (_27198_, _27197_, _27192_);
  or (_27199_, _27108_, _02303_);
  and (_27200_, _27199_, _01887_);
  and (_27201_, _27200_, _27198_);
  and (_27202_, _27135_, _01860_);
  or (_27203_, _27202_, _01537_);
  or (_27204_, _27203_, _27201_);
  and (_27205_, _11685_, _03693_);
  or (_27206_, _27103_, _01538_);
  or (_27208_, _27206_, _27205_);
  and (_27209_, _27208_, _38087_);
  and (_27210_, _27209_, _27204_);
  or (_27211_, _27210_, _27102_);
  and (_40313_, _27211_, _37580_);
  and (_27212_, _38088_, \oc8051_golden_model_1.TCON [6]);
  and (_27213_, _09335_, \oc8051_golden_model_1.TCON [6]);
  and (_27214_, _11709_, _03693_);
  or (_27215_, _27214_, _27213_);
  and (_27216_, _27215_, _02167_);
  nor (_27218_, _11730_, _09335_);
  or (_27219_, _27218_, _27213_);
  or (_27220_, _27219_, _02814_);
  and (_27221_, _03693_, \oc8051_golden_model_1.ACC [6]);
  or (_27222_, _27221_, _27213_);
  and (_27223_, _27222_, _02817_);
  and (_27224_, _02818_, \oc8051_golden_model_1.TCON [6]);
  or (_27225_, _27224_, _02001_);
  or (_27226_, _27225_, _27223_);
  and (_27227_, _27226_, _02024_);
  and (_27229_, _27227_, _27220_);
  and (_27230_, _09343_, \oc8051_golden_model_1.TCON [6]);
  and (_27231_, _11717_, _04315_);
  or (_27232_, _27231_, _27230_);
  and (_27233_, _27232_, _02007_);
  or (_27234_, _27233_, _01999_);
  or (_27235_, _27234_, _27229_);
  nor (_27236_, _03808_, _09335_);
  or (_27237_, _27236_, _27213_);
  or (_27238_, _27237_, _02840_);
  and (_27240_, _27238_, _27235_);
  or (_27241_, _27240_, _02006_);
  or (_27242_, _27222_, _02021_);
  and (_27243_, _27242_, _02025_);
  and (_27244_, _27243_, _27241_);
  and (_27245_, _11715_, _04315_);
  or (_27246_, _27245_, _27230_);
  and (_27247_, _27246_, _01997_);
  or (_27248_, _27247_, _01991_);
  or (_27249_, _27248_, _27244_);
  or (_27251_, _27230_, _11747_);
  and (_27252_, _27251_, _27232_);
  or (_27253_, _27252_, _02861_);
  and (_27254_, _27253_, _02408_);
  and (_27255_, _27254_, _27249_);
  nor (_27256_, _11713_, _09343_);
  or (_27257_, _27256_, _27230_);
  and (_27258_, _27257_, _01875_);
  or (_27259_, _27258_, _05994_);
  or (_27260_, _27259_, _27255_);
  or (_27261_, _27237_, _05249_);
  and (_27262_, _27261_, _27260_);
  or (_27263_, _27262_, _02528_);
  and (_27264_, _04861_, _03693_);
  or (_27265_, _27213_, _02888_);
  or (_27266_, _27265_, _27264_);
  and (_27267_, _27266_, _02043_);
  and (_27268_, _27267_, _27263_);
  nor (_27269_, _11820_, _09335_);
  or (_27270_, _27269_, _27213_);
  and (_27272_, _27270_, _01602_);
  or (_27273_, _27272_, _01869_);
  or (_27274_, _27273_, _27268_);
  and (_27275_, _09920_, _03693_);
  or (_27276_, _27275_, _27213_);
  or (_27277_, _27276_, _01870_);
  and (_27278_, _27277_, _27274_);
  or (_27279_, _27278_, _02079_);
  and (_27280_, _11835_, _03693_);
  or (_27281_, _27213_, _02166_);
  or (_27283_, _27281_, _27280_);
  and (_27284_, _27283_, _02912_);
  and (_27285_, _27284_, _27279_);
  or (_27286_, _27285_, _27216_);
  and (_27287_, _27286_, _02176_);
  or (_27288_, _27213_, _03863_);
  and (_27289_, _27276_, _02072_);
  and (_27290_, _27289_, _27288_);
  or (_27291_, _27290_, _27287_);
  and (_27292_, _27291_, _02907_);
  and (_27294_, _27222_, _02177_);
  and (_27295_, _27294_, _27288_);
  or (_27296_, _27295_, _02071_);
  or (_27297_, _27296_, _27292_);
  nor (_27298_, _11833_, _09335_);
  or (_27299_, _27213_, _04788_);
  or (_27300_, _27299_, _27298_);
  and (_27301_, _27300_, _04793_);
  and (_27302_, _27301_, _27297_);
  nor (_27303_, _11708_, _09335_);
  or (_27305_, _27303_, _27213_);
  and (_27306_, _27305_, _02173_);
  or (_27307_, _27306_, _02201_);
  or (_27308_, _27307_, _27302_);
  or (_27309_, _27219_, _02303_);
  and (_27310_, _27309_, _01887_);
  and (_27311_, _27310_, _27308_);
  and (_27312_, _27246_, _01860_);
  or (_27313_, _27312_, _01537_);
  or (_27314_, _27313_, _27311_);
  and (_27316_, _11887_, _03693_);
  or (_27317_, _27213_, _01538_);
  or (_27318_, _27317_, _27316_);
  and (_27319_, _27318_, _38087_);
  and (_27320_, _27319_, _27314_);
  or (_27321_, _27320_, _27212_);
  and (_40314_, _27321_, _37580_);
  and (_27322_, _38088_, \oc8051_golden_model_1.TH0 [0]);
  and (_27323_, _09439_, \oc8051_golden_model_1.TH0 [0]);
  nor (_27324_, _04106_, _09439_);
  or (_27326_, _27324_, _27323_);
  or (_27327_, _27326_, _02814_);
  and (_27328_, _03691_, \oc8051_golden_model_1.ACC [0]);
  or (_27329_, _27328_, _27323_);
  and (_27330_, _27329_, _02817_);
  and (_27331_, _02818_, \oc8051_golden_model_1.TH0 [0]);
  or (_27332_, _27331_, _02001_);
  or (_27333_, _27332_, _27330_);
  and (_27334_, _27333_, _02840_);
  and (_27335_, _27334_, _27327_);
  and (_27337_, _03691_, _03028_);
  or (_27338_, _27337_, _27323_);
  and (_27339_, _27338_, _01999_);
  or (_27340_, _27339_, _27335_);
  and (_27341_, _27340_, _02021_);
  and (_27342_, _27329_, _02006_);
  or (_27343_, _27342_, _05994_);
  or (_27344_, _27343_, _27341_);
  or (_27345_, _27338_, _05249_);
  and (_27346_, _27345_, _27344_);
  or (_27348_, _27346_, _02528_);
  and (_27349_, _04952_, _03691_);
  or (_27350_, _27323_, _02888_);
  or (_27351_, _27350_, _27349_);
  and (_27352_, _27351_, _27348_);
  or (_27353_, _27352_, _01602_);
  nor (_27354_, _10600_, _09439_);
  or (_27355_, _27354_, _27323_);
  or (_27356_, _27355_, _02043_);
  and (_27357_, _27356_, _01870_);
  and (_27359_, _27357_, _27353_);
  and (_27360_, _03691_, _04562_);
  or (_27361_, _27360_, _27323_);
  and (_27362_, _27361_, _01869_);
  or (_27363_, _27362_, _02079_);
  or (_27364_, _27363_, _27359_);
  and (_27365_, _10614_, _03691_);
  or (_27366_, _27365_, _27323_);
  or (_27367_, _27366_, _02166_);
  and (_27368_, _27367_, _27364_);
  or (_27370_, _27368_, _02167_);
  and (_27371_, _10620_, _03691_);
  or (_27372_, _27323_, _02912_);
  or (_27373_, _27372_, _27371_);
  and (_27374_, _27373_, _02176_);
  and (_27375_, _27374_, _27370_);
  nand (_27376_, _27361_, _02072_);
  nor (_27377_, _27376_, _27324_);
  or (_27378_, _27377_, _27375_);
  and (_27379_, _27378_, _02907_);
  or (_27381_, _27323_, _04106_);
  and (_27382_, _27329_, _02177_);
  and (_27383_, _27382_, _27381_);
  or (_27384_, _27383_, _02071_);
  or (_27385_, _27384_, _27379_);
  nor (_27386_, _10613_, _09439_);
  or (_27387_, _27323_, _04788_);
  or (_27388_, _27387_, _27386_);
  and (_27389_, _27388_, _04793_);
  and (_27390_, _27389_, _27385_);
  nor (_27392_, _10619_, _09439_);
  or (_27393_, _27392_, _27323_);
  and (_27394_, _27393_, _02173_);
  or (_27395_, _27394_, _15577_);
  or (_27396_, _27395_, _27390_);
  or (_27397_, _27326_, _02743_);
  and (_27398_, _27397_, _38087_);
  and (_27399_, _27398_, _27396_);
  or (_27400_, _27399_, _27322_);
  and (_40316_, _27400_, _37580_);
  and (_27402_, _38088_, \oc8051_golden_model_1.TH0 [1]);
  or (_27403_, _03691_, \oc8051_golden_model_1.TH0 [1]);
  and (_27404_, _10698_, _03691_);
  not (_27405_, _27404_);
  and (_27406_, _27405_, _27403_);
  or (_27407_, _27406_, _02814_);
  nand (_27408_, _03691_, _01613_);
  and (_27409_, _27408_, _27403_);
  and (_27410_, _27409_, _02817_);
  and (_27411_, _02818_, \oc8051_golden_model_1.TH0 [1]);
  or (_27413_, _27411_, _02001_);
  or (_27414_, _27413_, _27410_);
  and (_27415_, _27414_, _02840_);
  and (_27416_, _27415_, _27407_);
  nand (_27417_, _03691_, _02811_);
  and (_27418_, _27417_, _27403_);
  and (_27419_, _27418_, _01999_);
  or (_27420_, _27419_, _27416_);
  and (_27421_, _27420_, _02021_);
  and (_27422_, _27409_, _02006_);
  or (_27423_, _27422_, _05994_);
  or (_27424_, _27423_, _27421_);
  or (_27425_, _27418_, _05249_);
  and (_27426_, _27425_, _02888_);
  and (_27427_, _27426_, _27424_);
  or (_27428_, _04907_, _09439_);
  and (_27429_, _27403_, _02528_);
  and (_27430_, _27429_, _27428_);
  or (_27431_, _27430_, _27427_);
  and (_27432_, _27431_, _02043_);
  nand (_27434_, _10802_, _03691_);
  and (_27435_, _27403_, _01602_);
  and (_27436_, _27435_, _27434_);
  or (_27437_, _27436_, _27432_);
  and (_27438_, _27437_, _01870_);
  nand (_27439_, _03691_, _02687_);
  and (_27440_, _27403_, _01869_);
  and (_27441_, _27440_, _27439_);
  or (_27442_, _27441_, _27438_);
  and (_27443_, _27442_, _02166_);
  or (_27445_, _10816_, _09439_);
  and (_27446_, _27403_, _02079_);
  and (_27447_, _27446_, _27445_);
  or (_27448_, _27447_, _27443_);
  and (_27449_, _27448_, _02912_);
  or (_27450_, _10822_, _09439_);
  and (_27451_, _27403_, _02167_);
  and (_27452_, _27451_, _27450_);
  or (_27453_, _27452_, _27449_);
  and (_27454_, _27453_, _02176_);
  or (_27456_, _10692_, _09439_);
  and (_27457_, _27403_, _02072_);
  and (_27458_, _27457_, _27456_);
  or (_27459_, _27458_, _27454_);
  and (_27460_, _27459_, _02907_);
  and (_27461_, _09439_, \oc8051_golden_model_1.TH0 [1]);
  or (_27462_, _27461_, _04058_);
  and (_27463_, _27409_, _02177_);
  and (_27464_, _27463_, _27462_);
  or (_27465_, _27464_, _27460_);
  and (_27467_, _27465_, _02174_);
  or (_27468_, _27408_, _04058_);
  and (_27469_, _27403_, _02173_);
  and (_27470_, _27469_, _27468_);
  or (_27471_, _27470_, _02201_);
  or (_27472_, _27439_, _04058_);
  and (_27473_, _27403_, _02071_);
  and (_27474_, _27473_, _27472_);
  or (_27475_, _27474_, _27471_);
  or (_27476_, _27475_, _27467_);
  or (_27478_, _27406_, _02303_);
  and (_27479_, _27478_, _27476_);
  or (_27480_, _27479_, _01537_);
  or (_27481_, _27461_, _01538_);
  or (_27482_, _27481_, _27404_);
  and (_27483_, _27482_, _38087_);
  and (_27484_, _27483_, _27480_);
  or (_27485_, _27484_, _27402_);
  and (_40317_, _27485_, _37580_);
  and (_27486_, _38088_, \oc8051_golden_model_1.TH0 [2]);
  and (_27488_, _09439_, \oc8051_golden_model_1.TH0 [2]);
  nor (_27489_, _11019_, _09439_);
  or (_27490_, _27489_, _27488_);
  and (_27491_, _27490_, _02173_);
  or (_27492_, _27488_, _04156_);
  and (_27493_, _03691_, _04724_);
  or (_27494_, _27493_, _27488_);
  and (_27495_, _27494_, _02072_);
  and (_27496_, _27495_, _27492_);
  and (_27497_, _11020_, _03691_);
  or (_27499_, _27497_, _27488_);
  and (_27500_, _27499_, _02167_);
  nor (_27501_, _10905_, _09439_);
  or (_27502_, _27501_, _27488_);
  or (_27503_, _27502_, _02814_);
  and (_27504_, _03691_, \oc8051_golden_model_1.ACC [2]);
  or (_27505_, _27504_, _27488_);
  and (_27506_, _27505_, _02817_);
  and (_27507_, _02818_, \oc8051_golden_model_1.TH0 [2]);
  or (_27508_, _27507_, _02001_);
  or (_27510_, _27508_, _27506_);
  and (_27511_, _27510_, _02840_);
  and (_27512_, _27511_, _27503_);
  nor (_27513_, _09439_, _03455_);
  or (_27514_, _27513_, _27488_);
  and (_27515_, _27514_, _01999_);
  or (_27516_, _27515_, _27512_);
  and (_27517_, _27516_, _02021_);
  and (_27518_, _27505_, _02006_);
  or (_27519_, _27518_, _05994_);
  or (_27521_, _27519_, _27517_);
  or (_27522_, _27514_, _05249_);
  and (_27523_, _27522_, _27521_);
  or (_27524_, _27523_, _02528_);
  and (_27525_, _05043_, _03691_);
  or (_27526_, _27488_, _02888_);
  or (_27527_, _27526_, _27525_);
  and (_27528_, _27527_, _27524_);
  or (_27529_, _27528_, _01602_);
  nor (_27530_, _11000_, _09439_);
  or (_27532_, _27488_, _02043_);
  or (_27533_, _27532_, _27530_);
  and (_27534_, _27533_, _01870_);
  and (_27535_, _27534_, _27529_);
  and (_27536_, _27494_, _01869_);
  or (_27537_, _27536_, _02079_);
  or (_27538_, _27537_, _27535_);
  and (_27539_, _11014_, _03691_);
  or (_27540_, _27488_, _02166_);
  or (_27541_, _27540_, _27539_);
  and (_27543_, _27541_, _02912_);
  and (_27544_, _27543_, _27538_);
  or (_27545_, _27544_, _27500_);
  and (_27546_, _27545_, _02176_);
  or (_27547_, _27546_, _27496_);
  and (_27548_, _27547_, _02907_);
  and (_27549_, _27505_, _02177_);
  and (_27550_, _27549_, _27492_);
  or (_27551_, _27550_, _02071_);
  or (_27552_, _27551_, _27548_);
  nor (_27554_, _11013_, _09439_);
  or (_27555_, _27488_, _04788_);
  or (_27556_, _27555_, _27554_);
  and (_27557_, _27556_, _04793_);
  and (_27558_, _27557_, _27552_);
  or (_27559_, _27558_, _27491_);
  and (_27560_, _27559_, _02303_);
  and (_27561_, _27502_, _02201_);
  or (_27562_, _27561_, _01537_);
  or (_27563_, _27562_, _27560_);
  and (_27565_, _11072_, _03691_);
  or (_27566_, _27488_, _01538_);
  or (_27567_, _27566_, _27565_);
  and (_27568_, _27567_, _38087_);
  and (_27569_, _27568_, _27563_);
  or (_27570_, _27569_, _27486_);
  and (_40318_, _27570_, _37580_);
  or (_27571_, _38087_, \oc8051_golden_model_1.TH0 [3]);
  and (_27572_, _27571_, _37580_);
  and (_27573_, _09439_, \oc8051_golden_model_1.TH0 [3]);
  or (_27575_, _27573_, _04014_);
  and (_27576_, _03691_, _04678_);
  or (_27577_, _27576_, _27573_);
  and (_27578_, _27577_, _02072_);
  and (_27579_, _27578_, _27575_);
  and (_27580_, _11094_, _03691_);
  or (_27581_, _27580_, _27573_);
  and (_27582_, _27581_, _02167_);
  nor (_27583_, _11101_, _09439_);
  or (_27584_, _27583_, _27573_);
  or (_27586_, _27584_, _02814_);
  and (_27587_, _03691_, \oc8051_golden_model_1.ACC [3]);
  or (_27588_, _27587_, _27573_);
  and (_27589_, _27588_, _02817_);
  and (_27590_, _02818_, \oc8051_golden_model_1.TH0 [3]);
  or (_27591_, _27590_, _02001_);
  or (_27592_, _27591_, _27589_);
  and (_27593_, _27592_, _02840_);
  and (_27594_, _27593_, _27586_);
  nor (_27595_, _09439_, _03268_);
  or (_27596_, _27595_, _27573_);
  and (_27597_, _27596_, _01999_);
  or (_27598_, _27597_, _27594_);
  and (_27599_, _27598_, _02021_);
  and (_27600_, _27588_, _02006_);
  or (_27601_, _27600_, _05994_);
  or (_27602_, _27601_, _27599_);
  or (_27603_, _27596_, _05249_);
  and (_27604_, _27603_, _27602_);
  or (_27605_, _27604_, _02528_);
  and (_27607_, _04998_, _03691_);
  or (_27608_, _27573_, _02888_);
  or (_27609_, _27608_, _27607_);
  and (_27610_, _27609_, _02043_);
  and (_27611_, _27610_, _27605_);
  nor (_27612_, _11206_, _09439_);
  or (_27613_, _27612_, _27573_);
  and (_27614_, _27613_, _01602_);
  or (_27615_, _27614_, _01869_);
  or (_27616_, _27615_, _27611_);
  or (_27618_, _27577_, _01870_);
  and (_27619_, _27618_, _27616_);
  or (_27620_, _27619_, _02079_);
  and (_27621_, _11222_, _03691_);
  or (_27622_, _27573_, _02166_);
  or (_27623_, _27622_, _27621_);
  and (_27624_, _27623_, _02912_);
  and (_27625_, _27624_, _27620_);
  or (_27626_, _27625_, _27582_);
  and (_27627_, _27626_, _02176_);
  or (_27629_, _27627_, _27579_);
  and (_27630_, _27629_, _02907_);
  and (_27631_, _27588_, _02177_);
  and (_27632_, _27631_, _27575_);
  or (_27633_, _27632_, _02071_);
  or (_27634_, _27633_, _27630_);
  nor (_27635_, _11220_, _09439_);
  or (_27636_, _27573_, _04788_);
  or (_27637_, _27636_, _27635_);
  and (_27638_, _27637_, _04793_);
  and (_27640_, _27638_, _27634_);
  nor (_27641_, _11093_, _09439_);
  or (_27642_, _27641_, _27573_);
  and (_27643_, _27642_, _02173_);
  or (_27644_, _27643_, _02201_);
  or (_27645_, _27644_, _27640_);
  or (_27646_, _27584_, _02303_);
  and (_27647_, _27646_, _01538_);
  and (_27648_, _27647_, _27645_);
  and (_27649_, _11273_, _03691_);
  or (_27651_, _27649_, _27573_);
  and (_27652_, _27651_, _01537_);
  or (_27653_, _27652_, _38088_);
  or (_27654_, _27653_, _27648_);
  and (_40319_, _27654_, _27572_);
  or (_27655_, _38087_, \oc8051_golden_model_1.TH0 [4]);
  and (_27656_, _27655_, _37580_);
  and (_27657_, _09439_, \oc8051_golden_model_1.TH0 [4]);
  and (_27658_, _11431_, _03691_);
  or (_27659_, _27658_, _27657_);
  and (_27661_, _27659_, _02167_);
  nor (_27662_, _11317_, _09439_);
  or (_27663_, _27662_, _27657_);
  or (_27664_, _27663_, _02814_);
  and (_27665_, _03691_, \oc8051_golden_model_1.ACC [4]);
  or (_27666_, _27665_, _27657_);
  and (_27667_, _27666_, _02817_);
  and (_27668_, _02818_, \oc8051_golden_model_1.TH0 [4]);
  or (_27669_, _27668_, _02001_);
  or (_27670_, _27669_, _27667_);
  and (_27672_, _27670_, _02840_);
  and (_27673_, _27672_, _27664_);
  nor (_27674_, _04211_, _09439_);
  or (_27675_, _27674_, _27657_);
  and (_27676_, _27675_, _01999_);
  or (_27677_, _27676_, _27673_);
  and (_27678_, _27677_, _02021_);
  and (_27679_, _27666_, _02006_);
  or (_27680_, _27679_, _05994_);
  or (_27681_, _27680_, _27678_);
  or (_27683_, _27675_, _05249_);
  and (_27684_, _27683_, _27681_);
  or (_27685_, _27684_, _02528_);
  and (_27686_, _05135_, _03691_);
  or (_27687_, _27657_, _02888_);
  or (_27688_, _27687_, _27686_);
  and (_27689_, _27688_, _02043_);
  and (_27690_, _27689_, _27685_);
  nor (_27691_, _11411_, _09439_);
  or (_27692_, _27691_, _27657_);
  and (_27694_, _27692_, _01602_);
  or (_27695_, _27694_, _01869_);
  or (_27696_, _27695_, _27690_);
  and (_27697_, _04694_, _03691_);
  or (_27698_, _27697_, _27657_);
  or (_27699_, _27698_, _01870_);
  and (_27700_, _27699_, _27696_);
  or (_27701_, _27700_, _02079_);
  and (_27702_, _11425_, _03691_);
  or (_27703_, _27657_, _02166_);
  or (_27705_, _27703_, _27702_);
  and (_27706_, _27705_, _02912_);
  and (_27707_, _27706_, _27701_);
  or (_27708_, _27707_, _27661_);
  and (_27709_, _27708_, _02176_);
  or (_27710_, _27657_, _04258_);
  and (_27711_, _27698_, _02072_);
  and (_27712_, _27711_, _27710_);
  or (_27713_, _27712_, _27709_);
  and (_27714_, _27713_, _02907_);
  and (_27716_, _27666_, _02177_);
  and (_27717_, _27716_, _27710_);
  or (_27718_, _27717_, _02071_);
  or (_27719_, _27718_, _27714_);
  nor (_27720_, _11424_, _09439_);
  or (_27721_, _27657_, _04788_);
  or (_27722_, _27721_, _27720_);
  and (_27723_, _27722_, _04793_);
  and (_27724_, _27723_, _27719_);
  nor (_27725_, _11430_, _09439_);
  or (_27727_, _27725_, _27657_);
  and (_27728_, _27727_, _02173_);
  or (_27729_, _27728_, _02201_);
  or (_27730_, _27729_, _27724_);
  or (_27731_, _27663_, _02303_);
  and (_27732_, _27731_, _01538_);
  and (_27733_, _27732_, _27730_);
  and (_27734_, _11487_, _03691_);
  or (_27735_, _27734_, _27657_);
  and (_27736_, _27735_, _01537_);
  or (_27738_, _27736_, _38088_);
  or (_27739_, _27738_, _27733_);
  and (_40320_, _27739_, _27656_);
  or (_27740_, _38087_, \oc8051_golden_model_1.TH0 [5]);
  and (_27741_, _27740_, _37580_);
  and (_27742_, _09439_, \oc8051_golden_model_1.TH0 [5]);
  and (_27743_, _11635_, _03691_);
  or (_27744_, _27743_, _27742_);
  and (_27745_, _27744_, _02167_);
  nor (_27746_, _11525_, _09439_);
  or (_27748_, _27746_, _27742_);
  or (_27749_, _27748_, _02814_);
  and (_27750_, _03691_, \oc8051_golden_model_1.ACC [5]);
  or (_27751_, _27750_, _27742_);
  and (_27752_, _27751_, _02817_);
  and (_27753_, _02818_, \oc8051_golden_model_1.TH0 [5]);
  or (_27754_, _27753_, _02001_);
  or (_27755_, _27754_, _27752_);
  and (_27756_, _27755_, _02840_);
  and (_27757_, _27756_, _27749_);
  nor (_27759_, _03916_, _09439_);
  or (_27760_, _27759_, _27742_);
  and (_27761_, _27760_, _01999_);
  or (_27762_, _27761_, _27757_);
  and (_27763_, _27762_, _02021_);
  and (_27764_, _27751_, _02006_);
  or (_27765_, _27764_, _05994_);
  or (_27766_, _27765_, _27763_);
  or (_27767_, _27760_, _05249_);
  and (_27768_, _27767_, _27766_);
  or (_27770_, _27768_, _02528_);
  and (_27771_, _05090_, _03691_);
  or (_27772_, _27742_, _02888_);
  or (_27773_, _27772_, _27771_);
  and (_27774_, _27773_, _02043_);
  and (_27775_, _27774_, _27770_);
  nor (_27776_, _11615_, _09439_);
  or (_27777_, _27776_, _27742_);
  and (_27778_, _27777_, _01602_);
  or (_27779_, _27778_, _01869_);
  or (_27781_, _27779_, _27775_);
  and (_27782_, _04672_, _03691_);
  or (_27783_, _27782_, _27742_);
  or (_27784_, _27783_, _01870_);
  and (_27785_, _27784_, _27781_);
  or (_27786_, _27785_, _02079_);
  and (_27787_, _11629_, _03691_);
  or (_27788_, _27742_, _02166_);
  or (_27789_, _27788_, _27787_);
  and (_27790_, _27789_, _02912_);
  and (_27792_, _27790_, _27786_);
  or (_27793_, _27792_, _27745_);
  and (_27794_, _27793_, _02176_);
  or (_27795_, _27742_, _03965_);
  and (_27796_, _27783_, _02072_);
  and (_27797_, _27796_, _27795_);
  or (_27798_, _27797_, _27794_);
  and (_27799_, _27798_, _02907_);
  and (_27800_, _27751_, _02177_);
  and (_27801_, _27800_, _27795_);
  or (_27803_, _27801_, _02071_);
  or (_27804_, _27803_, _27799_);
  nor (_27805_, _11628_, _09439_);
  or (_27806_, _27742_, _04788_);
  or (_27807_, _27806_, _27805_);
  and (_27808_, _27807_, _04793_);
  and (_27809_, _27808_, _27804_);
  nor (_27810_, _11634_, _09439_);
  or (_27811_, _27810_, _27742_);
  and (_27812_, _27811_, _02173_);
  or (_27813_, _27812_, _02201_);
  or (_27814_, _27813_, _27809_);
  or (_27815_, _27748_, _02303_);
  and (_27816_, _27815_, _01538_);
  and (_27817_, _27816_, _27814_);
  and (_27818_, _11685_, _03691_);
  or (_27819_, _27818_, _27742_);
  and (_27820_, _27819_, _01537_);
  or (_27821_, _27820_, _38088_);
  or (_27822_, _27821_, _27817_);
  and (_40321_, _27822_, _27741_);
  or (_27824_, _38087_, \oc8051_golden_model_1.TH0 [6]);
  and (_27825_, _27824_, _37580_);
  and (_27826_, _09439_, \oc8051_golden_model_1.TH0 [6]);
  and (_27827_, _11709_, _03691_);
  or (_27828_, _27827_, _27826_);
  and (_27829_, _27828_, _02167_);
  nor (_27830_, _11730_, _09439_);
  or (_27831_, _27830_, _27826_);
  or (_27832_, _27831_, _02814_);
  and (_27834_, _03691_, \oc8051_golden_model_1.ACC [6]);
  or (_27835_, _27834_, _27826_);
  and (_27836_, _27835_, _02817_);
  and (_27837_, _02818_, \oc8051_golden_model_1.TH0 [6]);
  or (_27838_, _27837_, _02001_);
  or (_27839_, _27838_, _27836_);
  and (_27840_, _27839_, _02840_);
  and (_27841_, _27840_, _27832_);
  nor (_27842_, _03808_, _09439_);
  or (_27843_, _27842_, _27826_);
  and (_27845_, _27843_, _01999_);
  or (_27846_, _27845_, _27841_);
  and (_27847_, _27846_, _02021_);
  and (_27848_, _27835_, _02006_);
  or (_27849_, _27848_, _05994_);
  or (_27850_, _27849_, _27847_);
  or (_27851_, _27843_, _05249_);
  and (_27852_, _27851_, _27850_);
  or (_27853_, _27852_, _02528_);
  and (_27854_, _04861_, _03691_);
  or (_27856_, _27826_, _02888_);
  or (_27857_, _27856_, _27854_);
  and (_27858_, _27857_, _02043_);
  and (_27859_, _27858_, _27853_);
  nor (_27860_, _11820_, _09439_);
  or (_27861_, _27860_, _27826_);
  and (_27862_, _27861_, _01602_);
  or (_27863_, _27862_, _01869_);
  or (_27864_, _27863_, _27859_);
  and (_27865_, _09920_, _03691_);
  or (_27867_, _27865_, _27826_);
  or (_27868_, _27867_, _01870_);
  and (_27869_, _27868_, _27864_);
  or (_27870_, _27869_, _02079_);
  and (_27871_, _11835_, _03691_);
  or (_27872_, _27826_, _02166_);
  or (_27873_, _27872_, _27871_);
  and (_27874_, _27873_, _02912_);
  and (_27875_, _27874_, _27870_);
  or (_27876_, _27875_, _27829_);
  and (_27878_, _27876_, _02176_);
  or (_27879_, _27826_, _03863_);
  and (_27880_, _27867_, _02072_);
  and (_27881_, _27880_, _27879_);
  or (_27882_, _27881_, _27878_);
  and (_27883_, _27882_, _02907_);
  and (_27884_, _27835_, _02177_);
  and (_27885_, _27884_, _27879_);
  or (_27886_, _27885_, _02071_);
  or (_27887_, _27886_, _27883_);
  nor (_27889_, _11833_, _09439_);
  or (_27890_, _27826_, _04788_);
  or (_27891_, _27890_, _27889_);
  and (_27892_, _27891_, _04793_);
  and (_27893_, _27892_, _27887_);
  nor (_27894_, _11708_, _09439_);
  or (_27895_, _27894_, _27826_);
  and (_27896_, _27895_, _02173_);
  or (_27897_, _27896_, _02201_);
  or (_27898_, _27897_, _27893_);
  or (_27900_, _27831_, _02303_);
  and (_27901_, _27900_, _01538_);
  and (_27902_, _27901_, _27898_);
  and (_27903_, _11887_, _03691_);
  or (_27904_, _27903_, _27826_);
  and (_27905_, _27904_, _01537_);
  or (_27906_, _27905_, _38088_);
  or (_27907_, _27906_, _27902_);
  and (_40323_, _27907_, _27825_);
  and (_27908_, _38088_, \oc8051_golden_model_1.TH1 [0]);
  and (_27910_, _09517_, \oc8051_golden_model_1.TH1 [0]);
  and (_27911_, _03722_, _03028_);
  or (_27912_, _27911_, _27910_);
  or (_27913_, _27912_, _05249_);
  nor (_27914_, _04106_, _09517_);
  or (_27915_, _27914_, _27910_);
  or (_27916_, _27915_, _02814_);
  and (_27917_, _03722_, \oc8051_golden_model_1.ACC [0]);
  or (_27918_, _27917_, _27910_);
  and (_27919_, _27918_, _02817_);
  and (_27921_, _02818_, \oc8051_golden_model_1.TH1 [0]);
  or (_27922_, _27921_, _02001_);
  or (_27923_, _27922_, _27919_);
  and (_27924_, _27923_, _02840_);
  and (_27925_, _27924_, _27916_);
  and (_27926_, _27912_, _01999_);
  or (_27927_, _27926_, _27925_);
  and (_27928_, _27927_, _02021_);
  and (_27929_, _27918_, _02006_);
  or (_27930_, _27929_, _05994_);
  or (_27932_, _27930_, _27928_);
  and (_27933_, _27932_, _27913_);
  or (_27934_, _27933_, _02528_);
  and (_27935_, _04952_, _03722_);
  or (_27936_, _27910_, _02888_);
  or (_27937_, _27936_, _27935_);
  and (_27938_, _27937_, _27934_);
  or (_27939_, _27938_, _01602_);
  nor (_27940_, _10600_, _09517_);
  or (_27941_, _27940_, _27910_);
  or (_27943_, _27941_, _02043_);
  and (_27944_, _27943_, _01870_);
  and (_27945_, _27944_, _27939_);
  and (_27946_, _03722_, _04562_);
  or (_27947_, _27946_, _27910_);
  and (_27948_, _27947_, _01869_);
  or (_27949_, _27948_, _02079_);
  or (_27950_, _27949_, _27945_);
  and (_27951_, _10614_, _03722_);
  or (_27952_, _27951_, _27910_);
  or (_27954_, _27952_, _02166_);
  and (_27955_, _27954_, _27950_);
  or (_27956_, _27955_, _02167_);
  and (_27957_, _10620_, _03722_);
  or (_27958_, _27910_, _02912_);
  or (_27959_, _27958_, _27957_);
  and (_27960_, _27959_, _02176_);
  and (_27961_, _27960_, _27956_);
  nand (_27962_, _27947_, _02072_);
  nor (_27963_, _27962_, _27914_);
  or (_27965_, _27963_, _27961_);
  and (_27966_, _27965_, _02907_);
  or (_27967_, _27910_, _04106_);
  and (_27968_, _27918_, _02177_);
  and (_27969_, _27968_, _27967_);
  or (_27970_, _27969_, _02071_);
  or (_27971_, _27970_, _27966_);
  nor (_27972_, _10613_, _09517_);
  or (_27973_, _27910_, _04788_);
  or (_27974_, _27973_, _27972_);
  and (_27976_, _27974_, _04793_);
  and (_27977_, _27976_, _27971_);
  nor (_27978_, _10619_, _09517_);
  or (_27979_, _27978_, _27910_);
  and (_27980_, _27979_, _02173_);
  or (_27981_, _27980_, _15577_);
  or (_27982_, _27981_, _27977_);
  or (_27983_, _27915_, _02743_);
  and (_27984_, _27983_, _38087_);
  and (_27985_, _27984_, _27982_);
  or (_27987_, _27985_, _27908_);
  and (_40324_, _27987_, _37580_);
  and (_27988_, _38088_, \oc8051_golden_model_1.TH1 [1]);
  or (_27989_, _03722_, \oc8051_golden_model_1.TH1 [1]);
  and (_27990_, _10698_, _03722_);
  not (_27991_, _27990_);
  and (_27992_, _27991_, _27989_);
  or (_27993_, _27992_, _02814_);
  nand (_27994_, _03722_, _01613_);
  and (_27995_, _27994_, _27989_);
  and (_27997_, _27995_, _02817_);
  and (_27998_, _02818_, \oc8051_golden_model_1.TH1 [1]);
  or (_27999_, _27998_, _02001_);
  or (_28000_, _27999_, _27997_);
  and (_28001_, _28000_, _02840_);
  and (_28002_, _28001_, _27993_);
  nand (_28003_, _03722_, _02811_);
  and (_28004_, _28003_, _27989_);
  and (_28005_, _28004_, _01999_);
  or (_28006_, _28005_, _28002_);
  and (_28008_, _28006_, _02021_);
  and (_28009_, _27995_, _02006_);
  or (_28010_, _28009_, _05994_);
  or (_28011_, _28010_, _28008_);
  or (_28012_, _28004_, _05249_);
  and (_28013_, _28012_, _02888_);
  and (_28014_, _28013_, _28011_);
  or (_28015_, _04907_, _09517_);
  and (_28016_, _27989_, _02528_);
  and (_28017_, _28016_, _28015_);
  or (_28019_, _28017_, _28014_);
  and (_28020_, _28019_, _02043_);
  nand (_28021_, _10802_, _03722_);
  and (_28022_, _27989_, _01602_);
  and (_28023_, _28022_, _28021_);
  or (_28024_, _28023_, _28020_);
  and (_28025_, _28024_, _01870_);
  nand (_28026_, _03722_, _02687_);
  and (_28027_, _27989_, _01869_);
  and (_28028_, _28027_, _28026_);
  or (_28030_, _28028_, _28025_);
  and (_28031_, _28030_, _02166_);
  or (_28032_, _10816_, _09517_);
  and (_28033_, _27989_, _02079_);
  and (_28034_, _28033_, _28032_);
  or (_28035_, _28034_, _28031_);
  and (_28036_, _28035_, _02912_);
  or (_28037_, _10822_, _09517_);
  and (_28038_, _27989_, _02167_);
  and (_28039_, _28038_, _28037_);
  or (_28040_, _28039_, _28036_);
  and (_28041_, _28040_, _02176_);
  or (_28042_, _10692_, _09517_);
  and (_28043_, _27989_, _02072_);
  and (_28044_, _28043_, _28042_);
  or (_28045_, _28044_, _28041_);
  and (_28046_, _28045_, _02907_);
  and (_28047_, _09517_, \oc8051_golden_model_1.TH1 [1]);
  or (_28048_, _28047_, _04058_);
  and (_28049_, _27995_, _02177_);
  and (_28051_, _28049_, _28048_);
  or (_28052_, _28051_, _28046_);
  and (_28053_, _28052_, _02174_);
  or (_28054_, _27994_, _04058_);
  and (_28055_, _27989_, _02173_);
  and (_28056_, _28055_, _28054_);
  or (_28057_, _28056_, _02201_);
  or (_28058_, _28026_, _04058_);
  and (_28059_, _27989_, _02071_);
  and (_28060_, _28059_, _28058_);
  or (_28062_, _28060_, _28057_);
  or (_28063_, _28062_, _28053_);
  or (_28064_, _27992_, _02303_);
  and (_28065_, _28064_, _28063_);
  or (_28066_, _28065_, _01537_);
  or (_28067_, _28047_, _01538_);
  or (_28068_, _28067_, _27990_);
  and (_28069_, _28068_, _38087_);
  and (_28070_, _28069_, _28066_);
  or (_28071_, _28070_, _27988_);
  and (_40325_, _28071_, _37580_);
  and (_28073_, _38088_, \oc8051_golden_model_1.TH1 [2]);
  and (_28074_, _09517_, \oc8051_golden_model_1.TH1 [2]);
  nor (_28075_, _11019_, _09517_);
  or (_28076_, _28075_, _28074_);
  and (_28077_, _28076_, _02173_);
  and (_28078_, _11020_, _03722_);
  or (_28079_, _28078_, _28074_);
  and (_28080_, _28079_, _02167_);
  nor (_28081_, _10905_, _09517_);
  or (_28083_, _28081_, _28074_);
  or (_28084_, _28083_, _02814_);
  and (_28085_, _03722_, \oc8051_golden_model_1.ACC [2]);
  or (_28086_, _28085_, _28074_);
  and (_28087_, _28086_, _02817_);
  and (_28088_, _02818_, \oc8051_golden_model_1.TH1 [2]);
  or (_28089_, _28088_, _02001_);
  or (_28090_, _28089_, _28087_);
  and (_28091_, _28090_, _02840_);
  and (_28092_, _28091_, _28084_);
  nor (_28094_, _09517_, _03455_);
  or (_28095_, _28094_, _28074_);
  and (_28096_, _28095_, _01999_);
  or (_28097_, _28096_, _28092_);
  and (_28098_, _28097_, _02021_);
  and (_28099_, _28086_, _02006_);
  or (_28100_, _28099_, _05994_);
  or (_28101_, _28100_, _28098_);
  or (_28102_, _28095_, _05249_);
  and (_28103_, _28102_, _28101_);
  or (_28105_, _28103_, _02528_);
  and (_28106_, _05043_, _03722_);
  or (_28107_, _28074_, _02888_);
  or (_28108_, _28107_, _28106_);
  and (_28109_, _28108_, _28105_);
  or (_28110_, _28109_, _01602_);
  nor (_28111_, _11000_, _09517_);
  or (_28112_, _28074_, _02043_);
  or (_28113_, _28112_, _28111_);
  and (_28114_, _28113_, _01870_);
  and (_28116_, _28114_, _28110_);
  and (_28117_, _03722_, _04724_);
  or (_28118_, _28117_, _28074_);
  and (_28119_, _28118_, _01869_);
  or (_28120_, _28119_, _02079_);
  or (_28121_, _28120_, _28116_);
  and (_28122_, _11014_, _03722_);
  or (_28123_, _28074_, _02166_);
  or (_28124_, _28123_, _28122_);
  and (_28125_, _28124_, _02912_);
  and (_28127_, _28125_, _28121_);
  or (_28128_, _28127_, _28080_);
  and (_28129_, _28128_, _02176_);
  or (_28130_, _28074_, _04156_);
  and (_28131_, _28118_, _02072_);
  and (_28132_, _28131_, _28130_);
  or (_28133_, _28132_, _28129_);
  and (_28134_, _28133_, _02907_);
  and (_28135_, _28086_, _02177_);
  and (_28136_, _28135_, _28130_);
  or (_28138_, _28136_, _02071_);
  or (_28139_, _28138_, _28134_);
  nor (_28140_, _11013_, _09517_);
  or (_28141_, _28074_, _04788_);
  or (_28142_, _28141_, _28140_);
  and (_28143_, _28142_, _04793_);
  and (_28144_, _28143_, _28139_);
  or (_28145_, _28144_, _28077_);
  and (_28146_, _28145_, _02303_);
  and (_28147_, _28083_, _02201_);
  or (_28149_, _28147_, _01537_);
  or (_28150_, _28149_, _28146_);
  and (_28151_, _11072_, _03722_);
  or (_28152_, _28074_, _01538_);
  or (_28153_, _28152_, _28151_);
  and (_28154_, _28153_, _38087_);
  and (_28155_, _28154_, _28150_);
  or (_28156_, _28155_, _28073_);
  and (_40326_, _28156_, _37580_);
  or (_28157_, _38087_, \oc8051_golden_model_1.TH1 [3]);
  and (_28159_, _28157_, _37580_);
  and (_28160_, _09517_, \oc8051_golden_model_1.TH1 [3]);
  and (_28161_, _11094_, _03722_);
  or (_28162_, _28161_, _28160_);
  and (_28163_, _28162_, _02167_);
  nor (_28164_, _11101_, _09517_);
  or (_28165_, _28164_, _28160_);
  or (_28166_, _28165_, _02814_);
  and (_28167_, _03722_, \oc8051_golden_model_1.ACC [3]);
  or (_28168_, _28167_, _28160_);
  and (_28169_, _28168_, _02817_);
  and (_28170_, _02818_, \oc8051_golden_model_1.TH1 [3]);
  or (_28171_, _28170_, _02001_);
  or (_28172_, _28171_, _28169_);
  and (_28173_, _28172_, _02840_);
  and (_28174_, _28173_, _28166_);
  nor (_28175_, _09517_, _03268_);
  or (_28176_, _28175_, _28160_);
  and (_28177_, _28176_, _01999_);
  or (_28178_, _28177_, _28174_);
  and (_28180_, _28178_, _02021_);
  and (_28181_, _28168_, _02006_);
  or (_28182_, _28181_, _05994_);
  or (_28183_, _28182_, _28180_);
  or (_28184_, _28176_, _05249_);
  and (_28185_, _28184_, _28183_);
  or (_28186_, _28185_, _02528_);
  and (_28187_, _04998_, _03722_);
  or (_28188_, _28160_, _02888_);
  or (_28189_, _28188_, _28187_);
  and (_28191_, _28189_, _02043_);
  and (_28192_, _28191_, _28186_);
  nor (_28193_, _11206_, _09517_);
  or (_28194_, _28193_, _28160_);
  and (_28195_, _28194_, _01602_);
  or (_28196_, _28195_, _01869_);
  or (_28197_, _28196_, _28192_);
  and (_28198_, _03722_, _04678_);
  or (_28199_, _28198_, _28160_);
  or (_28200_, _28199_, _01870_);
  and (_28202_, _28200_, _28197_);
  or (_28203_, _28202_, _02079_);
  and (_28204_, _11222_, _03722_);
  or (_28205_, _28160_, _02166_);
  or (_28206_, _28205_, _28204_);
  and (_28207_, _28206_, _02912_);
  and (_28208_, _28207_, _28203_);
  or (_28209_, _28208_, _28163_);
  and (_28210_, _28209_, _02176_);
  or (_28211_, _28160_, _04014_);
  and (_28213_, _28199_, _02072_);
  and (_28214_, _28213_, _28211_);
  or (_28215_, _28214_, _28210_);
  and (_28216_, _28215_, _02907_);
  and (_28217_, _28168_, _02177_);
  and (_28218_, _28217_, _28211_);
  or (_28219_, _28218_, _02071_);
  or (_28220_, _28219_, _28216_);
  nor (_28221_, _11220_, _09517_);
  or (_28222_, _28160_, _04788_);
  or (_28224_, _28222_, _28221_);
  and (_28225_, _28224_, _04793_);
  and (_28226_, _28225_, _28220_);
  nor (_28227_, _11093_, _09517_);
  or (_28228_, _28227_, _28160_);
  and (_28229_, _28228_, _02173_);
  or (_28230_, _28229_, _02201_);
  or (_28231_, _28230_, _28226_);
  or (_28232_, _28165_, _02303_);
  and (_28233_, _28232_, _01538_);
  and (_28235_, _28233_, _28231_);
  and (_28236_, _11273_, _03722_);
  or (_28237_, _28236_, _28160_);
  and (_28238_, _28237_, _01537_);
  or (_28239_, _28238_, _38088_);
  or (_28240_, _28239_, _28235_);
  and (_40327_, _28240_, _28159_);
  or (_28241_, _38087_, \oc8051_golden_model_1.TH1 [4]);
  and (_28242_, _28241_, _37580_);
  and (_28243_, _09517_, \oc8051_golden_model_1.TH1 [4]);
  or (_28245_, _28243_, _04258_);
  and (_28246_, _04694_, _03722_);
  or (_28247_, _28246_, _28243_);
  and (_28248_, _28247_, _02072_);
  and (_28249_, _28248_, _28245_);
  and (_28250_, _11431_, _03722_);
  or (_28251_, _28250_, _28243_);
  and (_28252_, _28251_, _02167_);
  nor (_28253_, _11317_, _09517_);
  or (_28254_, _28253_, _28243_);
  or (_28256_, _28254_, _02814_);
  and (_28257_, _03722_, \oc8051_golden_model_1.ACC [4]);
  or (_28258_, _28257_, _28243_);
  and (_28259_, _28258_, _02817_);
  and (_28260_, _02818_, \oc8051_golden_model_1.TH1 [4]);
  or (_28261_, _28260_, _02001_);
  or (_28262_, _28261_, _28259_);
  and (_28263_, _28262_, _02840_);
  and (_28264_, _28263_, _28256_);
  nor (_28265_, _04211_, _09517_);
  or (_28267_, _28265_, _28243_);
  and (_28268_, _28267_, _01999_);
  or (_28269_, _28268_, _28264_);
  and (_28270_, _28269_, _02021_);
  and (_28271_, _28258_, _02006_);
  or (_28272_, _28271_, _05994_);
  or (_28273_, _28272_, _28270_);
  or (_28274_, _28267_, _05249_);
  and (_28275_, _28274_, _28273_);
  or (_28276_, _28275_, _02528_);
  and (_28278_, _05135_, _03722_);
  or (_28279_, _28243_, _02888_);
  or (_28280_, _28279_, _28278_);
  and (_28281_, _28280_, _02043_);
  and (_28282_, _28281_, _28276_);
  nor (_28283_, _11411_, _09517_);
  or (_28284_, _28283_, _28243_);
  and (_28285_, _28284_, _01602_);
  or (_28286_, _28285_, _01869_);
  or (_28287_, _28286_, _28282_);
  or (_28289_, _28247_, _01870_);
  and (_28290_, _28289_, _28287_);
  or (_28291_, _28290_, _02079_);
  and (_28292_, _11425_, _03722_);
  or (_28293_, _28243_, _02166_);
  or (_28294_, _28293_, _28292_);
  and (_28295_, _28294_, _02912_);
  and (_28296_, _28295_, _28291_);
  or (_28297_, _28296_, _28252_);
  and (_28298_, _28297_, _02176_);
  or (_28299_, _28298_, _28249_);
  and (_28300_, _28299_, _02907_);
  and (_28301_, _28258_, _02177_);
  and (_28302_, _28301_, _28245_);
  or (_28303_, _28302_, _02071_);
  or (_28304_, _28303_, _28300_);
  nor (_28305_, _11424_, _09517_);
  or (_28306_, _28243_, _04788_);
  or (_28307_, _28306_, _28305_);
  and (_28308_, _28307_, _04793_);
  and (_28310_, _28308_, _28304_);
  nor (_28311_, _11430_, _09517_);
  or (_28312_, _28311_, _28243_);
  and (_28313_, _28312_, _02173_);
  or (_28314_, _28313_, _02201_);
  or (_28315_, _28314_, _28310_);
  or (_28316_, _28254_, _02303_);
  and (_28317_, _28316_, _01538_);
  and (_28318_, _28317_, _28315_);
  and (_28319_, _11487_, _03722_);
  or (_28321_, _28319_, _28243_);
  and (_28322_, _28321_, _01537_);
  or (_28323_, _28322_, _38088_);
  or (_28324_, _28323_, _28318_);
  and (_40328_, _28324_, _28242_);
  or (_28325_, _38087_, \oc8051_golden_model_1.TH1 [5]);
  and (_28326_, _28325_, _37580_);
  and (_28327_, _09517_, \oc8051_golden_model_1.TH1 [5]);
  and (_28328_, _11635_, _03722_);
  or (_28329_, _28328_, _28327_);
  and (_28331_, _28329_, _02167_);
  nor (_28332_, _11525_, _09517_);
  or (_28333_, _28332_, _28327_);
  or (_28334_, _28333_, _02814_);
  and (_28335_, _03722_, \oc8051_golden_model_1.ACC [5]);
  or (_28336_, _28335_, _28327_);
  and (_28337_, _28336_, _02817_);
  and (_28338_, _02818_, \oc8051_golden_model_1.TH1 [5]);
  or (_28339_, _28338_, _02001_);
  or (_28340_, _28339_, _28337_);
  and (_28342_, _28340_, _02840_);
  and (_28343_, _28342_, _28334_);
  nor (_28344_, _03916_, _09517_);
  or (_28345_, _28344_, _28327_);
  and (_28346_, _28345_, _01999_);
  or (_28347_, _28346_, _28343_);
  and (_28348_, _28347_, _02021_);
  and (_28349_, _28336_, _02006_);
  or (_28350_, _28349_, _05994_);
  or (_28351_, _28350_, _28348_);
  or (_28353_, _28345_, _05249_);
  and (_28354_, _28353_, _28351_);
  or (_28355_, _28354_, _02528_);
  and (_28356_, _05090_, _03722_);
  or (_28357_, _28327_, _02888_);
  or (_28358_, _28357_, _28356_);
  and (_28359_, _28358_, _02043_);
  and (_28360_, _28359_, _28355_);
  nor (_28361_, _11615_, _09517_);
  or (_28362_, _28361_, _28327_);
  and (_28364_, _28362_, _01602_);
  or (_28365_, _28364_, _01869_);
  or (_28366_, _28365_, _28360_);
  and (_28367_, _04672_, _03722_);
  or (_28368_, _28367_, _28327_);
  or (_28369_, _28368_, _01870_);
  and (_28370_, _28369_, _28366_);
  or (_28371_, _28370_, _02079_);
  and (_28372_, _11629_, _03722_);
  or (_28373_, _28327_, _02166_);
  or (_28375_, _28373_, _28372_);
  and (_28376_, _28375_, _02912_);
  and (_28377_, _28376_, _28371_);
  or (_28378_, _28377_, _28331_);
  and (_28379_, _28378_, _02176_);
  or (_28380_, _28327_, _03965_);
  and (_28381_, _28368_, _02072_);
  and (_28382_, _28381_, _28380_);
  or (_28383_, _28382_, _28379_);
  and (_28384_, _28383_, _02907_);
  and (_28386_, _28336_, _02177_);
  and (_28387_, _28386_, _28380_);
  or (_28388_, _28387_, _02071_);
  or (_28389_, _28388_, _28384_);
  nor (_28390_, _11628_, _09517_);
  or (_28391_, _28327_, _04788_);
  or (_28392_, _28391_, _28390_);
  and (_28393_, _28392_, _04793_);
  and (_28394_, _28393_, _28389_);
  nor (_28395_, _11634_, _09517_);
  or (_28397_, _28395_, _28327_);
  and (_28398_, _28397_, _02173_);
  or (_28399_, _28398_, _02201_);
  or (_28400_, _28399_, _28394_);
  or (_28401_, _28333_, _02303_);
  and (_28402_, _28401_, _01538_);
  and (_28403_, _28402_, _28400_);
  and (_28404_, _11685_, _03722_);
  or (_28405_, _28404_, _28327_);
  and (_28406_, _28405_, _01537_);
  or (_28408_, _28406_, _38088_);
  or (_28409_, _28408_, _28403_);
  and (_40329_, _28409_, _28326_);
  or (_28410_, _38087_, \oc8051_golden_model_1.TH1 [6]);
  and (_28411_, _28410_, _37580_);
  and (_28412_, _09517_, \oc8051_golden_model_1.TH1 [6]);
  and (_28413_, _11709_, _03722_);
  or (_28414_, _28413_, _28412_);
  and (_28415_, _28414_, _02167_);
  nor (_28416_, _11730_, _09517_);
  or (_28418_, _28416_, _28412_);
  or (_28419_, _28418_, _02814_);
  and (_28420_, _03722_, \oc8051_golden_model_1.ACC [6]);
  or (_28421_, _28420_, _28412_);
  and (_28422_, _28421_, _02817_);
  and (_28423_, _02818_, \oc8051_golden_model_1.TH1 [6]);
  or (_28424_, _28423_, _02001_);
  or (_28425_, _28424_, _28422_);
  and (_28426_, _28425_, _02840_);
  and (_28427_, _28426_, _28419_);
  nor (_28429_, _03808_, _09517_);
  or (_28430_, _28429_, _28412_);
  and (_28431_, _28430_, _01999_);
  or (_28432_, _28431_, _28427_);
  and (_28433_, _28432_, _02021_);
  and (_28434_, _28421_, _02006_);
  or (_28435_, _28434_, _05994_);
  or (_28436_, _28435_, _28433_);
  or (_28437_, _28430_, _05249_);
  and (_28438_, _28437_, _28436_);
  or (_28440_, _28438_, _02528_);
  and (_28441_, _04861_, _03722_);
  or (_28442_, _28412_, _02888_);
  or (_28443_, _28442_, _28441_);
  and (_28444_, _28443_, _02043_);
  and (_28445_, _28444_, _28440_);
  nor (_28446_, _11820_, _09517_);
  or (_28447_, _28446_, _28412_);
  and (_28448_, _28447_, _01602_);
  or (_28449_, _28448_, _01869_);
  or (_28450_, _28449_, _28445_);
  and (_28451_, _09920_, _03722_);
  or (_28452_, _28451_, _28412_);
  or (_28453_, _28452_, _01870_);
  and (_28454_, _28453_, _28450_);
  or (_28455_, _28454_, _02079_);
  and (_28456_, _11835_, _03722_);
  or (_28457_, _28412_, _02166_);
  or (_28458_, _28457_, _28456_);
  and (_28459_, _28458_, _02912_);
  and (_28461_, _28459_, _28455_);
  or (_28462_, _28461_, _28415_);
  and (_28463_, _28462_, _02176_);
  or (_28464_, _28412_, _03863_);
  and (_28465_, _28452_, _02072_);
  and (_28466_, _28465_, _28464_);
  or (_28467_, _28466_, _28463_);
  and (_28468_, _28467_, _02907_);
  and (_28469_, _28421_, _02177_);
  and (_28470_, _28469_, _28464_);
  or (_28472_, _28470_, _02071_);
  or (_28473_, _28472_, _28468_);
  nor (_28474_, _11833_, _09517_);
  or (_28475_, _28412_, _04788_);
  or (_28476_, _28475_, _28474_);
  and (_28477_, _28476_, _04793_);
  and (_28478_, _28477_, _28473_);
  nor (_28479_, _11708_, _09517_);
  or (_28480_, _28479_, _28412_);
  and (_28481_, _28480_, _02173_);
  or (_28483_, _28481_, _02201_);
  or (_28484_, _28483_, _28478_);
  or (_28485_, _28418_, _02303_);
  and (_28486_, _28485_, _01538_);
  and (_28487_, _28486_, _28484_);
  and (_28488_, _11887_, _03722_);
  or (_28489_, _28488_, _28412_);
  and (_28490_, _28489_, _01537_);
  or (_28491_, _28490_, _38088_);
  or (_28492_, _28491_, _28487_);
  and (_40330_, _28492_, _28411_);
  not (_28494_, \oc8051_golden_model_1.TL0 [0]);
  nor (_28495_, _38087_, _28494_);
  nor (_28496_, _03730_, _28494_);
  and (_28497_, _03730_, _03028_);
  or (_28498_, _28497_, _28496_);
  or (_28499_, _28498_, _05249_);
  nor (_28500_, _04106_, _09595_);
  or (_28501_, _28500_, _28496_);
  or (_28502_, _28501_, _02814_);
  and (_28504_, _03730_, \oc8051_golden_model_1.ACC [0]);
  or (_28505_, _28504_, _28496_);
  and (_28506_, _28505_, _02817_);
  nor (_28507_, _02817_, _28494_);
  or (_28508_, _28507_, _02001_);
  or (_28509_, _28508_, _28506_);
  and (_28510_, _28509_, _02840_);
  and (_28511_, _28510_, _28502_);
  and (_28512_, _28498_, _01999_);
  or (_28513_, _28512_, _28511_);
  and (_28515_, _28513_, _02021_);
  and (_28516_, _28505_, _02006_);
  or (_28517_, _28516_, _05994_);
  or (_28518_, _28517_, _28515_);
  and (_28519_, _28518_, _28499_);
  or (_28520_, _28519_, _02528_);
  and (_28521_, _04952_, _03730_);
  or (_28522_, _28496_, _02888_);
  or (_28523_, _28522_, _28521_);
  and (_28524_, _28523_, _28520_);
  or (_28526_, _28524_, _01602_);
  nor (_28527_, _10600_, _09595_);
  or (_28528_, _28527_, _28496_);
  or (_28529_, _28528_, _02043_);
  and (_28530_, _28529_, _01870_);
  and (_28531_, _28530_, _28526_);
  and (_28532_, _03730_, _04562_);
  or (_28533_, _28532_, _28496_);
  and (_28534_, _28533_, _01869_);
  or (_28535_, _28534_, _02079_);
  or (_28537_, _28535_, _28531_);
  and (_28538_, _10614_, _03730_);
  or (_28539_, _28538_, _28496_);
  or (_28540_, _28539_, _02166_);
  and (_28541_, _28540_, _28537_);
  or (_28542_, _28541_, _02167_);
  and (_28543_, _10620_, _03730_);
  or (_28544_, _28496_, _02912_);
  or (_28545_, _28544_, _28543_);
  and (_28546_, _28545_, _02176_);
  and (_28548_, _28546_, _28542_);
  nand (_28549_, _28533_, _02072_);
  nor (_28550_, _28549_, _28500_);
  or (_28551_, _28550_, _28548_);
  and (_28552_, _28551_, _02907_);
  or (_28553_, _28496_, _04106_);
  and (_28554_, _28505_, _02177_);
  and (_28555_, _28554_, _28553_);
  or (_28556_, _28555_, _02071_);
  or (_28557_, _28556_, _28552_);
  nor (_28559_, _10613_, _09595_);
  or (_28560_, _28496_, _04788_);
  or (_28561_, _28560_, _28559_);
  and (_28562_, _28561_, _04793_);
  and (_28563_, _28562_, _28557_);
  nor (_28564_, _10619_, _09595_);
  or (_28565_, _28564_, _28496_);
  and (_28566_, _28565_, _02173_);
  or (_28567_, _28566_, _15577_);
  or (_28568_, _28567_, _28563_);
  or (_28570_, _28501_, _02743_);
  and (_28571_, _28570_, _38087_);
  and (_28572_, _28571_, _28568_);
  or (_28573_, _28572_, _28495_);
  and (_40332_, _28573_, _37580_);
  not (_28574_, \oc8051_golden_model_1.TL0 [1]);
  nor (_28575_, _38087_, _28574_);
  or (_28576_, _03730_, \oc8051_golden_model_1.TL0 [1]);
  and (_28577_, _10698_, _03730_);
  not (_28578_, _28577_);
  and (_28580_, _28578_, _28576_);
  or (_28581_, _28580_, _02814_);
  nand (_28582_, _03730_, _01613_);
  and (_28583_, _28582_, _28576_);
  and (_28584_, _28583_, _02817_);
  nor (_28585_, _02817_, _28574_);
  or (_28586_, _28585_, _02001_);
  or (_28587_, _28586_, _28584_);
  and (_28588_, _28587_, _02840_);
  and (_28589_, _28588_, _28581_);
  nand (_28590_, _03730_, _02811_);
  and (_28591_, _28590_, _28576_);
  and (_28592_, _28591_, _01999_);
  or (_28593_, _28592_, _28589_);
  and (_28594_, _28593_, _02021_);
  and (_28595_, _28583_, _02006_);
  or (_28596_, _28595_, _05994_);
  or (_28597_, _28596_, _28594_);
  or (_28598_, _28591_, _05249_);
  and (_28599_, _28598_, _02888_);
  and (_28601_, _28599_, _28597_);
  or (_28602_, _04907_, _09595_);
  and (_28603_, _28576_, _02528_);
  and (_28604_, _28603_, _28602_);
  or (_28605_, _28604_, _28601_);
  and (_28606_, _28605_, _02043_);
  nand (_28607_, _10802_, _03730_);
  and (_28608_, _28576_, _01602_);
  and (_28609_, _28608_, _28607_);
  or (_28610_, _28609_, _28606_);
  and (_28612_, _28610_, _01870_);
  nand (_28613_, _03730_, _02687_);
  and (_28614_, _28576_, _01869_);
  and (_28615_, _28614_, _28613_);
  or (_28616_, _28615_, _28612_);
  and (_28617_, _28616_, _02166_);
  or (_28618_, _10816_, _09595_);
  and (_28619_, _28576_, _02079_);
  and (_28620_, _28619_, _28618_);
  or (_28621_, _28620_, _28617_);
  and (_28623_, _28621_, _02912_);
  or (_28624_, _10822_, _09595_);
  and (_28625_, _28576_, _02167_);
  and (_28626_, _28625_, _28624_);
  or (_28627_, _28626_, _28623_);
  and (_28628_, _28627_, _02176_);
  or (_28629_, _10692_, _09595_);
  and (_28630_, _28576_, _02072_);
  and (_28631_, _28630_, _28629_);
  or (_28632_, _28631_, _28628_);
  and (_28634_, _28632_, _02907_);
  nor (_28635_, _03730_, _28574_);
  or (_28636_, _28635_, _04058_);
  and (_28637_, _28583_, _02177_);
  and (_28638_, _28637_, _28636_);
  or (_28639_, _28638_, _28634_);
  and (_28640_, _28639_, _02174_);
  or (_28641_, _28582_, _04058_);
  and (_28642_, _28576_, _02173_);
  and (_28643_, _28642_, _28641_);
  or (_28645_, _28643_, _02201_);
  or (_28646_, _28613_, _04058_);
  and (_28647_, _28576_, _02071_);
  and (_28648_, _28647_, _28646_);
  or (_28649_, _28648_, _28645_);
  or (_28650_, _28649_, _28640_);
  or (_28651_, _28580_, _02303_);
  and (_28652_, _28651_, _28650_);
  or (_28653_, _28652_, _01537_);
  or (_28654_, _28635_, _01538_);
  or (_28656_, _28654_, _28577_);
  and (_28657_, _28656_, _38087_);
  and (_28658_, _28657_, _28653_);
  or (_28659_, _28658_, _28575_);
  and (_40333_, _28659_, _37580_);
  not (_28660_, \oc8051_golden_model_1.TL0 [2]);
  nor (_28661_, _38087_, _28660_);
  nor (_28662_, _03730_, _28660_);
  nor (_28663_, _11019_, _09595_);
  or (_28664_, _28663_, _28662_);
  and (_28666_, _28664_, _02173_);
  and (_28667_, _11020_, _03730_);
  or (_28668_, _28667_, _28662_);
  and (_28669_, _28668_, _02167_);
  nor (_28670_, _10905_, _09595_);
  or (_28671_, _28670_, _28662_);
  or (_28672_, _28671_, _02814_);
  and (_28673_, _03730_, \oc8051_golden_model_1.ACC [2]);
  or (_28674_, _28673_, _28662_);
  and (_28675_, _28674_, _02817_);
  nor (_28677_, _02817_, _28660_);
  or (_28678_, _28677_, _02001_);
  or (_28679_, _28678_, _28675_);
  and (_28680_, _28679_, _02840_);
  and (_28681_, _28680_, _28672_);
  nor (_28682_, _09595_, _03455_);
  or (_28683_, _28682_, _28662_);
  and (_28684_, _28683_, _01999_);
  or (_28685_, _28684_, _28681_);
  and (_28686_, _28685_, _02021_);
  and (_28688_, _28674_, _02006_);
  or (_28689_, _28688_, _05994_);
  or (_28690_, _28689_, _28686_);
  or (_28691_, _28683_, _05249_);
  and (_28692_, _28691_, _28690_);
  or (_28693_, _28692_, _02528_);
  and (_28694_, _05043_, _03730_);
  or (_28695_, _28662_, _02888_);
  or (_28696_, _28695_, _28694_);
  and (_28697_, _28696_, _28693_);
  or (_28699_, _28697_, _01602_);
  nor (_28700_, _11000_, _09595_);
  or (_28701_, _28662_, _02043_);
  or (_28702_, _28701_, _28700_);
  and (_28703_, _28702_, _01870_);
  and (_28704_, _28703_, _28699_);
  and (_28705_, _03730_, _04724_);
  or (_28706_, _28705_, _28662_);
  and (_28707_, _28706_, _01869_);
  or (_28708_, _28707_, _02079_);
  or (_28710_, _28708_, _28704_);
  and (_28711_, _11014_, _03730_);
  or (_28712_, _28662_, _02166_);
  or (_28713_, _28712_, _28711_);
  and (_28714_, _28713_, _02912_);
  and (_28715_, _28714_, _28710_);
  or (_28716_, _28715_, _28669_);
  and (_28717_, _28716_, _02176_);
  or (_28718_, _28662_, _04156_);
  and (_28719_, _28706_, _02072_);
  and (_28721_, _28719_, _28718_);
  or (_28722_, _28721_, _28717_);
  and (_28723_, _28722_, _02907_);
  and (_28724_, _28674_, _02177_);
  and (_28725_, _28724_, _28718_);
  or (_28726_, _28725_, _02071_);
  or (_28727_, _28726_, _28723_);
  nor (_28728_, _11013_, _09595_);
  or (_28729_, _28662_, _04788_);
  or (_28730_, _28729_, _28728_);
  and (_28732_, _28730_, _04793_);
  and (_28733_, _28732_, _28727_);
  or (_28734_, _28733_, _28666_);
  and (_28735_, _28734_, _02303_);
  and (_28736_, _28671_, _02201_);
  or (_28737_, _28736_, _01537_);
  or (_28738_, _28737_, _28735_);
  and (_28739_, _11072_, _03730_);
  or (_28740_, _28662_, _01538_);
  or (_28741_, _28740_, _28739_);
  and (_28742_, _28741_, _38087_);
  and (_28743_, _28742_, _28738_);
  or (_28744_, _28743_, _28661_);
  and (_40334_, _28744_, _37580_);
  or (_28745_, _38087_, \oc8051_golden_model_1.TL0 [3]);
  and (_28746_, _28745_, _37580_);
  and (_28747_, _09595_, \oc8051_golden_model_1.TL0 [3]);
  and (_28748_, _11094_, _03730_);
  or (_28749_, _28748_, _28747_);
  and (_28750_, _28749_, _02167_);
  nor (_28752_, _11101_, _09595_);
  or (_28753_, _28752_, _28747_);
  or (_28754_, _28753_, _02814_);
  and (_28755_, _03730_, \oc8051_golden_model_1.ACC [3]);
  or (_28756_, _28755_, _28747_);
  and (_28757_, _28756_, _02817_);
  and (_28758_, _02818_, \oc8051_golden_model_1.TL0 [3]);
  or (_28759_, _28758_, _02001_);
  or (_28760_, _28759_, _28757_);
  and (_28761_, _28760_, _02840_);
  and (_28763_, _28761_, _28754_);
  nor (_28764_, _09595_, _03268_);
  or (_28765_, _28764_, _28747_);
  and (_28766_, _28765_, _01999_);
  or (_28767_, _28766_, _28763_);
  and (_28768_, _28767_, _02021_);
  and (_28769_, _28756_, _02006_);
  or (_28770_, _28769_, _05994_);
  or (_28771_, _28770_, _28768_);
  or (_28772_, _28765_, _05249_);
  and (_28774_, _28772_, _28771_);
  or (_28775_, _28774_, _02528_);
  and (_28776_, _04998_, _03730_);
  or (_28777_, _28747_, _02888_);
  or (_28778_, _28777_, _28776_);
  and (_28779_, _28778_, _02043_);
  and (_28780_, _28779_, _28775_);
  nor (_28781_, _11206_, _09595_);
  or (_28782_, _28781_, _28747_);
  and (_28783_, _28782_, _01602_);
  or (_28785_, _28783_, _01869_);
  or (_28786_, _28785_, _28780_);
  and (_28787_, _03730_, _04678_);
  or (_28788_, _28787_, _28747_);
  or (_28789_, _28788_, _01870_);
  and (_28790_, _28789_, _28786_);
  or (_28791_, _28790_, _02079_);
  and (_28792_, _11222_, _03730_);
  or (_28793_, _28747_, _02166_);
  or (_28794_, _28793_, _28792_);
  and (_28796_, _28794_, _02912_);
  and (_28797_, _28796_, _28791_);
  or (_28798_, _28797_, _28750_);
  and (_28799_, _28798_, _02176_);
  or (_28800_, _28747_, _04014_);
  and (_28801_, _28788_, _02072_);
  and (_28802_, _28801_, _28800_);
  or (_28803_, _28802_, _28799_);
  and (_28804_, _28803_, _02907_);
  and (_28805_, _28756_, _02177_);
  and (_28807_, _28805_, _28800_);
  or (_28808_, _28807_, _02071_);
  or (_28809_, _28808_, _28804_);
  nor (_28810_, _11220_, _09595_);
  or (_28811_, _28747_, _04788_);
  or (_28812_, _28811_, _28810_);
  and (_28813_, _28812_, _04793_);
  and (_28814_, _28813_, _28809_);
  nor (_28815_, _11093_, _09595_);
  or (_28816_, _28815_, _28747_);
  and (_28818_, _28816_, _02173_);
  or (_28819_, _28818_, _02201_);
  or (_28820_, _28819_, _28814_);
  or (_28821_, _28753_, _02303_);
  and (_28822_, _28821_, _01538_);
  and (_28823_, _28822_, _28820_);
  and (_28824_, _11273_, _03730_);
  or (_28825_, _28824_, _28747_);
  and (_28826_, _28825_, _01537_);
  or (_28827_, _28826_, _38088_);
  or (_28829_, _28827_, _28823_);
  and (_40335_, _28829_, _28746_);
  or (_28830_, _38087_, \oc8051_golden_model_1.TL0 [4]);
  and (_28831_, _28830_, _37580_);
  and (_28832_, _09595_, \oc8051_golden_model_1.TL0 [4]);
  and (_28833_, _11431_, _03730_);
  or (_28834_, _28833_, _28832_);
  and (_28835_, _28834_, _02167_);
  nor (_28836_, _04211_, _09595_);
  or (_28837_, _28836_, _28832_);
  or (_28839_, _28837_, _05249_);
  nor (_28840_, _11317_, _09595_);
  or (_28841_, _28840_, _28832_);
  or (_28842_, _28841_, _02814_);
  and (_28843_, _03730_, \oc8051_golden_model_1.ACC [4]);
  or (_28844_, _28843_, _28832_);
  and (_28845_, _28844_, _02817_);
  and (_28846_, _02818_, \oc8051_golden_model_1.TL0 [4]);
  or (_28847_, _28846_, _02001_);
  or (_28848_, _28847_, _28845_);
  and (_28850_, _28848_, _02840_);
  and (_28851_, _28850_, _28842_);
  and (_28852_, _28837_, _01999_);
  or (_28853_, _28852_, _28851_);
  and (_28854_, _28853_, _02021_);
  and (_28855_, _28844_, _02006_);
  or (_28856_, _28855_, _05994_);
  or (_28857_, _28856_, _28854_);
  and (_28858_, _28857_, _28839_);
  or (_28859_, _28858_, _02528_);
  and (_28861_, _05135_, _03730_);
  or (_28862_, _28832_, _02888_);
  or (_28863_, _28862_, _28861_);
  and (_28864_, _28863_, _02043_);
  and (_28865_, _28864_, _28859_);
  nor (_28866_, _11411_, _09595_);
  or (_28867_, _28866_, _28832_);
  and (_28868_, _28867_, _01602_);
  or (_28869_, _28868_, _01869_);
  or (_28870_, _28869_, _28865_);
  and (_28872_, _04694_, _03730_);
  or (_28873_, _28872_, _28832_);
  or (_28874_, _28873_, _01870_);
  and (_28875_, _28874_, _28870_);
  or (_28876_, _28875_, _02079_);
  and (_28877_, _11425_, _03730_);
  or (_28878_, _28832_, _02166_);
  or (_28879_, _28878_, _28877_);
  and (_28880_, _28879_, _02912_);
  and (_28881_, _28880_, _28876_);
  or (_28882_, _28881_, _28835_);
  and (_28883_, _28882_, _02176_);
  or (_28884_, _28832_, _04258_);
  and (_28885_, _28873_, _02072_);
  and (_28886_, _28885_, _28884_);
  or (_28887_, _28886_, _28883_);
  and (_28888_, _28887_, _02907_);
  and (_28889_, _28844_, _02177_);
  and (_28890_, _28889_, _28884_);
  or (_28891_, _28890_, _02071_);
  or (_28893_, _28891_, _28888_);
  nor (_28894_, _11424_, _09595_);
  or (_28895_, _28832_, _04788_);
  or (_28896_, _28895_, _28894_);
  and (_28897_, _28896_, _04793_);
  and (_28898_, _28897_, _28893_);
  nor (_28899_, _11430_, _09595_);
  or (_28900_, _28899_, _28832_);
  and (_28901_, _28900_, _02173_);
  or (_28902_, _28901_, _02201_);
  or (_28904_, _28902_, _28898_);
  or (_28905_, _28841_, _02303_);
  and (_28906_, _28905_, _01538_);
  and (_28907_, _28906_, _28904_);
  and (_28908_, _11487_, _03730_);
  or (_28909_, _28908_, _28832_);
  and (_28910_, _28909_, _01537_);
  or (_28911_, _28910_, _38088_);
  or (_28912_, _28911_, _28907_);
  and (_40336_, _28912_, _28831_);
  or (_28914_, _38087_, \oc8051_golden_model_1.TL0 [5]);
  and (_28915_, _28914_, _37580_);
  and (_28916_, _09595_, \oc8051_golden_model_1.TL0 [5]);
  and (_28917_, _11635_, _03730_);
  or (_28918_, _28917_, _28916_);
  and (_28919_, _28918_, _02167_);
  nor (_28920_, _03916_, _09595_);
  or (_28921_, _28920_, _28916_);
  or (_28922_, _28921_, _05249_);
  nor (_28923_, _11525_, _09595_);
  or (_28925_, _28923_, _28916_);
  or (_28926_, _28925_, _02814_);
  and (_28927_, _03730_, \oc8051_golden_model_1.ACC [5]);
  or (_28928_, _28927_, _28916_);
  and (_28929_, _28928_, _02817_);
  and (_28930_, _02818_, \oc8051_golden_model_1.TL0 [5]);
  or (_28931_, _28930_, _02001_);
  or (_28932_, _28931_, _28929_);
  and (_28933_, _28932_, _02840_);
  and (_28934_, _28933_, _28926_);
  and (_28936_, _28921_, _01999_);
  or (_28937_, _28936_, _28934_);
  and (_28938_, _28937_, _02021_);
  and (_28939_, _28928_, _02006_);
  or (_28940_, _28939_, _05994_);
  or (_28941_, _28940_, _28938_);
  and (_28942_, _28941_, _28922_);
  or (_28943_, _28942_, _02528_);
  and (_28944_, _05090_, _03730_);
  or (_28945_, _28916_, _02888_);
  or (_28947_, _28945_, _28944_);
  and (_28948_, _28947_, _02043_);
  and (_28949_, _28948_, _28943_);
  nor (_28950_, _11615_, _09595_);
  or (_28951_, _28950_, _28916_);
  and (_28952_, _28951_, _01602_);
  or (_28953_, _28952_, _01869_);
  or (_28954_, _28953_, _28949_);
  and (_28955_, _04672_, _03730_);
  or (_28956_, _28955_, _28916_);
  or (_28958_, _28956_, _01870_);
  and (_28959_, _28958_, _28954_);
  or (_28960_, _28959_, _02079_);
  and (_28961_, _11629_, _03730_);
  or (_28962_, _28916_, _02166_);
  or (_28963_, _28962_, _28961_);
  and (_28964_, _28963_, _02912_);
  and (_28965_, _28964_, _28960_);
  or (_28966_, _28965_, _28919_);
  and (_28967_, _28966_, _02176_);
  or (_28969_, _28916_, _03965_);
  and (_28970_, _28956_, _02072_);
  and (_28971_, _28970_, _28969_);
  or (_28972_, _28971_, _28967_);
  and (_28973_, _28972_, _02907_);
  and (_28974_, _28928_, _02177_);
  and (_28975_, _28974_, _28969_);
  or (_28976_, _28975_, _02071_);
  or (_28977_, _28976_, _28973_);
  nor (_28978_, _11628_, _09595_);
  or (_28980_, _28916_, _04788_);
  or (_28981_, _28980_, _28978_);
  and (_28982_, _28981_, _04793_);
  and (_28983_, _28982_, _28977_);
  nor (_28984_, _11634_, _09595_);
  or (_28985_, _28984_, _28916_);
  and (_28986_, _28985_, _02173_);
  or (_28987_, _28986_, _02201_);
  or (_28988_, _28987_, _28983_);
  or (_28989_, _28925_, _02303_);
  and (_28991_, _28989_, _01538_);
  and (_28992_, _28991_, _28988_);
  and (_28993_, _11685_, _03730_);
  or (_28994_, _28993_, _28916_);
  and (_28995_, _28994_, _01537_);
  or (_28996_, _28995_, _38088_);
  or (_28997_, _28996_, _28992_);
  and (_40337_, _28997_, _28915_);
  or (_28998_, _38087_, \oc8051_golden_model_1.TL0 [6]);
  and (_28999_, _28998_, _37580_);
  and (_29001_, _09595_, \oc8051_golden_model_1.TL0 [6]);
  and (_29002_, _11709_, _03730_);
  or (_29003_, _29002_, _29001_);
  and (_29004_, _29003_, _02167_);
  nor (_29005_, _03808_, _09595_);
  or (_29006_, _29005_, _29001_);
  or (_29007_, _29006_, _05249_);
  nor (_29008_, _11730_, _09595_);
  or (_29009_, _29008_, _29001_);
  or (_29010_, _29009_, _02814_);
  and (_29012_, _03730_, \oc8051_golden_model_1.ACC [6]);
  or (_29013_, _29012_, _29001_);
  and (_29014_, _29013_, _02817_);
  and (_29015_, _02818_, \oc8051_golden_model_1.TL0 [6]);
  or (_29016_, _29015_, _02001_);
  or (_29017_, _29016_, _29014_);
  and (_29018_, _29017_, _02840_);
  and (_29019_, _29018_, _29010_);
  and (_29020_, _29006_, _01999_);
  or (_29021_, _29020_, _29019_);
  and (_29023_, _29021_, _02021_);
  and (_29024_, _29013_, _02006_);
  or (_29025_, _29024_, _05994_);
  or (_29026_, _29025_, _29023_);
  and (_29027_, _29026_, _29007_);
  or (_29028_, _29027_, _02528_);
  and (_29029_, _04861_, _03730_);
  or (_29030_, _29001_, _02888_);
  or (_29031_, _29030_, _29029_);
  and (_29032_, _29031_, _02043_);
  and (_29033_, _29032_, _29028_);
  nor (_29034_, _11820_, _09595_);
  or (_29035_, _29034_, _29001_);
  and (_29036_, _29035_, _01602_);
  or (_29037_, _29036_, _01869_);
  or (_29038_, _29037_, _29033_);
  and (_29039_, _09920_, _03730_);
  or (_29040_, _29039_, _29001_);
  or (_29041_, _29040_, _01870_);
  and (_29042_, _29041_, _29038_);
  or (_29044_, _29042_, _02079_);
  and (_29045_, _11835_, _03730_);
  or (_29046_, _29001_, _02166_);
  or (_29047_, _29046_, _29045_);
  and (_29048_, _29047_, _02912_);
  and (_29049_, _29048_, _29044_);
  or (_29050_, _29049_, _29004_);
  and (_29051_, _29050_, _02176_);
  or (_29052_, _29001_, _03863_);
  and (_29053_, _29040_, _02072_);
  and (_29055_, _29053_, _29052_);
  or (_29056_, _29055_, _29051_);
  and (_29057_, _29056_, _02907_);
  and (_29058_, _29013_, _02177_);
  and (_29059_, _29058_, _29052_);
  or (_29060_, _29059_, _02071_);
  or (_29061_, _29060_, _29057_);
  nor (_29062_, _11833_, _09595_);
  or (_29063_, _29001_, _04788_);
  or (_29064_, _29063_, _29062_);
  and (_29066_, _29064_, _04793_);
  and (_29067_, _29066_, _29061_);
  nor (_29068_, _11708_, _09595_);
  or (_29069_, _29068_, _29001_);
  and (_29070_, _29069_, _02173_);
  or (_29071_, _29070_, _02201_);
  or (_29072_, _29071_, _29067_);
  or (_29073_, _29009_, _02303_);
  and (_29074_, _29073_, _01538_);
  and (_29075_, _29074_, _29072_);
  and (_29078_, _11887_, _03730_);
  or (_29079_, _29078_, _29001_);
  and (_29080_, _29079_, _01537_);
  or (_29081_, _29080_, _38088_);
  or (_29082_, _29081_, _29075_);
  and (_40338_, _29082_, _28999_);
  and (_29083_, _38088_, \oc8051_golden_model_1.TL1 [0]);
  and (_29084_, _09673_, \oc8051_golden_model_1.TL1 [0]);
  nor (_29085_, _04106_, _09678_);
  or (_29086_, _29085_, _29084_);
  or (_29088_, _29086_, _02814_);
  and (_29089_, _03708_, \oc8051_golden_model_1.ACC [0]);
  or (_29090_, _29089_, _29084_);
  and (_29091_, _29090_, _02817_);
  and (_29092_, _02818_, \oc8051_golden_model_1.TL1 [0]);
  or (_29093_, _29092_, _02001_);
  or (_29094_, _29093_, _29091_);
  and (_29095_, _29094_, _02840_);
  and (_29096_, _29095_, _29088_);
  and (_29097_, _03845_, _03028_);
  or (_29099_, _29097_, _29084_);
  and (_29100_, _29099_, _01999_);
  or (_29101_, _29100_, _29096_);
  and (_29102_, _29101_, _02021_);
  and (_29103_, _29090_, _02006_);
  or (_29104_, _29103_, _05994_);
  or (_29105_, _29104_, _29102_);
  or (_29106_, _29099_, _05249_);
  and (_29107_, _29106_, _29105_);
  or (_29108_, _29107_, _02528_);
  or (_29110_, _29084_, _02888_);
  and (_29111_, _04952_, _03708_);
  or (_29112_, _29111_, _29110_);
  and (_29113_, _29112_, _29108_);
  or (_29114_, _29113_, _01602_);
  nor (_29115_, _10600_, _09673_);
  or (_29116_, _29115_, _29084_);
  or (_29117_, _29116_, _02043_);
  and (_29118_, _29117_, _01870_);
  and (_29119_, _29118_, _29114_);
  and (_29121_, _03708_, _04562_);
  or (_29122_, _29121_, _29084_);
  and (_29123_, _29122_, _01869_);
  or (_29124_, _29123_, _02079_);
  or (_29125_, _29124_, _29119_);
  and (_29126_, _10614_, _03708_);
  or (_29127_, _29126_, _29084_);
  or (_29128_, _29127_, _02166_);
  and (_29129_, _29128_, _29125_);
  or (_29130_, _29129_, _02167_);
  and (_29132_, _10620_, _03845_);
  or (_29133_, _29084_, _02912_);
  or (_29134_, _29133_, _29132_);
  and (_29135_, _29134_, _02176_);
  and (_29136_, _29135_, _29130_);
  nand (_29137_, _29122_, _02072_);
  nor (_29138_, _29137_, _29085_);
  or (_29139_, _29138_, _29136_);
  and (_29140_, _29139_, _02907_);
  or (_29141_, _29084_, _04106_);
  and (_29143_, _29090_, _02177_);
  and (_29144_, _29143_, _29141_);
  or (_29145_, _29144_, _02071_);
  or (_29146_, _29145_, _29140_);
  nor (_29147_, _10613_, _09678_);
  or (_29148_, _29084_, _04788_);
  or (_29149_, _29148_, _29147_);
  and (_29150_, _29149_, _04793_);
  and (_29151_, _29150_, _29146_);
  nor (_29152_, _10619_, _09678_);
  or (_29154_, _29152_, _29084_);
  and (_29155_, _29154_, _02173_);
  or (_29156_, _29155_, _15577_);
  or (_29157_, _29156_, _29151_);
  or (_29158_, _29086_, _02743_);
  and (_29159_, _29158_, _38087_);
  and (_29160_, _29159_, _29157_);
  or (_29161_, _29160_, _29083_);
  and (_40340_, _29161_, _37580_);
  and (_29162_, _38088_, \oc8051_golden_model_1.TL1 [1]);
  or (_29163_, _03708_, \oc8051_golden_model_1.TL1 [1]);
  and (_29164_, _10698_, _03845_);
  not (_29165_, _29164_);
  and (_29166_, _29165_, _29163_);
  or (_29167_, _29166_, _02814_);
  nand (_29168_, _03845_, _01613_);
  and (_29169_, _29168_, _29163_);
  and (_29170_, _29169_, _02817_);
  and (_29171_, _02818_, \oc8051_golden_model_1.TL1 [1]);
  or (_29172_, _29171_, _02001_);
  or (_29174_, _29172_, _29170_);
  and (_29175_, _29174_, _02840_);
  and (_29176_, _29175_, _29167_);
  nand (_29177_, _03708_, _02811_);
  and (_29178_, _29177_, _29163_);
  and (_29179_, _29178_, _01999_);
  or (_29180_, _29179_, _29176_);
  and (_29181_, _29180_, _02021_);
  and (_29182_, _29169_, _02006_);
  or (_29183_, _29182_, _05994_);
  or (_29186_, _29183_, _29181_);
  or (_29187_, _29178_, _05249_);
  and (_29188_, _29187_, _02888_);
  and (_29189_, _29188_, _29186_);
  or (_29190_, _04907_, _09678_);
  and (_29191_, _29163_, _02528_);
  and (_29192_, _29191_, _29190_);
  or (_29193_, _29192_, _29189_);
  and (_29194_, _29193_, _02043_);
  nand (_29195_, _10802_, _03845_);
  and (_29197_, _29163_, _01602_);
  and (_29198_, _29197_, _29195_);
  or (_29199_, _29198_, _29194_);
  and (_29200_, _29199_, _01870_);
  and (_29201_, _29163_, _01869_);
  nand (_29202_, _03845_, _02687_);
  and (_29203_, _29202_, _29201_);
  or (_29204_, _29203_, _29200_);
  and (_29205_, _29204_, _02166_);
  or (_29206_, _10816_, _09678_);
  and (_29208_, _29163_, _02079_);
  and (_29209_, _29208_, _29206_);
  or (_29210_, _29209_, _29205_);
  and (_29211_, _29210_, _02912_);
  or (_29212_, _10822_, _09678_);
  and (_29213_, _29163_, _02167_);
  and (_29214_, _29213_, _29212_);
  or (_29215_, _29214_, _29211_);
  and (_29216_, _29215_, _02176_);
  or (_29217_, _10692_, _09678_);
  and (_29219_, _29163_, _02072_);
  and (_29220_, _29219_, _29217_);
  or (_29221_, _29220_, _29216_);
  and (_29222_, _29221_, _02907_);
  and (_29223_, _09673_, \oc8051_golden_model_1.TL1 [1]);
  or (_29224_, _29223_, _04058_);
  and (_29225_, _29169_, _02177_);
  and (_29226_, _29225_, _29224_);
  or (_29227_, _29226_, _29222_);
  and (_29228_, _29227_, _02174_);
  or (_29230_, _29168_, _04058_);
  and (_29231_, _29163_, _02173_);
  and (_29232_, _29231_, _29230_);
  or (_29233_, _29232_, _02201_);
  or (_29234_, _29202_, _04058_);
  and (_29235_, _29163_, _02071_);
  and (_29236_, _29235_, _29234_);
  or (_29237_, _29236_, _29233_);
  or (_29238_, _29237_, _29228_);
  or (_29239_, _29166_, _02303_);
  and (_29241_, _29239_, _29238_);
  or (_29242_, _29241_, _01537_);
  or (_29243_, _29223_, _01538_);
  or (_29244_, _29243_, _29164_);
  and (_29245_, _29244_, _38087_);
  and (_29246_, _29245_, _29242_);
  or (_29247_, _29246_, _29162_);
  and (_40341_, _29247_, _37580_);
  and (_29248_, _38088_, \oc8051_golden_model_1.TL1 [2]);
  and (_29249_, _09673_, \oc8051_golden_model_1.TL1 [2]);
  nor (_29251_, _11019_, _09678_);
  or (_29252_, _29251_, _29249_);
  and (_29253_, _29252_, _02173_);
  or (_29254_, _29249_, _04156_);
  and (_29255_, _03708_, _04724_);
  or (_29256_, _29255_, _29249_);
  and (_29257_, _29256_, _02072_);
  and (_29258_, _29257_, _29254_);
  and (_29259_, _05043_, _03708_);
  or (_29260_, _29259_, _29249_);
  and (_29262_, _29260_, _02528_);
  nor (_29263_, _10905_, _09678_);
  or (_29264_, _29263_, _29249_);
  or (_29265_, _29264_, _02814_);
  and (_29266_, _03708_, \oc8051_golden_model_1.ACC [2]);
  or (_29267_, _29266_, _29249_);
  and (_29268_, _29267_, _02817_);
  and (_29269_, _02818_, \oc8051_golden_model_1.TL1 [2]);
  or (_29270_, _29269_, _02001_);
  or (_29271_, _29270_, _29268_);
  and (_29273_, _29271_, _02840_);
  and (_29274_, _29273_, _29265_);
  nor (_29275_, _09678_, _03455_);
  or (_29276_, _29275_, _29249_);
  and (_29277_, _29276_, _01999_);
  or (_29278_, _29277_, _29274_);
  and (_29279_, _29278_, _02021_);
  and (_29280_, _29267_, _02006_);
  or (_29281_, _29280_, _05994_);
  or (_29282_, _29281_, _29279_);
  or (_29284_, _29276_, _05249_);
  and (_29285_, _29284_, _02888_);
  and (_29286_, _29285_, _29282_);
  or (_29287_, _29286_, _01602_);
  or (_29288_, _29287_, _29262_);
  nor (_29289_, _11000_, _09673_);
  or (_29290_, _29289_, _29249_);
  or (_29291_, _29290_, _02043_);
  and (_29292_, _29291_, _01870_);
  and (_29293_, _29292_, _29288_);
  and (_29296_, _29256_, _01869_);
  or (_29297_, _29296_, _02079_);
  or (_29298_, _29297_, _29293_);
  and (_29299_, _11014_, _03708_);
  or (_29300_, _29299_, _29249_);
  or (_29301_, _29300_, _02166_);
  and (_29302_, _29301_, _29298_);
  or (_29303_, _29302_, _02167_);
  and (_29304_, _11020_, _03845_);
  or (_29305_, _29249_, _02912_);
  or (_29306_, _29305_, _29304_);
  and (_29307_, _29306_, _02176_);
  and (_29308_, _29307_, _29303_);
  or (_29309_, _29308_, _29258_);
  and (_29310_, _29309_, _02907_);
  and (_29311_, _29267_, _02177_);
  and (_29312_, _29311_, _29254_);
  or (_29313_, _29312_, _02071_);
  or (_29314_, _29313_, _29310_);
  nor (_29315_, _11013_, _09678_);
  or (_29317_, _29249_, _04788_);
  or (_29318_, _29317_, _29315_);
  and (_29319_, _29318_, _04793_);
  and (_29320_, _29319_, _29314_);
  or (_29321_, _29320_, _29253_);
  and (_29322_, _29321_, _02303_);
  and (_29323_, _29264_, _02201_);
  or (_29324_, _29323_, _01537_);
  or (_29325_, _29324_, _29322_);
  and (_29326_, _11072_, _03845_);
  or (_29328_, _29249_, _01538_);
  or (_29329_, _29328_, _29326_);
  and (_29330_, _29329_, _38087_);
  and (_29331_, _29330_, _29325_);
  or (_29332_, _29331_, _29248_);
  and (_40342_, _29332_, _37580_);
  or (_29333_, _38087_, \oc8051_golden_model_1.TL1 [3]);
  and (_29334_, _29333_, _37580_);
  and (_29335_, _09673_, \oc8051_golden_model_1.TL1 [3]);
  or (_29336_, _29335_, _04014_);
  and (_29338_, _03708_, _04678_);
  or (_29339_, _29338_, _29335_);
  and (_29340_, _29339_, _02072_);
  and (_29341_, _29340_, _29336_);
  and (_29342_, _11094_, _03845_);
  or (_29343_, _29342_, _29335_);
  and (_29344_, _29343_, _02167_);
  nor (_29345_, _11101_, _09678_);
  or (_29346_, _29345_, _29335_);
  or (_29347_, _29346_, _02814_);
  and (_29349_, _03708_, \oc8051_golden_model_1.ACC [3]);
  or (_29350_, _29349_, _29335_);
  and (_29351_, _29350_, _02817_);
  and (_29352_, _02818_, \oc8051_golden_model_1.TL1 [3]);
  or (_29353_, _29352_, _02001_);
  or (_29354_, _29353_, _29351_);
  and (_29355_, _29354_, _02840_);
  and (_29356_, _29355_, _29347_);
  nor (_29357_, _09678_, _03268_);
  or (_29358_, _29357_, _29335_);
  and (_29360_, _29358_, _01999_);
  or (_29361_, _29360_, _29356_);
  and (_29362_, _29361_, _02021_);
  and (_29363_, _29350_, _02006_);
  or (_29364_, _29363_, _05994_);
  or (_29365_, _29364_, _29362_);
  or (_29366_, _29358_, _05249_);
  and (_29367_, _29366_, _29365_);
  or (_29368_, _29367_, _02528_);
  and (_29369_, _04998_, _03708_);
  or (_29371_, _29335_, _02888_);
  or (_29372_, _29371_, _29369_);
  and (_29373_, _29372_, _02043_);
  and (_29374_, _29373_, _29368_);
  nor (_29375_, _11206_, _09673_);
  or (_29376_, _29375_, _29335_);
  and (_29377_, _29376_, _01602_);
  or (_29378_, _29377_, _01869_);
  or (_29379_, _29378_, _29374_);
  or (_29380_, _29339_, _01870_);
  and (_29382_, _29380_, _29379_);
  or (_29383_, _29382_, _02079_);
  and (_29384_, _11222_, _03845_);
  or (_29385_, _29335_, _02166_);
  or (_29386_, _29385_, _29384_);
  and (_29387_, _29386_, _02912_);
  and (_29388_, _29387_, _29383_);
  or (_29389_, _29388_, _29344_);
  and (_29390_, _29389_, _02176_);
  or (_29391_, _29390_, _29341_);
  and (_29393_, _29391_, _02907_);
  and (_29394_, _29350_, _02177_);
  and (_29395_, _29394_, _29336_);
  or (_29396_, _29395_, _02071_);
  or (_29397_, _29396_, _29393_);
  nor (_29398_, _11220_, _09678_);
  or (_29399_, _29335_, _04788_);
  or (_29400_, _29399_, _29398_);
  and (_29401_, _29400_, _04793_);
  and (_29402_, _29401_, _29397_);
  nor (_29405_, _11093_, _09678_);
  or (_29406_, _29405_, _29335_);
  and (_29407_, _29406_, _02173_);
  or (_29408_, _29407_, _02201_);
  or (_29409_, _29408_, _29402_);
  or (_29410_, _29346_, _02303_);
  and (_29411_, _29410_, _01538_);
  and (_29412_, _29411_, _29409_);
  and (_29413_, _11273_, _03845_);
  or (_29414_, _29413_, _29335_);
  and (_29416_, _29414_, _01537_);
  or (_29417_, _29416_, _38088_);
  or (_29418_, _29417_, _29412_);
  and (_40343_, _29418_, _29334_);
  or (_29419_, _38087_, \oc8051_golden_model_1.TL1 [4]);
  and (_29420_, _29419_, _37580_);
  and (_29421_, _09673_, \oc8051_golden_model_1.TL1 [4]);
  and (_29422_, _11431_, _03845_);
  or (_29423_, _29422_, _29421_);
  and (_29424_, _29423_, _02167_);
  nor (_29426_, _11317_, _09678_);
  or (_29427_, _29426_, _29421_);
  or (_29428_, _29427_, _02814_);
  and (_29429_, _03708_, \oc8051_golden_model_1.ACC [4]);
  or (_29430_, _29429_, _29421_);
  and (_29431_, _29430_, _02817_);
  and (_29432_, _02818_, \oc8051_golden_model_1.TL1 [4]);
  or (_29433_, _29432_, _02001_);
  or (_29434_, _29433_, _29431_);
  and (_29435_, _29434_, _02840_);
  and (_29437_, _29435_, _29428_);
  nor (_29438_, _04211_, _09678_);
  or (_29439_, _29438_, _29421_);
  and (_29440_, _29439_, _01999_);
  or (_29441_, _29440_, _29437_);
  and (_29442_, _29441_, _02021_);
  and (_29443_, _29430_, _02006_);
  or (_29444_, _29443_, _05994_);
  or (_29445_, _29444_, _29442_);
  or (_29446_, _29439_, _05249_);
  and (_29447_, _29446_, _29445_);
  or (_29448_, _29447_, _02528_);
  or (_29449_, _29421_, _02888_);
  and (_29450_, _05135_, _03708_);
  or (_29451_, _29450_, _29449_);
  and (_29452_, _29451_, _02043_);
  and (_29453_, _29452_, _29448_);
  nor (_29454_, _11411_, _09673_);
  or (_29455_, _29454_, _29421_);
  and (_29456_, _29455_, _01602_);
  or (_29458_, _29456_, _01869_);
  or (_29459_, _29458_, _29453_);
  and (_29460_, _04694_, _03708_);
  or (_29461_, _29460_, _29421_);
  or (_29462_, _29461_, _01870_);
  and (_29463_, _29462_, _29459_);
  or (_29464_, _29463_, _02079_);
  and (_29465_, _11425_, _03845_);
  or (_29466_, _29421_, _02166_);
  or (_29467_, _29466_, _29465_);
  and (_29469_, _29467_, _02912_);
  and (_29470_, _29469_, _29464_);
  or (_29471_, _29470_, _29424_);
  and (_29472_, _29471_, _02176_);
  or (_29473_, _29421_, _04258_);
  and (_29474_, _29461_, _02072_);
  and (_29475_, _29474_, _29473_);
  or (_29476_, _29475_, _29472_);
  and (_29477_, _29476_, _02907_);
  and (_29478_, _29430_, _02177_);
  and (_29480_, _29478_, _29473_);
  or (_29481_, _29480_, _02071_);
  or (_29482_, _29481_, _29477_);
  nor (_29483_, _11424_, _09678_);
  or (_29484_, _29421_, _04788_);
  or (_29485_, _29484_, _29483_);
  and (_29486_, _29485_, _04793_);
  and (_29487_, _29486_, _29482_);
  nor (_29488_, _11430_, _09678_);
  or (_29489_, _29488_, _29421_);
  and (_29491_, _29489_, _02173_);
  or (_29492_, _29491_, _02201_);
  or (_29493_, _29492_, _29487_);
  or (_29494_, _29427_, _02303_);
  and (_29495_, _29494_, _01538_);
  and (_29496_, _29495_, _29493_);
  and (_29497_, _11487_, _03845_);
  or (_29498_, _29497_, _29421_);
  and (_29499_, _29498_, _01537_);
  or (_29500_, _29499_, _38088_);
  or (_29502_, _29500_, _29496_);
  and (_40345_, _29502_, _29420_);
  or (_29503_, _38087_, \oc8051_golden_model_1.TL1 [5]);
  and (_29504_, _29503_, _37580_);
  and (_29505_, _09673_, \oc8051_golden_model_1.TL1 [5]);
  and (_29506_, _11635_, _03845_);
  or (_29507_, _29506_, _29505_);
  and (_29508_, _29507_, _02167_);
  nor (_29509_, _11525_, _09678_);
  or (_29510_, _29509_, _29505_);
  or (_29513_, _29510_, _02814_);
  and (_29514_, _03708_, \oc8051_golden_model_1.ACC [5]);
  or (_29515_, _29514_, _29505_);
  and (_29516_, _29515_, _02817_);
  and (_29517_, _02818_, \oc8051_golden_model_1.TL1 [5]);
  or (_29518_, _29517_, _02001_);
  or (_29519_, _29518_, _29516_);
  and (_29520_, _29519_, _02840_);
  and (_29521_, _29520_, _29513_);
  nor (_29522_, _03916_, _09678_);
  or (_29524_, _29522_, _29505_);
  and (_29525_, _29524_, _01999_);
  or (_29526_, _29525_, _29521_);
  and (_29527_, _29526_, _02021_);
  and (_29528_, _29515_, _02006_);
  or (_29529_, _29528_, _05994_);
  or (_29530_, _29529_, _29527_);
  or (_29531_, _29524_, _05249_);
  and (_29532_, _29531_, _29530_);
  or (_29533_, _29532_, _02528_);
  or (_29535_, _29505_, _02888_);
  and (_29536_, _05090_, _03708_);
  or (_29537_, _29536_, _29535_);
  and (_29538_, _29537_, _02043_);
  and (_29539_, _29538_, _29533_);
  nor (_29540_, _11615_, _09673_);
  or (_29541_, _29540_, _29505_);
  and (_29542_, _29541_, _01602_);
  or (_29543_, _29542_, _01869_);
  or (_29544_, _29543_, _29539_);
  and (_29546_, _04672_, _03708_);
  or (_29547_, _29546_, _29505_);
  or (_29548_, _29547_, _01870_);
  and (_29549_, _29548_, _29544_);
  or (_29550_, _29549_, _02079_);
  and (_29551_, _11629_, _03845_);
  or (_29552_, _29505_, _02166_);
  or (_29553_, _29552_, _29551_);
  and (_29554_, _29553_, _02912_);
  and (_29555_, _29554_, _29550_);
  or (_29557_, _29555_, _29508_);
  and (_29558_, _29557_, _02176_);
  or (_29559_, _29505_, _03965_);
  and (_29560_, _29547_, _02072_);
  and (_29561_, _29560_, _29559_);
  or (_29562_, _29561_, _29558_);
  and (_29563_, _29562_, _02907_);
  and (_29564_, _29515_, _02177_);
  and (_29565_, _29564_, _29559_);
  or (_29566_, _29565_, _02071_);
  or (_29568_, _29566_, _29563_);
  nor (_29569_, _11628_, _09678_);
  or (_29570_, _29505_, _04788_);
  or (_29571_, _29570_, _29569_);
  and (_29572_, _29571_, _04793_);
  and (_29573_, _29572_, _29568_);
  nor (_29574_, _11634_, _09678_);
  or (_29575_, _29574_, _29505_);
  and (_29576_, _29575_, _02173_);
  or (_29577_, _29576_, _02201_);
  or (_29579_, _29577_, _29573_);
  or (_29580_, _29510_, _02303_);
  and (_29581_, _29580_, _01538_);
  and (_29582_, _29581_, _29579_);
  and (_29583_, _11685_, _03845_);
  or (_29584_, _29583_, _29505_);
  and (_29585_, _29584_, _01537_);
  or (_29586_, _29585_, _38088_);
  or (_29587_, _29586_, _29582_);
  and (_40346_, _29587_, _29504_);
  or (_29588_, _38087_, \oc8051_golden_model_1.TL1 [6]);
  and (_29589_, _29588_, _37580_);
  and (_29590_, _09673_, \oc8051_golden_model_1.TL1 [6]);
  and (_29591_, _11709_, _03845_);
  or (_29592_, _29591_, _29590_);
  and (_29593_, _29592_, _02167_);
  nor (_29594_, _03808_, _09678_);
  or (_29595_, _29594_, _29590_);
  or (_29596_, _29595_, _05249_);
  nor (_29597_, _11730_, _09678_);
  or (_29599_, _29597_, _29590_);
  or (_29600_, _29599_, _02814_);
  and (_29601_, _03708_, \oc8051_golden_model_1.ACC [6]);
  or (_29602_, _29601_, _29590_);
  and (_29603_, _29602_, _02817_);
  and (_29604_, _02818_, \oc8051_golden_model_1.TL1 [6]);
  or (_29605_, _29604_, _02001_);
  or (_29606_, _29605_, _29603_);
  and (_29607_, _29606_, _02840_);
  and (_29608_, _29607_, _29600_);
  and (_29610_, _29595_, _01999_);
  or (_29611_, _29610_, _29608_);
  and (_29612_, _29611_, _02021_);
  and (_29613_, _29602_, _02006_);
  or (_29614_, _29613_, _05994_);
  or (_29615_, _29614_, _29612_);
  and (_29616_, _29615_, _29596_);
  or (_29617_, _29616_, _02528_);
  or (_29618_, _29590_, _02888_);
  and (_29619_, _04861_, _03708_);
  or (_29622_, _29619_, _29618_);
  and (_29623_, _29622_, _02043_);
  and (_29624_, _29623_, _29617_);
  nor (_29625_, _11820_, _09673_);
  or (_29626_, _29625_, _29590_);
  and (_29627_, _29626_, _01602_);
  or (_29628_, _29627_, _01869_);
  or (_29629_, _29628_, _29624_);
  and (_29630_, _09920_, _03708_);
  or (_29631_, _29630_, _29590_);
  or (_29633_, _29631_, _01870_);
  and (_29634_, _29633_, _29629_);
  or (_29635_, _29634_, _02079_);
  and (_29636_, _11835_, _03845_);
  or (_29637_, _29590_, _02166_);
  or (_29638_, _29637_, _29636_);
  and (_29639_, _29638_, _02912_);
  and (_29640_, _29639_, _29635_);
  or (_29641_, _29640_, _29593_);
  and (_29642_, _29641_, _02176_);
  or (_29644_, _29590_, _03863_);
  and (_29645_, _29631_, _02072_);
  and (_29646_, _29645_, _29644_);
  or (_29647_, _29646_, _29642_);
  and (_29648_, _29647_, _02907_);
  and (_29649_, _29602_, _02177_);
  and (_29650_, _29649_, _29644_);
  or (_29651_, _29650_, _02071_);
  or (_29652_, _29651_, _29648_);
  nor (_29653_, _11833_, _09678_);
  or (_29655_, _29590_, _04788_);
  or (_29656_, _29655_, _29653_);
  and (_29657_, _29656_, _04793_);
  and (_29658_, _29657_, _29652_);
  nor (_29659_, _11708_, _09678_);
  or (_29660_, _29659_, _29590_);
  and (_29661_, _29660_, _02173_);
  or (_29662_, _29661_, _02201_);
  or (_29663_, _29662_, _29658_);
  or (_29664_, _29599_, _02303_);
  and (_29666_, _29664_, _01538_);
  and (_29667_, _29666_, _29663_);
  and (_29668_, _11887_, _03845_);
  or (_29669_, _29668_, _29590_);
  and (_29670_, _29669_, _01537_);
  or (_29671_, _29670_, _38088_);
  or (_29672_, _29671_, _29667_);
  and (_40347_, _29672_, _29589_);
  and (_29673_, _38088_, \oc8051_golden_model_1.TMOD [0]);
  nor (_29674_, _04106_, _09752_);
  and (_29676_, _09752_, \oc8051_golden_model_1.TMOD [0]);
  and (_29677_, _03726_, _04562_);
  or (_29678_, _29677_, _29676_);
  nand (_29679_, _29678_, _02072_);
  nor (_29680_, _29679_, _29674_);
  and (_29681_, _03726_, \oc8051_golden_model_1.ACC [0]);
  or (_29682_, _29681_, _29676_);
  and (_29683_, _29682_, _02006_);
  or (_29684_, _29683_, _05994_);
  or (_29685_, _29676_, _29674_);
  and (_29687_, _29685_, _02001_);
  and (_29688_, _02818_, \oc8051_golden_model_1.TMOD [0]);
  and (_29689_, _29682_, _02817_);
  or (_29690_, _29689_, _29688_);
  and (_29691_, _29690_, _02814_);
  or (_29692_, _29691_, _01999_);
  or (_29693_, _29692_, _29687_);
  and (_29694_, _29693_, _02021_);
  or (_29695_, _29694_, _29684_);
  and (_29696_, _03726_, _03028_);
  or (_29698_, _29676_, _23851_);
  or (_29699_, _29698_, _29696_);
  and (_29700_, _29699_, _29695_);
  or (_29701_, _29700_, _02528_);
  and (_29702_, _04952_, _03726_);
  or (_29703_, _29676_, _02888_);
  or (_29704_, _29703_, _29702_);
  and (_29705_, _29704_, _29701_);
  or (_29706_, _29705_, _01602_);
  nor (_29707_, _10600_, _09752_);
  or (_29709_, _29707_, _29676_);
  or (_29710_, _29709_, _02043_);
  and (_29711_, _29710_, _01870_);
  and (_29712_, _29711_, _29706_);
  and (_29713_, _29678_, _01869_);
  or (_29714_, _29713_, _02079_);
  or (_29715_, _29714_, _29712_);
  and (_29716_, _10614_, _03726_);
  or (_29717_, _29716_, _29676_);
  or (_29718_, _29717_, _02166_);
  and (_29720_, _29718_, _29715_);
  or (_29721_, _29720_, _02167_);
  and (_29722_, _10620_, _03726_);
  or (_29723_, _29676_, _02912_);
  or (_29724_, _29723_, _29722_);
  and (_29725_, _29724_, _02176_);
  and (_29726_, _29725_, _29721_);
  or (_29727_, _29726_, _29680_);
  and (_29728_, _29727_, _02907_);
  or (_29729_, _29676_, _04106_);
  and (_29731_, _29682_, _02177_);
  and (_29732_, _29731_, _29729_);
  or (_29733_, _29732_, _02071_);
  or (_29734_, _29733_, _29728_);
  nor (_29735_, _10613_, _09752_);
  or (_29736_, _29676_, _04788_);
  or (_29737_, _29736_, _29735_);
  and (_29738_, _29737_, _04793_);
  and (_29739_, _29738_, _29734_);
  nor (_29740_, _10619_, _09752_);
  or (_29742_, _29740_, _29676_);
  and (_29743_, _29742_, _02173_);
  or (_29744_, _29743_, _15577_);
  or (_29745_, _29744_, _29739_);
  or (_29746_, _29685_, _02743_);
  and (_29747_, _29746_, _38087_);
  and (_29748_, _29747_, _29745_);
  or (_29749_, _29748_, _29673_);
  and (_40349_, _29749_, _37580_);
  and (_29750_, _38088_, \oc8051_golden_model_1.TMOD [1]);
  or (_29752_, _03726_, \oc8051_golden_model_1.TMOD [1]);
  and (_29753_, _10698_, _03726_);
  not (_29754_, _29753_);
  and (_29755_, _29754_, _29752_);
  or (_29756_, _29755_, _02814_);
  nand (_29757_, _03726_, _01613_);
  and (_29758_, _29757_, _29752_);
  and (_29759_, _29758_, _02817_);
  and (_29760_, _02818_, \oc8051_golden_model_1.TMOD [1]);
  or (_29761_, _29760_, _02001_);
  or (_29763_, _29761_, _29759_);
  and (_29764_, _29763_, _02840_);
  and (_29765_, _29764_, _29756_);
  nand (_29766_, _03726_, _02811_);
  and (_29767_, _29766_, _29752_);
  and (_29768_, _29767_, _01999_);
  or (_29769_, _29768_, _29765_);
  and (_29770_, _29769_, _02021_);
  and (_29771_, _29758_, _02006_);
  or (_29772_, _29771_, _05994_);
  or (_29774_, _29772_, _29770_);
  or (_29775_, _29767_, _05249_);
  and (_29776_, _29775_, _02888_);
  and (_29777_, _29776_, _29774_);
  or (_29778_, _04907_, _09752_);
  and (_29779_, _29752_, _02528_);
  and (_29780_, _29779_, _29778_);
  or (_29781_, _29780_, _29777_);
  and (_29782_, _29781_, _02043_);
  nand (_29783_, _10802_, _03726_);
  and (_29785_, _29752_, _01602_);
  and (_29786_, _29785_, _29783_);
  or (_29787_, _29786_, _29782_);
  and (_29788_, _29787_, _01870_);
  nand (_29789_, _03726_, _02687_);
  and (_29790_, _29752_, _01869_);
  and (_29791_, _29790_, _29789_);
  or (_29792_, _29791_, _29788_);
  and (_29793_, _29792_, _02166_);
  or (_29794_, _10816_, _09752_);
  and (_29796_, _29752_, _02079_);
  and (_29797_, _29796_, _29794_);
  or (_29798_, _29797_, _29793_);
  and (_29799_, _29798_, _02912_);
  or (_29800_, _10822_, _09752_);
  and (_29801_, _29752_, _02167_);
  and (_29802_, _29801_, _29800_);
  or (_29803_, _29802_, _29799_);
  and (_29804_, _29803_, _02176_);
  or (_29805_, _10692_, _09752_);
  and (_29807_, _29752_, _02072_);
  and (_29808_, _29807_, _29805_);
  or (_29809_, _29808_, _29804_);
  and (_29810_, _29809_, _02907_);
  and (_29811_, _09752_, \oc8051_golden_model_1.TMOD [1]);
  or (_29812_, _29811_, _04058_);
  and (_29813_, _29758_, _02177_);
  and (_29814_, _29813_, _29812_);
  or (_29815_, _29814_, _29810_);
  and (_29816_, _29815_, _02174_);
  or (_29818_, _29757_, _04058_);
  and (_29819_, _29752_, _02173_);
  and (_29820_, _29819_, _29818_);
  or (_29821_, _29820_, _02201_);
  or (_29822_, _29789_, _04058_);
  and (_29823_, _29752_, _02071_);
  and (_29824_, _29823_, _29822_);
  or (_29825_, _29824_, _29821_);
  or (_29826_, _29825_, _29816_);
  or (_29827_, _29755_, _02303_);
  and (_29829_, _29827_, _29826_);
  or (_29830_, _29829_, _01537_);
  or (_29831_, _29811_, _01538_);
  or (_29832_, _29831_, _29753_);
  and (_29833_, _29832_, _38087_);
  and (_29834_, _29833_, _29830_);
  or (_29835_, _29834_, _29750_);
  and (_40350_, _29835_, _37580_);
  and (_29836_, _38088_, \oc8051_golden_model_1.TMOD [2]);
  and (_29837_, _09752_, \oc8051_golden_model_1.TMOD [2]);
  nor (_29839_, _11019_, _09752_);
  or (_29840_, _29839_, _29837_);
  and (_29841_, _29840_, _02173_);
  nor (_29842_, _09752_, _03455_);
  or (_29843_, _29842_, _29837_);
  or (_29844_, _29843_, _05249_);
  nor (_29845_, _10905_, _09752_);
  or (_29846_, _29845_, _29837_);
  and (_29847_, _29846_, _02001_);
  and (_29848_, _02818_, \oc8051_golden_model_1.TMOD [2]);
  and (_29850_, _03726_, \oc8051_golden_model_1.ACC [2]);
  or (_29851_, _29850_, _29837_);
  and (_29852_, _29851_, _02817_);
  or (_29853_, _29852_, _29848_);
  and (_29854_, _29853_, _02814_);
  or (_29855_, _29854_, _01999_);
  or (_29856_, _29855_, _29847_);
  or (_29857_, _29843_, _02840_);
  and (_29858_, _29857_, _02021_);
  and (_29859_, _29858_, _29856_);
  and (_29861_, _29851_, _02006_);
  or (_29862_, _29861_, _05994_);
  or (_29863_, _29862_, _29859_);
  and (_29864_, _29863_, _29844_);
  or (_29865_, _29864_, _02528_);
  and (_29866_, _05043_, _03726_);
  or (_29867_, _29837_, _02888_);
  or (_29868_, _29867_, _29866_);
  and (_29869_, _29868_, _29865_);
  or (_29870_, _29869_, _01602_);
  nor (_29871_, _11000_, _09752_);
  or (_29872_, _29871_, _29837_);
  or (_29873_, _29872_, _02043_);
  and (_29874_, _29873_, _01870_);
  and (_29875_, _29874_, _29870_);
  and (_29876_, _03726_, _04724_);
  or (_29877_, _29876_, _29837_);
  and (_29878_, _29877_, _01869_);
  or (_29879_, _29878_, _02079_);
  or (_29880_, _29879_, _29875_);
  and (_29882_, _11014_, _03726_);
  or (_29883_, _29882_, _29837_);
  or (_29884_, _29883_, _02166_);
  and (_29885_, _29884_, _29880_);
  or (_29886_, _29885_, _02167_);
  and (_29887_, _11020_, _03726_);
  or (_29888_, _29837_, _02912_);
  or (_29889_, _29888_, _29887_);
  and (_29890_, _29889_, _02176_);
  and (_29891_, _29890_, _29886_);
  or (_29893_, _29837_, _04156_);
  and (_29894_, _29877_, _02072_);
  and (_29895_, _29894_, _29893_);
  or (_29896_, _29895_, _29891_);
  and (_29897_, _29896_, _02907_);
  and (_29898_, _29851_, _02177_);
  and (_29899_, _29898_, _29893_);
  or (_29900_, _29899_, _02071_);
  or (_29901_, _29900_, _29897_);
  nor (_29902_, _11013_, _09752_);
  or (_29904_, _29837_, _04788_);
  or (_29905_, _29904_, _29902_);
  and (_29906_, _29905_, _04793_);
  and (_29907_, _29906_, _29901_);
  or (_29908_, _29907_, _29841_);
  and (_29909_, _29908_, _02303_);
  and (_29910_, _29846_, _02201_);
  or (_29911_, _29910_, _01537_);
  or (_29912_, _29911_, _29909_);
  and (_29913_, _11072_, _03726_);
  or (_29915_, _29837_, _01538_);
  or (_29916_, _29915_, _29913_);
  and (_29917_, _29916_, _38087_);
  and (_29918_, _29917_, _29912_);
  or (_29919_, _29918_, _29836_);
  and (_40351_, _29919_, _37580_);
  or (_29920_, _38087_, \oc8051_golden_model_1.TMOD [3]);
  and (_29921_, _29920_, _37580_);
  and (_29922_, _09752_, \oc8051_golden_model_1.TMOD [3]);
  and (_29923_, _11094_, _03726_);
  or (_29925_, _29923_, _29922_);
  and (_29926_, _29925_, _02167_);
  nor (_29927_, _11101_, _09752_);
  or (_29928_, _29927_, _29922_);
  or (_29929_, _29928_, _02814_);
  and (_29930_, _03726_, \oc8051_golden_model_1.ACC [3]);
  or (_29931_, _29930_, _29922_);
  and (_29932_, _29931_, _02817_);
  and (_29933_, _02818_, \oc8051_golden_model_1.TMOD [3]);
  or (_29934_, _29933_, _02001_);
  or (_29936_, _29934_, _29932_);
  and (_29937_, _29936_, _02840_);
  and (_29938_, _29937_, _29929_);
  nor (_29939_, _09752_, _03268_);
  or (_29940_, _29939_, _29922_);
  and (_29941_, _29940_, _01999_);
  or (_29942_, _29941_, _29938_);
  and (_29943_, _29942_, _02021_);
  and (_29944_, _29931_, _02006_);
  or (_29945_, _29944_, _05994_);
  or (_29947_, _29945_, _29943_);
  or (_29948_, _29940_, _05249_);
  and (_29949_, _29948_, _29947_);
  or (_29950_, _29949_, _02528_);
  and (_29951_, _04998_, _03726_);
  or (_29952_, _29922_, _02888_);
  or (_29953_, _29952_, _29951_);
  and (_29954_, _29953_, _02043_);
  and (_29955_, _29954_, _29950_);
  nor (_29956_, _11206_, _09752_);
  or (_29958_, _29956_, _29922_);
  and (_29959_, _29958_, _01602_);
  or (_29960_, _29959_, _01869_);
  or (_29961_, _29960_, _29955_);
  and (_29962_, _03726_, _04678_);
  or (_29963_, _29962_, _29922_);
  or (_29964_, _29963_, _01870_);
  and (_29965_, _29964_, _29961_);
  or (_29966_, _29965_, _02079_);
  and (_29967_, _11222_, _03726_);
  or (_29969_, _29922_, _02166_);
  or (_29970_, _29969_, _29967_);
  and (_29971_, _29970_, _02912_);
  and (_29972_, _29971_, _29966_);
  or (_29973_, _29972_, _29926_);
  and (_29974_, _29973_, _02176_);
  or (_29975_, _29922_, _04014_);
  and (_29976_, _29963_, _02072_);
  and (_29977_, _29976_, _29975_);
  or (_29978_, _29977_, _29974_);
  and (_29980_, _29978_, _02907_);
  and (_29981_, _29931_, _02177_);
  and (_29982_, _29981_, _29975_);
  or (_29983_, _29982_, _02071_);
  or (_29984_, _29983_, _29980_);
  nor (_29985_, _11220_, _09752_);
  or (_29986_, _29922_, _04788_);
  or (_29987_, _29986_, _29985_);
  and (_29988_, _29987_, _04793_);
  and (_29989_, _29988_, _29984_);
  nor (_29991_, _11093_, _09752_);
  or (_29992_, _29991_, _29922_);
  and (_29993_, _29992_, _02173_);
  or (_29994_, _29993_, _02201_);
  or (_29995_, _29994_, _29989_);
  or (_29996_, _29928_, _02303_);
  and (_29997_, _29996_, _01538_);
  and (_29998_, _29997_, _29995_);
  and (_29999_, _11273_, _03726_);
  or (_30000_, _29999_, _29922_);
  and (_30002_, _30000_, _01537_);
  or (_30003_, _30002_, _38088_);
  or (_30004_, _30003_, _29998_);
  and (_40352_, _30004_, _29921_);
  or (_30005_, _38087_, \oc8051_golden_model_1.TMOD [4]);
  and (_30006_, _30005_, _37580_);
  and (_30007_, _09752_, \oc8051_golden_model_1.TMOD [4]);
  and (_30008_, _11431_, _03726_);
  or (_30009_, _30008_, _30007_);
  and (_30010_, _30009_, _02167_);
  nor (_30011_, _04211_, _09752_);
  or (_30012_, _30011_, _30007_);
  or (_30013_, _30012_, _05249_);
  nor (_30014_, _11317_, _09752_);
  or (_30015_, _30014_, _30007_);
  or (_30016_, _30015_, _02814_);
  and (_30017_, _03726_, \oc8051_golden_model_1.ACC [4]);
  or (_30018_, _30017_, _30007_);
  and (_30019_, _30018_, _02817_);
  and (_30020_, _02818_, \oc8051_golden_model_1.TMOD [4]);
  or (_30022_, _30020_, _02001_);
  or (_30023_, _30022_, _30019_);
  and (_30024_, _30023_, _02840_);
  and (_30025_, _30024_, _30016_);
  and (_30026_, _30012_, _01999_);
  or (_30027_, _30026_, _30025_);
  and (_30028_, _30027_, _02021_);
  and (_30029_, _30018_, _02006_);
  or (_30030_, _30029_, _05994_);
  or (_30031_, _30030_, _30028_);
  and (_30033_, _30031_, _30013_);
  or (_30034_, _30033_, _02528_);
  and (_30035_, _05135_, _03726_);
  or (_30036_, _30007_, _02888_);
  or (_30037_, _30036_, _30035_);
  and (_30038_, _30037_, _02043_);
  and (_30039_, _30038_, _30034_);
  nor (_30040_, _11411_, _09752_);
  or (_30041_, _30040_, _30007_);
  and (_30042_, _30041_, _01602_);
  or (_30044_, _30042_, _01869_);
  or (_30045_, _30044_, _30039_);
  and (_30046_, _04694_, _03726_);
  or (_30047_, _30046_, _30007_);
  or (_30048_, _30047_, _01870_);
  and (_30049_, _30048_, _30045_);
  or (_30050_, _30049_, _02079_);
  and (_30051_, _11425_, _03726_);
  or (_30052_, _30007_, _02166_);
  or (_30053_, _30052_, _30051_);
  and (_30055_, _30053_, _02912_);
  and (_30056_, _30055_, _30050_);
  or (_30057_, _30056_, _30010_);
  and (_30058_, _30057_, _02176_);
  or (_30059_, _30007_, _04258_);
  and (_30060_, _30047_, _02072_);
  and (_30061_, _30060_, _30059_);
  or (_30062_, _30061_, _30058_);
  and (_30063_, _30062_, _02907_);
  and (_30064_, _30018_, _02177_);
  and (_30066_, _30064_, _30059_);
  or (_30067_, _30066_, _02071_);
  or (_30068_, _30067_, _30063_);
  nor (_30069_, _11424_, _09752_);
  or (_30070_, _30007_, _04788_);
  or (_30071_, _30070_, _30069_);
  and (_30072_, _30071_, _04793_);
  and (_30073_, _30072_, _30068_);
  nor (_30074_, _11430_, _09752_);
  or (_30075_, _30074_, _30007_);
  and (_30077_, _30075_, _02173_);
  or (_30078_, _30077_, _02201_);
  or (_30079_, _30078_, _30073_);
  or (_30080_, _30015_, _02303_);
  and (_30081_, _30080_, _01538_);
  and (_30082_, _30081_, _30079_);
  and (_30083_, _11487_, _03726_);
  or (_30084_, _30083_, _30007_);
  and (_30085_, _30084_, _01537_);
  or (_30086_, _30085_, _38088_);
  or (_30088_, _30086_, _30082_);
  and (_40353_, _30088_, _30006_);
  or (_30089_, _38087_, \oc8051_golden_model_1.TMOD [5]);
  and (_30090_, _30089_, _37580_);
  and (_30091_, _09752_, \oc8051_golden_model_1.TMOD [5]);
  and (_30092_, _11635_, _03726_);
  or (_30093_, _30092_, _30091_);
  and (_30094_, _30093_, _02167_);
  nor (_30095_, _03916_, _09752_);
  or (_30096_, _30095_, _30091_);
  or (_30098_, _30096_, _05249_);
  nor (_30099_, _11525_, _09752_);
  or (_30100_, _30099_, _30091_);
  or (_30101_, _30100_, _02814_);
  and (_30102_, _03726_, \oc8051_golden_model_1.ACC [5]);
  or (_30103_, _30102_, _30091_);
  and (_30104_, _30103_, _02817_);
  and (_30105_, _02818_, \oc8051_golden_model_1.TMOD [5]);
  or (_30106_, _30105_, _02001_);
  or (_30107_, _30106_, _30104_);
  and (_30109_, _30107_, _02840_);
  and (_30110_, _30109_, _30101_);
  and (_30111_, _30096_, _01999_);
  or (_30112_, _30111_, _30110_);
  and (_30113_, _30112_, _02021_);
  and (_30114_, _30103_, _02006_);
  or (_30115_, _30114_, _05994_);
  or (_30116_, _30115_, _30113_);
  and (_30117_, _30116_, _30098_);
  or (_30118_, _30117_, _02528_);
  and (_30120_, _05090_, _03726_);
  or (_30121_, _30091_, _02888_);
  or (_30122_, _30121_, _30120_);
  and (_30123_, _30122_, _02043_);
  and (_30124_, _30123_, _30118_);
  nor (_30125_, _11615_, _09752_);
  or (_30126_, _30125_, _30091_);
  and (_30127_, _30126_, _01602_);
  or (_30128_, _30127_, _01869_);
  or (_30129_, _30128_, _30124_);
  and (_30131_, _04672_, _03726_);
  or (_30132_, _30131_, _30091_);
  or (_30133_, _30132_, _01870_);
  and (_30134_, _30133_, _30129_);
  or (_30135_, _30134_, _02079_);
  and (_30136_, _11629_, _03726_);
  or (_30137_, _30091_, _02166_);
  or (_30138_, _30137_, _30136_);
  and (_30139_, _30138_, _02912_);
  and (_30140_, _30139_, _30135_);
  or (_30142_, _30140_, _30094_);
  and (_30143_, _30142_, _02176_);
  or (_30144_, _30091_, _03965_);
  and (_30145_, _30132_, _02072_);
  and (_30146_, _30145_, _30144_);
  or (_30147_, _30146_, _30143_);
  and (_30148_, _30147_, _02907_);
  and (_30149_, _30103_, _02177_);
  and (_30150_, _30149_, _30144_);
  or (_30151_, _30150_, _02071_);
  or (_30153_, _30151_, _30148_);
  nor (_30154_, _11628_, _09752_);
  or (_30155_, _30091_, _04788_);
  or (_30156_, _30155_, _30154_);
  and (_30157_, _30156_, _04793_);
  and (_30158_, _30157_, _30153_);
  nor (_30159_, _11634_, _09752_);
  or (_30160_, _30159_, _30091_);
  and (_30161_, _30160_, _02173_);
  or (_30162_, _30161_, _02201_);
  or (_30164_, _30162_, _30158_);
  or (_30165_, _30100_, _02303_);
  and (_30166_, _30165_, _01538_);
  and (_30167_, _30166_, _30164_);
  and (_30168_, _11685_, _03726_);
  or (_30169_, _30168_, _30091_);
  and (_30170_, _30169_, _01537_);
  or (_30171_, _30170_, _38088_);
  or (_30172_, _30171_, _30167_);
  and (_40354_, _30172_, _30090_);
  or (_30173_, _38087_, \oc8051_golden_model_1.TMOD [6]);
  and (_30174_, _30173_, _37580_);
  and (_30175_, _09752_, \oc8051_golden_model_1.TMOD [6]);
  and (_30176_, _11709_, _03726_);
  or (_30177_, _30176_, _30175_);
  and (_30178_, _30177_, _02167_);
  nor (_30179_, _11730_, _09752_);
  or (_30180_, _30179_, _30175_);
  or (_30181_, _30180_, _02814_);
  and (_30182_, _03726_, \oc8051_golden_model_1.ACC [6]);
  or (_30184_, _30182_, _30175_);
  and (_30185_, _30184_, _02817_);
  and (_30186_, _02818_, \oc8051_golden_model_1.TMOD [6]);
  or (_30187_, _30186_, _02001_);
  or (_30188_, _30187_, _30185_);
  and (_30189_, _30188_, _02840_);
  and (_30190_, _30189_, _30181_);
  nor (_30191_, _03808_, _09752_);
  or (_30192_, _30191_, _30175_);
  and (_30193_, _30192_, _01999_);
  or (_30195_, _30193_, _30190_);
  and (_30196_, _30195_, _02021_);
  and (_30197_, _30184_, _02006_);
  or (_30198_, _30197_, _05994_);
  or (_30199_, _30198_, _30196_);
  or (_30200_, _30192_, _05249_);
  and (_30201_, _30200_, _30199_);
  or (_30202_, _30201_, _02528_);
  and (_30203_, _04861_, _03726_);
  or (_30204_, _30175_, _02888_);
  or (_30206_, _30204_, _30203_);
  and (_30207_, _30206_, _02043_);
  and (_30208_, _30207_, _30202_);
  nor (_30209_, _11820_, _09752_);
  or (_30210_, _30209_, _30175_);
  and (_30211_, _30210_, _01602_);
  or (_30212_, _30211_, _01869_);
  or (_30213_, _30212_, _30208_);
  and (_30214_, _09920_, _03726_);
  or (_30215_, _30214_, _30175_);
  or (_30217_, _30215_, _01870_);
  and (_30218_, _30217_, _30213_);
  or (_30219_, _30218_, _02079_);
  and (_30220_, _11835_, _03726_);
  or (_30221_, _30175_, _02166_);
  or (_30222_, _30221_, _30220_);
  and (_30223_, _30222_, _02912_);
  and (_30224_, _30223_, _30219_);
  or (_30225_, _30224_, _30178_);
  and (_30226_, _30225_, _02176_);
  or (_30228_, _30175_, _03863_);
  and (_30229_, _30215_, _02072_);
  and (_30230_, _30229_, _30228_);
  or (_30231_, _30230_, _30226_);
  and (_30232_, _30231_, _02907_);
  and (_30233_, _30184_, _02177_);
  and (_30234_, _30233_, _30228_);
  or (_30235_, _30234_, _02071_);
  or (_30236_, _30235_, _30232_);
  nor (_30237_, _11833_, _09752_);
  or (_30239_, _30175_, _04788_);
  or (_30240_, _30239_, _30237_);
  and (_30241_, _30240_, _04793_);
  and (_30242_, _30241_, _30236_);
  nor (_30243_, _11708_, _09752_);
  or (_30244_, _30243_, _30175_);
  and (_30245_, _30244_, _02173_);
  or (_30246_, _30245_, _02201_);
  or (_30247_, _30246_, _30242_);
  or (_30248_, _30180_, _02303_);
  and (_30250_, _30248_, _01538_);
  and (_30251_, _30250_, _30247_);
  and (_30252_, _11887_, _03726_);
  or (_30253_, _30252_, _30175_);
  and (_30254_, _30253_, _01537_);
  or (_30255_, _30254_, _38088_);
  or (_30256_, _30255_, _30251_);
  and (_40355_, _30256_, _30174_);
  or (_30257_, _38087_, \oc8051_golden_model_1.PC [0]);
  and (_30258_, _30257_, _37580_);
  nand (_30260_, _08439_, \oc8051_golden_model_1.PC [0]);
  and (_30261_, _02568_, \oc8051_golden_model_1.PC [0]);
  nor (_30262_, _30261_, _09946_);
  or (_30263_, _30262_, _08439_);
  and (_30264_, _30263_, _30260_);
  and (_30265_, _30264_, _01860_);
  and (_30266_, _10438_, _10442_);
  or (_30267_, _30266_, _01280_);
  and (_30268_, _09844_, _07305_);
  or (_30269_, _30268_, _01280_);
  and (_30271_, _09846_, _07176_);
  not (_30272_, _01648_);
  nor (_30273_, _02568_, _30272_);
  and (_30274_, _09861_, _04788_);
  nor (_30275_, _02568_, _01633_);
  nand (_30276_, _02568_, _01638_);
  and (_30277_, _30276_, _10311_);
  and (_30278_, _08498_, _01280_);
  not (_30279_, _08498_);
  and (_30280_, _30262_, _30279_);
  or (_30282_, _30280_, _08494_);
  or (_30283_, _30282_, _30278_);
  and (_30284_, _01568_, _01562_);
  nor (_30285_, _30284_, _02568_);
  nor (_30286_, _06616_, _06629_);
  or (_30287_, _30286_, _01280_);
  and (_30288_, _30287_, _01568_);
  not (_30289_, _30286_);
  nor (_30290_, _21690_, _01280_);
  nand (_30291_, _21690_, _01280_);
  nand (_30293_, _30291_, _01562_);
  nor (_30294_, _30293_, _30290_);
  or (_30295_, _30294_, _30289_);
  and (_30296_, _30295_, _30288_);
  or (_30297_, _30296_, _04380_);
  or (_30298_, _30297_, _30285_);
  and (_30299_, _10107_, \oc8051_golden_model_1.PC [0]);
  and (_30300_, _02441_, _01280_);
  nor (_30301_, _30300_, _10055_);
  and (_30302_, _30301_, _10105_);
  or (_30304_, _30302_, _30299_);
  or (_30305_, _30304_, _04381_);
  and (_30306_, _30305_, _30298_);
  or (_30307_, _30306_, _01883_);
  nand (_30308_, _01883_, \oc8051_golden_model_1.PC [0]);
  and (_30309_, _30308_, _02814_);
  and (_30310_, _30309_, _30307_);
  not (_30311_, _09871_);
  or (_30312_, _09876_, _01280_);
  or (_30313_, _30262_, _09996_);
  and (_30315_, _30313_, _02001_);
  and (_30316_, _30315_, _30312_);
  or (_30317_, _30316_, _30311_);
  or (_30318_, _30317_, _30310_);
  or (_30319_, _09871_, _01280_);
  and (_30320_, _30319_, _01558_);
  and (_30321_, _30320_, _30318_);
  or (_30322_, _02568_, _01558_);
  and (_30323_, _10163_, _10156_);
  nand (_30324_, _30323_, _30322_);
  or (_30326_, _30324_, _30321_);
  or (_30327_, _30323_, _01280_);
  and (_30328_, _30327_, _01574_);
  and (_30329_, _30328_, _30326_);
  nor (_30330_, _02568_, _01574_);
  or (_30331_, _30330_, _08539_);
  or (_30332_, _30331_, _30329_);
  or (_30333_, _30262_, _08572_);
  nand (_30334_, _08572_, \oc8051_golden_model_1.PC [0]);
  and (_30335_, _30334_, _30333_);
  or (_30336_, _30335_, _08538_);
  and (_30337_, _30336_, _30332_);
  or (_30338_, _30337_, _08493_);
  and (_30339_, _30338_, _02444_);
  and (_30340_, _30339_, _30283_);
  and (_30341_, _08625_, _01280_);
  not (_30342_, _08625_);
  and (_30343_, _30262_, _30342_);
  or (_30344_, _30343_, _30341_);
  and (_30345_, _30344_, _01995_);
  or (_30347_, _30345_, _30340_);
  and (_30348_, _30347_, _02046_);
  nand (_30349_, _08664_, \oc8051_golden_model_1.PC [0]);
  or (_30350_, _30262_, _08664_);
  and (_30351_, _30350_, _02045_);
  and (_30352_, _30351_, _30349_);
  or (_30353_, _30352_, _08628_);
  or (_30354_, _30353_, _30348_);
  nand (_30355_, _08628_, \oc8051_golden_model_1.PC [0]);
  and (_30356_, _30355_, _01565_);
  and (_30358_, _30356_, _30354_);
  nor (_30359_, _02568_, _01565_);
  or (_30360_, _30359_, _10211_);
  or (_30361_, _30360_, _30358_);
  or (_30362_, _10207_, _01280_);
  and (_30363_, _30362_, _01572_);
  and (_30364_, _30363_, _30361_);
  or (_30365_, _02568_, _01572_);
  nor (_30366_, _10219_, _01549_);
  nand (_30367_, _30366_, _30365_);
  or (_30369_, _30367_, _30364_);
  or (_30370_, _30366_, _01280_);
  and (_30371_, _30370_, _04310_);
  and (_30372_, _30371_, _30369_);
  or (_30373_, _02568_, _04310_);
  nor (_30374_, _02080_, _01602_);
  and (_30375_, _30374_, _10245_);
  nand (_30376_, _30375_, _30373_);
  or (_30377_, _30376_, _30372_);
  not (_30378_, _01649_);
  or (_30380_, _30375_, _01280_);
  and (_30381_, _30380_, _30378_);
  and (_30382_, _30381_, _30377_);
  nor (_30383_, _02568_, _30378_);
  or (_30384_, _30383_, _10253_);
  or (_30385_, _30384_, _30382_);
  or (_30386_, _30301_, _10254_);
  and (_30387_, _30386_, _30385_);
  or (_30388_, _30387_, _01869_);
  nand (_30389_, _01869_, \oc8051_golden_model_1.PC [0]);
  and (_30391_, _10268_, _30389_);
  and (_30392_, _30391_, _30388_);
  and (_30393_, _10267_, _01703_);
  or (_30394_, _30393_, _01638_);
  or (_30395_, _30394_, _30392_);
  and (_30396_, _30395_, _30277_);
  and (_30397_, _10327_, _02166_);
  or (_30398_, _30301_, _07356_);
  nand (_30399_, _07356_, _01280_);
  and (_30400_, _30399_, _10310_);
  nand (_30402_, _30400_, _30398_);
  nand (_30403_, _30402_, _30397_);
  or (_30404_, _30403_, _30396_);
  or (_30405_, _30397_, _01280_);
  and (_30406_, _30405_, _22337_);
  and (_30407_, _30406_, _30404_);
  or (_30408_, _30301_, _10316_);
  or (_30409_, _07356_, \oc8051_golden_model_1.PC [0]);
  and (_30410_, _30409_, _10343_);
  and (_30411_, _30410_, _30408_);
  not (_30413_, _01645_);
  or (_30414_, _02568_, _30413_);
  nor (_30415_, _09863_, _02072_);
  nand (_30416_, _30415_, _30414_);
  or (_30417_, _30416_, _30411_);
  or (_30418_, _30417_, _30407_);
  or (_30419_, _30415_, _01280_);
  and (_30420_, _30419_, _01633_);
  and (_30421_, _30420_, _30418_);
  or (_30422_, _30421_, _30275_);
  and (_30424_, _30422_, _10364_);
  nor (_30425_, _06524_, _01280_);
  and (_30426_, _06524_, _01280_);
  or (_30427_, _30426_, _30425_);
  and (_30428_, _30427_, _10363_);
  nor (_30429_, _30428_, _30424_);
  nand (_30430_, _30429_, _30274_);
  or (_30431_, _30274_, _01280_);
  and (_30432_, _30431_, _30272_);
  and (_30433_, _30432_, _30430_);
  or (_30435_, _30433_, _30273_);
  and (_30436_, _30435_, _09849_);
  nor (_30437_, _06519_, _01280_);
  and (_30438_, _06519_, _01280_);
  or (_30439_, _30438_, _30437_);
  and (_30440_, _30439_, _09848_);
  nor (_30441_, _30440_, _30436_);
  nand (_30442_, _30441_, _30271_);
  or (_30443_, _30271_, _01280_);
  and (_30444_, _30443_, _09305_);
  and (_30446_, _30444_, _30442_);
  and (_30447_, _04952_, _02185_);
  or (_30448_, _30447_, _01636_);
  or (_30449_, _30448_, _30446_);
  nand (_30450_, _02568_, _01636_);
  and (_30451_, _30450_, _10403_);
  and (_30452_, _30451_, _30449_);
  or (_30453_, _30262_, _10408_);
  or (_30454_, _08439_, _01280_);
  and (_30455_, _30454_, _02083_);
  nand (_30457_, _30455_, _30453_);
  nand (_30458_, _30457_, _30268_);
  or (_30459_, _30458_, _30452_);
  and (_30460_, _30459_, _30269_);
  or (_30461_, _30460_, _01888_);
  or (_30462_, _04952_, _01889_);
  and (_30463_, _30462_, _10426_);
  and (_30464_, _30463_, _30461_);
  nor (_30465_, _02568_, _10426_);
  or (_30466_, _30465_, _30464_);
  and (_30468_, _30466_, _02202_);
  nand (_30469_, _30264_, _02082_);
  nand (_30470_, _30469_, _30266_);
  or (_30471_, _30470_, _30468_);
  and (_30472_, _30471_, _30267_);
  or (_30473_, _30472_, _03370_);
  nand (_30474_, _03370_, _02568_);
  and (_30475_, _30474_, _01887_);
  and (_30476_, _30475_, _30473_);
  or (_30477_, _30476_, _30265_);
  and (_30479_, _10461_, _10465_);
  and (_30480_, _30479_, _30477_);
  nor (_30481_, _02057_, _01651_);
  not (_30482_, _30481_);
  nor (_30483_, _30479_, \oc8051_golden_model_1.PC [0]);
  or (_30484_, _30483_, _30482_);
  or (_30485_, _30484_, _30480_);
  nand (_30486_, _30482_, _02568_);
  and (_30487_, _30486_, _10481_);
  and (_30488_, _30487_, _30485_);
  and (_30489_, _09829_, _01280_);
  or (_30490_, _30489_, _38088_);
  or (_30491_, _30490_, _30488_);
  and (_40358_, _30491_, _30258_);
  or (_30492_, _10465_, _01723_);
  nor (_30493_, _09948_, _09946_);
  nor (_30494_, _30493_, _09949_);
  or (_30495_, _30494_, _08439_);
  nand (_30496_, _08439_, _01723_);
  and (_30497_, _30496_, _30495_);
  and (_30499_, _30497_, _01860_);
  or (_30500_, _10442_, _01723_);
  not (_30501_, _02387_);
  nand (_30502_, _02718_, _01541_);
  and (_30503_, _30502_, _30501_);
  or (_30504_, _30503_, _01723_);
  and (_30505_, _02062_, _01652_);
  or (_30506_, _09861_, _01723_);
  nand (_30507_, _09863_, _01614_);
  or (_30508_, _10327_, _01723_);
  or (_30510_, _04757_, _01253_);
  nand (_30511_, _10219_, _01614_);
  nand (_30512_, _08628_, _01614_);
  or (_30513_, _30494_, _08572_);
  nand (_30514_, _08572_, _01723_);
  and (_30515_, _30514_, _30513_);
  or (_30516_, _30515_, _08538_);
  nor (_30517_, _02687_, _01574_);
  or (_30518_, _10163_, _01723_);
  nand (_30519_, _01883_, _01614_);
  or (_30521_, _10105_, _01253_);
  nor (_30522_, _10057_, _10055_);
  nor (_30523_, _30522_, _10058_);
  or (_30524_, _30523_, _10107_);
  and (_30525_, _30524_, _04380_);
  and (_30526_, _30525_, _30521_);
  nand (_30527_, _02687_, _02823_);
  nor (_30528_, _30290_, _02817_);
  or (_30529_, _30528_, _01253_);
  nand (_30530_, _30528_, _01253_);
  and (_30532_, _30530_, _30529_);
  nor (_30533_, _30532_, _02823_);
  nor (_30534_, _03122_, _01567_);
  or (_30535_, _30534_, _02353_);
  nor (_30536_, _30535_, _30533_);
  and (_30537_, _30536_, _30527_);
  nor (_30538_, _06620_, _02448_);
  nand (_30539_, _30535_, _01723_);
  nand (_30540_, _30539_, _30538_);
  or (_30541_, _30540_, _30537_);
  or (_30543_, _30538_, _01723_);
  and (_30544_, _30543_, _06618_);
  and (_30545_, _30544_, _30541_);
  and (_30546_, _02003_, _01253_);
  or (_30547_, _30546_, _06616_);
  or (_30548_, _30547_, _30545_);
  nand (_30549_, _06616_, _01614_);
  and (_30550_, _30549_, _30548_);
  or (_30551_, _30550_, _10140_);
  nand (_30552_, _02687_, _10140_);
  and (_30554_, _30552_, _04381_);
  and (_30555_, _30554_, _30551_);
  or (_30556_, _30555_, _01883_);
  or (_30557_, _30556_, _30526_);
  and (_30558_, _30557_, _30519_);
  or (_30559_, _30558_, _02001_);
  and (_30560_, _09996_, _01614_);
  and (_30561_, _30494_, _09876_);
  or (_30562_, _30561_, _30560_);
  or (_30563_, _30562_, _02814_);
  and (_30565_, _30563_, _30559_);
  or (_30566_, _30565_, _30311_);
  or (_30567_, _09871_, _01723_);
  and (_30568_, _30567_, _02024_);
  and (_30569_, _30568_, _30566_);
  and (_30570_, _02007_, _01253_);
  or (_30571_, _30570_, _03279_);
  or (_30572_, _30571_, _30569_);
  nand (_30573_, _02687_, _03279_);
  and (_30574_, _30573_, _02840_);
  and (_30576_, _30574_, _30572_);
  nand (_30577_, _01999_, _01253_);
  nand (_30578_, _30577_, _10156_);
  or (_30579_, _30578_, _30576_);
  or (_30580_, _10156_, _01723_);
  and (_30581_, _30580_, _02021_);
  and (_30582_, _30581_, _30579_);
  nand (_30583_, _02006_, _01253_);
  nand (_30584_, _30583_, _10163_);
  or (_30585_, _30584_, _30582_);
  and (_30587_, _30585_, _30518_);
  or (_30588_, _30587_, _01997_);
  nand (_30589_, _01997_, \oc8051_golden_model_1.PC [1]);
  and (_30590_, _30589_, _01574_);
  and (_30591_, _30590_, _30588_);
  or (_30592_, _30591_, _30517_);
  and (_30593_, _30592_, _01880_);
  nand (_30594_, _01878_, _01253_);
  nand (_30595_, _30594_, _08538_);
  or (_30596_, _30595_, _30593_);
  and (_30598_, _30596_, _30516_);
  or (_30599_, _30598_, _08493_);
  and (_30600_, _08498_, _01614_);
  and (_30601_, _30494_, _30279_);
  or (_30602_, _30601_, _08494_);
  or (_30603_, _30602_, _30600_);
  and (_30604_, _30603_, _30599_);
  or (_30605_, _30604_, _01995_);
  and (_30606_, _30494_, _30342_);
  and (_30607_, _08625_, _01614_);
  or (_30609_, _30607_, _02444_);
  or (_30610_, _30609_, _30606_);
  and (_30611_, _30610_, _02046_);
  and (_30612_, _30611_, _30605_);
  nand (_30613_, _08664_, _01723_);
  or (_30614_, _30494_, _08664_);
  and (_30615_, _30614_, _02045_);
  and (_30616_, _30615_, _30613_);
  or (_30617_, _30616_, _08628_);
  or (_30618_, _30617_, _30612_);
  and (_30620_, _30618_, _30512_);
  or (_30621_, _30620_, _01991_);
  nand (_30622_, _01991_, \oc8051_golden_model_1.PC [1]);
  and (_30623_, _30622_, _01565_);
  and (_30624_, _30623_, _30621_);
  nor (_30625_, _02687_, _01565_);
  and (_30626_, _02358_, _01965_);
  nor (_30627_, _30626_, _03489_);
  and (_30628_, _02340_, _01965_);
  nor (_30629_, _01992_, _30628_);
  and (_30631_, _30629_, _30627_);
  and (_30632_, _30631_, _04403_);
  not (_30633_, _30632_);
  or (_30634_, _30633_, _30625_);
  or (_30635_, _30634_, _30624_);
  or (_30636_, _30632_, _01253_);
  and (_30637_, _30636_, _10205_);
  and (_30638_, _30637_, _30635_);
  nand (_30639_, _10204_, _01723_);
  nand (_30640_, _30639_, _10206_);
  or (_30642_, _30640_, _30638_);
  or (_30643_, _10206_, _01723_);
  and (_30644_, _30643_, _08249_);
  and (_30645_, _30644_, _30642_);
  and (_30646_, _01967_, _01253_);
  or (_30647_, _30646_, _10213_);
  or (_30648_, _30647_, _30645_);
  nand (_30649_, _02687_, _10213_);
  and (_30650_, _30649_, _08248_);
  and (_30651_, _30650_, _30648_);
  and (_30652_, _01966_, _01253_);
  or (_30653_, _30652_, _10219_);
  or (_30654_, _30653_, _30651_);
  and (_30655_, _30654_, _30511_);
  or (_30656_, _30655_, _06776_);
  or (_30657_, _06775_, _01253_);
  and (_30658_, _30657_, _01550_);
  and (_30659_, _30658_, _30656_);
  and (_30660_, _01723_, _01549_);
  or (_30661_, _30660_, _01875_);
  or (_30663_, _30661_, _30659_);
  nand (_30664_, _01875_, \oc8051_golden_model_1.PC [1]);
  and (_30665_, _30664_, _30663_);
  or (_30666_, _30665_, _01604_);
  nand (_30667_, _02687_, _01604_);
  and (_30668_, _30667_, _07401_);
  and (_30669_, _30668_, _30666_);
  nand (_30670_, _02080_, _01614_);
  nand (_30671_, _30670_, _09211_);
  or (_30672_, _30671_, _30669_);
  or (_30674_, _09211_, _01253_);
  and (_30675_, _30674_, _02043_);
  and (_30676_, _30675_, _30672_);
  nand (_30677_, _01614_, _01602_);
  nand (_30678_, _30677_, _10245_);
  or (_30679_, _30678_, _30676_);
  not (_30680_, _01959_);
  or (_30681_, _10245_, _01723_);
  and (_30682_, _30681_, _30680_);
  and (_30683_, _30682_, _30679_);
  and (_30685_, _01959_, _01253_);
  or (_30686_, _30685_, _01649_);
  or (_30687_, _30686_, _30683_);
  nand (_30688_, _02687_, _01649_);
  and (_30689_, _30688_, _10254_);
  and (_30690_, _30689_, _30687_);
  and (_30691_, _30523_, _10253_);
  or (_30692_, _30691_, _04758_);
  or (_30693_, _30692_, _30690_);
  and (_30694_, _30693_, _30510_);
  or (_30696_, _30694_, _01869_);
  nand (_30697_, _01869_, _01723_);
  and (_30698_, _30697_, _06985_);
  and (_30699_, _30698_, _30696_);
  and (_30700_, _06984_, _01253_);
  or (_30701_, _30700_, _10267_);
  or (_30702_, _30701_, _30699_);
  or (_30703_, _10268_, _01721_);
  and (_30704_, _30703_, _02576_);
  and (_30705_, _30704_, _30702_);
  and (_30707_, _01958_, _01253_);
  or (_30708_, _30707_, _01638_);
  or (_30709_, _30708_, _30705_);
  nand (_30710_, _02687_, _01638_);
  and (_30711_, _30710_, _10311_);
  and (_30712_, _30711_, _30709_);
  or (_30713_, _30523_, _07356_);
  nand (_30714_, _07356_, \oc8051_golden_model_1.PC [1]);
  and (_30715_, _30714_, _10310_);
  and (_30716_, _30715_, _30713_);
  or (_30718_, _30716_, _10331_);
  or (_30719_, _30718_, _30712_);
  and (_30720_, _30719_, _30508_);
  or (_30721_, _30720_, _10330_);
  or (_30722_, _10329_, _01253_);
  and (_30723_, _30722_, _02166_);
  and (_30724_, _30723_, _30721_);
  and (_30725_, _02079_, _01614_);
  or (_30726_, _30725_, _02167_);
  or (_30727_, _30726_, _30724_);
  nand (_30729_, _02167_, \oc8051_golden_model_1.PC [1]);
  and (_30730_, _30729_, _30727_);
  or (_30731_, _30730_, _01645_);
  nand (_30732_, _02687_, _01645_);
  and (_30733_, _30732_, _10344_);
  and (_30734_, _30733_, _30731_);
  or (_30735_, _30523_, _10316_);
  or (_30736_, _07356_, _01253_);
  and (_30737_, _30736_, _10343_);
  and (_30738_, _30737_, _30735_);
  or (_30740_, _30738_, _09863_);
  or (_30741_, _30740_, _30734_);
  and (_30742_, _30741_, _30507_);
  or (_30743_, _30742_, _07042_);
  or (_30744_, _07041_, _01253_);
  and (_30745_, _30744_, _02176_);
  and (_30746_, _30745_, _30743_);
  and (_30747_, _02072_, _01614_);
  or (_30748_, _30747_, _02177_);
  or (_30749_, _30748_, _30746_);
  nand (_30751_, _02177_, \oc8051_golden_model_1.PC [1]);
  and (_30752_, _30751_, _30749_);
  or (_30753_, _30752_, _01632_);
  nand (_30754_, _02687_, _01632_);
  and (_30755_, _30754_, _10364_);
  and (_30756_, _30755_, _30753_);
  or (_30757_, _30523_, \oc8051_golden_model_1.PSW [7]);
  nand (_30758_, \oc8051_golden_model_1.PSW [7], \oc8051_golden_model_1.PC [1]);
  and (_30759_, _30758_, _10363_);
  and (_30760_, _30759_, _30757_);
  or (_30762_, _30760_, _10368_);
  or (_30763_, _30762_, _30756_);
  and (_30764_, _30763_, _30506_);
  or (_30765_, _30764_, _09854_);
  or (_30766_, _09853_, _01253_);
  and (_30767_, _30766_, _04788_);
  and (_30768_, _30767_, _30765_);
  and (_30769_, _02071_, _01614_);
  or (_30770_, _30769_, _02173_);
  or (_30771_, _30770_, _30768_);
  nand (_30773_, _02173_, \oc8051_golden_model_1.PC [1]);
  and (_30774_, _30773_, _30771_);
  or (_30775_, _30774_, _01648_);
  nand (_30776_, _02687_, _01648_);
  and (_30777_, _30776_, _09849_);
  and (_30778_, _30777_, _30775_);
  or (_30779_, _30523_, _06518_);
  or (_30780_, \oc8051_golden_model_1.PSW [7], _01253_);
  and (_30781_, _30780_, _09848_);
  and (_30782_, _30781_, _30779_);
  or (_30784_, _30782_, _30778_);
  and (_30785_, _30784_, _09846_);
  nor (_30786_, _09846_, _01614_);
  or (_30787_, _30786_, _07146_);
  or (_30788_, _30787_, _30785_);
  or (_30789_, _07145_, _01253_);
  and (_30790_, _30789_, _07176_);
  and (_30791_, _30790_, _30788_);
  and (_30792_, _07175_, _01723_);
  or (_30793_, _30792_, _02185_);
  or (_30795_, _30793_, _30791_);
  or (_30796_, _04907_, _09305_);
  and (_30797_, _30796_, _30795_);
  or (_30798_, _30797_, _01636_);
  nand (_30799_, _02687_, _01636_);
  and (_30800_, _30799_, _10403_);
  and (_30801_, _30800_, _30798_);
  nor (_30802_, _08439_, _01723_);
  and (_30803_, _30494_, _08439_);
  or (_30804_, _30803_, _30802_);
  and (_30806_, _30804_, _02083_);
  nor (_30807_, _30806_, _30801_);
  nor (_30808_, _30807_, _30505_);
  and (_30809_, _30505_, _01723_);
  or (_30810_, _02075_, _01975_);
  or (_30811_, _10321_, _02074_);
  or (_30812_, _30811_, _30810_);
  and (_30813_, _30812_, _01652_);
  or (_30814_, _30813_, _30809_);
  or (_30815_, _30814_, _30808_);
  and (_30816_, _30813_, _01614_);
  nor (_30817_, _30816_, _06455_);
  and (_30818_, _30817_, _30815_);
  nand (_30819_, _06455_, _01723_);
  and (_30820_, _02047_, _01652_);
  nor (_30821_, _30820_, _06450_);
  nand (_30822_, _30821_, _30819_);
  or (_30823_, _30822_, _30818_);
  nor (_30824_, _30821_, _01723_);
  and (_30825_, _07210_, _01434_);
  nor (_30827_, _30825_, _30824_);
  and (_30828_, _30827_, _30823_);
  and (_30829_, _30825_, _01723_);
  or (_30830_, _30829_, _07255_);
  or (_30831_, _30830_, _30828_);
  or (_30832_, _07254_, _01253_);
  and (_30833_, _30832_, _07305_);
  and (_30834_, _30833_, _30831_);
  and (_30835_, _07304_, _01723_);
  or (_30836_, _30835_, _01888_);
  or (_30838_, _30836_, _30834_);
  or (_30839_, _04907_, _01889_);
  and (_30840_, _30839_, _30838_);
  or (_30841_, _30840_, _01653_);
  nand (_30842_, _02687_, _01653_);
  and (_30843_, _30842_, _02202_);
  and (_30844_, _30843_, _30841_);
  nand (_30845_, _30497_, _02082_);
  nand (_30846_, _30845_, _30503_);
  or (_30847_, _30846_, _30844_);
  nand (_30849_, _30847_, _30504_);
  not (_30850_, _01542_);
  and (_30851_, _03521_, _30850_);
  nor (_30852_, _30851_, _02935_);
  nand (_30853_, _30852_, _30849_);
  or (_30854_, _30852_, _01723_);
  and (_30855_, _30854_, _02303_);
  and (_30856_, _30855_, _30853_);
  nand (_30857_, _02201_, _01253_);
  nand (_30858_, _30857_, _10442_);
  or (_30860_, _30858_, _30856_);
  and (_30861_, _30860_, _30500_);
  or (_30862_, _30861_, _03370_);
  nand (_30863_, _03370_, _02687_);
  and (_30864_, _30863_, _01887_);
  and (_30865_, _30864_, _30862_);
  or (_30866_, _30865_, _30499_);
  and (_30867_, _30866_, _05154_);
  or (_30868_, _05154_, _01614_);
  nor (_30869_, _02948_, _02952_);
  nand (_30871_, _30869_, _30868_);
  or (_30872_, _30871_, _30867_);
  or (_30873_, _30869_, _01723_);
  and (_30874_, _30873_, _01538_);
  and (_30875_, _30874_, _30872_);
  nand (_30876_, _01537_, _01253_);
  nand (_30877_, _30876_, _10465_);
  or (_30878_, _30877_, _30875_);
  and (_30879_, _30878_, _30492_);
  or (_30880_, _30879_, _30482_);
  nand (_30882_, _30482_, _02687_);
  and (_30883_, _30882_, _10481_);
  and (_30884_, _30883_, _30880_);
  and (_30885_, _09829_, _01723_);
  or (_30886_, _30885_, _38088_);
  or (_30887_, _30886_, _30884_);
  or (_30888_, _38087_, \oc8051_golden_model_1.PC [1]);
  and (_30889_, _30888_, _37580_);
  and (_40359_, _30889_, _30887_);
  and (_30890_, _01553_, _01537_);
  and (_30892_, _02201_, _01553_);
  or (_30893_, _09844_, _01582_);
  or (_30894_, _09846_, _01582_);
  or (_30895_, _09861_, _01582_);
  nand (_30896_, _09863_, _01583_);
  or (_30897_, _10327_, _01582_);
  nor (_30898_, _03140_, _02899_);
  and (_30899_, _30898_, _03138_);
  or (_30900_, _30899_, _01553_);
  and (_30901_, _02062_, _01637_);
  or (_30903_, _10245_, _01582_);
  and (_30904_, _02075_, _01601_);
  nand (_30905_, _10219_, _01583_);
  nand (_30906_, _08628_, _01583_);
  nor (_30907_, _09953_, _09951_);
  nor (_30908_, _30907_, _09954_);
  or (_30909_, _30908_, _08498_);
  nand (_30910_, _09943_, _08498_);
  and (_30911_, _30910_, _30909_);
  or (_30912_, _30911_, _08494_);
  or (_30914_, _30908_, _09996_);
  or (_30915_, _09876_, _09942_);
  and (_30916_, _30915_, _30914_);
  or (_30917_, _30916_, _02814_);
  and (_30918_, _10107_, _01553_);
  nor (_30919_, _10062_, _10060_);
  nor (_30920_, _30919_, _10063_);
  and (_30921_, _30920_, _10105_);
  or (_30922_, _30921_, _30918_);
  or (_30923_, _30922_, _04381_);
  nand (_30925_, _02338_, _02823_);
  and (_30926_, _21690_, _10129_);
  or (_30927_, _30926_, _01582_);
  nand (_30928_, _02817_, _01554_);
  or (_30929_, _02817_, \oc8051_golden_model_1.PC [2]);
  or (_30930_, _30929_, _10112_);
  and (_30931_, _30930_, _30928_);
  or (_30932_, _10125_, _06625_);
  or (_30933_, _30932_, _30931_);
  and (_30934_, _30933_, _06618_);
  and (_30936_, _30934_, _30927_);
  and (_30937_, _30936_, _30925_);
  and (_30938_, _02003_, _01553_);
  or (_30939_, _30938_, _06616_);
  or (_30940_, _30939_, _30937_);
  nand (_30941_, _06616_, _01583_);
  and (_30942_, _30941_, _01568_);
  and (_30943_, _30942_, _30940_);
  nor (_30944_, _02338_, _01568_);
  or (_30945_, _30944_, _04380_);
  or (_30947_, _30945_, _30943_);
  and (_30948_, _30947_, _04394_);
  and (_30949_, _30948_, _30923_);
  and (_30950_, _01883_, _01582_);
  or (_30951_, _30950_, _02001_);
  or (_30952_, _30951_, _30949_);
  and (_30953_, _30952_, _30917_);
  or (_30954_, _30953_, _30311_);
  or (_30955_, _09871_, _01582_);
  and (_30956_, _30955_, _02024_);
  and (_30958_, _30956_, _30954_);
  and (_30959_, _02007_, _01553_);
  or (_30960_, _30959_, _03279_);
  or (_30961_, _30960_, _30958_);
  nand (_30962_, _02338_, _03279_);
  and (_30963_, _30962_, _02840_);
  and (_30964_, _30963_, _30961_);
  nand (_30965_, _01999_, _01553_);
  nand (_30966_, _30965_, _10156_);
  or (_30967_, _30966_, _30964_);
  or (_30969_, _10156_, _01582_);
  and (_30970_, _30969_, _02021_);
  and (_30971_, _30970_, _30967_);
  nand (_30972_, _02006_, _01553_);
  nand (_30973_, _30972_, _10163_);
  or (_30974_, _30973_, _30971_);
  or (_30975_, _10163_, _01582_);
  and (_30976_, _30975_, _02025_);
  and (_30977_, _30976_, _30974_);
  and (_30978_, _01997_, _01553_);
  or (_30979_, _30978_, _10167_);
  or (_30980_, _30979_, _30977_);
  nand (_30981_, _02338_, _10167_);
  and (_30982_, _30981_, _01880_);
  and (_30983_, _30982_, _30980_);
  nand (_30984_, _01878_, _01553_);
  nand (_30985_, _30984_, _08538_);
  or (_30986_, _30985_, _30983_);
  or (_30987_, _30908_, _08572_);
  nand (_30988_, _09943_, _08572_);
  and (_30990_, _30988_, _30987_);
  or (_30991_, _30990_, _08538_);
  and (_30992_, _30991_, _30986_);
  or (_30993_, _30992_, _08493_);
  and (_30994_, _30993_, _30912_);
  or (_30995_, _30994_, _01995_);
  and (_30996_, _09942_, _08625_);
  and (_30997_, _30908_, _30342_);
  or (_30998_, _30997_, _02444_);
  or (_30999_, _30998_, _30996_);
  and (_31001_, _30999_, _02046_);
  and (_31002_, _31001_, _30995_);
  or (_31003_, _30908_, _08664_);
  nand (_31004_, _09943_, _08664_);
  and (_31005_, _31004_, _02045_);
  and (_31006_, _31005_, _31003_);
  or (_31007_, _31006_, _08628_);
  or (_31008_, _31007_, _31002_);
  and (_31009_, _31008_, _30906_);
  or (_31010_, _31009_, _01991_);
  nand (_31012_, _01991_, _01554_);
  and (_31013_, _31012_, _01565_);
  and (_31014_, _31013_, _31010_);
  nor (_31015_, _02338_, _01565_);
  nand (_31016_, _02047_, _01965_);
  nand (_31017_, _30631_, _31016_);
  or (_31018_, _31017_, _31015_);
  or (_31019_, _31018_, _31014_);
  nor (_31020_, _02508_, _01554_);
  or (_31021_, _31020_, _30632_);
  and (_31023_, _31021_, _31019_);
  nand (_31024_, _02508_, _01553_);
  nand (_31025_, _31024_, _10207_);
  or (_31026_, _31025_, _31023_);
  or (_31027_, _10207_, _01582_);
  and (_31028_, _31027_, _08249_);
  and (_31029_, _31028_, _31026_);
  and (_31030_, _01967_, _01553_);
  or (_31031_, _31030_, _10213_);
  or (_31032_, _31031_, _31029_);
  nand (_31034_, _02338_, _10213_);
  and (_31035_, _31034_, _08248_);
  and (_31036_, _31035_, _31032_);
  and (_31037_, _01966_, _01553_);
  or (_31038_, _31037_, _10219_);
  or (_31039_, _31038_, _31036_);
  and (_31040_, _31039_, _30905_);
  or (_31041_, _31040_, _06776_);
  or (_31042_, _06775_, _01553_);
  and (_31043_, _31042_, _01550_);
  and (_31045_, _31043_, _31041_);
  and (_31046_, _01582_, _01549_);
  or (_31047_, _31046_, _01875_);
  or (_31048_, _31047_, _31045_);
  nand (_31049_, _01875_, _01554_);
  and (_31050_, _31049_, _04310_);
  and (_31051_, _31050_, _31048_);
  nor (_31052_, _02338_, _04310_);
  or (_31053_, _31052_, _02080_);
  or (_31054_, _31053_, _31051_);
  and (_31056_, _02062_, _01601_);
  and (_31057_, _09943_, _02080_);
  nor (_31058_, _31057_, _31056_);
  and (_31059_, _31058_, _31054_);
  and (_31060_, _31056_, _01553_);
  nor (_31061_, _31060_, _31059_);
  nor (_31062_, _31061_, _30904_);
  nand (_31063_, _30904_, _01553_);
  nor (_31064_, _02049_, _02047_);
  nor (_31065_, _31064_, _02531_);
  not (_31067_, _31065_);
  not (_31068_, _05247_);
  nor (_31069_, _31068_, _02530_);
  and (_31070_, _31069_, _31067_);
  nand (_31071_, _31070_, _31063_);
  or (_31072_, _31071_, _31062_);
  or (_31073_, _31070_, _01553_);
  and (_31074_, _31073_, _02043_);
  and (_31075_, _31074_, _31072_);
  nand (_31076_, _09942_, _01602_);
  nand (_31078_, _31076_, _10245_);
  or (_31079_, _31078_, _31075_);
  and (_31080_, _31079_, _30903_);
  or (_31081_, _31080_, _01959_);
  nand (_31082_, _01959_, _01554_);
  and (_31083_, _31082_, _30378_);
  and (_31084_, _31083_, _31081_);
  nor (_31085_, _02338_, _30378_);
  or (_31086_, _31085_, _10253_);
  or (_31087_, _31086_, _31084_);
  or (_31089_, _30920_, _10254_);
  and (_31090_, _31089_, _31087_);
  or (_31091_, _31090_, _30901_);
  and (_31092_, _02075_, _01637_);
  and (_31093_, _30901_, _01554_);
  nor (_31094_, _31093_, _31092_);
  and (_31095_, _31094_, _31091_);
  nand (_31096_, _31092_, _01553_);
  nand (_31097_, _31096_, _30899_);
  or (_31098_, _31097_, _31095_);
  and (_31100_, _31098_, _30900_);
  or (_31101_, _31100_, _01869_);
  nand (_31102_, _09943_, _01869_);
  and (_31103_, _31102_, _06985_);
  and (_31104_, _31103_, _31101_);
  and (_31105_, _06984_, _01553_);
  or (_31106_, _31105_, _10267_);
  or (_31107_, _31106_, _31104_);
  or (_31108_, _10268_, _01599_);
  and (_31109_, _31108_, _02576_);
  and (_31111_, _31109_, _31107_);
  and (_31112_, _01958_, _01553_);
  or (_31113_, _31112_, _01638_);
  or (_31114_, _31113_, _31111_);
  nand (_31115_, _02338_, _01638_);
  and (_31116_, _31115_, _10311_);
  and (_31117_, _31116_, _31114_);
  or (_31118_, _30920_, _07356_);
  nand (_31119_, _07356_, _01554_);
  and (_31120_, _31119_, _10310_);
  and (_31122_, _31120_, _31118_);
  or (_31123_, _31122_, _10331_);
  or (_31124_, _31123_, _31117_);
  and (_31125_, _31124_, _30897_);
  or (_31126_, _31125_, _10330_);
  or (_31127_, _10329_, _01553_);
  and (_31128_, _31127_, _02166_);
  and (_31129_, _31128_, _31126_);
  and (_31130_, _09942_, _02079_);
  or (_31131_, _31130_, _02167_);
  or (_31133_, _31131_, _31129_);
  nand (_31134_, _02167_, _01554_);
  and (_31135_, _31134_, _31133_);
  or (_31136_, _31135_, _01645_);
  nand (_31137_, _02338_, _01645_);
  and (_31138_, _31137_, _10344_);
  and (_31139_, _31138_, _31136_);
  or (_31140_, _30920_, _10316_);
  or (_31141_, _07356_, _01553_);
  and (_31142_, _31141_, _10343_);
  and (_31143_, _31142_, _31140_);
  or (_31144_, _31143_, _09863_);
  or (_31145_, _31144_, _31139_);
  and (_31146_, _31145_, _30896_);
  or (_31147_, _31146_, _07042_);
  or (_31148_, _07041_, _01553_);
  and (_31149_, _31148_, _02176_);
  and (_31150_, _31149_, _31147_);
  and (_31151_, _09942_, _02072_);
  or (_31152_, _31151_, _02177_);
  or (_31154_, _31152_, _31150_);
  nand (_31155_, _02177_, _01554_);
  and (_31156_, _31155_, _31154_);
  or (_31157_, _31156_, _01632_);
  nand (_31158_, _02338_, _01632_);
  and (_31159_, _31158_, _10364_);
  and (_31160_, _31159_, _31157_);
  or (_31161_, _30920_, \oc8051_golden_model_1.PSW [7]);
  or (_31162_, _01553_, _06518_);
  and (_31163_, _31162_, _10363_);
  and (_31165_, _31163_, _31161_);
  or (_31166_, _31165_, _10368_);
  or (_31167_, _31166_, _31160_);
  and (_31168_, _31167_, _30895_);
  or (_31169_, _31168_, _09854_);
  or (_31170_, _09853_, _01553_);
  and (_31171_, _31170_, _04788_);
  and (_31172_, _31171_, _31169_);
  and (_31173_, _09942_, _02071_);
  or (_31174_, _31173_, _02173_);
  or (_31176_, _31174_, _31172_);
  nand (_31177_, _02173_, _01554_);
  and (_31178_, _31177_, _31176_);
  or (_31179_, _31178_, _01648_);
  nand (_31180_, _02338_, _01648_);
  and (_31181_, _31180_, _09849_);
  and (_31182_, _31181_, _31179_);
  or (_31183_, _30920_, _06518_);
  or (_31184_, _01553_, \oc8051_golden_model_1.PSW [7]);
  and (_31185_, _31184_, _09848_);
  and (_31187_, _31185_, _31183_);
  or (_31188_, _31187_, _10385_);
  or (_31189_, _31188_, _31182_);
  and (_31190_, _31189_, _30894_);
  or (_31191_, _31190_, _07146_);
  or (_31192_, _07145_, _01553_);
  and (_31193_, _31192_, _07176_);
  and (_31194_, _31193_, _31191_);
  and (_31195_, _07175_, _01582_);
  or (_31196_, _31195_, _02185_);
  or (_31198_, _31196_, _31194_);
  or (_31199_, _05043_, _09305_);
  and (_31200_, _31199_, _31198_);
  or (_31201_, _31200_, _01636_);
  nand (_31202_, _02338_, _01636_);
  and (_31203_, _31202_, _10403_);
  and (_31204_, _31203_, _31201_);
  or (_31205_, _30908_, _10408_);
  or (_31206_, _09942_, _08439_);
  and (_31207_, _31206_, _02083_);
  and (_31209_, _31207_, _31205_);
  or (_31210_, _31209_, _10407_);
  or (_31211_, _31210_, _31204_);
  and (_31212_, _31211_, _30893_);
  or (_31213_, _31212_, _07255_);
  or (_31214_, _07254_, _01553_);
  and (_31215_, _31214_, _07305_);
  and (_31216_, _31215_, _31213_);
  and (_31217_, _07304_, _01582_);
  or (_31218_, _31217_, _01888_);
  or (_31220_, _31218_, _31216_);
  or (_31221_, _05043_, _01889_);
  and (_31222_, _31221_, _31220_);
  or (_31223_, _31222_, _01653_);
  nand (_31224_, _02338_, _01653_);
  and (_31225_, _31224_, _02202_);
  and (_31226_, _31225_, _31223_);
  or (_31227_, _30908_, _08439_);
  nand (_31228_, _09943_, _08439_);
  and (_31229_, _31228_, _31227_);
  and (_31231_, _31229_, _02082_);
  or (_31232_, _31231_, _10435_);
  or (_31233_, _31232_, _31226_);
  nand (_31234_, _10435_, _01583_);
  and (_31235_, _31234_, _02303_);
  and (_31236_, _31235_, _31233_);
  or (_31237_, _31236_, _30892_);
  and (_31238_, _31237_, _10442_);
  nor (_31239_, _10442_, _01583_);
  or (_31240_, _31239_, _03370_);
  or (_31242_, _31240_, _31238_);
  nand (_31243_, _03370_, _02338_);
  and (_31244_, _31243_, _01887_);
  and (_31245_, _31244_, _31242_);
  and (_31246_, _31229_, _01860_);
  or (_31247_, _31246_, _10458_);
  or (_31248_, _31247_, _31245_);
  nand (_31249_, _10458_, _01583_);
  and (_31250_, _31249_, _01538_);
  and (_31251_, _31250_, _31248_);
  or (_31253_, _31251_, _30890_);
  and (_31254_, _31253_, _10465_);
  nor (_31255_, _10465_, _01583_);
  or (_31256_, _31255_, _30482_);
  or (_31257_, _31256_, _31254_);
  nand (_31258_, _30482_, _02338_);
  and (_31259_, _31258_, _10481_);
  and (_31260_, _31259_, _31257_);
  and (_31261_, _09829_, _01582_);
  or (_31262_, _31261_, _38088_);
  or (_31264_, _31262_, _31260_);
  or (_31265_, _38087_, \oc8051_golden_model_1.PC [2]);
  and (_31266_, _31265_, _37580_);
  and (_40360_, _31266_, _31264_);
  and (_31267_, _01682_, _01537_);
  or (_31268_, _09844_, _02103_);
  or (_31269_, _09846_, _02103_);
  or (_31270_, _09861_, _02103_);
  nand (_31271_, _09863_, _01675_);
  or (_31272_, _10327_, _02103_);
  or (_31274_, _04757_, _01682_);
  nand (_31275_, _01875_, _01683_);
  nand (_31276_, _10219_, _01675_);
  nand (_31277_, _08628_, _01675_);
  or (_31278_, _09940_, _09939_);
  nand (_31279_, _31278_, _09955_);
  or (_31280_, _31278_, _09955_);
  and (_31281_, _31280_, _31279_);
  or (_31282_, _31281_, _08498_);
  nand (_31283_, _09938_, _08498_);
  and (_31285_, _31283_, _31282_);
  or (_31286_, _31285_, _08494_);
  or (_31287_, _09876_, _09937_);
  or (_31288_, _31281_, _09996_);
  and (_31289_, _31288_, _31287_);
  or (_31290_, _31289_, _02814_);
  and (_31291_, _10107_, _01682_);
  or (_31292_, _10052_, _10051_);
  nand (_31293_, _31292_, _10064_);
  or (_31294_, _31292_, _10064_);
  and (_31295_, _31294_, _31293_);
  and (_31296_, _31295_, _10105_);
  or (_31297_, _31296_, _31291_);
  or (_31298_, _31297_, _04381_);
  nor (_31299_, _02159_, _01562_);
  nand (_31300_, _02817_, _01683_);
  and (_31301_, _31300_, _10121_);
  nor (_31302_, _10112_, _01249_);
  or (_31303_, _31302_, _02817_);
  and (_31304_, _31303_, _31301_);
  nor (_31306_, _21690_, _01675_);
  or (_31307_, _31306_, _06629_);
  or (_31308_, _31307_, _31304_);
  and (_31309_, _31308_, _01562_);
  or (_31310_, _31309_, _31299_);
  nand (_31311_, _06629_, _01675_);
  and (_31312_, _31311_, _06618_);
  and (_31313_, _31312_, _31310_);
  and (_31314_, _02003_, _01682_);
  or (_31315_, _31314_, _06616_);
  or (_31317_, _31315_, _31313_);
  nand (_31318_, _06616_, _01675_);
  and (_31319_, _31318_, _01568_);
  and (_31320_, _31319_, _31317_);
  nor (_31321_, _02159_, _01568_);
  or (_31322_, _31321_, _04380_);
  or (_31323_, _31322_, _31320_);
  and (_31324_, _31323_, _04394_);
  and (_31325_, _31324_, _31298_);
  and (_31326_, _01883_, _02103_);
  or (_31328_, _31326_, _02001_);
  or (_31329_, _31328_, _31325_);
  and (_31330_, _31329_, _31290_);
  or (_31331_, _31330_, _30311_);
  or (_31332_, _09871_, _02103_);
  and (_31333_, _31332_, _02024_);
  and (_31334_, _31333_, _31331_);
  and (_31335_, _02007_, _01682_);
  or (_31336_, _31335_, _03279_);
  or (_31337_, _31336_, _31334_);
  nand (_31339_, _02159_, _03279_);
  and (_31340_, _31339_, _02840_);
  and (_31341_, _31340_, _31337_);
  nand (_31342_, _01999_, _01682_);
  nand (_31343_, _31342_, _10156_);
  or (_31344_, _31343_, _31341_);
  or (_31345_, _10156_, _02103_);
  and (_31346_, _31345_, _02021_);
  and (_31347_, _31346_, _31344_);
  nand (_31348_, _02006_, _01682_);
  nand (_31350_, _31348_, _10163_);
  or (_31351_, _31350_, _31347_);
  or (_31352_, _10163_, _02103_);
  and (_31353_, _31352_, _02025_);
  and (_31354_, _31353_, _31351_);
  and (_31355_, _01997_, _01682_);
  or (_31356_, _31355_, _10167_);
  or (_31357_, _31356_, _31354_);
  nand (_31358_, _02159_, _10167_);
  and (_31359_, _31358_, _01880_);
  and (_31361_, _31359_, _31357_);
  nand (_31362_, _01878_, _01682_);
  nand (_31363_, _31362_, _08538_);
  or (_31364_, _31363_, _31361_);
  or (_31365_, _31281_, _08572_);
  nand (_31366_, _09938_, _08572_);
  and (_31367_, _31366_, _31365_);
  or (_31368_, _31367_, _08538_);
  and (_31369_, _31368_, _31364_);
  or (_31370_, _31369_, _08493_);
  and (_31372_, _31370_, _31286_);
  or (_31373_, _31372_, _01995_);
  and (_31374_, _31281_, _30342_);
  and (_31375_, _09937_, _08625_);
  or (_31376_, _31375_, _02444_);
  or (_31377_, _31376_, _31374_);
  and (_31378_, _31377_, _02046_);
  and (_31379_, _31378_, _31373_);
  nand (_31380_, _09938_, _08664_);
  or (_31381_, _31281_, _08664_);
  and (_31383_, _31381_, _02045_);
  and (_31384_, _31383_, _31380_);
  or (_31385_, _31384_, _08628_);
  or (_31386_, _31385_, _31379_);
  and (_31387_, _31386_, _31277_);
  or (_31388_, _31387_, _01991_);
  nand (_31389_, _01991_, _01683_);
  and (_31390_, _31389_, _01565_);
  and (_31391_, _31390_, _31388_);
  nor (_31392_, _02159_, _01565_);
  or (_31394_, _31392_, _30633_);
  or (_31395_, _31394_, _31391_);
  or (_31396_, _30632_, _01682_);
  and (_31397_, _31396_, _31395_);
  or (_31398_, _31397_, _10211_);
  or (_31399_, _10207_, _02103_);
  and (_31400_, _31399_, _08249_);
  and (_31401_, _31400_, _31398_);
  and (_31402_, _01967_, _01682_);
  or (_31403_, _31402_, _10213_);
  or (_31405_, _31403_, _31401_);
  nand (_31406_, _02159_, _10213_);
  and (_31407_, _31406_, _08248_);
  and (_31408_, _31407_, _31405_);
  and (_31409_, _01966_, _01682_);
  or (_31410_, _31409_, _10219_);
  or (_31411_, _31410_, _31408_);
  and (_31412_, _31411_, _31276_);
  or (_31413_, _31412_, _06776_);
  or (_31414_, _06775_, _01682_);
  and (_31416_, _31414_, _01550_);
  and (_31417_, _31416_, _31413_);
  and (_31418_, _01549_, _02103_);
  or (_31419_, _31418_, _01875_);
  or (_31420_, _31419_, _31417_);
  and (_31421_, _31420_, _31275_);
  or (_31422_, _31421_, _01604_);
  nand (_31423_, _02159_, _01604_);
  and (_31424_, _31423_, _07401_);
  and (_31425_, _31424_, _31422_);
  nand (_31427_, _09937_, _02080_);
  nand (_31428_, _31427_, _09211_);
  or (_31429_, _31428_, _31425_);
  or (_31430_, _09211_, _01682_);
  and (_31431_, _31430_, _02043_);
  and (_31432_, _31431_, _31429_);
  nand (_31433_, _09937_, _01602_);
  nand (_31434_, _31433_, _10245_);
  or (_31435_, _31434_, _31432_);
  or (_31436_, _10245_, _02103_);
  and (_31438_, _31436_, _30680_);
  and (_31439_, _31438_, _31435_);
  and (_31440_, _01959_, _01682_);
  or (_31441_, _31440_, _01649_);
  or (_31442_, _31441_, _31439_);
  nand (_31443_, _02159_, _01649_);
  and (_31444_, _31443_, _10254_);
  and (_31445_, _31444_, _31442_);
  and (_31446_, _31295_, _10253_);
  or (_31447_, _31446_, _04758_);
  or (_31448_, _31447_, _31445_);
  and (_31449_, _31448_, _31274_);
  or (_31450_, _31449_, _01869_);
  nand (_31451_, _09938_, _01869_);
  and (_31452_, _31451_, _06985_);
  and (_31453_, _31452_, _31450_);
  and (_31454_, _06984_, _01682_);
  or (_31455_, _31454_, _10267_);
  or (_31456_, _31455_, _31453_);
  or (_31457_, _10268_, _01671_);
  and (_31459_, _31457_, _02576_);
  and (_31460_, _31459_, _31456_);
  and (_31461_, _01958_, _01682_);
  or (_31462_, _31461_, _01638_);
  or (_31463_, _31462_, _31460_);
  nand (_31464_, _02159_, _01638_);
  and (_31465_, _31464_, _10311_);
  and (_31466_, _31465_, _31463_);
  or (_31467_, _31295_, _07356_);
  nand (_31468_, _07356_, _01683_);
  and (_31470_, _31468_, _10310_);
  and (_31471_, _31470_, _31467_);
  or (_31472_, _31471_, _10331_);
  or (_31473_, _31472_, _31466_);
  and (_31474_, _31473_, _31272_);
  or (_31475_, _31474_, _10330_);
  or (_31476_, _10329_, _01682_);
  and (_31477_, _31476_, _02166_);
  and (_31478_, _31477_, _31475_);
  and (_31479_, _09937_, _02079_);
  or (_31481_, _31479_, _02167_);
  or (_31482_, _31481_, _31478_);
  nand (_31483_, _02167_, _01683_);
  and (_31484_, _31483_, _31482_);
  or (_31485_, _31484_, _01645_);
  nand (_31486_, _02159_, _01645_);
  and (_31487_, _31486_, _10344_);
  and (_31488_, _31487_, _31485_);
  or (_31489_, _31295_, _10316_);
  or (_31490_, _07356_, _01682_);
  and (_31492_, _31490_, _10343_);
  and (_31493_, _31492_, _31489_);
  or (_31494_, _31493_, _09863_);
  or (_31495_, _31494_, _31488_);
  and (_31496_, _31495_, _31271_);
  or (_31497_, _31496_, _07042_);
  or (_31498_, _07041_, _01682_);
  and (_31499_, _31498_, _02176_);
  and (_31500_, _31499_, _31497_);
  and (_31501_, _09937_, _02072_);
  or (_31503_, _31501_, _02177_);
  or (_31504_, _31503_, _31500_);
  nand (_31505_, _02177_, _01683_);
  and (_31506_, _31505_, _31504_);
  or (_31507_, _31506_, _01632_);
  nand (_31508_, _02159_, _01632_);
  and (_31509_, _31508_, _10364_);
  and (_31510_, _31509_, _31507_);
  or (_31511_, _31295_, \oc8051_golden_model_1.PSW [7]);
  or (_31512_, _01682_, _06518_);
  and (_31514_, _31512_, _10363_);
  and (_31515_, _31514_, _31511_);
  or (_31516_, _31515_, _10368_);
  or (_31517_, _31516_, _31510_);
  and (_31518_, _31517_, _31270_);
  or (_31519_, _31518_, _09854_);
  or (_31520_, _09853_, _01682_);
  and (_31521_, _31520_, _04788_);
  and (_31522_, _31521_, _31519_);
  and (_31523_, _09937_, _02071_);
  or (_31525_, _31523_, _02173_);
  or (_31526_, _31525_, _31522_);
  nand (_31527_, _02173_, _01683_);
  and (_31528_, _31527_, _31526_);
  or (_31529_, _31528_, _01648_);
  nand (_31530_, _02159_, _01648_);
  and (_31531_, _31530_, _09849_);
  and (_31532_, _31531_, _31529_);
  or (_31533_, _31295_, _06518_);
  or (_31534_, _01682_, \oc8051_golden_model_1.PSW [7]);
  and (_31536_, _31534_, _09848_);
  and (_31537_, _31536_, _31533_);
  or (_31538_, _31537_, _10385_);
  or (_31539_, _31538_, _31532_);
  and (_31540_, _31539_, _31269_);
  or (_31541_, _31540_, _07146_);
  or (_31542_, _07145_, _01682_);
  and (_31543_, _31542_, _07176_);
  and (_31544_, _31543_, _31541_);
  and (_31545_, _07175_, _02103_);
  or (_31547_, _31545_, _02185_);
  or (_31548_, _31547_, _31544_);
  or (_31549_, _04998_, _09305_);
  and (_31550_, _31549_, _31548_);
  or (_31551_, _31550_, _01636_);
  nand (_31552_, _02159_, _01636_);
  and (_31553_, _31552_, _10403_);
  and (_31554_, _31553_, _31551_);
  or (_31555_, _31281_, _10408_);
  or (_31556_, _09937_, _08439_);
  and (_31558_, _31556_, _02083_);
  and (_31559_, _31558_, _31555_);
  or (_31560_, _31559_, _10407_);
  or (_31561_, _31560_, _31554_);
  and (_31562_, _31561_, _31268_);
  or (_31563_, _31562_, _07255_);
  or (_31564_, _07254_, _01682_);
  and (_31565_, _31564_, _07305_);
  and (_31566_, _31565_, _31563_);
  and (_31567_, _07304_, _02103_);
  or (_31569_, _31567_, _01888_);
  or (_31570_, _31569_, _31566_);
  or (_31571_, _04998_, _01889_);
  and (_31572_, _31571_, _31570_);
  or (_31573_, _31572_, _01653_);
  nand (_31574_, _02159_, _01653_);
  and (_31575_, _31574_, _02202_);
  and (_31576_, _31575_, _31573_);
  or (_31577_, _31281_, _08439_);
  nand (_31578_, _09938_, _08439_);
  and (_31580_, _31578_, _31577_);
  and (_31581_, _31580_, _02082_);
  or (_31582_, _31581_, _10435_);
  or (_31583_, _31582_, _31576_);
  nand (_31584_, _10435_, _01675_);
  and (_31585_, _31584_, _02303_);
  and (_31586_, _31585_, _31583_);
  nand (_31587_, _02201_, _01682_);
  nand (_31588_, _31587_, _10442_);
  or (_31589_, _31588_, _31586_);
  or (_31591_, _10442_, _02103_);
  and (_31592_, _31591_, _31589_);
  or (_31593_, _31592_, _03370_);
  nand (_31594_, _03370_, _02159_);
  and (_31595_, _31594_, _01887_);
  and (_31596_, _31595_, _31593_);
  and (_31597_, _31580_, _01860_);
  or (_31598_, _31597_, _10458_);
  or (_31599_, _31598_, _31596_);
  nand (_31600_, _10458_, _01675_);
  and (_31601_, _31600_, _01538_);
  and (_31602_, _31601_, _31599_);
  or (_31603_, _31602_, _31267_);
  and (_31604_, _31603_, _10465_);
  nor (_31605_, _10465_, _01675_);
  or (_31606_, _31605_, _30482_);
  or (_31607_, _31606_, _31604_);
  nand (_31608_, _30482_, _02159_);
  and (_31609_, _31608_, _10481_);
  and (_31610_, _31609_, _31607_);
  and (_31612_, _09829_, _02103_);
  or (_31613_, _31612_, _38088_);
  or (_31614_, _31613_, _31610_);
  or (_31615_, _38087_, \oc8051_golden_model_1.PC [3]);
  and (_31616_, _31615_, _37580_);
  and (_40361_, _31616_, _31614_);
  nand (_31617_, _04657_, _03370_);
  or (_31618_, _10068_, _10066_);
  and (_31619_, _31618_, _10069_);
  or (_31620_, _31619_, _06518_);
  or (_31622_, _10048_, \oc8051_golden_model_1.PSW [7]);
  and (_31623_, _31622_, _09848_);
  and (_31624_, _31623_, _31620_);
  or (_31625_, _31619_, _07356_);
  nand (_31626_, _10049_, _07356_);
  and (_31627_, _31626_, _10310_);
  and (_31628_, _31627_, _31625_);
  or (_31629_, _10048_, _04757_);
  nand (_31630_, _04657_, _10213_);
  and (_31631_, _09830_, \oc8051_golden_model_1.PC [4]);
  nor (_31633_, _09830_, \oc8051_golden_model_1.PC [4]);
  nor (_31634_, _31633_, _31631_);
  not (_31635_, _31634_);
  nand (_31636_, _31635_, _08628_);
  nand (_31637_, _10049_, _01997_);
  or (_31638_, _31634_, _10156_);
  and (_31639_, _31619_, _10105_);
  and (_31640_, _10107_, _10048_);
  or (_31641_, _31640_, _31639_);
  or (_31642_, _31641_, _04381_);
  nand (_31644_, _04657_, _02823_);
  nand (_31645_, _10049_, _02817_);
  and (_31646_, _31645_, _10121_);
  and (_31647_, _10113_, \oc8051_golden_model_1.PC [4]);
  or (_31648_, _31647_, _02817_);
  and (_31649_, _31648_, _31646_);
  nor (_31650_, _31635_, _21690_);
  or (_31651_, _31650_, _02823_);
  or (_31652_, _31651_, _31649_);
  and (_31653_, _31652_, _10129_);
  and (_31655_, _31653_, _31644_);
  and (_31656_, _31634_, _06629_);
  or (_31657_, _31656_, _02003_);
  or (_31658_, _31657_, _31655_);
  nand (_31659_, _10049_, _02003_);
  and (_31660_, _31659_, _31658_);
  or (_31661_, _31660_, _06616_);
  nand (_31662_, _31635_, _06616_);
  and (_31663_, _31662_, _01568_);
  and (_31664_, _31663_, _31661_);
  nor (_31666_, _04657_, _01568_);
  or (_31667_, _31666_, _04380_);
  or (_31668_, _31667_, _31664_);
  and (_31669_, _31668_, _31642_);
  or (_31670_, _31669_, _01883_);
  nand (_31671_, _31635_, _01883_);
  and (_31672_, _31671_, _02814_);
  and (_31673_, _31672_, _31670_);
  or (_31674_, _09876_, _09934_);
  or (_31675_, _09959_, _09957_);
  and (_31677_, _31675_, _09960_);
  or (_31678_, _31677_, _09996_);
  and (_31679_, _31678_, _02001_);
  and (_31680_, _31679_, _31674_);
  or (_31681_, _31680_, _30311_);
  or (_31682_, _31681_, _31673_);
  or (_31683_, _31634_, _09871_);
  and (_31684_, _31683_, _31682_);
  or (_31685_, _31684_, _02007_);
  nand (_31686_, _10049_, _02007_);
  and (_31688_, _31686_, _01558_);
  and (_31689_, _31688_, _31685_);
  nor (_31690_, _04657_, _01558_);
  or (_31691_, _31690_, _01999_);
  or (_31692_, _31691_, _31689_);
  nand (_31693_, _10049_, _01999_);
  and (_31694_, _31693_, _31692_);
  or (_31695_, _31694_, _10157_);
  and (_31696_, _31695_, _31638_);
  or (_31697_, _31696_, _02006_);
  nand (_31699_, _10049_, _02006_);
  and (_31700_, _31699_, _10163_);
  and (_31701_, _31700_, _31697_);
  nor (_31702_, _31635_, _10163_);
  or (_31703_, _31702_, _01997_);
  or (_31704_, _31703_, _31701_);
  and (_31705_, _31704_, _31637_);
  or (_31706_, _31705_, _10167_);
  nand (_31707_, _04657_, _10167_);
  and (_31708_, _31707_, _01880_);
  and (_31710_, _31708_, _31706_);
  nand (_31711_, _10048_, _01878_);
  nand (_31712_, _31711_, _08538_);
  or (_31713_, _31712_, _31710_);
  and (_31714_, _09934_, _08572_);
  and (_31715_, _31677_, _08573_);
  or (_31716_, _31715_, _31714_);
  or (_31717_, _31716_, _08538_);
  and (_31718_, _31717_, _31713_);
  or (_31719_, _31718_, _08493_);
  and (_31721_, _09934_, _08498_);
  and (_31722_, _31677_, _30279_);
  or (_31723_, _31722_, _31721_);
  or (_31724_, _31723_, _08494_);
  and (_31725_, _31724_, _31719_);
  or (_31726_, _31725_, _01995_);
  and (_31727_, _31677_, _30342_);
  and (_31728_, _09934_, _08625_);
  or (_31729_, _31728_, _02444_);
  or (_31730_, _31729_, _31727_);
  and (_31732_, _31730_, _02046_);
  and (_31733_, _31732_, _31726_);
  or (_31734_, _31677_, _08664_);
  not (_31735_, _08664_);
  or (_31736_, _09934_, _31735_);
  and (_31737_, _31736_, _02045_);
  and (_31738_, _31737_, _31734_);
  or (_31739_, _31738_, _08628_);
  or (_31740_, _31739_, _31733_);
  and (_31741_, _31740_, _31636_);
  or (_31743_, _31741_, _01991_);
  nand (_31744_, _10049_, _01991_);
  and (_31745_, _31744_, _01565_);
  and (_31746_, _31745_, _31743_);
  nor (_31747_, _04657_, _01565_);
  or (_31748_, _31747_, _30633_);
  or (_31749_, _31748_, _31746_);
  or (_31750_, _30632_, _10048_);
  and (_31751_, _31750_, _10207_);
  and (_31752_, _31751_, _31749_);
  nor (_31753_, _31635_, _10207_);
  or (_31754_, _31753_, _01967_);
  or (_31755_, _31754_, _31752_);
  nand (_31756_, _10049_, _01967_);
  and (_31757_, _31756_, _31755_);
  or (_31758_, _31757_, _10213_);
  and (_31759_, _31758_, _31630_);
  or (_31760_, _31759_, _01966_);
  and (_31761_, _10049_, _01966_);
  nor (_31762_, _31761_, _10219_);
  and (_31764_, _31762_, _31760_);
  and (_31765_, _31634_, _10219_);
  or (_31766_, _31765_, _06776_);
  or (_31767_, _31766_, _31764_);
  or (_31768_, _10048_, _06775_);
  and (_31769_, _31768_, _01550_);
  and (_31770_, _31769_, _31767_);
  and (_31771_, _31634_, _01549_);
  or (_31772_, _31771_, _01875_);
  or (_31773_, _31772_, _31770_);
  nand (_31775_, _10049_, _01875_);
  and (_31776_, _31775_, _31773_);
  or (_31777_, _31776_, _01604_);
  nand (_31778_, _04657_, _01604_);
  and (_31779_, _31778_, _07401_);
  and (_31780_, _31779_, _31777_);
  nand (_31781_, _09934_, _02080_);
  nand (_31782_, _31781_, _09211_);
  or (_31783_, _31782_, _31780_);
  or (_31784_, _10048_, _09211_);
  and (_31786_, _31784_, _02043_);
  and (_31787_, _31786_, _31783_);
  nand (_31788_, _09934_, _01602_);
  nand (_31789_, _31788_, _10245_);
  or (_31790_, _31789_, _31787_);
  or (_31791_, _31634_, _10245_);
  and (_31792_, _31791_, _30680_);
  and (_31793_, _31792_, _31790_);
  and (_31794_, _10048_, _01959_);
  or (_31795_, _31794_, _01649_);
  or (_31797_, _31795_, _31793_);
  nand (_31798_, _04657_, _01649_);
  and (_31799_, _31798_, _10254_);
  and (_31800_, _31799_, _31797_);
  and (_31801_, _31619_, _10253_);
  or (_31802_, _31801_, _04758_);
  or (_31803_, _31802_, _31800_);
  and (_31804_, _31803_, _31629_);
  or (_31805_, _31804_, _01869_);
  or (_31806_, _09934_, _01870_);
  and (_31808_, _31806_, _06985_);
  and (_31809_, _31808_, _31805_);
  and (_31810_, _10048_, _06984_);
  or (_31811_, _31810_, _10267_);
  or (_31812_, _31811_, _31809_);
  nor (_31813_, _10285_, _10283_);
  nor (_31814_, _31813_, _10286_);
  or (_31815_, _31814_, _10268_);
  and (_31816_, _31815_, _02576_);
  and (_31817_, _31816_, _31812_);
  and (_31819_, _10048_, _01958_);
  or (_31820_, _31819_, _01638_);
  or (_31821_, _31820_, _31817_);
  nand (_31822_, _04657_, _01638_);
  and (_31823_, _31822_, _10311_);
  and (_31824_, _31823_, _31821_);
  or (_31825_, _31824_, _31628_);
  and (_31826_, _31825_, _10327_);
  nor (_31827_, _31635_, _10327_);
  or (_31828_, _31827_, _10330_);
  or (_31830_, _31828_, _31826_);
  or (_31831_, _10048_, _10329_);
  and (_31832_, _31831_, _02166_);
  and (_31833_, _31832_, _31830_);
  and (_31834_, _09934_, _02079_);
  or (_31835_, _31834_, _02167_);
  or (_31836_, _31835_, _31833_);
  nand (_31837_, _10049_, _02167_);
  and (_31838_, _31837_, _31836_);
  or (_31839_, _31838_, _01645_);
  nand (_31841_, _04657_, _01645_);
  and (_31842_, _31841_, _10344_);
  and (_31843_, _31842_, _31839_);
  or (_31844_, _31619_, _10316_);
  or (_31845_, _10048_, _07356_);
  and (_31846_, _31845_, _10343_);
  and (_31847_, _31846_, _31844_);
  or (_31848_, _31847_, _31843_);
  and (_31849_, _31848_, _09864_);
  and (_31850_, _31634_, _09863_);
  or (_31852_, _31850_, _07042_);
  or (_31853_, _31852_, _31849_);
  or (_31854_, _10048_, _07041_);
  and (_31855_, _31854_, _02176_);
  and (_31856_, _31855_, _31853_);
  and (_31857_, _09934_, _02072_);
  or (_31858_, _31857_, _02177_);
  or (_31859_, _31858_, _31856_);
  nand (_31860_, _10049_, _02177_);
  and (_31861_, _31860_, _31859_);
  or (_31863_, _31861_, _01632_);
  nand (_31864_, _04657_, _01632_);
  and (_31865_, _31864_, _10364_);
  and (_31866_, _31865_, _31863_);
  or (_31867_, _31619_, \oc8051_golden_model_1.PSW [7]);
  or (_31868_, _10048_, _06518_);
  and (_31869_, _31868_, _10363_);
  and (_31870_, _31869_, _31867_);
  or (_31871_, _31870_, _31866_);
  and (_31872_, _31871_, _09861_);
  nor (_31874_, _31635_, _09861_);
  or (_31875_, _31874_, _09854_);
  or (_31876_, _31875_, _31872_);
  or (_31877_, _10048_, _09853_);
  and (_31878_, _31877_, _04788_);
  and (_31879_, _31878_, _31876_);
  and (_31880_, _09934_, _02071_);
  or (_31881_, _31880_, _02173_);
  or (_31882_, _31881_, _31879_);
  nand (_31883_, _10049_, _02173_);
  and (_31885_, _31883_, _31882_);
  or (_31886_, _31885_, _01648_);
  nand (_31887_, _04657_, _01648_);
  and (_31888_, _31887_, _09849_);
  and (_31889_, _31888_, _31886_);
  or (_31890_, _31889_, _31624_);
  and (_31891_, _31890_, _09846_);
  nor (_31892_, _31635_, _09846_);
  or (_31893_, _31892_, _07146_);
  or (_31894_, _31893_, _31891_);
  or (_31896_, _10048_, _07145_);
  and (_31897_, _31896_, _07176_);
  and (_31898_, _31897_, _31894_);
  and (_31899_, _31634_, _07175_);
  or (_31900_, _31899_, _02185_);
  or (_31901_, _31900_, _31898_);
  or (_31902_, _05135_, _09305_);
  and (_31903_, _31902_, _31901_);
  or (_31904_, _31903_, _01636_);
  nand (_31905_, _04657_, _01636_);
  and (_31906_, _31905_, _10403_);
  and (_31907_, _31906_, _31904_);
  or (_31908_, _31677_, _10408_);
  or (_31909_, _09934_, _08439_);
  and (_31910_, _31909_, _02083_);
  and (_31911_, _31910_, _31908_);
  or (_31912_, _31911_, _31907_);
  and (_31913_, _31912_, _09844_);
  nor (_31914_, _31635_, _09844_);
  or (_31915_, _31914_, _07255_);
  or (_31917_, _31915_, _31913_);
  or (_31918_, _10048_, _07254_);
  and (_31919_, _31918_, _07305_);
  and (_31920_, _31919_, _31917_);
  and (_31921_, _31634_, _07304_);
  or (_31922_, _31921_, _01888_);
  or (_31923_, _31922_, _31920_);
  or (_31924_, _05135_, _01889_);
  and (_31925_, _31924_, _10426_);
  and (_31926_, _31925_, _31923_);
  nor (_31928_, _04657_, _10426_);
  or (_31929_, _31928_, _02082_);
  or (_31930_, _31929_, _31926_);
  or (_31931_, _31677_, _08439_);
  or (_31932_, _09934_, _10408_);
  and (_31933_, _31932_, _31931_);
  or (_31934_, _31933_, _02202_);
  and (_31935_, _31934_, _10438_);
  and (_31936_, _31935_, _31930_);
  and (_31937_, _31634_, _10435_);
  or (_31939_, _31937_, _02201_);
  or (_31940_, _31939_, _31936_);
  nand (_31941_, _10049_, _02201_);
  and (_31942_, _31941_, _10442_);
  and (_31943_, _31942_, _31940_);
  nor (_31944_, _31635_, _10442_);
  or (_31945_, _31944_, _03370_);
  or (_31946_, _31945_, _31943_);
  and (_31947_, _31946_, _31617_);
  or (_31948_, _31947_, _01860_);
  or (_31950_, _31933_, _01887_);
  and (_31951_, _31950_, _10461_);
  and (_31952_, _31951_, _31948_);
  and (_31953_, _31634_, _10458_);
  or (_31954_, _31953_, _01537_);
  or (_31955_, _31954_, _31952_);
  nand (_31956_, _10049_, _01537_);
  and (_31957_, _31956_, _10465_);
  and (_31958_, _31957_, _31955_);
  nor (_31959_, _31635_, _10465_);
  or (_31961_, _31959_, _30482_);
  or (_31962_, _31961_, _31958_);
  nand (_31963_, _30482_, _04657_);
  and (_31964_, _31963_, _10481_);
  and (_31965_, _31964_, _31962_);
  and (_31966_, _31634_, _09829_);
  or (_31967_, _31966_, _38088_);
  or (_31968_, _31967_, _31965_);
  or (_31969_, _38087_, \oc8051_golden_model_1.PC [4]);
  and (_31970_, _31969_, _37580_);
  and (_40362_, _31970_, _31968_);
  or (_31972_, _38087_, \oc8051_golden_model_1.PC [5]);
  and (_31973_, _31972_, _37580_);
  and (_31974_, _10043_, _01537_);
  nor (_31975_, \oc8051_golden_model_1.PC [5], \oc8051_golden_model_1.PC [0]);
  nor (_31976_, _10043_, _01280_);
  nor (_31977_, _31976_, _31975_);
  or (_31978_, _31977_, _10442_);
  or (_31979_, _05090_, _01889_);
  or (_31980_, _31977_, _09844_);
  or (_31982_, _31977_, _09846_);
  or (_31983_, _31977_, _09861_);
  not (_31984_, _31977_);
  nand (_31985_, _31984_, _09863_);
  or (_31986_, _31977_, _10327_);
  or (_31987_, _10043_, _04757_);
  nand (_31988_, _10044_, _01875_);
  nand (_31989_, _31984_, _10219_);
  nand (_31990_, _31984_, _08628_);
  or (_31991_, _09932_, _09931_);
  nand (_31993_, _31991_, _09961_);
  or (_31994_, _31991_, _09961_);
  and (_31995_, _31994_, _31993_);
  or (_31996_, _31995_, _08498_);
  nand (_31997_, _09930_, _08498_);
  and (_31998_, _31997_, _31996_);
  or (_31999_, _31998_, _08494_);
  or (_32000_, _31995_, _09996_);
  or (_32001_, _09876_, _09929_);
  and (_32002_, _32001_, _32000_);
  or (_32004_, _32002_, _02814_);
  and (_32005_, _10107_, _10043_);
  or (_32006_, _10046_, _10045_);
  nand (_32007_, _32006_, _10070_);
  or (_32008_, _32006_, _10070_);
  and (_32009_, _32008_, _32007_);
  and (_32010_, _32009_, _10105_);
  or (_32011_, _32010_, _32005_);
  or (_32012_, _32011_, _04381_);
  nor (_32013_, _04626_, _01562_);
  nand (_32015_, _10044_, _02817_);
  and (_32016_, _32015_, _10121_);
  and (_32017_, _10113_, \oc8051_golden_model_1.PC [5]);
  or (_32018_, _32017_, _02817_);
  and (_32019_, _32018_, _32016_);
  nor (_32020_, _31984_, _21690_);
  or (_32021_, _32020_, _06629_);
  or (_32022_, _32021_, _32019_);
  and (_32023_, _32022_, _01562_);
  or (_32024_, _32023_, _32013_);
  nand (_32026_, _31984_, _06629_);
  and (_32027_, _32026_, _06618_);
  and (_32028_, _32027_, _32024_);
  and (_32029_, _10043_, _02003_);
  or (_32030_, _32029_, _06616_);
  or (_32031_, _32030_, _32028_);
  nand (_32032_, _31984_, _06616_);
  and (_32033_, _32032_, _01568_);
  and (_32034_, _32033_, _32031_);
  nor (_32035_, _04626_, _01568_);
  or (_32037_, _32035_, _04380_);
  or (_32038_, _32037_, _32034_);
  and (_32039_, _32038_, _04394_);
  and (_32040_, _32039_, _32012_);
  and (_32041_, _31977_, _01883_);
  or (_32042_, _32041_, _02001_);
  or (_32043_, _32042_, _32040_);
  and (_32044_, _32043_, _32004_);
  or (_32045_, _32044_, _30311_);
  or (_32046_, _31977_, _09871_);
  and (_32048_, _32046_, _02024_);
  and (_32049_, _32048_, _32045_);
  and (_32050_, _10043_, _02007_);
  or (_32051_, _32050_, _03279_);
  or (_32052_, _32051_, _32049_);
  nand (_32053_, _04626_, _03279_);
  and (_32054_, _32053_, _02840_);
  and (_32055_, _32054_, _32052_);
  nand (_32056_, _10043_, _01999_);
  nand (_32057_, _32056_, _10156_);
  or (_32058_, _32057_, _32055_);
  or (_32059_, _31977_, _10156_);
  and (_32060_, _32059_, _02021_);
  and (_32061_, _32060_, _32058_);
  nand (_32062_, _10043_, _02006_);
  nand (_32063_, _32062_, _10163_);
  or (_32064_, _32063_, _32061_);
  or (_32065_, _31977_, _10163_);
  and (_32066_, _32065_, _02025_);
  and (_32067_, _32066_, _32064_);
  and (_32069_, _10043_, _01997_);
  or (_32070_, _32069_, _10167_);
  or (_32071_, _32070_, _32067_);
  nand (_32072_, _04626_, _10167_);
  and (_32073_, _32072_, _01880_);
  and (_32074_, _32073_, _32071_);
  nand (_32075_, _10043_, _01878_);
  nand (_32076_, _32075_, _08538_);
  or (_32077_, _32076_, _32074_);
  or (_32078_, _31995_, _08572_);
  nand (_32080_, _09930_, _08572_);
  and (_32081_, _32080_, _32078_);
  or (_32082_, _32081_, _08538_);
  and (_32083_, _32082_, _32077_);
  or (_32084_, _32083_, _08493_);
  and (_32085_, _32084_, _31999_);
  or (_32086_, _32085_, _01995_);
  and (_32087_, _09929_, _08625_);
  and (_32088_, _31995_, _30342_);
  or (_32089_, _32088_, _02444_);
  or (_32091_, _32089_, _32087_);
  and (_32092_, _32091_, _02046_);
  and (_32093_, _32092_, _32086_);
  or (_32094_, _31995_, _08664_);
  nand (_32095_, _09930_, _08664_);
  and (_32096_, _32095_, _02045_);
  and (_32097_, _32096_, _32094_);
  or (_32098_, _32097_, _08628_);
  or (_32099_, _32098_, _32093_);
  and (_32100_, _32099_, _31990_);
  or (_32102_, _32100_, _01991_);
  nand (_32103_, _10044_, _01991_);
  and (_32104_, _32103_, _01565_);
  and (_32105_, _32104_, _32102_);
  nor (_32106_, _04626_, _01565_);
  or (_32107_, _32106_, _30633_);
  or (_32108_, _32107_, _32105_);
  or (_32109_, _30632_, _10043_);
  and (_32110_, _32109_, _32108_);
  or (_32111_, _32110_, _10211_);
  or (_32113_, _31977_, _10207_);
  and (_32114_, _32113_, _08249_);
  and (_32115_, _32114_, _32111_);
  and (_32116_, _10043_, _01967_);
  or (_32117_, _32116_, _10213_);
  or (_32118_, _32117_, _32115_);
  nand (_32119_, _04626_, _10213_);
  and (_32120_, _32119_, _08248_);
  and (_32121_, _32120_, _32118_);
  and (_32122_, _10043_, _01966_);
  or (_32124_, _32122_, _10219_);
  or (_32125_, _32124_, _32121_);
  and (_32126_, _32125_, _31989_);
  or (_32127_, _32126_, _06776_);
  or (_32128_, _10043_, _06775_);
  and (_32129_, _32128_, _01550_);
  and (_32130_, _32129_, _32127_);
  and (_32131_, _31977_, _01549_);
  or (_32132_, _32131_, _01875_);
  or (_32133_, _32132_, _32130_);
  and (_32135_, _32133_, _31988_);
  or (_32136_, _32135_, _01604_);
  nand (_32137_, _04626_, _01604_);
  and (_32138_, _32137_, _07401_);
  and (_32139_, _32138_, _32136_);
  nand (_32140_, _09929_, _02080_);
  nand (_32141_, _32140_, _09211_);
  or (_32142_, _32141_, _32139_);
  or (_32143_, _10043_, _09211_);
  and (_32144_, _32143_, _02043_);
  and (_32146_, _32144_, _32142_);
  nand (_32147_, _09929_, _01602_);
  nand (_32148_, _32147_, _10245_);
  or (_32149_, _32148_, _32146_);
  or (_32150_, _31977_, _10245_);
  and (_32151_, _32150_, _30680_);
  and (_32152_, _32151_, _32149_);
  nor (_32153_, _10043_, _01649_);
  nor (_32154_, _32153_, _10247_);
  or (_32155_, _32154_, _32152_);
  nand (_32157_, _04626_, _01649_);
  and (_32158_, _32157_, _10254_);
  and (_32159_, _32158_, _32155_);
  and (_32160_, _32009_, _10253_);
  or (_32161_, _32160_, _04758_);
  or (_32162_, _32161_, _32159_);
  and (_32163_, _32162_, _31987_);
  or (_32164_, _32163_, _01869_);
  nand (_32165_, _09930_, _01869_);
  and (_32166_, _32165_, _06985_);
  and (_32168_, _32166_, _32164_);
  and (_32169_, _10043_, _06984_);
  or (_32170_, _32169_, _10267_);
  or (_32171_, _32170_, _32168_);
  nor (_32172_, _10288_, _10280_);
  nor (_32173_, _32172_, _10289_);
  or (_32174_, _32173_, _10268_);
  and (_32175_, _32174_, _02576_);
  and (_32176_, _32175_, _32171_);
  and (_32177_, _10043_, _01958_);
  or (_32179_, _32177_, _01638_);
  or (_32180_, _32179_, _32176_);
  nand (_32181_, _04626_, _01638_);
  and (_32182_, _32181_, _10311_);
  and (_32183_, _32182_, _32180_);
  or (_32184_, _32009_, _07356_);
  or (_32185_, _10043_, _10316_);
  and (_32186_, _32185_, _10310_);
  and (_32187_, _32186_, _32184_);
  or (_32188_, _32187_, _10331_);
  or (_32190_, _32188_, _32183_);
  and (_32191_, _32190_, _31986_);
  or (_32192_, _32191_, _10330_);
  or (_32193_, _10043_, _10329_);
  and (_32194_, _32193_, _02166_);
  and (_32195_, _32194_, _32192_);
  and (_32196_, _09929_, _02079_);
  or (_32197_, _32196_, _02167_);
  or (_32198_, _32197_, _32195_);
  nand (_32199_, _10044_, _02167_);
  and (_32201_, _32199_, _32198_);
  or (_32202_, _32201_, _01645_);
  nand (_32203_, _04626_, _01645_);
  and (_32204_, _32203_, _10344_);
  and (_32205_, _32204_, _32202_);
  or (_32206_, _32009_, _10316_);
  or (_32207_, _10043_, _07356_);
  and (_32208_, _32207_, _10343_);
  and (_32209_, _32208_, _32206_);
  or (_32210_, _32209_, _09863_);
  or (_32211_, _32210_, _32205_);
  and (_32212_, _32211_, _31985_);
  or (_32213_, _32212_, _07042_);
  or (_32214_, _10043_, _07041_);
  and (_32215_, _32214_, _02176_);
  and (_32216_, _32215_, _32213_);
  and (_32217_, _09929_, _02072_);
  or (_32218_, _32217_, _02177_);
  or (_32219_, _32218_, _32216_);
  nand (_32220_, _10044_, _02177_);
  and (_32222_, _32220_, _32219_);
  or (_32223_, _32222_, _01632_);
  nand (_32224_, _04626_, _01632_);
  and (_32225_, _32224_, _10364_);
  and (_32226_, _32225_, _32223_);
  or (_32227_, _32009_, \oc8051_golden_model_1.PSW [7]);
  or (_32228_, _10043_, _06518_);
  and (_32229_, _32228_, _10363_);
  and (_32230_, _32229_, _32227_);
  or (_32231_, _32230_, _10368_);
  or (_32233_, _32231_, _32226_);
  and (_32234_, _32233_, _31983_);
  or (_32235_, _32234_, _09854_);
  or (_32236_, _10043_, _09853_);
  and (_32237_, _32236_, _04788_);
  and (_32238_, _32237_, _32235_);
  and (_32239_, _09929_, _02071_);
  or (_32240_, _32239_, _02173_);
  or (_32241_, _32240_, _32238_);
  nand (_32242_, _10044_, _02173_);
  and (_32244_, _32242_, _32241_);
  or (_32245_, _32244_, _01648_);
  nand (_32246_, _04626_, _01648_);
  and (_32247_, _32246_, _09849_);
  and (_32248_, _32247_, _32245_);
  or (_32249_, _32009_, _06518_);
  or (_32250_, _10043_, \oc8051_golden_model_1.PSW [7]);
  and (_32251_, _32250_, _09848_);
  and (_32252_, _32251_, _32249_);
  or (_32253_, _32252_, _10385_);
  or (_32255_, _32253_, _32248_);
  and (_32256_, _32255_, _31982_);
  or (_32257_, _32256_, _07146_);
  or (_32258_, _10043_, _07145_);
  and (_32259_, _32258_, _07176_);
  and (_32260_, _32259_, _32257_);
  and (_32261_, _31977_, _07175_);
  or (_32262_, _32261_, _02185_);
  or (_32263_, _32262_, _32260_);
  or (_32264_, _05090_, _09305_);
  and (_32266_, _32264_, _32263_);
  or (_32267_, _32266_, _01636_);
  nand (_32268_, _04626_, _01636_);
  and (_32269_, _32268_, _10403_);
  and (_32270_, _32269_, _32267_);
  or (_32271_, _31995_, _10408_);
  or (_32272_, _09929_, _08439_);
  and (_32273_, _32272_, _02083_);
  and (_32274_, _32273_, _32271_);
  or (_32275_, _32274_, _10407_);
  or (_32277_, _32275_, _32270_);
  and (_32278_, _32277_, _31980_);
  or (_32279_, _32278_, _07255_);
  or (_32280_, _10043_, _07254_);
  and (_32281_, _32280_, _07305_);
  and (_32282_, _32281_, _32279_);
  and (_32283_, _31977_, _07304_);
  or (_32284_, _32283_, _01888_);
  or (_32285_, _32284_, _32282_);
  and (_32286_, _32285_, _31979_);
  or (_32288_, _32286_, _01653_);
  nand (_32289_, _04626_, _01653_);
  and (_32290_, _32289_, _02202_);
  and (_32291_, _32290_, _32288_);
  or (_32292_, _31995_, _08439_);
  nand (_32293_, _09930_, _08439_);
  and (_32294_, _32293_, _32292_);
  and (_32295_, _32294_, _02082_);
  or (_32296_, _32295_, _10435_);
  or (_32297_, _32296_, _32291_);
  nand (_32299_, _31984_, _10435_);
  and (_32300_, _32299_, _02303_);
  and (_32301_, _32300_, _32297_);
  nand (_32302_, _10043_, _02201_);
  nand (_32303_, _32302_, _10442_);
  or (_32304_, _32303_, _32301_);
  and (_32305_, _32304_, _31978_);
  or (_32306_, _32305_, _03370_);
  nand (_32307_, _04626_, _03370_);
  and (_32308_, _32307_, _01887_);
  and (_32310_, _32308_, _32306_);
  and (_32311_, _32294_, _01860_);
  or (_32312_, _32311_, _10458_);
  or (_32313_, _32312_, _32310_);
  nand (_32314_, _31984_, _10458_);
  and (_32315_, _32314_, _01538_);
  and (_32316_, _32315_, _32313_);
  or (_32317_, _32316_, _31974_);
  and (_32318_, _32317_, _10465_);
  nor (_32319_, _31984_, _10465_);
  or (_32321_, _32319_, _30482_);
  or (_32322_, _32321_, _32318_);
  nand (_32323_, _30482_, _04626_);
  and (_32324_, _32323_, _10481_);
  and (_32325_, _32324_, _32322_);
  and (_32326_, _31977_, _09829_);
  or (_32327_, _32326_, _38088_);
  or (_32328_, _32327_, _32325_);
  and (_40363_, _32328_, _31973_);
  or (_32329_, _38087_, \oc8051_golden_model_1.PC [6]);
  and (_32331_, _32329_, _37580_);
  nand (_32332_, _04594_, _03370_);
  nor (_32333_, _09831_, \oc8051_golden_model_1.PC [6]);
  nor (_32334_, _32333_, _09832_);
  not (_32335_, _32334_);
  nand (_32336_, _32335_, _07304_);
  or (_32337_, _09923_, _04788_);
  or (_32338_, _09923_, _02176_);
  or (_32339_, _09923_, _02166_);
  nand (_32340_, _10037_, _01958_);
  or (_32341_, _10072_, _10040_);
  and (_32342_, _32341_, _10073_);
  and (_32343_, _32342_, _10253_);
  nand (_32344_, _32335_, _08628_);
  or (_32345_, _09923_, _30342_);
  or (_32346_, _09963_, _09926_);
  and (_32347_, _32346_, _09964_);
  or (_32348_, _32347_, _08625_);
  and (_32349_, _32348_, _01995_);
  and (_32350_, _32349_, _32345_);
  and (_32352_, _09923_, _08498_);
  and (_32353_, _32347_, _30279_);
  or (_32354_, _32353_, _32352_);
  and (_32355_, _32354_, _08493_);
  nand (_32356_, _10037_, _01997_);
  or (_32357_, _32334_, _10150_);
  not (_32358_, _10144_);
  nand (_32359_, _04594_, _02823_);
  nand (_32360_, _10037_, _02817_);
  and (_32361_, _32360_, _10121_);
  not (_32363_, \oc8051_golden_model_1.PC [6]);
  nor (_32364_, _10112_, _32363_);
  or (_32365_, _32364_, _02817_);
  and (_32366_, _32365_, _32361_);
  nor (_32367_, _32335_, _21690_);
  or (_32368_, _32367_, _02823_);
  or (_32369_, _32368_, _32366_);
  and (_32370_, _32369_, _10129_);
  and (_32371_, _32370_, _32359_);
  and (_32372_, _32334_, _06629_);
  or (_32374_, _32372_, _02003_);
  or (_32375_, _32374_, _32371_);
  nand (_32376_, _10037_, _02003_);
  and (_32377_, _32376_, _32375_);
  or (_32378_, _32377_, _06616_);
  nand (_32379_, _32335_, _06616_);
  and (_32380_, _32379_, _01568_);
  and (_32381_, _32380_, _32378_);
  nor (_32382_, _04594_, _01568_);
  or (_32383_, _32382_, _04380_);
  or (_32385_, _32383_, _32381_);
  and (_32386_, _32342_, _10105_);
  and (_32387_, _10107_, _10036_);
  or (_32388_, _32387_, _04381_);
  or (_32389_, _32388_, _32386_);
  and (_32390_, _32389_, _32385_);
  or (_32391_, _32390_, _32358_);
  and (_32392_, _32347_, _09876_);
  and (_32393_, _09996_, _09923_);
  or (_32394_, _32393_, _02814_);
  or (_32396_, _32394_, _32392_);
  and (_32397_, _32396_, _32391_);
  or (_32398_, _32397_, _30311_);
  and (_32399_, _32398_, _32357_);
  or (_32400_, _32399_, _02007_);
  nand (_32401_, _10037_, _02007_);
  and (_32402_, _32401_, _01558_);
  and (_32403_, _32402_, _32400_);
  nor (_32404_, _04594_, _01558_);
  or (_32405_, _32404_, _01999_);
  or (_32407_, _32405_, _32403_);
  nand (_32408_, _10037_, _01999_);
  and (_32409_, _32408_, _32407_);
  or (_32410_, _32409_, _10157_);
  or (_32411_, _32334_, _10156_);
  and (_32412_, _32411_, _32410_);
  or (_32413_, _32412_, _02006_);
  nand (_32414_, _10037_, _02006_);
  and (_32415_, _32414_, _10163_);
  and (_32416_, _32415_, _32413_);
  nor (_32418_, _32335_, _10163_);
  or (_32419_, _32418_, _01997_);
  or (_32420_, _32419_, _32416_);
  and (_32421_, _32420_, _32356_);
  or (_32422_, _32421_, _10167_);
  nand (_32423_, _04594_, _10167_);
  and (_32424_, _32423_, _01880_);
  and (_32425_, _32424_, _32422_);
  nand (_32426_, _10036_, _01878_);
  nand (_32427_, _32426_, _08538_);
  or (_32429_, _32427_, _32425_);
  and (_32430_, _09923_, _08572_);
  and (_32431_, _32347_, _08573_);
  or (_32432_, _32431_, _32430_);
  or (_32433_, _32432_, _08538_);
  and (_32434_, _32433_, _08494_);
  and (_32435_, _32434_, _32429_);
  or (_32436_, _32435_, _32355_);
  and (_32437_, _32436_, _02444_);
  or (_32438_, _32437_, _32350_);
  and (_32440_, _32438_, _02046_);
  and (_32441_, _09923_, _08664_);
  and (_32442_, _32347_, _31735_);
  or (_32443_, _32442_, _32441_);
  and (_32444_, _32443_, _02045_);
  or (_32445_, _32444_, _08628_);
  or (_32446_, _32445_, _32440_);
  and (_32447_, _32446_, _32344_);
  or (_32448_, _32447_, _01991_);
  nand (_32449_, _10037_, _01991_);
  and (_32451_, _32449_, _01565_);
  and (_32452_, _32451_, _32448_);
  nor (_32453_, _04594_, _01565_);
  or (_32454_, _32453_, _30633_);
  or (_32455_, _32454_, _32452_);
  or (_32456_, _30632_, _10036_);
  and (_32457_, _32456_, _32455_);
  or (_32458_, _32457_, _10211_);
  or (_32459_, _32334_, _10207_);
  and (_32460_, _32459_, _08249_);
  and (_32462_, _32460_, _32458_);
  and (_32463_, _10036_, _01967_);
  or (_32464_, _32463_, _10213_);
  or (_32465_, _32464_, _32462_);
  nand (_32466_, _04594_, _10213_);
  and (_32467_, _32466_, _08248_);
  and (_32468_, _32467_, _32465_);
  and (_32469_, _10036_, _01966_);
  or (_32470_, _32469_, _10219_);
  or (_32471_, _32470_, _32468_);
  nand (_32473_, _32335_, _10219_);
  and (_32474_, _32473_, _06775_);
  and (_32475_, _32474_, _32471_);
  nor (_32476_, _10037_, _06775_);
  or (_32477_, _32476_, _01549_);
  or (_32478_, _32477_, _32475_);
  nand (_32479_, _32335_, _01549_);
  and (_32480_, _32479_, _32478_);
  or (_32481_, _32480_, _01875_);
  nand (_32482_, _10037_, _01875_);
  and (_32483_, _32482_, _04310_);
  and (_32484_, _32483_, _32481_);
  nor (_32485_, _04594_, _04310_);
  or (_32486_, _32485_, _02080_);
  or (_32487_, _32486_, _32484_);
  or (_32488_, _09923_, _07401_);
  and (_32489_, _32488_, _32487_);
  or (_32490_, _32489_, _09212_);
  or (_32491_, _10036_, _09211_);
  and (_32492_, _32491_, _32490_);
  or (_32493_, _32492_, _01602_);
  or (_32494_, _09923_, _02043_);
  and (_32495_, _32494_, _10245_);
  and (_32496_, _32495_, _32493_);
  nor (_32497_, _32335_, _10245_);
  or (_32498_, _32497_, _01959_);
  or (_32499_, _32498_, _32496_);
  nand (_32500_, _10037_, _01959_);
  and (_32501_, _32500_, _30378_);
  and (_32502_, _32501_, _32499_);
  nor (_32503_, _04594_, _30378_);
  or (_32504_, _32503_, _32502_);
  and (_32505_, _32504_, _10254_);
  or (_32506_, _32505_, _32343_);
  and (_32507_, _32506_, _04757_);
  nor (_32508_, _10037_, _04757_);
  or (_32509_, _32508_, _01869_);
  or (_32510_, _32509_, _32507_);
  or (_32511_, _09923_, _01870_);
  and (_32512_, _32511_, _06985_);
  and (_32514_, _32512_, _32510_);
  and (_32515_, _10036_, _06984_);
  or (_32516_, _32515_, _10267_);
  or (_32517_, _32516_, _32514_);
  or (_32518_, _10290_, _10277_);
  and (_32519_, _32518_, _10291_);
  or (_32520_, _32519_, _10268_);
  and (_32521_, _32520_, _32517_);
  or (_32522_, _32521_, _01958_);
  and (_32523_, _32522_, _32340_);
  or (_32525_, _32523_, _01638_);
  nand (_32526_, _04594_, _01638_);
  and (_32527_, _32526_, _10311_);
  and (_32528_, _32527_, _32525_);
  or (_32529_, _32342_, _07356_);
  or (_32530_, _10036_, _10316_);
  and (_32531_, _32530_, _10310_);
  and (_32532_, _32531_, _32529_);
  or (_32533_, _32532_, _10331_);
  or (_32534_, _32533_, _32528_);
  or (_32535_, _32334_, _10327_);
  and (_32536_, _32535_, _10329_);
  and (_32537_, _32536_, _32534_);
  nor (_32538_, _10037_, _10329_);
  or (_32539_, _32538_, _02079_);
  or (_32540_, _32539_, _32537_);
  and (_32541_, _32540_, _32339_);
  or (_32542_, _32541_, _02167_);
  nand (_32543_, _10037_, _02167_);
  and (_32544_, _32543_, _30413_);
  and (_32546_, _32544_, _32542_);
  nor (_32547_, _04594_, _30413_);
  or (_32548_, _32547_, _32546_);
  and (_32549_, _32548_, _10344_);
  or (_32550_, _32342_, _10316_);
  or (_32551_, _10036_, _07356_);
  and (_32552_, _32551_, _10343_);
  and (_32553_, _32552_, _32550_);
  or (_32554_, _32553_, _09863_);
  or (_32555_, _32554_, _32549_);
  nand (_32557_, _32335_, _09863_);
  and (_32558_, _32557_, _07041_);
  and (_32559_, _32558_, _32555_);
  nor (_32560_, _10037_, _07041_);
  or (_32561_, _32560_, _02072_);
  or (_32562_, _32561_, _32559_);
  and (_32563_, _32562_, _32338_);
  or (_32564_, _32563_, _02177_);
  nand (_32565_, _10037_, _02177_);
  and (_32566_, _32565_, _01633_);
  and (_32568_, _32566_, _32564_);
  nor (_32569_, _04594_, _01633_);
  or (_32570_, _32569_, _32568_);
  and (_32571_, _32570_, _10364_);
  or (_32572_, _32342_, \oc8051_golden_model_1.PSW [7]);
  or (_32573_, _10036_, _06518_);
  and (_32574_, _32573_, _10363_);
  and (_32575_, _32574_, _32572_);
  or (_32576_, _32575_, _10368_);
  or (_32577_, _32576_, _32571_);
  or (_32579_, _32334_, _09861_);
  and (_32580_, _32579_, _09853_);
  and (_32581_, _32580_, _32577_);
  nor (_32582_, _10037_, _09853_);
  or (_32583_, _32582_, _02071_);
  or (_32584_, _32583_, _32581_);
  and (_32585_, _32584_, _32337_);
  or (_32586_, _32585_, _02173_);
  nand (_32587_, _10037_, _02173_);
  and (_32588_, _32587_, _30272_);
  and (_32590_, _32588_, _32586_);
  nor (_32591_, _04594_, _30272_);
  or (_32592_, _32591_, _32590_);
  and (_32593_, _32592_, _09849_);
  or (_32594_, _32342_, _06518_);
  or (_32595_, _10036_, \oc8051_golden_model_1.PSW [7]);
  and (_32596_, _32595_, _09848_);
  and (_32597_, _32596_, _32594_);
  or (_32598_, _32597_, _10385_);
  or (_32599_, _32598_, _32593_);
  or (_32601_, _32334_, _09846_);
  and (_32602_, _32601_, _07145_);
  and (_32603_, _32602_, _32599_);
  nor (_32604_, _10037_, _07145_);
  or (_32605_, _32604_, _07175_);
  or (_32606_, _32605_, _32603_);
  nand (_32607_, _32335_, _07175_);
  and (_32608_, _32607_, _09305_);
  and (_32609_, _32608_, _32606_);
  and (_32610_, _04861_, _02185_);
  or (_32612_, _32610_, _01636_);
  or (_32613_, _32612_, _32609_);
  nand (_32614_, _04594_, _01636_);
  and (_32615_, _32614_, _10403_);
  and (_32616_, _32615_, _32613_);
  or (_32617_, _32347_, _10408_);
  or (_32618_, _09923_, _08439_);
  and (_32619_, _32618_, _02083_);
  and (_32620_, _32619_, _32617_);
  or (_32621_, _32620_, _10407_);
  or (_32623_, _32621_, _32616_);
  or (_32624_, _32334_, _09844_);
  and (_32625_, _32624_, _07254_);
  and (_32626_, _32625_, _32623_);
  nor (_32627_, _10037_, _07254_);
  or (_32628_, _32627_, _07304_);
  or (_32629_, _32628_, _32626_);
  and (_32630_, _32629_, _32336_);
  or (_32631_, _32630_, _01888_);
  or (_32632_, _04861_, _01889_);
  and (_32634_, _32632_, _10426_);
  and (_32635_, _32634_, _32631_);
  nor (_32636_, _04594_, _10426_);
  or (_32637_, _32636_, _02082_);
  or (_32638_, _32637_, _32635_);
  or (_32639_, _09923_, _10408_);
  or (_32640_, _32347_, _08439_);
  and (_32641_, _32640_, _32639_);
  or (_32642_, _32641_, _02202_);
  and (_32643_, _32642_, _32638_);
  or (_32645_, _32643_, _10435_);
  nand (_32646_, _32335_, _10435_);
  and (_32647_, _32646_, _32645_);
  or (_32648_, _32647_, _02201_);
  nand (_32649_, _10037_, _02201_);
  and (_32650_, _32649_, _10442_);
  and (_32651_, _32650_, _32648_);
  nor (_32652_, _32335_, _10442_);
  or (_32653_, _32652_, _03370_);
  or (_32654_, _32653_, _32651_);
  and (_32656_, _32654_, _32332_);
  or (_32657_, _32656_, _01860_);
  or (_32658_, _32641_, _01887_);
  and (_32659_, _32658_, _10461_);
  and (_32660_, _32659_, _32657_);
  and (_32661_, _32334_, _10458_);
  or (_32662_, _32661_, _01537_);
  or (_32663_, _32662_, _32660_);
  nand (_32664_, _10037_, _01537_);
  and (_32665_, _32664_, _10465_);
  and (_32667_, _32665_, _32663_);
  nor (_32668_, _32335_, _10465_);
  or (_32669_, _32668_, _30482_);
  or (_32670_, _32669_, _32667_);
  nand (_32671_, _30482_, _04594_);
  and (_32672_, _32671_, _10481_);
  and (_32673_, _32672_, _32670_);
  and (_32674_, _32334_, _09829_);
  or (_32675_, _32674_, _38088_);
  or (_32676_, _32675_, _32673_);
  and (_40364_, _32676_, _32331_);
  and (_32678_, _04387_, _01537_);
  and (_32679_, _04387_, _02201_);
  and (_32680_, _04269_, _09830_);
  and (_32681_, _32680_, \oc8051_golden_model_1.PC [7]);
  nor (_32682_, _32680_, \oc8051_golden_model_1.PC [7]);
  nor (_32683_, _32682_, _32681_);
  or (_32684_, _32683_, _09844_);
  or (_32685_, _32683_, _09846_);
  or (_32686_, _32683_, _09861_);
  not (_32688_, _32683_);
  nand (_32689_, _32688_, _09863_);
  or (_32690_, _32683_, _10327_);
  or (_32691_, _04757_, _04387_);
  nand (_32692_, _04388_, _01875_);
  nand (_32693_, _32688_, _10219_);
  nand (_32694_, _32688_, _08628_);
  or (_32695_, _09918_, _09919_);
  nand (_32696_, _32695_, _09965_);
  or (_32697_, _32695_, _09965_);
  and (_32699_, _32697_, _32696_);
  or (_32700_, _32699_, _08498_);
  nand (_32701_, _08498_, _04275_);
  and (_32702_, _32701_, _32700_);
  or (_32703_, _32702_, _08494_);
  or (_32704_, _09876_, _04274_);
  or (_32705_, _32699_, _09996_);
  and (_32706_, _32705_, _32704_);
  or (_32707_, _32706_, _02814_);
  and (_32708_, _10107_, _04387_);
  or (_32710_, _10032_, _10033_);
  nand (_32711_, _32710_, _10074_);
  or (_32712_, _32710_, _10074_);
  and (_32713_, _32712_, _32711_);
  and (_32714_, _32713_, _10105_);
  or (_32715_, _32714_, _32708_);
  or (_32716_, _32715_, _04381_);
  nor (_32717_, _04307_, _01562_);
  nand (_32718_, _04388_, _02817_);
  and (_32719_, _32718_, _10121_);
  and (_32721_, _10113_, \oc8051_golden_model_1.PC [7]);
  or (_32722_, _32721_, _02817_);
  and (_32723_, _32722_, _32719_);
  nor (_32724_, _32688_, _21690_);
  or (_32725_, _32724_, _06629_);
  or (_32726_, _32725_, _32723_);
  and (_32727_, _32726_, _01562_);
  or (_32728_, _32727_, _32717_);
  nand (_32729_, _32688_, _06629_);
  and (_32730_, _32729_, _06618_);
  and (_32732_, _32730_, _32728_);
  and (_32733_, _04387_, _02003_);
  or (_32734_, _32733_, _06616_);
  or (_32735_, _32734_, _32732_);
  nand (_32736_, _32688_, _06616_);
  and (_32737_, _32736_, _01568_);
  and (_32738_, _32737_, _32735_);
  nor (_32739_, _04307_, _01568_);
  or (_32740_, _32739_, _04380_);
  or (_32741_, _32740_, _32738_);
  and (_32743_, _32741_, _04394_);
  and (_32744_, _32743_, _32716_);
  and (_32745_, _32683_, _01883_);
  or (_32746_, _32745_, _02001_);
  or (_32747_, _32746_, _32744_);
  and (_32748_, _32747_, _32707_);
  or (_32749_, _32748_, _30311_);
  or (_32750_, _32683_, _09871_);
  and (_32751_, _32750_, _02024_);
  and (_32752_, _32751_, _32749_);
  and (_32754_, _04387_, _02007_);
  or (_32755_, _32754_, _03279_);
  or (_32756_, _32755_, _32752_);
  nand (_32757_, _04307_, _03279_);
  and (_32758_, _32757_, _02840_);
  and (_32759_, _32758_, _32756_);
  nand (_32760_, _04387_, _01999_);
  nand (_32761_, _32760_, _10156_);
  or (_32762_, _32761_, _32759_);
  or (_32763_, _32683_, _10156_);
  and (_32765_, _32763_, _02021_);
  and (_32766_, _32765_, _32762_);
  nand (_32767_, _04387_, _02006_);
  nand (_32768_, _32767_, _10163_);
  or (_32769_, _32768_, _32766_);
  or (_32770_, _32683_, _10163_);
  and (_32771_, _32770_, _02025_);
  and (_32772_, _32771_, _32769_);
  and (_32773_, _04387_, _01997_);
  or (_32774_, _32773_, _10167_);
  or (_32776_, _32774_, _32772_);
  nand (_32777_, _04307_, _10167_);
  and (_32778_, _32777_, _01880_);
  and (_32779_, _32778_, _32776_);
  nand (_32780_, _04387_, _01878_);
  nand (_32781_, _32780_, _08538_);
  or (_32782_, _32781_, _32779_);
  or (_32783_, _32699_, _08572_);
  nand (_32784_, _08572_, _04275_);
  and (_32785_, _32784_, _32783_);
  or (_32787_, _32785_, _08538_);
  and (_32788_, _32787_, _32782_);
  or (_32789_, _32788_, _08493_);
  and (_32790_, _32789_, _32703_);
  or (_32791_, _32790_, _01995_);
  and (_32792_, _32699_, _30342_);
  and (_32793_, _08625_, _04274_);
  or (_32794_, _32793_, _02444_);
  or (_32795_, _32794_, _32792_);
  and (_32796_, _32795_, _02046_);
  and (_32798_, _32796_, _32791_);
  or (_32799_, _32699_, _08664_);
  nand (_32800_, _08664_, _04275_);
  and (_32801_, _32800_, _02045_);
  and (_32802_, _32801_, _32799_);
  or (_32803_, _32802_, _08628_);
  or (_32804_, _32803_, _32798_);
  and (_32805_, _32804_, _32694_);
  or (_32806_, _32805_, _01991_);
  nand (_32807_, _04388_, _01991_);
  and (_32809_, _32807_, _01565_);
  and (_32810_, _32809_, _32806_);
  nor (_32811_, _04307_, _01565_);
  or (_32812_, _32811_, _30633_);
  or (_32813_, _32812_, _32810_);
  or (_32814_, _30632_, _04387_);
  and (_32815_, _32814_, _32813_);
  or (_32816_, _32815_, _10211_);
  or (_32817_, _32683_, _10207_);
  and (_32818_, _32817_, _08249_);
  and (_32820_, _32818_, _32816_);
  and (_32821_, _04387_, _01967_);
  or (_32822_, _32821_, _10213_);
  or (_32823_, _32822_, _32820_);
  nand (_32824_, _04307_, _10213_);
  and (_32825_, _32824_, _08248_);
  and (_32826_, _32825_, _32823_);
  and (_32827_, _04387_, _01966_);
  or (_32828_, _32827_, _10219_);
  or (_32829_, _32828_, _32826_);
  and (_32831_, _32829_, _32693_);
  or (_32832_, _32831_, _06776_);
  or (_32833_, _06775_, _04387_);
  and (_32834_, _32833_, _01550_);
  and (_32835_, _32834_, _32832_);
  and (_32836_, _32683_, _01549_);
  or (_32837_, _32836_, _01875_);
  or (_32838_, _32837_, _32835_);
  and (_32839_, _32838_, _32692_);
  or (_32840_, _32839_, _01604_);
  nand (_32842_, _04307_, _01604_);
  and (_32843_, _32842_, _07401_);
  and (_32844_, _32843_, _32840_);
  nand (_32845_, _04274_, _02080_);
  nand (_32846_, _32845_, _09211_);
  or (_32847_, _32846_, _32844_);
  or (_32848_, _09211_, _04387_);
  and (_32849_, _32848_, _02043_);
  and (_32850_, _32849_, _32847_);
  nand (_32851_, _04274_, _01602_);
  nand (_32853_, _32851_, _10245_);
  or (_32854_, _32853_, _32850_);
  or (_32855_, _32683_, _10245_);
  and (_32856_, _32855_, _30680_);
  and (_32857_, _32856_, _32854_);
  nor (_32858_, _04387_, _01649_);
  nor (_32859_, _32858_, _10247_);
  or (_32860_, _32859_, _32857_);
  nand (_32861_, _04307_, _01649_);
  and (_32862_, _32861_, _10254_);
  and (_32864_, _32862_, _32860_);
  and (_32865_, _32713_, _10253_);
  or (_32866_, _32865_, _04758_);
  or (_32867_, _32866_, _32864_);
  and (_32868_, _32867_, _32691_);
  or (_32869_, _32868_, _01869_);
  nand (_32870_, _04275_, _01869_);
  and (_32871_, _32870_, _06985_);
  and (_32872_, _32871_, _32869_);
  and (_32873_, _06984_, _04387_);
  or (_32875_, _32873_, _10267_);
  or (_32876_, _32875_, _32872_);
  or (_32877_, _10273_, _10274_);
  nand (_32878_, _32877_, _10292_);
  or (_32879_, _32877_, _10292_);
  and (_32880_, _32879_, _32878_);
  or (_32881_, _32880_, _10268_);
  and (_32882_, _32881_, _02576_);
  and (_32883_, _32882_, _32876_);
  and (_32884_, _04387_, _01958_);
  or (_32886_, _32884_, _01638_);
  or (_32887_, _32886_, _32883_);
  nand (_32888_, _04307_, _01638_);
  and (_32889_, _32888_, _10311_);
  and (_32890_, _32889_, _32887_);
  or (_32891_, _32713_, _07356_);
  or (_32892_, _10316_, _04387_);
  and (_32893_, _32892_, _10310_);
  and (_32894_, _32893_, _32891_);
  or (_32895_, _32894_, _10331_);
  or (_32896_, _32895_, _32890_);
  and (_32897_, _32896_, _32690_);
  or (_32898_, _32897_, _10330_);
  or (_32899_, _10329_, _04387_);
  and (_32900_, _32899_, _02166_);
  and (_32901_, _32900_, _32898_);
  and (_32902_, _04274_, _02079_);
  or (_32903_, _32902_, _02167_);
  or (_32904_, _32903_, _32901_);
  nand (_32905_, _04388_, _02167_);
  and (_32907_, _32905_, _32904_);
  or (_32908_, _32907_, _01645_);
  nand (_32909_, _04307_, _01645_);
  and (_32910_, _32909_, _10344_);
  and (_32911_, _32910_, _32908_);
  or (_32912_, _32713_, _10316_);
  or (_32913_, _07356_, _04387_);
  and (_32914_, _32913_, _10343_);
  and (_32915_, _32914_, _32912_);
  or (_32916_, _32915_, _09863_);
  or (_32918_, _32916_, _32911_);
  and (_32919_, _32918_, _32689_);
  or (_32920_, _32919_, _07042_);
  or (_32921_, _07041_, _04387_);
  and (_32922_, _32921_, _02176_);
  and (_32923_, _32922_, _32920_);
  and (_32924_, _04274_, _02072_);
  or (_32925_, _32924_, _02177_);
  or (_32926_, _32925_, _32923_);
  nand (_32927_, _04388_, _02177_);
  and (_32929_, _32927_, _32926_);
  or (_32930_, _32929_, _01632_);
  nand (_32931_, _04307_, _01632_);
  and (_32932_, _32931_, _10364_);
  and (_32933_, _32932_, _32930_);
  or (_32934_, _32713_, \oc8051_golden_model_1.PSW [7]);
  or (_32935_, _04387_, _06518_);
  and (_32936_, _32935_, _10363_);
  and (_32937_, _32936_, _32934_);
  or (_32938_, _32937_, _10368_);
  or (_32940_, _32938_, _32933_);
  and (_32941_, _32940_, _32686_);
  or (_32942_, _32941_, _09854_);
  or (_32943_, _09853_, _04387_);
  and (_32944_, _32943_, _04788_);
  and (_32945_, _32944_, _32942_);
  and (_32946_, _04274_, _02071_);
  or (_32947_, _32946_, _02173_);
  or (_32948_, _32947_, _32945_);
  nand (_32949_, _04388_, _02173_);
  and (_32951_, _32949_, _32948_);
  or (_32952_, _32951_, _01648_);
  nand (_32953_, _04307_, _01648_);
  and (_32954_, _32953_, _09849_);
  and (_32955_, _32954_, _32952_);
  or (_32956_, _32713_, _06518_);
  or (_32957_, _04387_, \oc8051_golden_model_1.PSW [7]);
  and (_32958_, _32957_, _09848_);
  and (_32959_, _32958_, _32956_);
  or (_32960_, _32959_, _10385_);
  or (_32962_, _32960_, _32955_);
  and (_32963_, _32962_, _32685_);
  or (_32964_, _32963_, _07146_);
  or (_32965_, _07145_, _04387_);
  and (_32966_, _32965_, _07176_);
  and (_32967_, _32966_, _32964_);
  and (_32968_, _32683_, _07175_);
  or (_32969_, _32968_, _02185_);
  or (_32970_, _32969_, _32967_);
  or (_32971_, _04483_, _09305_);
  and (_32973_, _32971_, _32970_);
  or (_32974_, _32973_, _01636_);
  nand (_32975_, _04307_, _01636_);
  and (_32976_, _32975_, _10403_);
  and (_32977_, _32976_, _32974_);
  or (_32978_, _32699_, _10408_);
  or (_32979_, _08439_, _04274_);
  and (_32980_, _32979_, _02083_);
  and (_32981_, _32980_, _32978_);
  or (_32982_, _32981_, _10407_);
  or (_32984_, _32982_, _32977_);
  and (_32985_, _32984_, _32684_);
  or (_32986_, _32985_, _07255_);
  or (_32987_, _07254_, _04387_);
  and (_32988_, _32987_, _07305_);
  and (_32989_, _32988_, _32986_);
  and (_32990_, _32683_, _07304_);
  or (_32991_, _32990_, _01888_);
  or (_32992_, _32991_, _32989_);
  or (_32993_, _04483_, _01889_);
  and (_32995_, _32993_, _32992_);
  or (_32996_, _32995_, _01653_);
  nand (_32997_, _04307_, _01653_);
  and (_32998_, _32997_, _02202_);
  and (_32999_, _32998_, _32996_);
  nand (_33000_, _08439_, _04275_);
  or (_33001_, _32699_, _08439_);
  and (_33002_, _33001_, _33000_);
  and (_33003_, _33002_, _02082_);
  or (_33004_, _33003_, _10435_);
  or (_33006_, _33004_, _32999_);
  nand (_33007_, _32688_, _10435_);
  and (_33008_, _33007_, _02303_);
  and (_33009_, _33008_, _33006_);
  or (_33010_, _33009_, _32679_);
  and (_33011_, _33010_, _10442_);
  nor (_33012_, _32688_, _10442_);
  or (_33013_, _33012_, _03370_);
  or (_33014_, _33013_, _33011_);
  nand (_33015_, _04307_, _03370_);
  and (_33017_, _33015_, _01887_);
  and (_33018_, _33017_, _33014_);
  and (_33019_, _33002_, _01860_);
  or (_33020_, _33019_, _10458_);
  or (_33021_, _33020_, _33018_);
  nand (_33022_, _32688_, _10458_);
  and (_33023_, _33022_, _01538_);
  and (_33024_, _33023_, _33021_);
  or (_33025_, _33024_, _32678_);
  and (_33026_, _33025_, _10465_);
  nor (_33028_, _32688_, _10465_);
  or (_33029_, _33028_, _30482_);
  or (_33030_, _33029_, _33026_);
  nand (_33031_, _30482_, _04307_);
  and (_33032_, _33031_, _10481_);
  and (_33033_, _33032_, _33030_);
  and (_33034_, _32683_, _09829_);
  or (_33035_, _33034_, _38088_);
  or (_33036_, _33035_, _33033_);
  or (_33037_, _38087_, \oc8051_golden_model_1.PC [7]);
  and (_33039_, _33037_, _37580_);
  and (_40365_, _33039_, _33036_);
  or (_33040_, _38087_, \oc8051_golden_model_1.PC [8]);
  and (_33041_, _33040_, _37580_);
  nor (_33042_, _02441_, _10470_);
  nor (_33043_, _02441_, _05195_);
  nor (_33044_, _09848_, _01648_);
  or (_33045_, _09969_, _02176_);
  or (_33046_, _10030_, _04757_);
  nor (_33047_, _10253_, _01649_);
  and (_33049_, _10030_, _01959_);
  nor (_33050_, _32681_, \oc8051_golden_model_1.PC [8]);
  and (_33051_, _32681_, \oc8051_golden_model_1.PC [8]);
  nor (_33052_, _33051_, _33050_);
  not (_33053_, _33052_);
  nand (_33054_, _33053_, _01549_);
  or (_33055_, _09972_, _09967_);
  and (_33056_, _33055_, _09973_);
  or (_33057_, _33056_, _08498_);
  or (_33058_, _09969_, _30279_);
  and (_33060_, _33058_, _33057_);
  or (_33061_, _33060_, _08494_);
  and (_33062_, _10030_, _01997_);
  nor (_33063_, _01999_, _03279_);
  and (_33064_, _10030_, _02007_);
  or (_33065_, _09876_, _09969_);
  or (_33066_, _33056_, _09996_);
  and (_33067_, _33066_, _33065_);
  or (_33068_, _33067_, _02814_);
  and (_33069_, _10107_, _10030_);
  or (_33071_, _10078_, _10076_);
  and (_33072_, _33071_, _10079_);
  and (_33073_, _33072_, _10105_);
  or (_33074_, _33073_, _33069_);
  or (_33075_, _33074_, _04381_);
  or (_33076_, _33052_, _30286_);
  and (_33077_, _10030_, _02817_);
  and (_33078_, _02818_, \oc8051_golden_model_1.PC [8]);
  and (_33079_, _33078_, _21690_);
  or (_33080_, _33079_, _10125_);
  and (_33082_, _33080_, _06618_);
  or (_33083_, _33082_, _33077_);
  and (_33084_, _33083_, _33076_);
  nand (_33085_, _21690_, _10136_);
  and (_33086_, _33085_, _33052_);
  nand (_33087_, _10030_, _02003_);
  nand (_33088_, _33087_, _21702_);
  or (_33089_, _33088_, _33086_);
  or (_33090_, _33089_, _33084_);
  and (_33091_, _33090_, _04394_);
  and (_33093_, _33091_, _33075_);
  and (_33094_, _33052_, _01883_);
  or (_33095_, _33094_, _02001_);
  or (_33096_, _33095_, _33093_);
  and (_33097_, _33096_, _33068_);
  or (_33098_, _33097_, _30311_);
  or (_33099_, _33052_, _09871_);
  and (_33100_, _33099_, _02024_);
  and (_33101_, _33100_, _33098_);
  or (_33102_, _33101_, _33064_);
  and (_33104_, _33102_, _33063_);
  nand (_33105_, _10030_, _01999_);
  nand (_33106_, _33105_, _10156_);
  or (_33107_, _33106_, _33104_);
  or (_33108_, _33052_, _10156_);
  and (_33109_, _33108_, _02021_);
  and (_33110_, _33109_, _33107_);
  nand (_33111_, _10030_, _02006_);
  nand (_33112_, _33111_, _10163_);
  or (_33113_, _33112_, _33110_);
  or (_33115_, _33052_, _10163_);
  and (_33116_, _33115_, _02025_);
  and (_33117_, _33116_, _33113_);
  or (_33118_, _33117_, _33062_);
  and (_33119_, _33118_, _10168_);
  nand (_33120_, _10030_, _01878_);
  nand (_33121_, _33120_, _08538_);
  or (_33122_, _33121_, _33119_);
  and (_33123_, _09969_, _08572_);
  and (_33124_, _33056_, _08573_);
  or (_33126_, _33124_, _33123_);
  or (_33127_, _33126_, _08538_);
  and (_33128_, _33127_, _33122_);
  or (_33129_, _33128_, _08493_);
  and (_33130_, _33129_, _33061_);
  or (_33131_, _33130_, _01995_);
  and (_33132_, _09969_, _08625_);
  and (_33133_, _33056_, _30342_);
  or (_33134_, _33133_, _02444_);
  or (_33135_, _33134_, _33132_);
  and (_33137_, _33135_, _02046_);
  and (_33138_, _33137_, _33131_);
  or (_33139_, _33056_, _08664_);
  or (_33140_, _09969_, _31735_);
  and (_33141_, _33140_, _02045_);
  and (_33142_, _33141_, _33139_);
  or (_33143_, _33142_, _08628_);
  or (_33144_, _33143_, _33138_);
  nand (_33145_, _33053_, _08628_);
  and (_33146_, _33145_, _02861_);
  and (_33148_, _33146_, _33144_);
  and (_33149_, _10030_, _01991_);
  or (_33150_, _33149_, _03131_);
  or (_33151_, _33150_, _33148_);
  and (_33152_, _33151_, _30632_);
  nor (_33153_, _30632_, _10685_);
  or (_33154_, _33153_, _10211_);
  or (_33155_, _33154_, _33152_);
  or (_33156_, _33052_, _10207_);
  and (_33157_, _33156_, _08249_);
  and (_33159_, _33157_, _33155_);
  and (_33160_, _10030_, _01967_);
  or (_33161_, _33160_, _10213_);
  or (_33162_, _33161_, _33159_);
  and (_33163_, _33162_, _08248_);
  and (_33164_, _10030_, _01966_);
  or (_33165_, _33164_, _10219_);
  or (_33166_, _33165_, _33163_);
  nand (_33167_, _33053_, _10219_);
  and (_33168_, _33167_, _06775_);
  and (_33170_, _33168_, _33166_);
  nor (_33171_, _10685_, _06775_);
  or (_33172_, _33171_, _01549_);
  or (_33173_, _33172_, _33170_);
  and (_33174_, _33173_, _33054_);
  or (_33175_, _33174_, _01875_);
  nand (_33176_, _10685_, _01875_);
  and (_33177_, _33176_, _22053_);
  and (_33178_, _33177_, _33175_);
  nand (_33179_, _09969_, _02080_);
  nand (_33181_, _33179_, _09211_);
  or (_33182_, _33181_, _33178_);
  or (_33183_, _10030_, _09211_);
  and (_33184_, _33183_, _02043_);
  and (_33185_, _33184_, _33182_);
  nand (_33186_, _09969_, _01602_);
  nand (_33187_, _33186_, _10245_);
  or (_33188_, _33187_, _33185_);
  or (_33189_, _33052_, _10245_);
  and (_33190_, _33189_, _30680_);
  and (_33192_, _33190_, _33188_);
  or (_33193_, _33192_, _33049_);
  and (_33194_, _33193_, _33047_);
  and (_33195_, _33072_, _10253_);
  or (_33196_, _33195_, _04758_);
  or (_33197_, _33196_, _33194_);
  and (_33198_, _33197_, _33046_);
  or (_33199_, _33198_, _01869_);
  or (_33200_, _09969_, _01870_);
  and (_33201_, _33200_, _06985_);
  and (_33203_, _33201_, _33199_);
  and (_33204_, _10030_, _06984_);
  or (_33205_, _33204_, _10267_);
  or (_33206_, _33205_, _33203_);
  nor (_33207_, _10294_, \oc8051_golden_model_1.DPH [0]);
  nor (_33208_, _33207_, _10295_);
  or (_33209_, _33208_, _10268_);
  and (_33210_, _33209_, _02576_);
  and (_33211_, _33210_, _33206_);
  and (_33212_, _10030_, _01958_);
  or (_33214_, _33212_, _01638_);
  or (_33215_, _33214_, _33211_);
  and (_33216_, _33215_, _10311_);
  or (_33217_, _33072_, _07356_);
  or (_33218_, _10030_, _10316_);
  and (_33219_, _33218_, _10310_);
  and (_33220_, _33219_, _33217_);
  or (_33221_, _33220_, _10331_);
  or (_33222_, _33221_, _33216_);
  or (_33223_, _33052_, _10327_);
  and (_33225_, _33223_, _10329_);
  and (_33226_, _33225_, _33222_);
  nor (_33227_, _10685_, _10329_);
  or (_33228_, _33227_, _02079_);
  or (_33229_, _33228_, _33226_);
  or (_33230_, _09969_, _02166_);
  and (_33231_, _33230_, _02912_);
  and (_33232_, _33231_, _33229_);
  and (_33233_, _10030_, _02167_);
  or (_33234_, _33233_, _01645_);
  or (_33236_, _33234_, _33232_);
  and (_33237_, _33236_, _10344_);
  or (_33238_, _33072_, _10316_);
  or (_33239_, _10030_, _07356_);
  and (_33240_, _33239_, _10343_);
  and (_33241_, _33240_, _33238_);
  or (_33242_, _33241_, _09863_);
  or (_33243_, _33242_, _33237_);
  nand (_33244_, _33053_, _09863_);
  and (_33245_, _33244_, _07041_);
  and (_33247_, _33245_, _33243_);
  nor (_33248_, _10685_, _07041_);
  or (_33249_, _33248_, _02072_);
  or (_33250_, _33249_, _33247_);
  and (_33251_, _33250_, _33045_);
  or (_33252_, _33251_, _02177_);
  nor (_33253_, _10363_, _01632_);
  nand (_33254_, _10685_, _02177_);
  and (_33255_, _33254_, _33253_);
  and (_33256_, _33255_, _33252_);
  or (_33258_, _33072_, \oc8051_golden_model_1.PSW [7]);
  or (_33259_, _10030_, _06518_);
  and (_33260_, _33259_, _10363_);
  and (_33261_, _33260_, _33258_);
  or (_33262_, _33261_, _10368_);
  or (_33263_, _33262_, _33256_);
  or (_33264_, _33052_, _09861_);
  and (_33265_, _33264_, _09853_);
  and (_33266_, _33265_, _33263_);
  nor (_33267_, _10685_, _09853_);
  or (_33268_, _33267_, _02071_);
  or (_33269_, _33268_, _33266_);
  or (_33270_, _09969_, _04788_);
  and (_33271_, _33270_, _04793_);
  and (_33272_, _33271_, _33269_);
  and (_33273_, _10030_, _02173_);
  or (_33274_, _33273_, _33272_);
  and (_33275_, _33274_, _33044_);
  or (_33276_, _33072_, _06518_);
  or (_33277_, _10030_, \oc8051_golden_model_1.PSW [7]);
  and (_33279_, _33277_, _09848_);
  and (_33280_, _33279_, _33276_);
  or (_33281_, _33280_, _10385_);
  or (_33282_, _33281_, _33275_);
  or (_33283_, _33052_, _09846_);
  and (_33284_, _33283_, _07145_);
  and (_33285_, _33284_, _33282_);
  nor (_33286_, _10685_, _07145_);
  or (_33287_, _33286_, _07175_);
  or (_33288_, _33287_, _33285_);
  nand (_33290_, _33053_, _07175_);
  and (_33291_, _33290_, _09305_);
  and (_33292_, _33291_, _33288_);
  and (_33293_, _03028_, _02185_);
  or (_33294_, _33293_, _01636_);
  or (_33295_, _33294_, _33292_);
  and (_33296_, _33295_, _10403_);
  or (_33297_, _33056_, _10408_);
  or (_33298_, _09969_, _08439_);
  and (_33299_, _33298_, _02083_);
  and (_33301_, _33299_, _33297_);
  or (_33302_, _33301_, _10407_);
  or (_33303_, _33302_, _33296_);
  or (_33304_, _33052_, _09844_);
  and (_33305_, _33304_, _07254_);
  and (_33306_, _33305_, _33303_);
  nor (_33307_, _10685_, _07254_);
  or (_33308_, _33307_, _07304_);
  or (_33309_, _33308_, _33306_);
  nand (_33310_, _33053_, _07304_);
  and (_33312_, _33310_, _01889_);
  and (_33313_, _33312_, _33309_);
  and (_33314_, _03028_, _01888_);
  or (_33315_, _33314_, _01653_);
  or (_33316_, _33315_, _33313_);
  and (_33317_, _33316_, _02202_);
  or (_33318_, _09969_, _10408_);
  or (_33319_, _33056_, _08439_);
  and (_33320_, _33319_, _33318_);
  and (_33321_, _33320_, _02082_);
  or (_33323_, _33321_, _10435_);
  or (_33324_, _33323_, _33317_);
  nand (_33325_, _33053_, _10435_);
  and (_33326_, _33325_, _02303_);
  and (_33327_, _33326_, _33324_);
  nand (_33328_, _10030_, _02201_);
  nand (_33329_, _33328_, _10442_);
  or (_33330_, _33329_, _33327_);
  or (_33331_, _33052_, _10442_);
  and (_33332_, _33331_, _05195_);
  and (_33334_, _33332_, _33330_);
  or (_33335_, _33334_, _33043_);
  nor (_33336_, _01860_, _01642_);
  and (_33337_, _33336_, _33335_);
  and (_33338_, _33320_, _01860_);
  or (_33339_, _33338_, _10458_);
  or (_33340_, _33339_, _33337_);
  nand (_33341_, _33053_, _10458_);
  and (_33342_, _33341_, _01538_);
  and (_33343_, _33342_, _33340_);
  nand (_33345_, _10030_, _01537_);
  nand (_33346_, _33345_, _10465_);
  or (_33347_, _33346_, _33343_);
  or (_33348_, _33052_, _10465_);
  and (_33349_, _33348_, _10470_);
  and (_33350_, _33349_, _33347_);
  or (_33351_, _33350_, _33042_);
  and (_33352_, _33351_, _22954_);
  and (_33353_, _33052_, _09829_);
  or (_33354_, _33353_, _38088_);
  or (_33356_, _33354_, _33352_);
  and (_40367_, _33356_, _33041_);
  or (_33357_, _38087_, \oc8051_golden_model_1.PC [9]);
  and (_33358_, _33357_, _37580_);
  nor (_33359_, _10470_, _01822_);
  nor (_33360_, _05195_, _01822_);
  not (_33361_, \oc8051_golden_model_1.PC [9]);
  and (_33362_, _04270_, _09830_);
  and (_33363_, _33362_, \oc8051_golden_model_1.PC [8]);
  nor (_33364_, _33363_, _33361_);
  and (_33366_, _33363_, _33361_);
  or (_33367_, _33366_, _33364_);
  or (_33368_, _33367_, _09844_);
  or (_33369_, _33367_, _09846_);
  and (_33370_, _09912_, _02071_);
  or (_33371_, _33367_, _09861_);
  and (_33372_, _09912_, _02072_);
  not (_33373_, _33367_);
  nand (_33374_, _33373_, _09863_);
  and (_33375_, _09912_, _02079_);
  or (_33377_, _33367_, _10327_);
  or (_33378_, _10026_, _04757_);
  and (_33379_, _10026_, _01959_);
  nand (_33380_, _33373_, _10219_);
  or (_33381_, _33367_, _10207_);
  nand (_33382_, _33373_, _08628_);
  nand (_33383_, _33373_, _06629_);
  and (_33384_, _10026_, _02817_);
  nor (_33385_, _02817_, _33361_);
  and (_33386_, _33385_, _21690_);
  or (_33388_, _33386_, _10125_);
  and (_33389_, _33388_, _06618_);
  or (_33390_, _33389_, _33384_);
  and (_33391_, _33390_, _33383_);
  and (_33392_, _10026_, _02003_);
  nor (_33393_, _33373_, _21690_);
  or (_33394_, _33393_, _33392_);
  or (_33395_, _33394_, _33391_);
  and (_33396_, _33395_, _10136_);
  nand (_33397_, _33367_, _06616_);
  nand (_33399_, _33397_, _21702_);
  or (_33400_, _33399_, _33396_);
  and (_33401_, _10107_, _10026_);
  or (_33402_, _10028_, _10027_);
  nand (_33403_, _33402_, _10080_);
  or (_33404_, _33402_, _10080_);
  and (_33405_, _33404_, _33403_);
  and (_33406_, _33405_, _10105_);
  or (_33407_, _33406_, _33401_);
  or (_33408_, _33407_, _04381_);
  and (_33410_, _33408_, _33400_);
  or (_33411_, _33410_, _01883_);
  nand (_33412_, _33373_, _01883_);
  and (_33413_, _33412_, _02814_);
  and (_33414_, _33413_, _33411_);
  not (_33415_, _09970_);
  and (_33416_, _09973_, _33415_);
  and (_33417_, _33416_, _09916_);
  nor (_33418_, _33416_, _09916_);
  or (_33419_, _33418_, _33417_);
  or (_33421_, _33419_, _09996_);
  or (_33422_, _09876_, _09912_);
  and (_33423_, _33422_, _02001_);
  and (_33424_, _33423_, _33421_);
  or (_33425_, _33424_, _30311_);
  or (_33426_, _33425_, _33414_);
  or (_33427_, _33367_, _09871_);
  and (_33428_, _33427_, _02024_);
  and (_33429_, _33428_, _33426_);
  and (_33430_, _10026_, _02007_);
  or (_33432_, _33430_, _03279_);
  or (_33433_, _33432_, _33429_);
  and (_33434_, _33433_, _02840_);
  nand (_33435_, _10026_, _01999_);
  nand (_33436_, _33435_, _10156_);
  or (_33437_, _33436_, _33434_);
  or (_33438_, _33367_, _10156_);
  and (_33439_, _33438_, _02021_);
  and (_33440_, _33439_, _33437_);
  nand (_33441_, _10026_, _02006_);
  nand (_33443_, _33441_, _10163_);
  or (_33444_, _33443_, _33440_);
  or (_33445_, _33367_, _10163_);
  and (_33446_, _33445_, _02025_);
  and (_33447_, _33446_, _33444_);
  and (_33448_, _10026_, _01997_);
  or (_33449_, _33448_, _10167_);
  or (_33450_, _33449_, _33447_);
  and (_33451_, _33450_, _01880_);
  nand (_33452_, _10026_, _01878_);
  nand (_33454_, _33452_, _08538_);
  or (_33455_, _33454_, _33451_);
  or (_33456_, _33419_, _08572_);
  nand (_33457_, _09913_, _08572_);
  and (_33458_, _33457_, _33456_);
  or (_33459_, _33458_, _08538_);
  and (_33460_, _33459_, _33455_);
  or (_33461_, _33460_, _08493_);
  nand (_33462_, _09913_, _08498_);
  or (_33463_, _33419_, _08498_);
  and (_33465_, _33463_, _33462_);
  or (_33466_, _33465_, _08494_);
  and (_33467_, _33466_, _33461_);
  or (_33468_, _33467_, _01995_);
  and (_33469_, _09912_, _08625_);
  and (_33470_, _33419_, _30342_);
  or (_33471_, _33470_, _02444_);
  or (_33472_, _33471_, _33469_);
  and (_33473_, _33472_, _02046_);
  and (_33474_, _33473_, _33468_);
  or (_33476_, _33419_, _08664_);
  nand (_33477_, _09913_, _08664_);
  and (_33478_, _33477_, _02045_);
  and (_33479_, _33478_, _33476_);
  or (_33480_, _33479_, _08628_);
  or (_33481_, _33480_, _33474_);
  and (_33482_, _33481_, _33382_);
  or (_33483_, _33482_, _01991_);
  or (_33484_, _10026_, _02861_);
  nor (_33485_, _02871_, _30628_);
  and (_33487_, _33485_, _21871_);
  and (_33488_, _33487_, _30627_);
  and (_33489_, _33488_, _33484_);
  and (_33490_, _33489_, _33483_);
  and (_33491_, _30633_, _10026_);
  or (_33492_, _33491_, _10211_);
  or (_33493_, _33492_, _33490_);
  and (_33494_, _33493_, _33381_);
  or (_33495_, _33494_, _01967_);
  or (_33496_, _10026_, _08249_);
  and (_33498_, _33496_, _10214_);
  and (_33499_, _33498_, _33495_);
  and (_33500_, _10026_, _01966_);
  or (_33501_, _33500_, _10219_);
  or (_33502_, _33501_, _33499_);
  and (_33503_, _33502_, _33380_);
  or (_33504_, _33503_, _06776_);
  or (_33505_, _10026_, _06775_);
  and (_33506_, _33505_, _01550_);
  and (_33507_, _33506_, _33504_);
  and (_33509_, _33367_, _01549_);
  or (_33510_, _33509_, _01875_);
  or (_33511_, _33510_, _33507_);
  or (_33512_, _10026_, _02408_);
  and (_33513_, _33512_, _22053_);
  and (_33514_, _33513_, _33511_);
  nand (_33515_, _09912_, _02080_);
  nand (_33516_, _33515_, _09211_);
  or (_33517_, _33516_, _33514_);
  or (_33518_, _10026_, _09211_);
  and (_33520_, _33518_, _02043_);
  and (_33521_, _33520_, _33517_);
  nand (_33522_, _09912_, _01602_);
  nand (_33523_, _33522_, _10245_);
  or (_33524_, _33523_, _33521_);
  or (_33525_, _33367_, _10245_);
  and (_33526_, _33525_, _30680_);
  and (_33527_, _33526_, _33524_);
  or (_33528_, _33527_, _33379_);
  and (_33529_, _33528_, _33047_);
  and (_33531_, _33405_, _10253_);
  or (_33532_, _33531_, _04758_);
  or (_33533_, _33532_, _33529_);
  and (_33534_, _33533_, _33378_);
  or (_33535_, _33534_, _01869_);
  nand (_33536_, _09913_, _01869_);
  and (_33537_, _33536_, _06985_);
  and (_33538_, _33537_, _33535_);
  and (_33539_, _10026_, _06984_);
  or (_33540_, _33539_, _10267_);
  or (_33541_, _33540_, _33538_);
  nor (_33542_, _10295_, \oc8051_golden_model_1.DPH [1]);
  nor (_33543_, _33542_, _10296_);
  or (_33544_, _33543_, _10268_);
  and (_33545_, _33544_, _02576_);
  and (_33546_, _33545_, _33541_);
  and (_33547_, _10026_, _01958_);
  or (_33548_, _33547_, _01638_);
  or (_33549_, _33548_, _33546_);
  and (_33550_, _33549_, _10311_);
  or (_33552_, _33405_, _07356_);
  or (_33553_, _10026_, _10316_);
  and (_33554_, _33553_, _10310_);
  and (_33555_, _33554_, _33552_);
  or (_33556_, _33555_, _10331_);
  or (_33557_, _33556_, _33550_);
  and (_33558_, _33557_, _33377_);
  or (_33559_, _33558_, _10330_);
  or (_33560_, _10026_, _10329_);
  and (_33561_, _33560_, _02166_);
  and (_33563_, _33561_, _33559_);
  or (_33564_, _33563_, _33375_);
  and (_33565_, _33564_, _02912_);
  and (_33566_, _10026_, _02167_);
  or (_33567_, _33566_, _01645_);
  or (_33568_, _33567_, _33565_);
  and (_33569_, _33568_, _10344_);
  or (_33570_, _33405_, _10316_);
  or (_33571_, _10026_, _07356_);
  and (_33572_, _33571_, _10343_);
  and (_33574_, _33572_, _33570_);
  or (_33575_, _33574_, _09863_);
  or (_33576_, _33575_, _33569_);
  and (_33577_, _33576_, _33374_);
  or (_33578_, _33577_, _07042_);
  or (_33579_, _10026_, _07041_);
  and (_33580_, _33579_, _02176_);
  and (_33581_, _33580_, _33578_);
  or (_33582_, _33581_, _33372_);
  and (_33583_, _33582_, _02907_);
  and (_33585_, _10026_, _02177_);
  or (_33586_, _33585_, _01632_);
  or (_33587_, _33586_, _33583_);
  and (_33588_, _33587_, _10364_);
  or (_33589_, _33405_, \oc8051_golden_model_1.PSW [7]);
  or (_33590_, _10026_, _06518_);
  and (_33591_, _33590_, _10363_);
  and (_33592_, _33591_, _33589_);
  or (_33593_, _33592_, _10368_);
  or (_33594_, _33593_, _33588_);
  and (_33596_, _33594_, _33371_);
  or (_33597_, _33596_, _09854_);
  or (_33598_, _10026_, _09853_);
  and (_33599_, _33598_, _04788_);
  and (_33600_, _33599_, _33597_);
  or (_33601_, _33600_, _33370_);
  and (_33602_, _33601_, _04793_);
  and (_33603_, _10026_, _02173_);
  or (_33604_, _33603_, _01648_);
  or (_33605_, _33604_, _33602_);
  and (_33607_, _33605_, _09849_);
  or (_33608_, _33405_, _06518_);
  or (_33609_, _10026_, \oc8051_golden_model_1.PSW [7]);
  and (_33610_, _33609_, _09848_);
  and (_33611_, _33610_, _33608_);
  or (_33612_, _33611_, _10385_);
  or (_33613_, _33612_, _33607_);
  and (_33614_, _33613_, _33369_);
  or (_33615_, _33614_, _07146_);
  or (_33616_, _10026_, _07145_);
  and (_33618_, _33616_, _07176_);
  and (_33619_, _33618_, _33615_);
  and (_33620_, _33367_, _07175_);
  or (_33621_, _33620_, _02185_);
  or (_33622_, _33621_, _33619_);
  nor (_33623_, _02083_, _01636_);
  nand (_33624_, _02811_, _02185_);
  and (_33625_, _33624_, _33623_);
  and (_33626_, _33625_, _33622_);
  or (_33627_, _33419_, _10408_);
  or (_33629_, _09912_, _08439_);
  and (_33630_, _33629_, _02083_);
  and (_33631_, _33630_, _33627_);
  or (_33632_, _33631_, _10407_);
  or (_33633_, _33632_, _33626_);
  and (_33634_, _33633_, _33368_);
  or (_33635_, _33634_, _07255_);
  or (_33636_, _10026_, _07254_);
  and (_33637_, _33636_, _07305_);
  and (_33638_, _33637_, _33635_);
  and (_33640_, _33367_, _07304_);
  or (_33641_, _33640_, _01888_);
  or (_33642_, _33641_, _33638_);
  nand (_33643_, _02811_, _01888_);
  and (_33644_, _33643_, _22866_);
  and (_33645_, _33644_, _33642_);
  or (_33646_, _33419_, _08439_);
  nand (_33647_, _09913_, _08439_);
  and (_33648_, _33647_, _33646_);
  and (_33649_, _33648_, _02082_);
  or (_33651_, _33649_, _10435_);
  or (_33652_, _33651_, _33645_);
  nand (_33653_, _33373_, _10435_);
  and (_33654_, _33653_, _02303_);
  and (_33655_, _33654_, _33652_);
  nand (_33656_, _10026_, _02201_);
  nand (_33657_, _33656_, _10442_);
  or (_33658_, _33657_, _33655_);
  or (_33659_, _33367_, _10442_);
  and (_33660_, _33659_, _05195_);
  and (_33662_, _33660_, _33658_);
  or (_33663_, _33662_, _33360_);
  and (_33664_, _33663_, _33336_);
  and (_33665_, _33648_, _01860_);
  or (_33666_, _33665_, _10458_);
  or (_33667_, _33666_, _33664_);
  nand (_33668_, _33373_, _10458_);
  and (_33669_, _33668_, _01538_);
  and (_33670_, _33669_, _33667_);
  nand (_33671_, _10026_, _01537_);
  nand (_33673_, _33671_, _10465_);
  or (_33674_, _33673_, _33670_);
  or (_33675_, _33367_, _10465_);
  and (_33676_, _33675_, _10470_);
  and (_33677_, _33676_, _33674_);
  or (_33678_, _33677_, _33359_);
  and (_33679_, _33678_, _22954_);
  and (_33680_, _33367_, _09829_);
  or (_33681_, _33680_, _38088_);
  or (_33682_, _33681_, _33679_);
  and (_40368_, _33682_, _33358_);
  nor (_33684_, _09835_, \oc8051_golden_model_1.PC [10]);
  nor (_33685_, _33684_, _09836_);
  not (_33686_, _33685_);
  nand (_33687_, _33686_, _10458_);
  nand (_33688_, _33686_, _10435_);
  nand (_33689_, _33686_, _07175_);
  or (_33690_, _09906_, _04788_);
  or (_33691_, _09906_, _02176_);
  or (_33692_, _09906_, _02166_);
  nor (_33694_, _33686_, _10163_);
  or (_33695_, _33685_, _10156_);
  nor (_33696_, _33686_, _10150_);
  or (_33697_, _09976_, _09974_);
  and (_33698_, _33697_, _09909_);
  nor (_33699_, _33697_, _09909_);
  nor (_33700_, _33699_, _33698_);
  or (_33701_, _33700_, _09996_);
  or (_33702_, _09876_, _09906_);
  and (_33703_, _33702_, _02001_);
  and (_33704_, _33703_, _33701_);
  and (_33705_, _10107_, _10021_);
  or (_33706_, _10082_, _10024_);
  and (_33707_, _33706_, _10083_);
  and (_33708_, _33707_, _10105_);
  or (_33709_, _33708_, _04381_);
  or (_33710_, _33709_, _33705_);
  or (_33711_, _10112_, \oc8051_golden_model_1.PC [10]);
  nand (_33712_, _33686_, _10112_);
  and (_33713_, _33712_, _33711_);
  or (_33715_, _33713_, _02817_);
  nand (_33716_, _11080_, _02817_);
  and (_33717_, _33716_, _10121_);
  and (_33718_, _33717_, _33715_);
  and (_33719_, _33685_, _06625_);
  or (_33720_, _33719_, _02823_);
  or (_33721_, _33720_, _06629_);
  or (_33722_, _33721_, _33718_);
  nand (_33723_, _33686_, _06629_);
  and (_33724_, _33723_, _33722_);
  or (_33726_, _33724_, _02003_);
  nand (_33727_, _11080_, _02003_);
  and (_33728_, _33727_, _10136_);
  and (_33729_, _33728_, _33726_);
  nand (_33730_, _33685_, _06616_);
  nand (_33731_, _33730_, _21702_);
  or (_33732_, _33731_, _33729_);
  and (_33733_, _33732_, _10144_);
  and (_33734_, _33733_, _33710_);
  or (_33735_, _33734_, _33704_);
  and (_33737_, _33735_, _09871_);
  or (_33738_, _33737_, _33696_);
  and (_33739_, _33738_, _02008_);
  nor (_33740_, _11080_, _02008_);
  nor (_33741_, _33740_, _03279_);
  nand (_33742_, _33741_, _10156_);
  or (_33743_, _33742_, _33739_);
  and (_33744_, _33743_, _33695_);
  or (_33745_, _33744_, _02006_);
  nand (_33746_, _11080_, _02006_);
  and (_33748_, _33746_, _10163_);
  and (_33749_, _33748_, _33745_);
  or (_33750_, _33749_, _33694_);
  and (_33751_, _33750_, _02025_);
  and (_33752_, _10021_, _01997_);
  or (_33753_, _33752_, _10167_);
  or (_33754_, _33753_, _33751_);
  and (_33755_, _33754_, _01880_);
  nand (_33756_, _10021_, _01878_);
  nand (_33757_, _33756_, _08538_);
  or (_33759_, _33757_, _33755_);
  and (_33760_, _09906_, _08572_);
  and (_33761_, _33700_, _08573_);
  or (_33762_, _33761_, _33760_);
  or (_33763_, _33762_, _08538_);
  and (_33764_, _33763_, _33759_);
  or (_33765_, _33764_, _08493_);
  and (_33766_, _33700_, _30279_);
  and (_33767_, _09906_, _08498_);
  or (_33768_, _33767_, _08494_);
  or (_33770_, _33768_, _33766_);
  and (_33771_, _33770_, _33765_);
  or (_33772_, _33771_, _01995_);
  and (_33773_, _09906_, _08625_);
  and (_33774_, _33700_, _30342_);
  or (_33775_, _33774_, _02444_);
  or (_33776_, _33775_, _33773_);
  and (_33777_, _33776_, _02046_);
  and (_33778_, _33777_, _33772_);
  or (_33779_, _33700_, _08664_);
  or (_33781_, _09906_, _31735_);
  and (_33782_, _33781_, _02045_);
  and (_33783_, _33782_, _33779_);
  or (_33784_, _33783_, _08628_);
  or (_33785_, _33784_, _33778_);
  nand (_33786_, _33686_, _08628_);
  and (_33787_, _30632_, _02861_);
  and (_33788_, _33787_, _33786_);
  and (_33789_, _33788_, _33785_);
  nor (_33790_, _33787_, _11080_);
  nand (_33792_, _10207_, _01565_);
  or (_33793_, _33792_, _33790_);
  or (_33794_, _33793_, _33789_);
  or (_33795_, _33685_, _10207_);
  and (_33796_, _33795_, _08249_);
  and (_33797_, _33796_, _33794_);
  or (_33798_, _33797_, _10213_);
  and (_33799_, _33798_, _08248_);
  nor (_33800_, _11080_, _01968_);
  or (_33801_, _33800_, _10219_);
  or (_33803_, _33801_, _33799_);
  nand (_33804_, _33686_, _10219_);
  and (_33805_, _33804_, _06775_);
  and (_33806_, _33805_, _33803_);
  nor (_33807_, _11080_, _06775_);
  or (_33808_, _33807_, _01549_);
  or (_33809_, _33808_, _33806_);
  nand (_33810_, _33686_, _01549_);
  and (_33811_, _33810_, _02408_);
  and (_33812_, _33811_, _33809_);
  nand (_33814_, _10021_, _01875_);
  nand (_33815_, _33814_, _22053_);
  or (_33816_, _33815_, _33812_);
  or (_33817_, _09906_, _07401_);
  and (_33818_, _33817_, _09211_);
  and (_33819_, _33818_, _33816_);
  nor (_33820_, _11080_, _09211_);
  or (_33821_, _33820_, _01602_);
  or (_33822_, _33821_, _33819_);
  or (_33823_, _09906_, _02043_);
  and (_33825_, _33823_, _10245_);
  and (_33826_, _33825_, _33822_);
  nor (_33827_, _33686_, _10245_);
  or (_33828_, _33827_, _33826_);
  and (_33829_, _33828_, _30680_);
  nand (_33830_, _10021_, _01959_);
  nand (_33831_, _33830_, _33047_);
  or (_33832_, _33831_, _33829_);
  or (_33833_, _33707_, _10254_);
  and (_33834_, _33833_, _04757_);
  and (_33835_, _33834_, _33832_);
  nor (_33836_, _11080_, _04757_);
  or (_33837_, _33836_, _01869_);
  or (_33838_, _33837_, _33835_);
  or (_33839_, _09906_, _01870_);
  and (_33840_, _33839_, _06985_);
  and (_33841_, _33840_, _33838_);
  and (_33842_, _10021_, _06984_);
  or (_33843_, _33842_, _10267_);
  or (_33844_, _33843_, _33841_);
  nor (_33846_, _10296_, \oc8051_golden_model_1.DPH [2]);
  nor (_33847_, _33846_, _10297_);
  or (_33848_, _33847_, _10268_);
  and (_33849_, _33848_, _33844_);
  or (_33850_, _33849_, _01958_);
  nor (_33851_, _10310_, _01638_);
  nand (_33852_, _11080_, _01958_);
  and (_33853_, _33852_, _33851_);
  and (_33854_, _33853_, _33850_);
  or (_33855_, _33707_, _07356_);
  or (_33857_, _10021_, _10316_);
  and (_33858_, _33857_, _10310_);
  and (_33859_, _33858_, _33855_);
  or (_33860_, _33859_, _10331_);
  or (_33861_, _33860_, _33854_);
  or (_33862_, _33685_, _10327_);
  and (_33863_, _33862_, _10329_);
  and (_33864_, _33863_, _33861_);
  nor (_33865_, _11080_, _10329_);
  or (_33866_, _33865_, _02079_);
  or (_33868_, _33866_, _33864_);
  and (_33869_, _33868_, _33692_);
  or (_33870_, _33869_, _02167_);
  nand (_33871_, _11080_, _02167_);
  and (_33872_, _33871_, _22337_);
  and (_33873_, _33872_, _33870_);
  or (_33874_, _33707_, _10316_);
  or (_33875_, _10021_, _07356_);
  and (_33876_, _33875_, _10343_);
  and (_33877_, _33876_, _33874_);
  or (_33879_, _33877_, _09863_);
  or (_33880_, _33879_, _33873_);
  nand (_33881_, _33686_, _09863_);
  and (_33882_, _33881_, _07041_);
  and (_33883_, _33882_, _33880_);
  nor (_33884_, _11080_, _07041_);
  or (_33885_, _33884_, _02072_);
  or (_33886_, _33885_, _33883_);
  and (_33887_, _33886_, _33691_);
  or (_33888_, _33887_, _02177_);
  nand (_33890_, _11080_, _02177_);
  and (_33891_, _33890_, _33253_);
  and (_33892_, _33891_, _33888_);
  or (_33893_, _33707_, \oc8051_golden_model_1.PSW [7]);
  or (_33894_, _10021_, _06518_);
  and (_33895_, _33894_, _10363_);
  and (_33896_, _33895_, _33893_);
  or (_33897_, _33896_, _10368_);
  or (_33898_, _33897_, _33892_);
  or (_33899_, _33685_, _09861_);
  and (_33901_, _33899_, _09853_);
  and (_33902_, _33901_, _33898_);
  nor (_33903_, _11080_, _09853_);
  or (_33904_, _33903_, _02071_);
  or (_33905_, _33904_, _33902_);
  and (_33906_, _33905_, _33690_);
  or (_33907_, _33906_, _02173_);
  nand (_33908_, _11080_, _02173_);
  and (_33909_, _33908_, _33044_);
  and (_33910_, _33909_, _33907_);
  or (_33912_, _33707_, _06518_);
  or (_33913_, _10021_, \oc8051_golden_model_1.PSW [7]);
  and (_33914_, _33913_, _09848_);
  and (_33915_, _33914_, _33912_);
  or (_33916_, _33915_, _10385_);
  or (_33917_, _33916_, _33910_);
  or (_33918_, _33685_, _09846_);
  and (_33919_, _33918_, _07145_);
  and (_33920_, _33919_, _33917_);
  nor (_33921_, _11080_, _07145_);
  or (_33923_, _33921_, _07175_);
  or (_33924_, _33923_, _33920_);
  and (_33925_, _33924_, _33689_);
  or (_33926_, _33925_, _02185_);
  nand (_33927_, _03455_, _02185_);
  and (_33928_, _33927_, _33623_);
  and (_33929_, _33928_, _33926_);
  or (_33930_, _33700_, _10408_);
  or (_33931_, _09906_, _08439_);
  and (_33932_, _33931_, _02083_);
  and (_33934_, _33932_, _33930_);
  or (_33935_, _33934_, _10407_);
  or (_33936_, _33935_, _33929_);
  or (_33937_, _33685_, _09844_);
  and (_33938_, _33937_, _07254_);
  and (_33939_, _33938_, _33936_);
  nor (_33940_, _11080_, _07254_);
  or (_33941_, _33940_, _07304_);
  or (_33942_, _33941_, _33939_);
  nand (_33943_, _33686_, _07304_);
  and (_33945_, _33943_, _33942_);
  or (_33946_, _33945_, _01888_);
  nand (_33947_, _03455_, _01888_);
  and (_33948_, _33947_, _22866_);
  and (_33949_, _33948_, _33946_);
  or (_33950_, _09906_, _10408_);
  or (_33951_, _33700_, _08439_);
  and (_33952_, _33951_, _33950_);
  and (_33953_, _33952_, _02082_);
  or (_33954_, _33953_, _10435_);
  or (_33955_, _33954_, _33949_);
  and (_33956_, _33955_, _33688_);
  or (_33957_, _33956_, _02201_);
  nand (_33958_, _11080_, _02201_);
  and (_33959_, _33958_, _10442_);
  and (_33960_, _33959_, _33957_);
  nor (_33961_, _33686_, _10442_);
  or (_33962_, _33961_, _02058_);
  or (_33963_, _33962_, _33960_);
  nand (_33964_, _02294_, _02058_);
  and (_33966_, _33964_, _33336_);
  and (_33967_, _33966_, _33963_);
  and (_33968_, _33952_, _01860_);
  or (_33969_, _33968_, _10458_);
  or (_33970_, _33969_, _33967_);
  and (_33971_, _33970_, _33687_);
  or (_33972_, _33971_, _01537_);
  nand (_33973_, _11080_, _01537_);
  and (_33974_, _33973_, _10465_);
  and (_33975_, _33974_, _33972_);
  nor (_33977_, _33686_, _10465_);
  or (_33978_, _33977_, _02057_);
  or (_33979_, _33978_, _33975_);
  nand (_33980_, _02294_, _02057_);
  and (_33981_, _33980_, _22954_);
  and (_33982_, _33981_, _33979_);
  and (_33983_, _33685_, _09829_);
  or (_33984_, _33983_, _38088_);
  or (_33985_, _33984_, _33982_);
  or (_33986_, _38087_, \oc8051_golden_model_1.PC [10]);
  and (_33988_, _33986_, _37580_);
  and (_40369_, _33988_, _33985_);
  nor (_33989_, _38087_, _09897_);
  and (_33990_, _32681_, _05197_);
  nor (_33991_, _33990_, _09897_);
  and (_33992_, _33990_, _09897_);
  or (_33993_, _33992_, _33991_);
  or (_33994_, _33993_, _09844_);
  or (_33995_, _33993_, _09846_);
  or (_33996_, _33993_, _09861_);
  not (_33998_, _33993_);
  nand (_33999_, _33998_, _09863_);
  or (_34000_, _10018_, _10019_);
  nand (_34001_, _34000_, _10084_);
  or (_34002_, _34000_, _10084_);
  and (_34003_, _34002_, _34001_);
  or (_34004_, _34003_, _07356_);
  or (_34005_, _10017_, _10316_);
  and (_34006_, _34005_, _10310_);
  and (_34007_, _34006_, _34004_);
  or (_34009_, _10017_, _04757_);
  or (_34010_, _33993_, _10245_);
  and (_34011_, _10017_, _02006_);
  or (_34012_, _09869_, _10017_);
  or (_34013_, _09876_, _09900_);
  nor (_34014_, _33698_, _09907_);
  and (_34015_, _34014_, _09904_);
  nor (_34016_, _34014_, _09904_);
  or (_34017_, _34016_, _34015_);
  or (_34018_, _34017_, _09996_);
  and (_34020_, _34018_, _02001_);
  and (_34021_, _34020_, _34013_);
  and (_34022_, _10107_, _10017_);
  and (_34023_, _34003_, _10105_);
  or (_34024_, _34023_, _04381_);
  or (_34025_, _34024_, _34022_);
  or (_34026_, _33993_, _30926_);
  nand (_34027_, _11281_, _02817_);
  or (_34028_, _02817_, \oc8051_golden_model_1.PC [11]);
  or (_34029_, _34028_, _10112_);
  and (_34031_, _34029_, _34027_);
  or (_34032_, _34031_, _30932_);
  nor (_34033_, _10017_, _01562_);
  nor (_34034_, _34033_, _02003_);
  and (_34035_, _34034_, _34032_);
  and (_34036_, _34035_, _34026_);
  and (_34037_, _10017_, _02003_);
  or (_34038_, _34037_, _06616_);
  or (_34039_, _34038_, _34036_);
  nand (_34040_, _33998_, _06616_);
  and (_34041_, _34040_, _01568_);
  and (_34042_, _34041_, _34039_);
  nor (_34043_, _11281_, _01568_);
  or (_34044_, _34043_, _04380_);
  or (_34045_, _34044_, _34042_);
  and (_34046_, _34045_, _10144_);
  and (_34047_, _34046_, _34025_);
  or (_34048_, _34047_, _34021_);
  and (_34049_, _34048_, _09871_);
  nor (_34050_, _33998_, _10150_);
  or (_34052_, _34050_, _10149_);
  or (_34053_, _34052_, _34049_);
  and (_34054_, _34053_, _34012_);
  or (_34055_, _34054_, _10157_);
  or (_34056_, _33993_, _10156_);
  and (_34057_, _34056_, _02021_);
  and (_34058_, _34057_, _34055_);
  or (_34059_, _34058_, _34011_);
  and (_34060_, _34059_, _10163_);
  or (_34061_, _33998_, _10163_);
  nand (_34063_, _34061_, _10169_);
  or (_34064_, _34063_, _34060_);
  or (_34065_, _10169_, _10017_);
  and (_34066_, _34065_, _34064_);
  or (_34067_, _34066_, _08539_);
  or (_34068_, _34017_, _08572_);
  nand (_34069_, _09901_, _08572_);
  and (_34070_, _34069_, _34068_);
  or (_34071_, _34070_, _08538_);
  and (_34072_, _34071_, _34067_);
  or (_34074_, _34072_, _08493_);
  nand (_34075_, _09901_, _08498_);
  or (_34076_, _34017_, _08498_);
  and (_34077_, _34076_, _34075_);
  or (_34078_, _34077_, _08494_);
  and (_34079_, _34078_, _34074_);
  and (_34080_, _34079_, _08441_);
  or (_34081_, _34017_, _08664_);
  nand (_34082_, _09901_, _08664_);
  and (_34083_, _34082_, _02045_);
  and (_34085_, _34083_, _34081_);
  nand (_34086_, _09901_, _08625_);
  or (_34087_, _34017_, _08625_);
  and (_34088_, _34087_, _01995_);
  and (_34089_, _34088_, _34086_);
  or (_34090_, _34089_, _34085_);
  or (_34091_, _34090_, _34080_);
  and (_34092_, _34091_, _09867_);
  nand (_34093_, _33993_, _08628_);
  nand (_34094_, _34093_, _10201_);
  or (_34096_, _34094_, _34092_);
  or (_34097_, _10201_, _10017_);
  and (_34098_, _34097_, _10207_);
  and (_34099_, _34098_, _34096_);
  nor (_34100_, _33998_, _10207_);
  or (_34101_, _34100_, _10216_);
  or (_34102_, _34101_, _34099_);
  or (_34103_, _10215_, _10017_);
  and (_34104_, _34103_, _10220_);
  and (_34105_, _34104_, _34102_);
  and (_34107_, _33993_, _10219_);
  or (_34108_, _34107_, _06776_);
  or (_34109_, _34108_, _34105_);
  or (_34110_, _10017_, _06775_);
  and (_34111_, _34110_, _01550_);
  and (_34112_, _34111_, _34109_);
  nand (_34113_, _33993_, _01549_);
  nand (_34114_, _34113_, _10231_);
  or (_34115_, _34114_, _34112_);
  or (_34116_, _10231_, _10017_);
  and (_34118_, _34116_, _07401_);
  and (_34119_, _34118_, _34115_);
  nand (_34120_, _09900_, _02080_);
  nand (_34121_, _34120_, _09211_);
  or (_34122_, _34121_, _34119_);
  or (_34123_, _10017_, _09211_);
  and (_34124_, _34123_, _02043_);
  and (_34125_, _34124_, _34122_);
  nand (_34126_, _09900_, _01602_);
  nand (_34127_, _34126_, _10245_);
  or (_34129_, _34127_, _34125_);
  and (_34130_, _34129_, _34010_);
  or (_34131_, _34130_, _10248_);
  or (_34132_, _10247_, _10017_);
  and (_34133_, _34132_, _10254_);
  and (_34134_, _34133_, _34131_);
  and (_34135_, _34003_, _10253_);
  or (_34136_, _34135_, _04758_);
  or (_34137_, _34136_, _34134_);
  and (_34138_, _34137_, _34009_);
  or (_34140_, _34138_, _01869_);
  nand (_34141_, _09901_, _01869_);
  and (_34142_, _34141_, _06985_);
  and (_34143_, _34142_, _34140_);
  and (_34144_, _10017_, _06984_);
  or (_34145_, _34144_, _34143_);
  and (_34146_, _34145_, _10268_);
  nor (_34147_, _10297_, \oc8051_golden_model_1.DPH [3]);
  nor (_34148_, _34147_, _10298_);
  and (_34149_, _34148_, _10267_);
  or (_34150_, _34149_, _10307_);
  or (_34151_, _34150_, _34146_);
  or (_34152_, _10306_, _10017_);
  and (_34153_, _34152_, _10311_);
  and (_34154_, _34153_, _34151_);
  or (_34155_, _34154_, _34007_);
  and (_34156_, _34155_, _10327_);
  nor (_34157_, _33998_, _10327_);
  or (_34158_, _34157_, _10330_);
  or (_34159_, _34158_, _34156_);
  or (_34161_, _10017_, _10329_);
  and (_34162_, _34161_, _02166_);
  and (_34163_, _34162_, _34159_);
  nand (_34164_, _09900_, _02079_);
  nand (_34165_, _34164_, _10339_);
  or (_34166_, _34165_, _34163_);
  or (_34167_, _10339_, _10017_);
  and (_34168_, _34167_, _10344_);
  and (_34169_, _34168_, _34166_);
  or (_34170_, _34003_, _10316_);
  or (_34172_, _10017_, _07356_);
  and (_34173_, _34172_, _10343_);
  and (_34174_, _34173_, _34170_);
  or (_34175_, _34174_, _09863_);
  or (_34176_, _34175_, _34169_);
  and (_34177_, _34176_, _33999_);
  or (_34178_, _34177_, _07042_);
  or (_34179_, _10017_, _07041_);
  and (_34180_, _34179_, _02176_);
  and (_34181_, _34180_, _34178_);
  nand (_34183_, _09900_, _02072_);
  nand (_34184_, _34183_, _09292_);
  or (_34185_, _34184_, _34181_);
  nor (_34186_, _10363_, _11281_);
  or (_34187_, _34186_, _22459_);
  and (_34188_, _34187_, _34185_);
  or (_34189_, _34003_, \oc8051_golden_model_1.PSW [7]);
  or (_34190_, _10017_, _06518_);
  and (_34191_, _34190_, _10363_);
  and (_34192_, _34191_, _34189_);
  or (_34194_, _34192_, _10368_);
  or (_34195_, _34194_, _34188_);
  and (_34196_, _34195_, _33996_);
  or (_34197_, _34196_, _09854_);
  or (_34198_, _10017_, _09853_);
  and (_34199_, _34198_, _04788_);
  and (_34200_, _34199_, _34197_);
  nand (_34201_, _09900_, _02071_);
  nand (_34202_, _34201_, _09850_);
  or (_34203_, _34202_, _34200_);
  nor (_34205_, _11281_, _09848_);
  or (_34206_, _34205_, _22602_);
  and (_34207_, _34206_, _34203_);
  or (_34208_, _34003_, _06518_);
  or (_34209_, _10017_, \oc8051_golden_model_1.PSW [7]);
  and (_34210_, _34209_, _09848_);
  and (_34211_, _34210_, _34208_);
  or (_34212_, _34211_, _10385_);
  or (_34213_, _34212_, _34207_);
  and (_34214_, _34213_, _33995_);
  or (_34216_, _34214_, _07146_);
  or (_34217_, _10017_, _07145_);
  and (_34218_, _34217_, _07176_);
  and (_34219_, _34218_, _34216_);
  and (_34220_, _33993_, _07175_);
  or (_34221_, _34220_, _02185_);
  or (_34222_, _34221_, _34219_);
  nand (_34223_, _03268_, _02185_);
  and (_34224_, _34223_, _34222_);
  or (_34225_, _34224_, _01636_);
  nand (_34227_, _11281_, _01636_);
  and (_34228_, _34227_, _10403_);
  and (_34229_, _34228_, _34225_);
  or (_34230_, _34017_, _10408_);
  or (_34231_, _09900_, _08439_);
  and (_34232_, _34231_, _02083_);
  and (_34233_, _34232_, _34230_);
  or (_34234_, _34233_, _10407_);
  or (_34235_, _34234_, _34229_);
  and (_34236_, _34235_, _33994_);
  or (_34238_, _34236_, _07255_);
  or (_34239_, _10017_, _07254_);
  and (_34240_, _34239_, _07305_);
  and (_34241_, _34240_, _34238_);
  and (_34242_, _33993_, _07304_);
  or (_34243_, _34242_, _01888_);
  or (_34244_, _34243_, _34241_);
  nand (_34245_, _03268_, _01888_);
  and (_34246_, _34245_, _34244_);
  or (_34247_, _34246_, _01653_);
  nand (_34249_, _11281_, _01653_);
  and (_34250_, _34249_, _02202_);
  and (_34251_, _34250_, _34247_);
  or (_34252_, _34017_, _08439_);
  nand (_34253_, _09901_, _08439_);
  and (_34254_, _34253_, _34252_);
  and (_34255_, _34254_, _02082_);
  or (_34256_, _34255_, _10435_);
  or (_34257_, _34256_, _34251_);
  nand (_34258_, _33998_, _10435_);
  and (_34260_, _34258_, _02303_);
  and (_34261_, _34260_, _34257_);
  nand (_34262_, _10017_, _02201_);
  nand (_34263_, _34262_, _10442_);
  or (_34264_, _34263_, _34261_);
  or (_34265_, _33993_, _10442_);
  and (_34266_, _34265_, _05195_);
  and (_34267_, _34266_, _34264_);
  nor (_34268_, _05195_, _01954_);
  or (_34269_, _34268_, _01642_);
  or (_34271_, _34269_, _34267_);
  nand (_34272_, _11281_, _01642_);
  and (_34273_, _34272_, _01887_);
  and (_34274_, _34273_, _34271_);
  and (_34275_, _34254_, _01860_);
  or (_34276_, _34275_, _10458_);
  or (_34277_, _34276_, _34274_);
  nand (_34278_, _33998_, _10458_);
  and (_34279_, _34278_, _01538_);
  and (_34280_, _34279_, _34277_);
  nand (_34282_, _10017_, _01537_);
  nand (_34283_, _34282_, _10465_);
  or (_34284_, _34283_, _34280_);
  or (_34285_, _33993_, _10465_);
  and (_34286_, _34285_, _10470_);
  and (_34287_, _34286_, _34284_);
  nor (_34288_, _10470_, _01954_);
  or (_34289_, _34288_, _01651_);
  or (_34290_, _34289_, _34287_);
  nand (_34291_, _11281_, _01651_);
  and (_34293_, _34291_, _34290_);
  or (_34294_, _34293_, _09829_);
  nand (_34295_, _33998_, _09829_);
  and (_34296_, _34295_, _38087_);
  and (_34297_, _34296_, _34294_);
  or (_34298_, _34297_, _33989_);
  and (_40370_, _34298_, _37580_);
  or (_34299_, _38087_, \oc8051_golden_model_1.PC [12]);
  and (_34300_, _34299_, _37580_);
  and (_34301_, _33990_, \oc8051_golden_model_1.PC [11]);
  and (_34303_, _34301_, \oc8051_golden_model_1.PC [12]);
  nor (_34304_, _34301_, \oc8051_golden_model_1.PC [12]);
  nor (_34305_, _34304_, _34303_);
  not (_34306_, _34305_);
  nand (_34307_, _34306_, _07304_);
  and (_34308_, _10013_, _10380_);
  and (_34309_, _10013_, _10359_);
  and (_34310_, _10340_, _10013_);
  and (_34311_, _10307_, _10013_);
  or (_34312_, _10088_, _10086_);
  and (_34314_, _34312_, _10089_);
  and (_34315_, _34314_, _10253_);
  and (_34316_, _34305_, _10219_);
  or (_34317_, _09982_, _09980_);
  and (_34318_, _34317_, _09983_);
  or (_34319_, _34318_, _08498_);
  or (_34320_, _09895_, _30279_);
  and (_34321_, _34320_, _34319_);
  or (_34322_, _34321_, _08494_);
  or (_34323_, _34305_, _10150_);
  nand (_34325_, _34306_, _06629_);
  or (_34326_, _34305_, _21690_);
  nor (_34327_, _02817_, \oc8051_golden_model_1.PC [12]);
  nand (_34328_, _34327_, _21690_);
  or (_34329_, _34328_, _30289_);
  and (_34330_, _34329_, _34326_);
  or (_34331_, _34330_, _02823_);
  and (_34332_, _34331_, _34325_);
  or (_34333_, _34332_, _02003_);
  nand (_34334_, _34306_, _06616_);
  and (_34336_, _34334_, _34333_);
  or (_34337_, _34336_, _10140_);
  and (_34338_, _09224_, _06618_);
  and (_34339_, _34338_, _01568_);
  or (_34340_, _34339_, _10013_);
  and (_34341_, _34340_, _34337_);
  or (_34342_, _34341_, _04380_);
  and (_34343_, _34314_, _10105_);
  and (_34344_, _10107_, _10013_);
  or (_34345_, _34344_, _04381_);
  or (_34347_, _34345_, _34343_);
  and (_34348_, _34347_, _34342_);
  or (_34349_, _34348_, _32358_);
  and (_34350_, _34318_, _09876_);
  and (_34351_, _09996_, _09895_);
  or (_34352_, _34351_, _02814_);
  or (_34353_, _34352_, _34350_);
  and (_34354_, _34353_, _34349_);
  or (_34355_, _34354_, _30311_);
  and (_34356_, _34355_, _34323_);
  or (_34358_, _34356_, _10149_);
  or (_34359_, _09869_, _10013_);
  and (_34360_, _34359_, _10156_);
  and (_34361_, _34360_, _34358_);
  nor (_34362_, _34306_, _10156_);
  or (_34363_, _34362_, _02006_);
  or (_34364_, _34363_, _34361_);
  not (_34365_, _10013_);
  nand (_34366_, _34365_, _02006_);
  and (_34367_, _34366_, _10163_);
  and (_34369_, _34367_, _34364_);
  or (_34370_, _34306_, _10163_);
  nand (_34371_, _34370_, _10169_);
  or (_34372_, _34371_, _34369_);
  or (_34373_, _10169_, _10013_);
  and (_34374_, _34373_, _08538_);
  and (_34375_, _34374_, _34372_);
  and (_34376_, _09895_, _08572_);
  and (_34377_, _34318_, _08573_);
  or (_34378_, _34377_, _34376_);
  and (_34379_, _34378_, _08539_);
  or (_34380_, _34379_, _08493_);
  or (_34381_, _34380_, _34375_);
  and (_34382_, _34381_, _08441_);
  and (_34383_, _34382_, _34322_);
  or (_34384_, _09895_, _30342_);
  or (_34385_, _34318_, _08625_);
  and (_34386_, _34385_, _01995_);
  and (_34387_, _34386_, _34384_);
  or (_34388_, _34318_, _08664_);
  or (_34390_, _09895_, _31735_);
  and (_34391_, _34390_, _02045_);
  and (_34392_, _34391_, _34388_);
  or (_34393_, _34392_, _08628_);
  or (_34394_, _34393_, _34387_);
  or (_34395_, _34394_, _34383_);
  nand (_34396_, _34306_, _08628_);
  and (_34397_, _34396_, _10201_);
  and (_34398_, _34397_, _34395_);
  nor (_34399_, _10201_, _34365_);
  or (_34401_, _34399_, _10211_);
  or (_34402_, _34401_, _34398_);
  or (_34403_, _34305_, _10207_);
  and (_34404_, _34403_, _34402_);
  or (_34405_, _34404_, _10216_);
  or (_34406_, _10215_, _10013_);
  and (_34407_, _34406_, _10220_);
  and (_34408_, _34407_, _34405_);
  or (_34409_, _34408_, _34316_);
  and (_34410_, _34409_, _06775_);
  nor (_34412_, _34365_, _06775_);
  or (_34413_, _34412_, _01549_);
  or (_34414_, _34413_, _34410_);
  nand (_34415_, _34306_, _01549_);
  and (_34416_, _34415_, _10231_);
  and (_34417_, _34416_, _34414_);
  nor (_34418_, _10231_, _34365_);
  or (_34419_, _34418_, _02080_);
  or (_34420_, _34419_, _34417_);
  or (_34421_, _09895_, _07401_);
  and (_34423_, _34421_, _09211_);
  and (_34424_, _34423_, _34420_);
  nor (_34425_, _34365_, _09211_);
  or (_34426_, _34425_, _01602_);
  or (_34427_, _34426_, _34424_);
  or (_34428_, _09895_, _02043_);
  and (_34429_, _34428_, _10245_);
  and (_34430_, _34429_, _34427_);
  nor (_34431_, _34306_, _10245_);
  or (_34432_, _34431_, _10248_);
  or (_34434_, _34432_, _34430_);
  or (_34435_, _10247_, _10013_);
  and (_34436_, _34435_, _10254_);
  and (_34437_, _34436_, _34434_);
  or (_34438_, _34437_, _34315_);
  and (_34439_, _34438_, _04757_);
  nor (_34440_, _34365_, _04757_);
  or (_34441_, _34440_, _01869_);
  or (_34442_, _34441_, _34439_);
  or (_34443_, _09895_, _01870_);
  and (_34444_, _34443_, _06985_);
  and (_34445_, _34444_, _34442_);
  and (_34446_, _10013_, _06984_);
  or (_34447_, _34446_, _10267_);
  or (_34448_, _34447_, _34445_);
  nor (_34449_, _10298_, \oc8051_golden_model_1.DPH [4]);
  nor (_34450_, _34449_, _10299_);
  or (_34451_, _34450_, _10268_);
  and (_34452_, _34451_, _10306_);
  and (_34453_, _34452_, _34448_);
  or (_34455_, _34453_, _34311_);
  and (_34456_, _34455_, _10311_);
  or (_34457_, _34314_, _07356_);
  or (_34458_, _10013_, _10316_);
  and (_34459_, _34458_, _10310_);
  and (_34460_, _34459_, _34457_);
  or (_34461_, _34460_, _10331_);
  or (_34462_, _34461_, _34456_);
  or (_34463_, _34305_, _10327_);
  and (_34464_, _34463_, _10329_);
  and (_34466_, _34464_, _34462_);
  nor (_34467_, _34365_, _10329_);
  or (_34468_, _34467_, _02079_);
  or (_34469_, _34468_, _34466_);
  or (_34470_, _09895_, _02166_);
  and (_34471_, _34470_, _10339_);
  and (_34472_, _34471_, _34469_);
  or (_34473_, _34472_, _34310_);
  and (_34474_, _34473_, _10344_);
  or (_34475_, _34314_, _10316_);
  or (_34477_, _10013_, _07356_);
  and (_34478_, _34477_, _10343_);
  and (_34479_, _34478_, _34475_);
  or (_34480_, _34479_, _09863_);
  or (_34481_, _34480_, _34474_);
  nand (_34482_, _34306_, _09863_);
  and (_34483_, _34482_, _07041_);
  and (_34484_, _34483_, _34481_);
  nor (_34485_, _34365_, _07041_);
  or (_34486_, _34485_, _02072_);
  or (_34488_, _34486_, _34484_);
  or (_34489_, _09895_, _02176_);
  and (_34490_, _34489_, _09292_);
  and (_34491_, _34490_, _34488_);
  or (_34492_, _34491_, _34309_);
  and (_34493_, _34492_, _10364_);
  or (_34494_, _34314_, \oc8051_golden_model_1.PSW [7]);
  or (_34495_, _10013_, _06518_);
  and (_34496_, _34495_, _10363_);
  and (_34497_, _34496_, _34494_);
  or (_34499_, _34497_, _10368_);
  or (_34500_, _34499_, _34493_);
  or (_34501_, _34305_, _09861_);
  and (_34502_, _34501_, _09853_);
  and (_34503_, _34502_, _34500_);
  nor (_34504_, _34365_, _09853_);
  or (_34505_, _34504_, _02071_);
  or (_34506_, _34505_, _34503_);
  or (_34507_, _09895_, _04788_);
  and (_34508_, _34507_, _09850_);
  and (_34509_, _34508_, _34506_);
  or (_34510_, _34509_, _34308_);
  and (_34511_, _34510_, _09849_);
  or (_34512_, _34314_, _06518_);
  or (_34513_, _10013_, \oc8051_golden_model_1.PSW [7]);
  and (_34514_, _34513_, _09848_);
  and (_34515_, _34514_, _34512_);
  or (_34516_, _34515_, _10385_);
  or (_34517_, _34516_, _34511_);
  or (_34518_, _34305_, _09846_);
  and (_34519_, _34518_, _07145_);
  and (_34520_, _34519_, _34517_);
  nor (_34521_, _34365_, _07145_);
  or (_34522_, _34521_, _07175_);
  or (_34523_, _34522_, _34520_);
  nand (_34524_, _34306_, _07175_);
  and (_34525_, _34524_, _09305_);
  and (_34526_, _34525_, _34523_);
  nor (_34527_, _04211_, _09305_);
  or (_34528_, _34527_, _01636_);
  or (_34530_, _34528_, _34526_);
  nand (_34531_, _34365_, _01636_);
  and (_34532_, _34531_, _10403_);
  and (_34533_, _34532_, _34530_);
  or (_34534_, _34318_, _10408_);
  or (_34535_, _09895_, _08439_);
  and (_34536_, _34535_, _02083_);
  and (_34537_, _34536_, _34534_);
  or (_34538_, _34537_, _10407_);
  or (_34539_, _34538_, _34533_);
  or (_34541_, _34305_, _09844_);
  and (_34542_, _34541_, _07254_);
  and (_34543_, _34542_, _34539_);
  nor (_34544_, _34365_, _07254_);
  or (_34545_, _34544_, _07304_);
  or (_34546_, _34545_, _34543_);
  and (_34547_, _34546_, _34307_);
  or (_34548_, _34547_, _01888_);
  nand (_34549_, _04211_, _01888_);
  and (_34550_, _34549_, _10426_);
  and (_34552_, _34550_, _34548_);
  and (_34553_, _10013_, _01653_);
  or (_34554_, _34553_, _02082_);
  or (_34555_, _34554_, _34552_);
  or (_34556_, _09895_, _10408_);
  or (_34557_, _34318_, _08439_);
  and (_34558_, _34557_, _34556_);
  or (_34559_, _34558_, _02202_);
  and (_34560_, _34559_, _34555_);
  or (_34561_, _34560_, _10435_);
  nand (_34562_, _34306_, _10435_);
  and (_34563_, _34562_, _34561_);
  or (_34564_, _34563_, _02201_);
  nand (_34565_, _34365_, _02201_);
  and (_34566_, _34565_, _10442_);
  and (_34567_, _34566_, _34564_);
  nor (_34568_, _34306_, _10442_);
  or (_34569_, _34568_, _02058_);
  or (_34570_, _34569_, _34567_);
  nand (_34571_, _02058_, _01855_);
  and (_34573_, _34571_, _10453_);
  and (_34574_, _34573_, _34570_);
  and (_34575_, _10013_, _01642_);
  or (_34576_, _34575_, _01860_);
  or (_34577_, _34576_, _34574_);
  or (_34578_, _34558_, _01887_);
  and (_34579_, _34578_, _10461_);
  and (_34580_, _34579_, _34577_);
  and (_34581_, _34305_, _10458_);
  or (_34582_, _34581_, _01537_);
  or (_34584_, _34582_, _34580_);
  nand (_34585_, _34365_, _01537_);
  and (_34586_, _34585_, _10465_);
  and (_34587_, _34586_, _34584_);
  nor (_34588_, _34306_, _10465_);
  or (_34589_, _34588_, _02057_);
  or (_34590_, _34589_, _34587_);
  nand (_34591_, _02057_, _01855_);
  and (_34592_, _34591_, _34590_);
  or (_34593_, _34592_, _01651_);
  nand (_34594_, _34365_, _01651_);
  and (_34595_, _34594_, _10481_);
  and (_34596_, _34595_, _34593_);
  and (_34597_, _34305_, _09829_);
  or (_34598_, _34597_, _38088_);
  or (_34599_, _34598_, _34596_);
  and (_40371_, _34599_, _34300_);
  nor (_34600_, _38087_, _09883_);
  nand (_34601_, _03916_, _01888_);
  and (_34602_, _33362_, _09885_);
  and (_34604_, _34602_, \oc8051_golden_model_1.PC [12]);
  nor (_34605_, _34604_, _09883_);
  and (_34606_, _34604_, _09883_);
  or (_34607_, _34606_, _34605_);
  or (_34608_, _34607_, _09844_);
  or (_34609_, _34607_, _09846_);
  or (_34610_, _34607_, _09861_);
  or (_34611_, _10011_, _10010_);
  nand (_34612_, _34611_, _10090_);
  or (_34613_, _34611_, _10090_);
  and (_34614_, _34613_, _34612_);
  or (_34615_, _34614_, _10316_);
  or (_34616_, _10009_, _07356_);
  and (_34617_, _34616_, _10343_);
  and (_34618_, _34617_, _34615_);
  or (_34619_, _10009_, _04757_);
  or (_34620_, _34607_, _10245_);
  nand (_34621_, _09891_, _08498_);
  or (_34622_, _09893_, _09892_);
  nand (_34623_, _34622_, _09984_);
  or (_34625_, _34622_, _09984_);
  and (_34626_, _34625_, _34623_);
  or (_34627_, _34626_, _08498_);
  and (_34628_, _34627_, _34621_);
  or (_34629_, _34628_, _08494_);
  and (_34630_, _10009_, _02006_);
  or (_34631_, _09869_, _10009_);
  or (_34632_, _09876_, _09890_);
  or (_34633_, _34626_, _09996_);
  and (_34634_, _34633_, _02001_);
  and (_34636_, _34634_, _34632_);
  and (_34637_, _10107_, _10009_);
  and (_34638_, _34614_, _10105_);
  or (_34639_, _34638_, _04381_);
  or (_34640_, _34639_, _34637_);
  not (_34641_, _34607_);
  nand (_34642_, _34641_, _06616_);
  nand (_34643_, _34641_, _06629_);
  or (_34644_, _34607_, _21690_);
  nor (_34645_, _02817_, \oc8051_golden_model_1.PC [13]);
  nand (_34647_, _34645_, _21690_);
  or (_34648_, _34647_, _30289_);
  and (_34649_, _34648_, _34644_);
  or (_34650_, _34649_, _02823_);
  and (_34651_, _34650_, _34643_);
  or (_34652_, _34651_, _02003_);
  nand (_34653_, _34652_, _34642_);
  and (_34654_, _34653_, _01568_);
  nor (_34655_, _34339_, _10009_);
  or (_34656_, _34655_, _34654_);
  nand (_34658_, _34656_, _04381_);
  and (_34659_, _34658_, _10144_);
  and (_34660_, _34659_, _34640_);
  or (_34661_, _34660_, _34636_);
  and (_34662_, _34661_, _09871_);
  nor (_34663_, _34641_, _10150_);
  or (_34664_, _34663_, _10149_);
  or (_34665_, _34664_, _34662_);
  and (_34666_, _34665_, _34631_);
  or (_34667_, _34666_, _10157_);
  or (_34669_, _34607_, _10156_);
  and (_34670_, _34669_, _02021_);
  and (_34671_, _34670_, _34667_);
  or (_34672_, _34671_, _34630_);
  and (_34673_, _34672_, _10163_);
  or (_34674_, _34641_, _10163_);
  nand (_34675_, _34674_, _10169_);
  or (_34676_, _34675_, _34673_);
  or (_34677_, _10169_, _10009_);
  and (_34678_, _34677_, _08538_);
  and (_34680_, _34678_, _34676_);
  nand (_34681_, _09891_, _08572_);
  or (_34682_, _34626_, _08572_);
  and (_34683_, _34682_, _08539_);
  and (_34684_, _34683_, _34681_);
  or (_34685_, _34684_, _08493_);
  or (_34686_, _34685_, _34680_);
  and (_34687_, _34686_, _34629_);
  or (_34688_, _34687_, _01995_);
  and (_34689_, _09890_, _08625_);
  and (_34691_, _34626_, _30342_);
  or (_34692_, _34691_, _02444_);
  or (_34693_, _34692_, _34689_);
  and (_34694_, _34693_, _02046_);
  and (_34695_, _34694_, _34688_);
  or (_34696_, _34626_, _08664_);
  nand (_34697_, _09891_, _08664_);
  and (_34698_, _34697_, _02045_);
  and (_34699_, _34698_, _34696_);
  or (_34700_, _34699_, _34695_);
  and (_34702_, _34700_, _09867_);
  nand (_34703_, _34607_, _08628_);
  nand (_34704_, _34703_, _10201_);
  or (_34705_, _34704_, _34702_);
  or (_34706_, _10201_, _10009_);
  and (_34707_, _34706_, _10207_);
  and (_34708_, _34707_, _34705_);
  nor (_34709_, _34641_, _10207_);
  or (_34710_, _34709_, _10216_);
  or (_34711_, _34710_, _34708_);
  or (_34713_, _10215_, _10009_);
  and (_34714_, _34713_, _10220_);
  and (_34715_, _34714_, _34711_);
  and (_34716_, _34607_, _10219_);
  or (_34717_, _34716_, _06776_);
  or (_34718_, _34717_, _34715_);
  or (_34719_, _10009_, _06775_);
  and (_34720_, _34719_, _01550_);
  and (_34721_, _34720_, _34718_);
  nand (_34722_, _34607_, _01549_);
  nand (_34724_, _34722_, _10231_);
  or (_34725_, _34724_, _34721_);
  or (_34726_, _10231_, _10009_);
  and (_34727_, _34726_, _07401_);
  and (_34728_, _34727_, _34725_);
  nand (_34729_, _09890_, _02080_);
  nand (_34730_, _34729_, _09211_);
  or (_34731_, _34730_, _34728_);
  or (_34732_, _10009_, _09211_);
  and (_34733_, _34732_, _02043_);
  and (_34735_, _34733_, _34731_);
  nand (_34736_, _09890_, _01602_);
  nand (_34737_, _34736_, _10245_);
  or (_34738_, _34737_, _34735_);
  and (_34739_, _34738_, _34620_);
  or (_34740_, _34739_, _10248_);
  or (_34741_, _10247_, _10009_);
  and (_34742_, _34741_, _10254_);
  and (_34743_, _34742_, _34740_);
  and (_34744_, _34614_, _10253_);
  or (_34746_, _34744_, _04758_);
  or (_34747_, _34746_, _34743_);
  and (_34748_, _34747_, _34619_);
  or (_34749_, _34748_, _01869_);
  nand (_34750_, _09891_, _01869_);
  and (_34751_, _34750_, _06985_);
  and (_34752_, _34751_, _34749_);
  and (_34753_, _10009_, _06984_);
  or (_34754_, _34753_, _34752_);
  and (_34755_, _34754_, _10268_);
  or (_34757_, _10299_, \oc8051_golden_model_1.DPH [5]);
  and (_34758_, _34757_, _10300_);
  and (_34759_, _34758_, _10267_);
  or (_34760_, _34759_, _10307_);
  or (_34761_, _34760_, _34755_);
  or (_34762_, _10306_, _10009_);
  and (_34763_, _34762_, _10311_);
  and (_34764_, _34763_, _34761_);
  or (_34765_, _34614_, _07356_);
  or (_34766_, _10009_, _10316_);
  and (_34768_, _34766_, _10310_);
  and (_34769_, _34768_, _34765_);
  or (_34770_, _34769_, _34764_);
  and (_34771_, _34770_, _10327_);
  nor (_34772_, _34641_, _10327_);
  or (_34773_, _34772_, _10330_);
  or (_34774_, _34773_, _34771_);
  or (_34775_, _10009_, _10329_);
  and (_34776_, _34775_, _02166_);
  and (_34777_, _34776_, _34774_);
  nand (_34779_, _09890_, _02079_);
  nand (_34780_, _34779_, _10339_);
  or (_34781_, _34780_, _34777_);
  or (_34782_, _10339_, _10009_);
  and (_34783_, _34782_, _10344_);
  and (_34784_, _34783_, _34781_);
  or (_34785_, _34784_, _34618_);
  and (_34786_, _34785_, _09864_);
  and (_34787_, _34607_, _09863_);
  or (_34788_, _34787_, _07042_);
  or (_34790_, _34788_, _34786_);
  or (_34791_, _10009_, _07041_);
  and (_34792_, _34791_, _02176_);
  and (_34793_, _34792_, _34790_);
  nand (_34794_, _09890_, _02072_);
  nand (_34795_, _34794_, _09292_);
  or (_34796_, _34795_, _34793_);
  nor (_34797_, _10363_, _11694_);
  or (_34798_, _34797_, _22459_);
  and (_34799_, _34798_, _34796_);
  or (_34800_, _34614_, \oc8051_golden_model_1.PSW [7]);
  or (_34801_, _10009_, _06518_);
  and (_34802_, _34801_, _10363_);
  and (_34803_, _34802_, _34800_);
  or (_34804_, _34803_, _10368_);
  or (_34805_, _34804_, _34799_);
  and (_34806_, _34805_, _34610_);
  or (_34807_, _34806_, _09854_);
  or (_34808_, _10009_, _09853_);
  and (_34809_, _34808_, _04788_);
  and (_34811_, _34809_, _34807_);
  nand (_34812_, _09890_, _02071_);
  nand (_34813_, _34812_, _09850_);
  or (_34814_, _34813_, _34811_);
  nor (_34815_, _11694_, _09848_);
  or (_34816_, _34815_, _22602_);
  and (_34817_, _34816_, _34814_);
  or (_34818_, _34614_, _06518_);
  or (_34819_, _10009_, \oc8051_golden_model_1.PSW [7]);
  and (_34820_, _34819_, _09848_);
  and (_34822_, _34820_, _34818_);
  or (_34823_, _34822_, _10385_);
  or (_34824_, _34823_, _34817_);
  and (_34825_, _34824_, _34609_);
  or (_34826_, _34825_, _07146_);
  or (_34827_, _10009_, _07145_);
  and (_34828_, _34827_, _07176_);
  and (_34829_, _34828_, _34826_);
  and (_34830_, _34607_, _07175_);
  or (_34831_, _34830_, _02185_);
  or (_34833_, _34831_, _34829_);
  nand (_34834_, _03916_, _02185_);
  and (_34835_, _34834_, _34833_);
  or (_34836_, _34835_, _01636_);
  nand (_34837_, _11694_, _01636_);
  and (_34838_, _34837_, _10403_);
  and (_34839_, _34838_, _34836_);
  or (_34840_, _34626_, _10408_);
  or (_34841_, _09890_, _08439_);
  and (_34842_, _34841_, _02083_);
  and (_34844_, _34842_, _34840_);
  or (_34845_, _34844_, _10407_);
  or (_34846_, _34845_, _34839_);
  and (_34847_, _34846_, _34608_);
  or (_34848_, _34847_, _07255_);
  or (_34849_, _10009_, _07254_);
  and (_34850_, _34849_, _07305_);
  and (_34851_, _34850_, _34848_);
  and (_34852_, _34607_, _07304_);
  or (_34853_, _34852_, _01888_);
  or (_34855_, _34853_, _34851_);
  and (_34856_, _34855_, _34601_);
  or (_34857_, _34856_, _01653_);
  nand (_34858_, _11694_, _01653_);
  and (_34859_, _34858_, _02202_);
  and (_34860_, _34859_, _34857_);
  or (_34861_, _34626_, _08439_);
  nand (_34862_, _09891_, _08439_);
  and (_34863_, _34862_, _34861_);
  and (_34864_, _34863_, _02082_);
  or (_34866_, _34864_, _10435_);
  or (_34867_, _34866_, _34860_);
  nand (_34868_, _34641_, _10435_);
  and (_34869_, _34868_, _02303_);
  and (_34870_, _34869_, _34867_);
  nand (_34871_, _10009_, _02201_);
  nand (_34872_, _34871_, _10442_);
  or (_34873_, _34872_, _34870_);
  or (_34874_, _34607_, _10442_);
  and (_34875_, _34874_, _05195_);
  and (_34877_, _34875_, _34873_);
  nor (_34878_, _02252_, _05195_);
  or (_34879_, _34878_, _01642_);
  or (_34880_, _34879_, _34877_);
  nand (_34881_, _11694_, _01642_);
  and (_34882_, _34881_, _01887_);
  and (_34883_, _34882_, _34880_);
  and (_34884_, _34863_, _01860_);
  or (_34885_, _34884_, _10458_);
  or (_34886_, _34885_, _34883_);
  nand (_34888_, _34641_, _10458_);
  and (_34889_, _34888_, _01538_);
  and (_34890_, _34889_, _34886_);
  nand (_34891_, _10009_, _01537_);
  nand (_34892_, _34891_, _10465_);
  or (_34893_, _34892_, _34890_);
  or (_34894_, _34607_, _10465_);
  and (_34895_, _34894_, _10470_);
  and (_34896_, _34895_, _34893_);
  nor (_34897_, _02252_, _10470_);
  or (_34899_, _34897_, _01651_);
  or (_34900_, _34899_, _34896_);
  nand (_34901_, _11694_, _01651_);
  and (_34902_, _34901_, _34900_);
  or (_34903_, _34902_, _09829_);
  nand (_34904_, _34641_, _09829_);
  and (_34905_, _34904_, _38087_);
  and (_34906_, _34905_, _34903_);
  or (_34907_, _34906_, _34600_);
  and (_40372_, _34907_, _37580_);
  or (_34909_, _38087_, \oc8051_golden_model_1.PC [14]);
  and (_34910_, _34909_, _37580_);
  nor (_34911_, _09839_, \oc8051_golden_model_1.PC [14]);
  nor (_34912_, _34911_, _09840_);
  or (_34913_, _34912_, _07305_);
  nor (_34914_, _11895_, _09850_);
  nor (_34915_, _11895_, _09292_);
  nor (_34916_, _10339_, _11895_);
  nor (_34917_, _10306_, _11895_);
  and (_34918_, _34912_, _10219_);
  or (_34919_, _34912_, _10207_);
  or (_34920_, _09986_, _09882_);
  and (_34921_, _34920_, _09987_);
  and (_34922_, _34921_, _30279_);
  and (_34923_, _09879_, _08498_);
  or (_34924_, _34923_, _34922_);
  and (_34925_, _34924_, _08493_);
  and (_34926_, _34912_, _10165_);
  or (_34927_, _34912_, _10156_);
  and (_34928_, _34921_, _09876_);
  and (_34930_, _09996_, _09879_);
  or (_34931_, _34930_, _02814_);
  or (_34932_, _34931_, _34928_);
  or (_34933_, _10092_, _10004_);
  and (_34934_, _34933_, _10093_);
  and (_34935_, _34934_, _10105_);
  and (_34936_, _10107_, _10001_);
  or (_34937_, _34936_, _04381_);
  or (_34938_, _34937_, _34935_);
  and (_34939_, _34912_, _06616_);
  and (_34940_, _34912_, _06625_);
  and (_34941_, _34912_, _10112_);
  and (_34942_, _10136_, \oc8051_golden_model_1.PC [14]);
  and (_34943_, _34942_, _10129_);
  and (_34944_, _34943_, _21690_);
  or (_34945_, _34944_, _34941_);
  and (_34946_, _34945_, _02818_);
  or (_34947_, _34946_, _34940_);
  and (_34948_, _34947_, _01562_);
  and (_34949_, _34912_, _06629_);
  or (_34951_, _34949_, _34948_);
  and (_34952_, _34951_, _06618_);
  or (_34953_, _34952_, _34939_);
  and (_34954_, _34953_, _01568_);
  nor (_34955_, _34339_, _11895_);
  or (_34956_, _34955_, _04380_);
  or (_34957_, _34956_, _34954_);
  and (_34958_, _34957_, _04394_);
  and (_34959_, _34958_, _34938_);
  and (_34960_, _34912_, _01883_);
  or (_34961_, _34960_, _02001_);
  or (_34962_, _34961_, _34959_);
  and (_34963_, _34962_, _34932_);
  or (_34964_, _34963_, _30311_);
  or (_34965_, _34912_, _09871_);
  and (_34966_, _34965_, _09869_);
  and (_34967_, _34966_, _34964_);
  or (_34968_, _09869_, _11895_);
  nand (_34969_, _34968_, _10156_);
  or (_34970_, _34969_, _34967_);
  and (_34972_, _34970_, _34927_);
  or (_34973_, _34972_, _02006_);
  nand (_34974_, _11895_, _02006_);
  and (_34975_, _34974_, _10163_);
  and (_34976_, _34975_, _34973_);
  or (_34977_, _34976_, _34926_);
  and (_34978_, _34977_, _10169_);
  or (_34979_, _10169_, _11895_);
  nand (_34980_, _34979_, _08538_);
  or (_34981_, _34980_, _34978_);
  and (_34983_, _09879_, _08572_);
  and (_34984_, _34921_, _08573_);
  or (_34985_, _34984_, _34983_);
  or (_34986_, _34985_, _08538_);
  and (_34987_, _34986_, _08494_);
  and (_34988_, _34987_, _34981_);
  or (_34989_, _34988_, _01995_);
  or (_34990_, _34989_, _34925_);
  and (_34991_, _34921_, _30342_);
  and (_34992_, _09879_, _08625_);
  or (_34994_, _34992_, _02444_);
  or (_34995_, _34994_, _34991_);
  and (_34996_, _34995_, _02046_);
  and (_34997_, _34996_, _34990_);
  or (_34998_, _34921_, _08664_);
  or (_34999_, _09879_, _31735_);
  and (_35000_, _34999_, _02045_);
  and (_35001_, _35000_, _34998_);
  or (_35002_, _35001_, _08628_);
  or (_35003_, _35002_, _34997_);
  or (_35005_, _34912_, _09867_);
  and (_35006_, _35005_, _10201_);
  and (_35007_, _35006_, _35003_);
  nor (_35008_, _10201_, _11895_);
  or (_35009_, _35008_, _10211_);
  or (_35010_, _35009_, _35007_);
  and (_35011_, _35010_, _34919_);
  or (_35012_, _35011_, _10216_);
  or (_35013_, _10215_, _10001_);
  and (_35014_, _35013_, _10220_);
  and (_35015_, _35014_, _35012_);
  or (_35016_, _35015_, _34918_);
  and (_35017_, _35016_, _06775_);
  nor (_35018_, _11895_, _06775_);
  or (_35019_, _35018_, _01549_);
  or (_35020_, _35019_, _35017_);
  or (_35021_, _34912_, _01550_);
  and (_35022_, _35021_, _10231_);
  and (_35023_, _35022_, _35020_);
  nor (_35024_, _10231_, _11895_);
  or (_35026_, _35024_, _02080_);
  or (_35027_, _35026_, _35023_);
  or (_35028_, _09879_, _07401_);
  and (_35029_, _35028_, _09211_);
  and (_35030_, _35029_, _35027_);
  nor (_35031_, _11895_, _09211_);
  or (_35032_, _35031_, _01602_);
  or (_35033_, _35032_, _35030_);
  or (_35034_, _09879_, _02043_);
  and (_35035_, _35034_, _10245_);
  and (_35037_, _35035_, _35033_);
  and (_35038_, _34912_, _10249_);
  or (_35039_, _35038_, _10248_);
  or (_35040_, _35039_, _35037_);
  or (_35041_, _10247_, _10001_);
  and (_35042_, _35041_, _10254_);
  and (_35043_, _35042_, _35040_);
  and (_35044_, _34934_, _10253_);
  or (_35045_, _35044_, _35043_);
  and (_35046_, _35045_, _04757_);
  nor (_35048_, _11895_, _04757_);
  or (_35049_, _35048_, _01869_);
  or (_35050_, _35049_, _35046_);
  or (_35051_, _09879_, _01870_);
  and (_35052_, _35051_, _06985_);
  and (_35053_, _35052_, _35050_);
  and (_35054_, _10001_, _06984_);
  or (_35055_, _35054_, _10267_);
  or (_35056_, _35055_, _35053_);
  and (_35057_, _10300_, _10272_);
  nor (_35059_, _35057_, _10301_);
  or (_35060_, _35059_, _10268_);
  and (_35061_, _35060_, _10306_);
  and (_35062_, _35061_, _35056_);
  or (_35063_, _35062_, _34917_);
  and (_35064_, _35063_, _10311_);
  or (_35065_, _34934_, _07356_);
  or (_35066_, _10001_, _10316_);
  and (_35067_, _35066_, _10310_);
  and (_35068_, _35067_, _35065_);
  or (_35070_, _35068_, _10331_);
  or (_35071_, _35070_, _35064_);
  or (_35072_, _34912_, _10327_);
  and (_35073_, _35072_, _10329_);
  and (_35074_, _35073_, _35071_);
  nor (_35075_, _11895_, _10329_);
  or (_35076_, _35075_, _02079_);
  or (_35077_, _35076_, _35074_);
  or (_35078_, _09879_, _02166_);
  and (_35079_, _35078_, _10339_);
  and (_35081_, _35079_, _35077_);
  or (_35082_, _35081_, _34916_);
  and (_35083_, _35082_, _10344_);
  or (_35084_, _34934_, _10316_);
  or (_35085_, _10001_, _07356_);
  and (_35086_, _35085_, _10343_);
  and (_35087_, _35086_, _35084_);
  or (_35088_, _35087_, _09863_);
  or (_35089_, _35088_, _35083_);
  or (_35090_, _34912_, _09864_);
  and (_35092_, _35090_, _07041_);
  and (_35093_, _35092_, _35089_);
  nor (_35094_, _11895_, _07041_);
  or (_35095_, _35094_, _02072_);
  or (_35096_, _35095_, _35093_);
  or (_35097_, _09879_, _02176_);
  and (_35098_, _35097_, _09292_);
  and (_35099_, _35098_, _35096_);
  or (_35100_, _35099_, _34915_);
  and (_35101_, _35100_, _10364_);
  or (_35103_, _34934_, \oc8051_golden_model_1.PSW [7]);
  or (_35104_, _10001_, _06518_);
  and (_35105_, _35104_, _10363_);
  and (_35106_, _35105_, _35103_);
  or (_35107_, _35106_, _10368_);
  or (_35108_, _35107_, _35101_);
  or (_35109_, _34912_, _09861_);
  and (_35110_, _35109_, _09853_);
  and (_35111_, _35110_, _35108_);
  nor (_35112_, _11895_, _09853_);
  or (_35114_, _35112_, _02071_);
  or (_35115_, _35114_, _35111_);
  or (_35116_, _09879_, _04788_);
  and (_35117_, _35116_, _09850_);
  and (_35118_, _35117_, _35115_);
  or (_35119_, _35118_, _34914_);
  and (_35120_, _35119_, _09849_);
  or (_35121_, _34934_, _06518_);
  or (_35122_, _10001_, \oc8051_golden_model_1.PSW [7]);
  and (_35123_, _35122_, _09848_);
  and (_35125_, _35123_, _35121_);
  or (_35126_, _35125_, _10385_);
  or (_35127_, _35126_, _35120_);
  or (_35128_, _34912_, _09846_);
  and (_35129_, _35128_, _07145_);
  and (_35130_, _35129_, _35127_);
  nor (_35131_, _11895_, _07145_);
  or (_35132_, _35131_, _07175_);
  or (_35133_, _35132_, _35130_);
  or (_35134_, _34912_, _07176_);
  and (_35136_, _35134_, _09305_);
  and (_35137_, _35136_, _35133_);
  nor (_35138_, _03808_, _09305_);
  or (_35139_, _35138_, _01636_);
  or (_35140_, _35139_, _35137_);
  nand (_35141_, _11895_, _01636_);
  and (_35142_, _35141_, _10403_);
  and (_35143_, _35142_, _35140_);
  or (_35144_, _34921_, _10408_);
  or (_35145_, _09879_, _08439_);
  and (_35147_, _35145_, _02083_);
  and (_35148_, _35147_, _35144_);
  or (_35149_, _35148_, _10407_);
  or (_35150_, _35149_, _35143_);
  or (_35151_, _34912_, _09844_);
  and (_35152_, _35151_, _07254_);
  and (_35153_, _35152_, _35150_);
  nor (_35154_, _11895_, _07254_);
  or (_35155_, _35154_, _07304_);
  or (_35156_, _35155_, _35153_);
  and (_35158_, _35156_, _34913_);
  or (_35159_, _35158_, _01888_);
  nand (_35160_, _03808_, _01888_);
  and (_35161_, _35160_, _10426_);
  and (_35162_, _35161_, _35159_);
  and (_35163_, _10001_, _01653_);
  or (_35164_, _35163_, _02082_);
  or (_35165_, _35164_, _35162_);
  or (_35166_, _09879_, _10408_);
  or (_35167_, _34921_, _08439_);
  and (_35169_, _35167_, _35166_);
  or (_35170_, _35169_, _02202_);
  and (_35171_, _35170_, _35165_);
  or (_35172_, _35171_, _10435_);
  or (_35173_, _34912_, _10438_);
  and (_35174_, _35173_, _35172_);
  or (_35175_, _35174_, _02201_);
  nand (_35176_, _11895_, _02201_);
  and (_35177_, _35176_, _10442_);
  and (_35178_, _35177_, _35175_);
  and (_35180_, _34912_, _10443_);
  or (_35181_, _35180_, _02058_);
  or (_35182_, _35181_, _35178_);
  nand (_35183_, _02058_, _01922_);
  and (_35184_, _35183_, _10453_);
  and (_35185_, _35184_, _35182_);
  and (_35186_, _10001_, _01642_);
  or (_35187_, _35186_, _01860_);
  or (_35188_, _35187_, _35185_);
  or (_35189_, _35169_, _01887_);
  and (_35191_, _35189_, _10461_);
  and (_35192_, _35191_, _35188_);
  and (_35193_, _34912_, _10458_);
  or (_35194_, _35193_, _01537_);
  or (_35195_, _35194_, _35192_);
  nand (_35196_, _11895_, _01537_);
  and (_35197_, _35196_, _10465_);
  and (_35198_, _35197_, _35195_);
  and (_35199_, _34912_, _10466_);
  or (_35200_, _35199_, _02057_);
  or (_35202_, _35200_, _35198_);
  nand (_35203_, _02057_, _01922_);
  and (_35204_, _35203_, _35202_);
  or (_35205_, _35204_, _01651_);
  nand (_35206_, _11895_, _01651_);
  and (_35207_, _35206_, _10481_);
  and (_35208_, _35207_, _35205_);
  and (_35209_, _34912_, _09829_);
  or (_35210_, _35209_, _38088_);
  or (_35211_, _35210_, _35208_);
  and (_40373_, _35211_, _34910_);
  and (_35213_, _38088_, \oc8051_golden_model_1.P0INREG [0]);
  or (_35214_, _35213_, _38455_);
  and (_40374_, _35214_, _37580_);
  and (_35215_, _38088_, \oc8051_golden_model_1.P0INREG [1]);
  or (_35216_, _35215_, _38448_);
  and (_40375_, _35216_, _37580_);
  and (_35217_, _38088_, \oc8051_golden_model_1.P0INREG [2]);
  or (_35218_, _35217_, _38440_);
  and (_40376_, _35218_, _37580_);
  and (_35220_, _38088_, \oc8051_golden_model_1.P0INREG [3]);
  or (_35221_, _35220_, _38433_);
  and (_40377_, _35221_, _37580_);
  and (_35222_, _38088_, \oc8051_golden_model_1.P0INREG [4]);
  or (_35223_, _35222_, _38487_);
  and (_40378_, _35223_, _37580_);
  and (_35224_, _38088_, \oc8051_golden_model_1.P0INREG [5]);
  or (_35225_, _35224_, _38480_);
  and (_40379_, _35225_, _37580_);
  and (_35226_, _38088_, \oc8051_golden_model_1.P0INREG [6]);
  or (_35228_, _35226_, _38472_);
  and (_40381_, _35228_, _37580_);
  and (_35229_, _38088_, \oc8051_golden_model_1.P1INREG [0]);
  or (_35230_, _35229_, _38161_);
  and (_40382_, _35230_, _37580_);
  and (_35231_, _38088_, \oc8051_golden_model_1.P1INREG [1]);
  or (_35232_, _35231_, _38154_);
  and (_40383_, _35232_, _37580_);
  and (_35233_, _38088_, \oc8051_golden_model_1.P1INREG [2]);
  or (_35234_, _35233_, _38146_);
  and (_40385_, _35234_, _37580_);
  and (_35236_, _38088_, \oc8051_golden_model_1.P1INREG [3]);
  or (_35237_, _35236_, _38139_);
  and (_40386_, _35237_, _37580_);
  and (_35238_, _38088_, \oc8051_golden_model_1.P1INREG [4]);
  or (_35239_, _35238_, _38262_);
  and (_40387_, _35239_, _37580_);
  and (_35240_, _38088_, \oc8051_golden_model_1.P1INREG [5]);
  or (_35241_, _35240_, _38255_);
  and (_40388_, _35241_, _37580_);
  and (_35243_, _38088_, \oc8051_golden_model_1.P1INREG [6]);
  or (_35244_, _35243_, _38247_);
  and (_40389_, _35244_, _37580_);
  and (_35245_, _38088_, \oc8051_golden_model_1.P2INREG [0]);
  or (_35246_, _35245_, _38117_);
  and (_40391_, _35246_, _37580_);
  and (_35247_, _38088_, \oc8051_golden_model_1.P2INREG [1]);
  or (_35248_, _35247_, _38109_);
  and (_40392_, _35248_, _37580_);
  and (_35249_, _38088_, \oc8051_golden_model_1.P2INREG [2]);
  or (_35251_, _35249_, _38100_);
  and (_40393_, _35251_, _37580_);
  and (_35252_, _38088_, \oc8051_golden_model_1.P2INREG [3]);
  or (_35253_, _35252_, _38090_);
  and (_40394_, _35253_, _37580_);
  and (_35254_, _38088_, \oc8051_golden_model_1.P2INREG [4]);
  or (_35255_, _35254_, _38221_);
  and (_40395_, _35255_, _37580_);
  and (_35256_, _38088_, \oc8051_golden_model_1.P2INREG [5]);
  or (_35257_, _35256_, _38214_);
  and (_40396_, _35257_, _37580_);
  and (_35260_, _38088_, \oc8051_golden_model_1.P2INREG [6]);
  or (_35261_, _35260_, _38206_);
  and (_40397_, _35261_, _37580_);
  and (_35262_, _38088_, \oc8051_golden_model_1.P3INREG [0]);
  or (_35263_, _35262_, _38381_);
  and (_40399_, _35263_, _37580_);
  and (_35264_, _38088_, \oc8051_golden_model_1.P3INREG [1]);
  or (_35265_, _35264_, _38373_);
  and (_40400_, _35265_, _37580_);
  and (_35267_, _38088_, \oc8051_golden_model_1.P3INREG [2]);
  or (_35268_, _35267_, _38366_);
  and (_40401_, _35268_, _37580_);
  and (_35269_, _38088_, \oc8051_golden_model_1.P3INREG [3]);
  or (_35270_, _35269_, _38388_);
  and (_40402_, _35270_, _37580_);
  and (_35271_, _38088_, \oc8051_golden_model_1.P3INREG [4]);
  or (_35272_, _35271_, _38413_);
  and (_40404_, _35272_, _37580_);
  and (_35273_, _38088_, \oc8051_golden_model_1.P3INREG [5]);
  or (_35275_, _35273_, _38405_);
  and (_40405_, _35275_, _37580_);
  and (_35276_, _38088_, \oc8051_golden_model_1.P3INREG [6]);
  or (_35277_, _35276_, _38398_);
  and (_40406_, _35277_, _37580_);
  and (_00003_[6], _38399_, _37580_);
  and (_00003_[5], _38406_, _37580_);
  and (_00003_[4], _38414_, _37580_);
  and (_00003_[3], _38389_, _37580_);
  and (_00003_[2], _38367_, _37580_);
  and (_00003_[1], _38374_, _37580_);
  and (_00003_[0], _38382_, _37580_);
  and (_00002_[6], _38207_, _37580_);
  and (_00002_[5], _38215_, _37580_);
  and (_00002_[4], _38222_, _37580_);
  and (_00002_[3], _38091_, _37580_);
  and (_00002_[2], _38101_, _37580_);
  and (_00002_[1], _38110_, _37580_);
  and (_00002_[0], _38118_, _37580_);
  and (_00001_[6], _38248_, _37580_);
  and (_00001_[5], _38256_, _37580_);
  and (_00001_[4], _38263_, _37580_);
  and (_00001_[3], _38140_, _37580_);
  and (_00001_[2], _38147_, _37580_);
  and (_00001_[1], _38155_, _37580_);
  and (_00001_[0], _38162_, _37580_);
  and (_00000_[6], _38473_, _37580_);
  and (_00000_[5], _38481_, _37580_);
  and (_00000_[4], _38488_, _37580_);
  and (_00000_[3], _38434_, _37580_);
  and (_00000_[2], _38441_, _37580_);
  and (_00000_[1], _38449_, _37580_);
  and (_00000_[0], _38456_, _37580_);
  not (_35281_, _37932_);
  nor (_35282_, _02338_, _35281_);
  and (_35283_, _02338_, _35281_);
  or (_35284_, _35283_, _35282_);
  not (_35285_, _37949_);
  nor (_35286_, _02159_, _35285_);
  and (_35287_, _02159_, _35285_);
  or (_35288_, _35287_, _35286_);
  or (_35289_, _35288_, _35284_);
  not (_35290_, _37966_);
  nor (_35291_, _04657_, _35290_);
  and (_35292_, _04657_, _35290_);
  or (_35293_, _35292_, _35291_);
  not (_35294_, _37983_);
  nor (_35295_, _04626_, _35294_);
  and (_35296_, _04626_, _35294_);
  or (_35297_, _35296_, _35295_);
  or (_35299_, _35297_, _35293_);
  or (_35300_, _35299_, _35289_);
  or (_35301_, _02687_, _37915_);
  nand (_35302_, _02687_, _37915_);
  and (_35303_, _35302_, _35301_);
  nand (_35304_, _02568_, _37898_);
  or (_35305_, _02568_, _37898_);
  and (_35306_, _35305_, _35304_);
  or (_35307_, _35306_, _35303_);
  nand (_35308_, _04594_, _38000_);
  or (_35310_, _04594_, _38000_);
  and (_35311_, _35310_, _35308_);
  nor (_35312_, _04560_, _37881_);
  and (_35313_, _04560_, _37881_);
  or (_35314_, _35313_, _35312_);
  or (_35315_, _35314_, _35311_);
  or (_35316_, _35315_, _35307_);
  or (_35317_, _35316_, _35300_);
  nand (_35318_, _02095_, _39673_);
  or (_35319_, _02095_, _39673_);
  and (_35321_, _35319_, _35318_);
  or (_35322_, _01559_, _20640_);
  nand (_35323_, _01559_, _20640_);
  and (_35324_, _35323_, _35322_);
  or (_35325_, _01544_, _19887_);
  or (_35326_, _01369_, _19898_);
  and (_35327_, _35326_, _35325_);
  or (_35328_, _35327_, _35324_);
  or (_35329_, _01434_, _19648_);
  nand (_35330_, _01434_, _19648_);
  and (_35332_, _35330_, _35329_);
  and (_35333_, _01465_, _19408_);
  nor (_35334_, _01465_, _19408_);
  or (_35335_, _35334_, _35333_);
  or (_35336_, _35335_, _35332_);
  or (_35337_, _35336_, _35328_);
  nor (_35338_, _01533_, _19131_);
  and (_35339_, _01533_, _19131_);
  or (_35340_, _35339_, _35338_);
  nor (_35341_, _01498_, _18869_);
  and (_35343_, _01498_, _18869_);
  or (_35344_, _35343_, _35341_);
  or (_35345_, _35344_, _35340_);
  or (_35346_, _01306_, _20400_);
  nand (_35347_, _01306_, _20400_);
  and (_35348_, _35347_, _35346_);
  not (_35349_, _01337_);
  and (_35350_, _35349_, _20160_);
  nor (_35351_, _35349_, _20160_);
  or (_35352_, _35351_, _35350_);
  or (_35354_, _35352_, _35348_);
  or (_35355_, _35354_, _35345_);
  or (_35356_, _35355_, _35337_);
  nor (_35357_, \oc8051_golden_model_1.PC [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_35358_, \oc8051_golden_model_1.PC [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  or (_35359_, _35358_, _35357_);
  nor (_35360_, \oc8051_golden_model_1.PC [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_35361_, \oc8051_golden_model_1.PC [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  or (_35362_, _35361_, _35360_);
  and (_35363_, _35362_, _35359_);
  or (_35365_, \oc8051_golden_model_1.PC [12], _39711_);
  nand (_35366_, \oc8051_golden_model_1.PC [12], _39711_);
  and (_35367_, _35366_, _35365_);
  or (_35368_, _09883_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  or (_35369_, \oc8051_golden_model_1.PC [13], _39715_);
  and (_35370_, _35369_, _35368_);
  and (_35371_, _35370_, _35367_);
  and (_35372_, _35371_, _35363_);
  and (_35373_, \oc8051_golden_model_1.PC [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_35374_, \oc8051_golden_model_1.PC [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  or (_35376_, _35374_, _35373_);
  nor (_35377_, \oc8051_golden_model_1.PC [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_35378_, \oc8051_golden_model_1.PC [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  or (_35379_, _35378_, _35377_);
  and (_35380_, _35379_, _35376_);
  and (_35381_, \oc8051_golden_model_1.PC [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor (_35382_, \oc8051_golden_model_1.PC [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  or (_35383_, _35382_, _35381_);
  nor (_35384_, \oc8051_golden_model_1.PC [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_35385_, \oc8051_golden_model_1.PC [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  or (_35387_, _35385_, _35384_);
  and (_35388_, _35387_, _35383_);
  and (_35389_, _35388_, _35380_);
  and (_35390_, _35389_, _35372_);
  or (_35391_, \oc8051_golden_model_1.PC [1], _39673_);
  or (_35392_, _01253_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_35393_, _35392_, _35391_);
  nor (_35394_, \oc8051_golden_model_1.PC [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_35395_, \oc8051_golden_model_1.PC [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  or (_35396_, _35395_, _35394_);
  and (_35398_, _35396_, _35393_);
  and (_35399_, \oc8051_golden_model_1.PC [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nor (_35400_, \oc8051_golden_model_1.PC [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  or (_35401_, _35400_, _35399_);
  or (_35402_, _01249_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  or (_35403_, \oc8051_golden_model_1.PC [3], _39681_);
  and (_35404_, _35403_, _35402_);
  and (_35405_, _35404_, _35401_);
  and (_35406_, _35405_, _35398_);
  nor (_35407_, \oc8051_golden_model_1.PC [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_35409_, \oc8051_golden_model_1.PC [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  or (_35410_, _35409_, _35407_);
  nor (_35411_, \oc8051_golden_model_1.PC [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_35412_, \oc8051_golden_model_1.PC [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  or (_35413_, _35412_, _35411_);
  and (_35414_, _35413_, _35410_);
  and (_35415_, \oc8051_golden_model_1.PC [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor (_35416_, \oc8051_golden_model_1.PC [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  or (_35417_, _35416_, _35415_);
  or (_35418_, \oc8051_golden_model_1.PC [6], _39691_);
  or (_35420_, _32363_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_35421_, _35420_, _35418_);
  and (_35422_, _35421_, _35417_);
  and (_35423_, _35422_, _35414_);
  and (_35424_, _35423_, _35406_);
  and (_35425_, _35424_, _35390_);
  and (_35426_, _35425_, _38087_);
  and (_35427_, _35426_, _35356_);
  and (_35428_, _35427_, _35321_);
  and (_35429_, _39045_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_35431_, \oc8051_top_1.oc8051_memory_interface1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor (_35432_, _35431_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nor (_35433_, _35432_, _35429_);
  nand (_35434_, _35433_, _01662_);
  or (_35435_, _35433_, _01662_);
  and (_35436_, _35435_, _35434_);
  and (_35437_, _35436_, _35428_);
  or (_35438_, _01718_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_35439_, _31634_, \oc8051_golden_model_1.ACC [4]);
  nor (_35440_, _31634_, \oc8051_golden_model_1.ACC [4]);
  nor (_35443_, _35440_, _35439_);
  nor (_35444_, _01691_, _01688_);
  nor (_35445_, _35444_, _01690_);
  nor (_35446_, _35445_, _35443_);
  and (_35447_, _35445_, _35443_);
  or (_35448_, _35447_, _35446_);
  or (_35449_, _35448_, _01609_);
  nor (_35450_, _31814_, _01550_);
  nor (_35451_, _31634_, _01549_);
  and (_35452_, _35451_, _01577_);
  or (_35454_, _35452_, _35450_);
  nand (_35455_, _35454_, _01708_);
  and (_35456_, _35455_, _35449_);
  or (_35457_, _35456_, _01658_);
  or (_35458_, _10048_, _01716_);
  and (_35459_, _35458_, _35457_);
  or (_35460_, _39046_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_35461_, _35460_, _39047_);
  or (_35462_, _35461_, _39669_);
  or (_35463_, \oc8051_top_1.oc8051_memory_interface1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_35465_, _35463_, _35462_);
  nor (_35466_, _35465_, _35459_);
  and (_35467_, _35465_, _35459_);
  or (_35468_, _35467_, _35466_);
  and (_35469_, _35468_, _35438_);
  nor (_35470_, _39053_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  nor (_35471_, _35470_, _39054_);
  not (_35472_, _35471_);
  nor (_35473_, _10021_, _02089_);
  and (_35474_, _33686_, _02089_);
  nor (_35476_, _35474_, _35473_);
  nand (_35477_, _35476_, _35472_);
  nor (_35478_, _10001_, _02089_);
  not (_35479_, _34912_);
  and (_35480_, _35479_, _02089_);
  or (_35481_, _35480_, _35478_);
  or (_35482_, _35481_, _40164_);
  and (_35483_, _35482_, _35477_);
  or (_35484_, _10013_, _02089_);
  nand (_35485_, _34306_, _02089_);
  nand (_35487_, _35485_, _35484_);
  nand (_35488_, _35487_, _40119_);
  nor (_35489_, _39050_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor (_35490_, _35489_, _39051_);
  nor (_35491_, _04388_, _02089_);
  and (_35492_, _32683_, _02089_);
  nor (_35493_, _35492_, _35491_);
  nand (_35494_, _35493_, _35490_);
  and (_35495_, _35494_, _35488_);
  and (_35496_, _35495_, _35483_);
  nor (_35498_, _39049_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_35499_, _35498_, _39050_);
  nor (_35500_, _10036_, _02089_);
  and (_35501_, _32335_, _02089_);
  nor (_35502_, _35501_, _35500_);
  not (_35503_, _35502_);
  nand (_35504_, _35503_, _35499_);
  or (_35505_, _02092_, _39669_);
  and (_35506_, _35505_, _35504_);
  and (_35507_, _39051_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor (_35509_, _39051_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor (_35510_, _35509_, _35507_);
  nor (_35511_, _10030_, _02089_);
  and (_35512_, _33053_, _02089_);
  or (_35513_, _35512_, _35511_);
  or (_35514_, _35513_, _35510_);
  or (_35515_, _35476_, _35472_);
  and (_35516_, _35515_, _35514_);
  and (_35517_, _35516_, _35506_);
  and (_35518_, _35517_, _35496_);
  and (_35520_, _34607_, _02089_);
  nor (_35521_, _11694_, _02089_);
  nor (_35522_, _35521_, _35520_);
  nand (_35523_, _35522_, _40143_);
  or (_35524_, _35503_, _35499_);
  or (_35525_, _35522_, _40143_);
  and (_35526_, _35525_, _35524_);
  and (_35527_, _35526_, _35523_);
  or (_35528_, _35493_, _35490_);
  nor (_35529_, _39045_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nor (_35531_, _35529_, _39046_);
  or (_35532_, _35531_, _02105_);
  and (_35533_, _35532_, _35528_);
  nor (_35534_, _35507_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  or (_35535_, _35534_, _39053_);
  and (_35536_, _33367_, _02089_);
  not (_35537_, _10026_);
  nor (_35538_, _35537_, _02089_);
  or (_35539_, _35538_, _35536_);
  or (_35540_, _35539_, _35535_);
  or (_35542_, _10049_, _02089_);
  nand (_35543_, _31634_, _02089_);
  and (_35544_, _35543_, _35542_);
  or (_35545_, _35544_, _35461_);
  and (_35546_, _35545_, _35540_);
  and (_35547_, _35546_, _35533_);
  and (_35548_, _35547_, _35527_);
  and (_35549_, _35548_, _35518_);
  and (_35550_, _35549_, _35469_);
  and (_35551_, _35550_, _35437_);
  and (_35552_, _35551_, _35317_);
  nor (_35553_, _11895_, _01657_);
  nor (_35554_, _35059_, _01550_);
  nor (_35555_, _34912_, _01579_);
  and (_35556_, _11895_, _01579_);
  nor (_35557_, _35556_, _35555_);
  nor (_35558_, _35557_, _01549_);
  nor (_35559_, _35558_, _01663_);
  not (_35560_, _35559_);
  nor (_35561_, _35560_, _35554_);
  nor (_35563_, _11895_, _01605_);
  or (_35564_, _35563_, _01608_);
  nor (_35565_, _35564_, _35561_);
  and (_35566_, _32683_, \oc8051_golden_model_1.ACC [7]);
  nor (_35567_, _32683_, \oc8051_golden_model_1.ACC [7]);
  nor (_35568_, _35567_, _35566_);
  and (_35569_, _32334_, \oc8051_golden_model_1.ACC [6]);
  nor (_35570_, _32334_, \oc8051_golden_model_1.ACC [6]);
  nor (_35571_, _35570_, _35569_);
  and (_35572_, _31977_, \oc8051_golden_model_1.ACC [5]);
  nor (_35574_, _31977_, \oc8051_golden_model_1.ACC [5]);
  nor (_35575_, _35574_, _35572_);
  and (_35576_, _35575_, _35439_);
  nor (_35577_, _35576_, _35572_);
  not (_35578_, _35445_);
  and (_35579_, _35575_, _35443_);
  nand (_35580_, _35579_, _35578_);
  nand (_35581_, _35580_, _35577_);
  and (_35582_, _35581_, _35571_);
  or (_35583_, _35582_, _35569_);
  and (_35585_, _35583_, _35568_);
  nor (_35586_, _35585_, _35566_);
  and (_35587_, _33367_, _33052_);
  and (_35588_, _33993_, _33685_);
  and (_35589_, _35588_, _35587_);
  not (_35590_, _35589_);
  nor (_35591_, _35590_, _35586_);
  and (_35592_, _34607_, _34305_);
  and (_35593_, _35592_, _35591_);
  and (_35594_, _35593_, _34912_);
  nor (_35596_, _35593_, _34912_);
  nor (_35597_, _35596_, _35594_);
  nor (_35598_, _35597_, _01609_);
  nor (_35599_, _35598_, _01658_);
  not (_35600_, _35599_);
  nor (_35601_, _35600_, _35565_);
  nor (_35602_, _35601_, _35553_);
  and (_35603_, \oc8051_top_1.oc8051_memory_interface1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_35604_, _39051_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_35605_, _35604_, _39164_);
  and (_35607_, _35605_, _35603_);
  and (_35608_, _35607_, _39076_);
  nor (_35609_, _35607_, _39076_);
  or (_35610_, _35609_, _35608_);
  nand (_35611_, _35610_, _35602_);
  or (_35612_, _35610_, _35602_);
  and (_35613_, _35612_, _35611_);
  and (_35614_, _02584_, _36057_);
  nor (_35615_, _02584_, _36057_);
  or (_35616_, _35615_, _35614_);
  not (_35618_, _36175_);
  nor (_35619_, _01822_, _35618_);
  and (_35620_, _01822_, _35618_);
  or (_35621_, _35620_, _35619_);
  or (_35622_, _35621_, _35616_);
  nand (_35623_, _02252_, _35921_);
  or (_35624_, _02252_, _35921_);
  and (_35625_, _35624_, _35623_);
  and (_35626_, _01790_, _35844_);
  nor (_35627_, _01790_, _35844_);
  or (_35629_, _35627_, _35626_);
  or (_35630_, _35629_, _35625_);
  or (_35631_, _35630_, _35622_);
  nand (_35632_, _02294_, _35976_);
  or (_35633_, _02294_, _35976_);
  and (_35634_, _35633_, _35632_);
  and (_35635_, _01955_, _36020_);
  nor (_35636_, _01955_, _36020_);
  or (_35637_, _35636_, _35635_);
  or (_35638_, _35637_, _35634_);
  or (_35640_, _01855_, _36151_);
  nand (_35641_, _01855_, _36151_);
  and (_35642_, _35641_, _35640_);
  nor (_35643_, _03379_, _36088_);
  and (_35644_, _03379_, _36088_);
  or (_35645_, _35644_, _35643_);
  or (_35646_, _35645_, _35642_);
  or (_35647_, _35646_, _35638_);
  or (_35648_, _35647_, _35631_);
  and (_35649_, _35648_, _35613_);
  and (property_invalid_rom_pc, _35649_, _35552_);
  and (_00000_[7], _38466_, _37580_);
  and (_00001_[7], _38241_, _37580_);
  and (_00002_[7], _38200_, _37580_);
  and (_00003_[7], _38421_, _37580_);
  buf (_00065_, _37580_);
  buf (_00116_, _37580_);
  buf (_00168_, _37580_);
  buf (_00220_, _37580_);
  buf (_00272_, _37580_);
  buf (_00324_, _37580_);
  buf (_00376_, _37580_);
  buf (_00428_, _37580_);
  buf (_00480_, _37580_);
  buf (_00532_, _37580_);
  buf (_00584_, _37580_);
  buf (_00636_, _37580_);
  buf (_00687_, _37580_);
  buf (_00739_, _37580_);
  buf (_00790_, _37580_);
  buf (_00842_, _37580_);
  buf (_03175_, _00918_);
  buf (_03178_, _00922_);
  buf (_03212_, _00918_);
  buf (_03215_, _00922_);
  buf (_05689_, _01063_);
  buf (_05691_, _01066_);
  buf (_05693_, _01069_);
  buf (_05695_, _01072_);
  buf (_05697_, _01075_);
  buf (_05699_, _01078_);
  buf (_05701_, _01081_);
  buf (_05703_, _01084_);
  buf (_05705_, _01087_);
  buf (_05707_, _01090_);
  buf (_05709_, _01093_);
  buf (_05711_, _01095_);
  buf (_05713_, _01098_);
  buf (_05715_, _01101_);
  buf (_05809_, _01063_);
  buf (_05811_, _01066_);
  buf (_05813_, _01069_);
  buf (_05815_, _01072_);
  buf (_05817_, _01075_);
  buf (_05819_, _01078_);
  buf (_05821_, _01081_);
  buf (_05823_, _01084_);
  buf (_05825_, _01087_);
  buf (_05827_, _01090_);
  buf (_05829_, _01093_);
  buf (_05831_, _01095_);
  buf (_05833_, _01098_);
  buf (_05835_, _01101_);
  buf (_08208_, _01528_);
  buf (_08311_, _01528_);
  dff (p0in_reg[0], _00000_[0]);
  dff (p0in_reg[1], _00000_[1]);
  dff (p0in_reg[2], _00000_[2]);
  dff (p0in_reg[3], _00000_[3]);
  dff (p0in_reg[4], _00000_[4]);
  dff (p0in_reg[5], _00000_[5]);
  dff (p0in_reg[6], _00000_[6]);
  dff (p0in_reg[7], _00000_[7]);
  dff (p1in_reg[0], _00001_[0]);
  dff (p1in_reg[1], _00001_[1]);
  dff (p1in_reg[2], _00001_[2]);
  dff (p1in_reg[3], _00001_[3]);
  dff (p1in_reg[4], _00001_[4]);
  dff (p1in_reg[5], _00001_[5]);
  dff (p1in_reg[6], _00001_[6]);
  dff (p1in_reg[7], _00001_[7]);
  dff (p2in_reg[0], _00002_[0]);
  dff (p2in_reg[1], _00002_[1]);
  dff (p2in_reg[2], _00002_[2]);
  dff (p2in_reg[3], _00002_[3]);
  dff (p2in_reg[4], _00002_[4]);
  dff (p2in_reg[5], _00002_[5]);
  dff (p2in_reg[6], _00002_[6]);
  dff (p2in_reg[7], _00002_[7]);
  dff (p3in_reg[0], _00003_[0]);
  dff (p3in_reg[1], _00003_[1]);
  dff (p3in_reg[2], _00003_[2]);
  dff (p3in_reg[3], _00003_[3]);
  dff (p3in_reg[4], _00003_[4]);
  dff (p3in_reg[5], _00003_[5]);
  dff (p3in_reg[6], _00003_[6]);
  dff (p3in_reg[7], _00003_[7]);
  dff (\oc8051_gm_cxrom_1.cell0.data [0], _00094_);
  dff (\oc8051_gm_cxrom_1.cell0.data [1], _00096_);
  dff (\oc8051_gm_cxrom_1.cell0.data [2], _00098_);
  dff (\oc8051_gm_cxrom_1.cell0.data [3], _00100_);
  dff (\oc8051_gm_cxrom_1.cell0.data [4], _00102_);
  dff (\oc8051_gm_cxrom_1.cell0.data [5], _00104_);
  dff (\oc8051_gm_cxrom_1.cell0.data [6], _00106_);
  dff (\oc8051_gm_cxrom_1.cell0.data [7], _00062_);
  dff (\oc8051_gm_cxrom_1.cell0.valid , _00065_);
  dff (\oc8051_gm_cxrom_1.cell1.data [0], _00145_);
  dff (\oc8051_gm_cxrom_1.cell1.data [1], _00147_);
  dff (\oc8051_gm_cxrom_1.cell1.data [2], _00149_);
  dff (\oc8051_gm_cxrom_1.cell1.data [3], _00151_);
  dff (\oc8051_gm_cxrom_1.cell1.data [4], _00153_);
  dff (\oc8051_gm_cxrom_1.cell1.data [5], _00155_);
  dff (\oc8051_gm_cxrom_1.cell1.data [6], _00157_);
  dff (\oc8051_gm_cxrom_1.cell1.data [7], _00113_);
  dff (\oc8051_gm_cxrom_1.cell1.valid , _00116_);
  dff (\oc8051_gm_cxrom_1.cell10.data [0], _00613_);
  dff (\oc8051_gm_cxrom_1.cell10.data [1], _00615_);
  dff (\oc8051_gm_cxrom_1.cell10.data [2], _00617_);
  dff (\oc8051_gm_cxrom_1.cell10.data [3], _00619_);
  dff (\oc8051_gm_cxrom_1.cell10.data [4], _00621_);
  dff (\oc8051_gm_cxrom_1.cell10.data [5], _00623_);
  dff (\oc8051_gm_cxrom_1.cell10.data [6], _00625_);
  dff (\oc8051_gm_cxrom_1.cell10.data [7], _00581_);
  dff (\oc8051_gm_cxrom_1.cell10.valid , _00584_);
  dff (\oc8051_gm_cxrom_1.cell11.data [0], _00665_);
  dff (\oc8051_gm_cxrom_1.cell11.data [1], _00667_);
  dff (\oc8051_gm_cxrom_1.cell11.data [2], _00669_);
  dff (\oc8051_gm_cxrom_1.cell11.data [3], _00671_);
  dff (\oc8051_gm_cxrom_1.cell11.data [4], _00673_);
  dff (\oc8051_gm_cxrom_1.cell11.data [5], _00675_);
  dff (\oc8051_gm_cxrom_1.cell11.data [6], _00677_);
  dff (\oc8051_gm_cxrom_1.cell11.data [7], _00633_);
  dff (\oc8051_gm_cxrom_1.cell11.valid , _00636_);
  dff (\oc8051_gm_cxrom_1.cell12.data [0], _00716_);
  dff (\oc8051_gm_cxrom_1.cell12.data [1], _00718_);
  dff (\oc8051_gm_cxrom_1.cell12.data [2], _00720_);
  dff (\oc8051_gm_cxrom_1.cell12.data [3], _00722_);
  dff (\oc8051_gm_cxrom_1.cell12.data [4], _00724_);
  dff (\oc8051_gm_cxrom_1.cell12.data [5], _00726_);
  dff (\oc8051_gm_cxrom_1.cell12.data [6], _00728_);
  dff (\oc8051_gm_cxrom_1.cell12.data [7], _00684_);
  dff (\oc8051_gm_cxrom_1.cell12.valid , _00687_);
  dff (\oc8051_gm_cxrom_1.cell13.data [0], _00768_);
  dff (\oc8051_gm_cxrom_1.cell13.data [1], _00770_);
  dff (\oc8051_gm_cxrom_1.cell13.data [2], _00772_);
  dff (\oc8051_gm_cxrom_1.cell13.data [3], _00774_);
  dff (\oc8051_gm_cxrom_1.cell13.data [4], _00776_);
  dff (\oc8051_gm_cxrom_1.cell13.data [5], _00778_);
  dff (\oc8051_gm_cxrom_1.cell13.data [6], _00780_);
  dff (\oc8051_gm_cxrom_1.cell13.data [7], _00736_);
  dff (\oc8051_gm_cxrom_1.cell13.valid , _00739_);
  dff (\oc8051_gm_cxrom_1.cell14.data [0], _00819_);
  dff (\oc8051_gm_cxrom_1.cell14.data [1], _00821_);
  dff (\oc8051_gm_cxrom_1.cell14.data [2], _00823_);
  dff (\oc8051_gm_cxrom_1.cell14.data [3], _00825_);
  dff (\oc8051_gm_cxrom_1.cell14.data [4], _00827_);
  dff (\oc8051_gm_cxrom_1.cell14.data [5], _00829_);
  dff (\oc8051_gm_cxrom_1.cell14.data [6], _00831_);
  dff (\oc8051_gm_cxrom_1.cell14.data [7], _00787_);
  dff (\oc8051_gm_cxrom_1.cell14.valid , _00790_);
  dff (\oc8051_gm_cxrom_1.cell15.data [0], _00871_);
  dff (\oc8051_gm_cxrom_1.cell15.data [1], _00873_);
  dff (\oc8051_gm_cxrom_1.cell15.data [2], _00875_);
  dff (\oc8051_gm_cxrom_1.cell15.data [3], _00877_);
  dff (\oc8051_gm_cxrom_1.cell15.data [4], _00879_);
  dff (\oc8051_gm_cxrom_1.cell15.data [5], _00881_);
  dff (\oc8051_gm_cxrom_1.cell15.data [6], _00883_);
  dff (\oc8051_gm_cxrom_1.cell15.data [7], _00839_);
  dff (\oc8051_gm_cxrom_1.cell15.valid , _00842_);
  dff (\oc8051_gm_cxrom_1.cell2.data [0], _00197_);
  dff (\oc8051_gm_cxrom_1.cell2.data [1], _00199_);
  dff (\oc8051_gm_cxrom_1.cell2.data [2], _00201_);
  dff (\oc8051_gm_cxrom_1.cell2.data [3], _00203_);
  dff (\oc8051_gm_cxrom_1.cell2.data [4], _00205_);
  dff (\oc8051_gm_cxrom_1.cell2.data [5], _00207_);
  dff (\oc8051_gm_cxrom_1.cell2.data [6], _00209_);
  dff (\oc8051_gm_cxrom_1.cell2.data [7], _00165_);
  dff (\oc8051_gm_cxrom_1.cell2.valid , _00168_);
  dff (\oc8051_gm_cxrom_1.cell3.data [0], _00249_);
  dff (\oc8051_gm_cxrom_1.cell3.data [1], _00251_);
  dff (\oc8051_gm_cxrom_1.cell3.data [2], _00253_);
  dff (\oc8051_gm_cxrom_1.cell3.data [3], _00255_);
  dff (\oc8051_gm_cxrom_1.cell3.data [4], _00257_);
  dff (\oc8051_gm_cxrom_1.cell3.data [5], _00259_);
  dff (\oc8051_gm_cxrom_1.cell3.data [6], _00261_);
  dff (\oc8051_gm_cxrom_1.cell3.data [7], _00217_);
  dff (\oc8051_gm_cxrom_1.cell3.valid , _00220_);
  dff (\oc8051_gm_cxrom_1.cell4.data [0], _00302_);
  dff (\oc8051_gm_cxrom_1.cell4.data [1], _00304_);
  dff (\oc8051_gm_cxrom_1.cell4.data [2], _00306_);
  dff (\oc8051_gm_cxrom_1.cell4.data [3], _00307_);
  dff (\oc8051_gm_cxrom_1.cell4.data [4], _00309_);
  dff (\oc8051_gm_cxrom_1.cell4.data [5], _00311_);
  dff (\oc8051_gm_cxrom_1.cell4.data [6], _00313_);
  dff (\oc8051_gm_cxrom_1.cell4.data [7], _00269_);
  dff (\oc8051_gm_cxrom_1.cell4.valid , _00272_);
  dff (\oc8051_gm_cxrom_1.cell5.data [0], _00354_);
  dff (\oc8051_gm_cxrom_1.cell5.data [1], _00356_);
  dff (\oc8051_gm_cxrom_1.cell5.data [2], _00358_);
  dff (\oc8051_gm_cxrom_1.cell5.data [3], _00360_);
  dff (\oc8051_gm_cxrom_1.cell5.data [4], _00362_);
  dff (\oc8051_gm_cxrom_1.cell5.data [5], _00364_);
  dff (\oc8051_gm_cxrom_1.cell5.data [6], _00365_);
  dff (\oc8051_gm_cxrom_1.cell5.data [7], _00321_);
  dff (\oc8051_gm_cxrom_1.cell5.valid , _00324_);
  dff (\oc8051_gm_cxrom_1.cell6.data [0], _00406_);
  dff (\oc8051_gm_cxrom_1.cell6.data [1], _00408_);
  dff (\oc8051_gm_cxrom_1.cell6.data [2], _00410_);
  dff (\oc8051_gm_cxrom_1.cell6.data [3], _00412_);
  dff (\oc8051_gm_cxrom_1.cell6.data [4], _00414_);
  dff (\oc8051_gm_cxrom_1.cell6.data [5], _00416_);
  dff (\oc8051_gm_cxrom_1.cell6.data [6], _00418_);
  dff (\oc8051_gm_cxrom_1.cell6.data [7], _00373_);
  dff (\oc8051_gm_cxrom_1.cell6.valid , _00376_);
  dff (\oc8051_gm_cxrom_1.cell7.data [0], _00458_);
  dff (\oc8051_gm_cxrom_1.cell7.data [1], _00460_);
  dff (\oc8051_gm_cxrom_1.cell7.data [2], _00462_);
  dff (\oc8051_gm_cxrom_1.cell7.data [3], _00464_);
  dff (\oc8051_gm_cxrom_1.cell7.data [4], _00466_);
  dff (\oc8051_gm_cxrom_1.cell7.data [5], _00468_);
  dff (\oc8051_gm_cxrom_1.cell7.data [6], _00470_);
  dff (\oc8051_gm_cxrom_1.cell7.data [7], _00425_);
  dff (\oc8051_gm_cxrom_1.cell7.valid , _00428_);
  dff (\oc8051_gm_cxrom_1.cell8.data [0], _00510_);
  dff (\oc8051_gm_cxrom_1.cell8.data [1], _00512_);
  dff (\oc8051_gm_cxrom_1.cell8.data [2], _00514_);
  dff (\oc8051_gm_cxrom_1.cell8.data [3], _00516_);
  dff (\oc8051_gm_cxrom_1.cell8.data [4], _00518_);
  dff (\oc8051_gm_cxrom_1.cell8.data [5], _00520_);
  dff (\oc8051_gm_cxrom_1.cell8.data [6], _00522_);
  dff (\oc8051_gm_cxrom_1.cell8.data [7], _00477_);
  dff (\oc8051_gm_cxrom_1.cell8.valid , _00480_);
  dff (\oc8051_gm_cxrom_1.cell9.data [0], _00562_);
  dff (\oc8051_gm_cxrom_1.cell9.data [1], _00564_);
  dff (\oc8051_gm_cxrom_1.cell9.data [2], _00565_);
  dff (\oc8051_gm_cxrom_1.cell9.data [3], _00567_);
  dff (\oc8051_gm_cxrom_1.cell9.data [4], _00569_);
  dff (\oc8051_gm_cxrom_1.cell9.data [5], _00571_);
  dff (\oc8051_gm_cxrom_1.cell9.data [6], _00573_);
  dff (\oc8051_gm_cxrom_1.cell9.data [7], _00530_);
  dff (\oc8051_gm_cxrom_1.cell9.valid , _00532_);
  dff (\oc8051_golden_model_1.IRAM[15] [0], _37373_);
  dff (\oc8051_golden_model_1.IRAM[15] [1], _37374_);
  dff (\oc8051_golden_model_1.IRAM[15] [2], _37375_);
  dff (\oc8051_golden_model_1.IRAM[15] [3], _37377_);
  dff (\oc8051_golden_model_1.IRAM[15] [4], _37378_);
  dff (\oc8051_golden_model_1.IRAM[15] [5], _37379_);
  dff (\oc8051_golden_model_1.IRAM[15] [6], _37380_);
  dff (\oc8051_golden_model_1.IRAM[15] [7], _37136_);
  dff (\oc8051_golden_model_1.IRAM[14] [0], _37362_);
  dff (\oc8051_golden_model_1.IRAM[14] [1], _37363_);
  dff (\oc8051_golden_model_1.IRAM[14] [2], _37364_);
  dff (\oc8051_golden_model_1.IRAM[14] [3], _37366_);
  dff (\oc8051_golden_model_1.IRAM[14] [4], _37367_);
  dff (\oc8051_golden_model_1.IRAM[14] [5], _37368_);
  dff (\oc8051_golden_model_1.IRAM[14] [6], _37369_);
  dff (\oc8051_golden_model_1.IRAM[14] [7], _37370_);
  dff (\oc8051_golden_model_1.IRAM[13] [0], _37351_);
  dff (\oc8051_golden_model_1.IRAM[13] [1], _37352_);
  dff (\oc8051_golden_model_1.IRAM[13] [2], _37353_);
  dff (\oc8051_golden_model_1.IRAM[13] [3], _37354_);
  dff (\oc8051_golden_model_1.IRAM[13] [4], _37355_);
  dff (\oc8051_golden_model_1.IRAM[13] [5], _37356_);
  dff (\oc8051_golden_model_1.IRAM[13] [6], _37357_);
  dff (\oc8051_golden_model_1.IRAM[13] [7], _37358_);
  dff (\oc8051_golden_model_1.IRAM[12] [0], _37339_);
  dff (\oc8051_golden_model_1.IRAM[12] [1], _37340_);
  dff (\oc8051_golden_model_1.IRAM[12] [2], _37341_);
  dff (\oc8051_golden_model_1.IRAM[12] [3], _37342_);
  dff (\oc8051_golden_model_1.IRAM[12] [4], _37344_);
  dff (\oc8051_golden_model_1.IRAM[12] [5], _37345_);
  dff (\oc8051_golden_model_1.IRAM[12] [6], _37346_);
  dff (\oc8051_golden_model_1.IRAM[12] [7], _37347_);
  dff (\oc8051_golden_model_1.IRAM[11] [0], _37327_);
  dff (\oc8051_golden_model_1.IRAM[11] [1], _37329_);
  dff (\oc8051_golden_model_1.IRAM[11] [2], _37330_);
  dff (\oc8051_golden_model_1.IRAM[11] [3], _37331_);
  dff (\oc8051_golden_model_1.IRAM[11] [4], _37332_);
  dff (\oc8051_golden_model_1.IRAM[11] [5], _37333_);
  dff (\oc8051_golden_model_1.IRAM[11] [6], _37335_);
  dff (\oc8051_golden_model_1.IRAM[11] [7], _37336_);
  dff (\oc8051_golden_model_1.IRAM[10] [0], _37316_);
  dff (\oc8051_golden_model_1.IRAM[10] [1], _37317_);
  dff (\oc8051_golden_model_1.IRAM[10] [2], _37318_);
  dff (\oc8051_golden_model_1.IRAM[10] [3], _37319_);
  dff (\oc8051_golden_model_1.IRAM[10] [4], _37320_);
  dff (\oc8051_golden_model_1.IRAM[10] [5], _37321_);
  dff (\oc8051_golden_model_1.IRAM[10] [6], _37323_);
  dff (\oc8051_golden_model_1.IRAM[10] [7], _37324_);
  dff (\oc8051_golden_model_1.IRAM[9] [0], _37304_);
  dff (\oc8051_golden_model_1.IRAM[9] [1], _37305_);
  dff (\oc8051_golden_model_1.IRAM[9] [2], _37307_);
  dff (\oc8051_golden_model_1.IRAM[9] [3], _37308_);
  dff (\oc8051_golden_model_1.IRAM[9] [4], _37309_);
  dff (\oc8051_golden_model_1.IRAM[9] [5], _37310_);
  dff (\oc8051_golden_model_1.IRAM[9] [6], _37311_);
  dff (\oc8051_golden_model_1.IRAM[9] [7], _37313_);
  dff (\oc8051_golden_model_1.IRAM[8] [0], _37293_);
  dff (\oc8051_golden_model_1.IRAM[8] [1], _37294_);
  dff (\oc8051_golden_model_1.IRAM[8] [2], _37296_);
  dff (\oc8051_golden_model_1.IRAM[8] [3], _37297_);
  dff (\oc8051_golden_model_1.IRAM[8] [4], _37298_);
  dff (\oc8051_golden_model_1.IRAM[8] [5], _37299_);
  dff (\oc8051_golden_model_1.IRAM[8] [6], _37300_);
  dff (\oc8051_golden_model_1.IRAM[8] [7], _37302_);
  dff (\oc8051_golden_model_1.IRAM[7] [0], _37281_);
  dff (\oc8051_golden_model_1.IRAM[7] [1], _37283_);
  dff (\oc8051_golden_model_1.IRAM[7] [2], _37284_);
  dff (\oc8051_golden_model_1.IRAM[7] [3], _37285_);
  dff (\oc8051_golden_model_1.IRAM[7] [4], _37286_);
  dff (\oc8051_golden_model_1.IRAM[7] [5], _37287_);
  dff (\oc8051_golden_model_1.IRAM[7] [6], _37288_);
  dff (\oc8051_golden_model_1.IRAM[7] [7], _37289_);
  dff (\oc8051_golden_model_1.IRAM[6] [0], _37269_);
  dff (\oc8051_golden_model_1.IRAM[6] [1], _37271_);
  dff (\oc8051_golden_model_1.IRAM[6] [2], _37272_);
  dff (\oc8051_golden_model_1.IRAM[6] [3], _37273_);
  dff (\oc8051_golden_model_1.IRAM[6] [4], _37274_);
  dff (\oc8051_golden_model_1.IRAM[6] [5], _37275_);
  dff (\oc8051_golden_model_1.IRAM[6] [6], _37277_);
  dff (\oc8051_golden_model_1.IRAM[6] [7], _37278_);
  dff (\oc8051_golden_model_1.IRAM[5] [0], _37258_);
  dff (\oc8051_golden_model_1.IRAM[5] [1], _37259_);
  dff (\oc8051_golden_model_1.IRAM[5] [2], _37261_);
  dff (\oc8051_golden_model_1.IRAM[5] [3], _37262_);
  dff (\oc8051_golden_model_1.IRAM[5] [4], _37263_);
  dff (\oc8051_golden_model_1.IRAM[5] [5], _37264_);
  dff (\oc8051_golden_model_1.IRAM[5] [6], _37265_);
  dff (\oc8051_golden_model_1.IRAM[5] [7], _37267_);
  dff (\oc8051_golden_model_1.IRAM[4] [0], _37247_);
  dff (\oc8051_golden_model_1.IRAM[4] [1], _37248_);
  dff (\oc8051_golden_model_1.IRAM[4] [2], _37250_);
  dff (\oc8051_golden_model_1.IRAM[4] [3], _37251_);
  dff (\oc8051_golden_model_1.IRAM[4] [4], _37252_);
  dff (\oc8051_golden_model_1.IRAM[4] [5], _37253_);
  dff (\oc8051_golden_model_1.IRAM[4] [6], _37254_);
  dff (\oc8051_golden_model_1.IRAM[4] [7], _37255_);
  dff (\oc8051_golden_model_1.IRAM[3] [0], _37235_);
  dff (\oc8051_golden_model_1.IRAM[3] [1], _37236_);
  dff (\oc8051_golden_model_1.IRAM[3] [2], _37237_);
  dff (\oc8051_golden_model_1.IRAM[3] [3], _37238_);
  dff (\oc8051_golden_model_1.IRAM[3] [4], _37239_);
  dff (\oc8051_golden_model_1.IRAM[3] [5], _37240_);
  dff (\oc8051_golden_model_1.IRAM[3] [6], _37242_);
  dff (\oc8051_golden_model_1.IRAM[3] [7], _37243_);
  dff (\oc8051_golden_model_1.IRAM[2] [0], _37223_);
  dff (\oc8051_golden_model_1.IRAM[2] [1], _37224_);
  dff (\oc8051_golden_model_1.IRAM[2] [2], _37226_);
  dff (\oc8051_golden_model_1.IRAM[2] [3], _37227_);
  dff (\oc8051_golden_model_1.IRAM[2] [4], _37228_);
  dff (\oc8051_golden_model_1.IRAM[2] [5], _37229_);
  dff (\oc8051_golden_model_1.IRAM[2] [6], _37230_);
  dff (\oc8051_golden_model_1.IRAM[2] [7], _37232_);
  dff (\oc8051_golden_model_1.IRAM[1] [0], _37211_);
  dff (\oc8051_golden_model_1.IRAM[1] [1], _37213_);
  dff (\oc8051_golden_model_1.IRAM[1] [2], _37214_);
  dff (\oc8051_golden_model_1.IRAM[1] [3], _37215_);
  dff (\oc8051_golden_model_1.IRAM[1] [4], _37216_);
  dff (\oc8051_golden_model_1.IRAM[1] [5], _37217_);
  dff (\oc8051_golden_model_1.IRAM[1] [6], _37219_);
  dff (\oc8051_golden_model_1.IRAM[1] [7], _37220_);
  dff (\oc8051_golden_model_1.IRAM[0] [0], _37199_);
  dff (\oc8051_golden_model_1.IRAM[0] [1], _37200_);
  dff (\oc8051_golden_model_1.IRAM[0] [2], _37201_);
  dff (\oc8051_golden_model_1.IRAM[0] [3], _37203_);
  dff (\oc8051_golden_model_1.IRAM[0] [4], _37204_);
  dff (\oc8051_golden_model_1.IRAM[0] [5], _37206_);
  dff (\oc8051_golden_model_1.IRAM[0] [6], _37207_);
  dff (\oc8051_golden_model_1.IRAM[0] [7], _37208_);
  dff (\oc8051_golden_model_1.B [0], _40184_);
  dff (\oc8051_golden_model_1.B [1], _40185_);
  dff (\oc8051_golden_model_1.B [2], _40186_);
  dff (\oc8051_golden_model_1.B [3], _40187_);
  dff (\oc8051_golden_model_1.B [4], _40188_);
  dff (\oc8051_golden_model_1.B [5], _40189_);
  dff (\oc8051_golden_model_1.B [6], _40190_);
  dff (\oc8051_golden_model_1.B [7], _37137_);
  dff (\oc8051_golden_model_1.ACC [0], _40192_);
  dff (\oc8051_golden_model_1.ACC [1], _40193_);
  dff (\oc8051_golden_model_1.ACC [2], _40194_);
  dff (\oc8051_golden_model_1.ACC [3], _40195_);
  dff (\oc8051_golden_model_1.ACC [4], _40196_);
  dff (\oc8051_golden_model_1.ACC [5], _40197_);
  dff (\oc8051_golden_model_1.ACC [6], _40199_);
  dff (\oc8051_golden_model_1.ACC [7], _37139_);
  dff (\oc8051_golden_model_1.DPL [0], _40200_);
  dff (\oc8051_golden_model_1.DPL [1], _40201_);
  dff (\oc8051_golden_model_1.DPL [2], _40203_);
  dff (\oc8051_golden_model_1.DPL [3], _40204_);
  dff (\oc8051_golden_model_1.DPL [4], _40205_);
  dff (\oc8051_golden_model_1.DPL [5], _40206_);
  dff (\oc8051_golden_model_1.DPL [6], _40207_);
  dff (\oc8051_golden_model_1.DPL [7], _37140_);
  dff (\oc8051_golden_model_1.DPH [0], _40209_);
  dff (\oc8051_golden_model_1.DPH [1], _40210_);
  dff (\oc8051_golden_model_1.DPH [2], _40211_);
  dff (\oc8051_golden_model_1.DPH [3], _40212_);
  dff (\oc8051_golden_model_1.DPH [4], _40213_);
  dff (\oc8051_golden_model_1.DPH [5], _40214_);
  dff (\oc8051_golden_model_1.DPH [6], _40215_);
  dff (\oc8051_golden_model_1.DPH [7], _37141_);
  dff (\oc8051_golden_model_1.IE [0], _40217_);
  dff (\oc8051_golden_model_1.IE [1], _40218_);
  dff (\oc8051_golden_model_1.IE [2], _40219_);
  dff (\oc8051_golden_model_1.IE [3], _40220_);
  dff (\oc8051_golden_model_1.IE [4], _40222_);
  dff (\oc8051_golden_model_1.IE [5], _40223_);
  dff (\oc8051_golden_model_1.IE [6], _40224_);
  dff (\oc8051_golden_model_1.IE [7], _37142_);
  dff (\oc8051_golden_model_1.IP [0], _40225_);
  dff (\oc8051_golden_model_1.IP [1], _40226_);
  dff (\oc8051_golden_model_1.IP [2], _40227_);
  dff (\oc8051_golden_model_1.IP [3], _40228_);
  dff (\oc8051_golden_model_1.IP [4], _40229_);
  dff (\oc8051_golden_model_1.IP [5], _40230_);
  dff (\oc8051_golden_model_1.IP [6], _40231_);
  dff (\oc8051_golden_model_1.IP [7], _37143_);
  dff (\oc8051_golden_model_1.P0 [0], _40233_);
  dff (\oc8051_golden_model_1.P0 [1], _40234_);
  dff (\oc8051_golden_model_1.P0 [2], _40235_);
  dff (\oc8051_golden_model_1.P0 [3], _40236_);
  dff (\oc8051_golden_model_1.P0 [4], _40237_);
  dff (\oc8051_golden_model_1.P0 [5], _40238_);
  dff (\oc8051_golden_model_1.P0 [6], _40240_);
  dff (\oc8051_golden_model_1.P0 [7], _37145_);
  dff (\oc8051_golden_model_1.P1 [0], _40241_);
  dff (\oc8051_golden_model_1.P1 [1], _40242_);
  dff (\oc8051_golden_model_1.P1 [2], _40244_);
  dff (\oc8051_golden_model_1.P1 [3], _40245_);
  dff (\oc8051_golden_model_1.P1 [4], _40246_);
  dff (\oc8051_golden_model_1.P1 [5], _40247_);
  dff (\oc8051_golden_model_1.P1 [6], _40248_);
  dff (\oc8051_golden_model_1.P1 [7], _37146_);
  dff (\oc8051_golden_model_1.P2 [0], _40250_);
  dff (\oc8051_golden_model_1.P2 [1], _40251_);
  dff (\oc8051_golden_model_1.P2 [2], _40252_);
  dff (\oc8051_golden_model_1.P2 [3], _40253_);
  dff (\oc8051_golden_model_1.P2 [4], _40254_);
  dff (\oc8051_golden_model_1.P2 [5], _40255_);
  dff (\oc8051_golden_model_1.P2 [6], _40256_);
  dff (\oc8051_golden_model_1.P2 [7], _37147_);
  dff (\oc8051_golden_model_1.P3 [0], _40258_);
  dff (\oc8051_golden_model_1.P3 [1], _40259_);
  dff (\oc8051_golden_model_1.P3 [2], _40260_);
  dff (\oc8051_golden_model_1.P3 [3], _40261_);
  dff (\oc8051_golden_model_1.P3 [4], _40263_);
  dff (\oc8051_golden_model_1.P3 [5], _40264_);
  dff (\oc8051_golden_model_1.P3 [6], _40265_);
  dff (\oc8051_golden_model_1.P3 [7], _37148_);
  dff (\oc8051_golden_model_1.PSW [0], _40267_);
  dff (\oc8051_golden_model_1.PSW [1], _40268_);
  dff (\oc8051_golden_model_1.PSW [2], _40269_);
  dff (\oc8051_golden_model_1.PSW [3], _40270_);
  dff (\oc8051_golden_model_1.PSW [4], _40271_);
  dff (\oc8051_golden_model_1.PSW [5], _40272_);
  dff (\oc8051_golden_model_1.PSW [6], _40273_);
  dff (\oc8051_golden_model_1.PSW [7], _37149_);
  dff (\oc8051_golden_model_1.PCON [0], _40274_);
  dff (\oc8051_golden_model_1.PCON [1], _40275_);
  dff (\oc8051_golden_model_1.PCON [2], _40276_);
  dff (\oc8051_golden_model_1.PCON [3], _40277_);
  dff (\oc8051_golden_model_1.PCON [4], _40278_);
  dff (\oc8051_golden_model_1.PCON [5], _40279_);
  dff (\oc8051_golden_model_1.PCON [6], _40281_);
  dff (\oc8051_golden_model_1.PCON [7], _37150_);
  dff (\oc8051_golden_model_1.SBUF [0], _40282_);
  dff (\oc8051_golden_model_1.SBUF [1], _40283_);
  dff (\oc8051_golden_model_1.SBUF [2], _40285_);
  dff (\oc8051_golden_model_1.SBUF [3], _40286_);
  dff (\oc8051_golden_model_1.SBUF [4], _40287_);
  dff (\oc8051_golden_model_1.SBUF [5], _40288_);
  dff (\oc8051_golden_model_1.SBUF [6], _40289_);
  dff (\oc8051_golden_model_1.SBUF [7], _37151_);
  dff (\oc8051_golden_model_1.SCON [0], _40291_);
  dff (\oc8051_golden_model_1.SCON [1], _40292_);
  dff (\oc8051_golden_model_1.SCON [2], _40293_);
  dff (\oc8051_golden_model_1.SCON [3], _40294_);
  dff (\oc8051_golden_model_1.SCON [4], _40295_);
  dff (\oc8051_golden_model_1.SCON [5], _40296_);
  dff (\oc8051_golden_model_1.SCON [6], _40297_);
  dff (\oc8051_golden_model_1.SCON [7], _37152_);
  dff (\oc8051_golden_model_1.SP [0], _40299_);
  dff (\oc8051_golden_model_1.SP [1], _40300_);
  dff (\oc8051_golden_model_1.SP [2], _40301_);
  dff (\oc8051_golden_model_1.SP [3], _40302_);
  dff (\oc8051_golden_model_1.SP [4], _40304_);
  dff (\oc8051_golden_model_1.SP [5], _40305_);
  dff (\oc8051_golden_model_1.SP [6], _40306_);
  dff (\oc8051_golden_model_1.SP [7], _37153_);
  dff (\oc8051_golden_model_1.TCON [0], _40308_);
  dff (\oc8051_golden_model_1.TCON [1], _40309_);
  dff (\oc8051_golden_model_1.TCON [2], _40310_);
  dff (\oc8051_golden_model_1.TCON [3], _40311_);
  dff (\oc8051_golden_model_1.TCON [4], _40312_);
  dff (\oc8051_golden_model_1.TCON [5], _40313_);
  dff (\oc8051_golden_model_1.TCON [6], _40314_);
  dff (\oc8051_golden_model_1.TCON [7], _37154_);
  dff (\oc8051_golden_model_1.TH0 [0], _40316_);
  dff (\oc8051_golden_model_1.TH0 [1], _40317_);
  dff (\oc8051_golden_model_1.TH0 [2], _40318_);
  dff (\oc8051_golden_model_1.TH0 [3], _40319_);
  dff (\oc8051_golden_model_1.TH0 [4], _40320_);
  dff (\oc8051_golden_model_1.TH0 [5], _40321_);
  dff (\oc8051_golden_model_1.TH0 [6], _40323_);
  dff (\oc8051_golden_model_1.TH0 [7], _37156_);
  dff (\oc8051_golden_model_1.TH1 [0], _40324_);
  dff (\oc8051_golden_model_1.TH1 [1], _40325_);
  dff (\oc8051_golden_model_1.TH1 [2], _40326_);
  dff (\oc8051_golden_model_1.TH1 [3], _40327_);
  dff (\oc8051_golden_model_1.TH1 [4], _40328_);
  dff (\oc8051_golden_model_1.TH1 [5], _40329_);
  dff (\oc8051_golden_model_1.TH1 [6], _40330_);
  dff (\oc8051_golden_model_1.TH1 [7], _37157_);
  dff (\oc8051_golden_model_1.TL0 [0], _40332_);
  dff (\oc8051_golden_model_1.TL0 [1], _40333_);
  dff (\oc8051_golden_model_1.TL0 [2], _40334_);
  dff (\oc8051_golden_model_1.TL0 [3], _40335_);
  dff (\oc8051_golden_model_1.TL0 [4], _40336_);
  dff (\oc8051_golden_model_1.TL0 [5], _40337_);
  dff (\oc8051_golden_model_1.TL0 [6], _40338_);
  dff (\oc8051_golden_model_1.TL0 [7], _37158_);
  dff (\oc8051_golden_model_1.TL1 [0], _40340_);
  dff (\oc8051_golden_model_1.TL1 [1], _40341_);
  dff (\oc8051_golden_model_1.TL1 [2], _40342_);
  dff (\oc8051_golden_model_1.TL1 [3], _40343_);
  dff (\oc8051_golden_model_1.TL1 [4], _40345_);
  dff (\oc8051_golden_model_1.TL1 [5], _40346_);
  dff (\oc8051_golden_model_1.TL1 [6], _40347_);
  dff (\oc8051_golden_model_1.TL1 [7], _37159_);
  dff (\oc8051_golden_model_1.TMOD [0], _40349_);
  dff (\oc8051_golden_model_1.TMOD [1], _40350_);
  dff (\oc8051_golden_model_1.TMOD [2], _40351_);
  dff (\oc8051_golden_model_1.TMOD [3], _40352_);
  dff (\oc8051_golden_model_1.TMOD [4], _40353_);
  dff (\oc8051_golden_model_1.TMOD [5], _40354_);
  dff (\oc8051_golden_model_1.TMOD [6], _40355_);
  dff (\oc8051_golden_model_1.TMOD [7], _37160_);
  dff (\oc8051_golden_model_1.PC [0], _40358_);
  dff (\oc8051_golden_model_1.PC [1], _40359_);
  dff (\oc8051_golden_model_1.PC [2], _40360_);
  dff (\oc8051_golden_model_1.PC [3], _40361_);
  dff (\oc8051_golden_model_1.PC [4], _40362_);
  dff (\oc8051_golden_model_1.PC [5], _40363_);
  dff (\oc8051_golden_model_1.PC [6], _40364_);
  dff (\oc8051_golden_model_1.PC [7], _40365_);
  dff (\oc8051_golden_model_1.PC [8], _40367_);
  dff (\oc8051_golden_model_1.PC [9], _40368_);
  dff (\oc8051_golden_model_1.PC [10], _40369_);
  dff (\oc8051_golden_model_1.PC [11], _40370_);
  dff (\oc8051_golden_model_1.PC [12], _40371_);
  dff (\oc8051_golden_model_1.PC [13], _40372_);
  dff (\oc8051_golden_model_1.PC [14], _40373_);
  dff (\oc8051_golden_model_1.PC [15], _37162_);
  dff (\oc8051_golden_model_1.P0INREG [0], _40374_);
  dff (\oc8051_golden_model_1.P0INREG [1], _40375_);
  dff (\oc8051_golden_model_1.P0INREG [2], _40376_);
  dff (\oc8051_golden_model_1.P0INREG [3], _40377_);
  dff (\oc8051_golden_model_1.P0INREG [4], _40378_);
  dff (\oc8051_golden_model_1.P0INREG [5], _40379_);
  dff (\oc8051_golden_model_1.P0INREG [6], _40381_);
  dff (\oc8051_golden_model_1.P0INREG [7], _37163_);
  dff (\oc8051_golden_model_1.P1INREG [0], _40382_);
  dff (\oc8051_golden_model_1.P1INREG [1], _40383_);
  dff (\oc8051_golden_model_1.P1INREG [2], _40385_);
  dff (\oc8051_golden_model_1.P1INREG [3], _40386_);
  dff (\oc8051_golden_model_1.P1INREG [4], _40387_);
  dff (\oc8051_golden_model_1.P1INREG [5], _40388_);
  dff (\oc8051_golden_model_1.P1INREG [6], _40389_);
  dff (\oc8051_golden_model_1.P1INREG [7], _37164_);
  dff (\oc8051_golden_model_1.P2INREG [0], _40391_);
  dff (\oc8051_golden_model_1.P2INREG [1], _40392_);
  dff (\oc8051_golden_model_1.P2INREG [2], _40393_);
  dff (\oc8051_golden_model_1.P2INREG [3], _40394_);
  dff (\oc8051_golden_model_1.P2INREG [4], _40395_);
  dff (\oc8051_golden_model_1.P2INREG [5], _40396_);
  dff (\oc8051_golden_model_1.P2INREG [6], _40397_);
  dff (\oc8051_golden_model_1.P2INREG [7], _37165_);
  dff (\oc8051_golden_model_1.P3INREG [0], _40399_);
  dff (\oc8051_golden_model_1.P3INREG [1], _40400_);
  dff (\oc8051_golden_model_1.P3INREG [2], _40401_);
  dff (\oc8051_golden_model_1.P3INREG [3], _40402_);
  dff (\oc8051_golden_model_1.P3INREG [4], _40404_);
  dff (\oc8051_golden_model_1.P3INREG [5], _40405_);
  dff (\oc8051_golden_model_1.P3INREG [6], _40406_);
  dff (\oc8051_golden_model_1.P3INREG [7], _37166_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [0], _01043_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [1], _01046_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [2], _01049_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [3], _01051_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [4], _01054_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [5], _01057_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [6], _01060_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [7], _00914_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [0], _01063_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [1], _01066_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [2], _01069_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [3], _01072_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [4], _01075_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [5], _01078_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [6], _01081_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [7], _00918_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [0], _01084_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [1], _01087_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [2], _01090_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [3], _01093_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [4], _01095_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [5], _01098_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [6], _01101_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [7], _00922_);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [0], _35781_);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [1], _12280_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [0], _35782_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [1], _12283_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _35783_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _35784_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], _12285_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [0], _35785_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [1], _35786_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [2], _12288_);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [0], _35787_);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [1], _12291_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [0], _35788_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [1], _35789_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [2], _35790_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [3], _12293_);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [0], _35792_);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [1], _12296_);
  dff (\oc8051_top_1.oc8051_decoder1.wr , _12299_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], _12341_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], _12343_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], _12267_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [0], _12345_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [1], _12348_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [2], _12269_);
  dff (\oc8051_top_1.oc8051_decoder1.state [0], _12351_);
  dff (\oc8051_top_1.oc8051_decoder1.state [1], _12272_);
  dff (\oc8051_top_1.oc8051_decoder1.op [0], _12353_);
  dff (\oc8051_top_1.oc8051_decoder1.op [1], _12356_);
  dff (\oc8051_top_1.oc8051_decoder1.op [2], _12359_);
  dff (\oc8051_top_1.oc8051_decoder1.op [3], _12362_);
  dff (\oc8051_top_1.oc8051_decoder1.op [4], _12365_);
  dff (\oc8051_top_1.oc8051_decoder1.op [5], _12367_);
  dff (\oc8051_top_1.oc8051_decoder1.op [6], _12370_);
  dff (\oc8051_top_1.oc8051_decoder1.op [7], _12275_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel3 , _12277_);
  dff (\oc8051_top_1.oc8051_indi_addr1.wr_bit_r , _08208_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [0], _03635_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [1], _03637_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [2], _03639_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [3], _03641_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [4], _03643_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [5], _03645_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [6], _03647_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [7], _03649_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [8], _03651_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [9], _03653_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [10], _03655_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [11], _03657_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [12], _03659_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [13], _03661_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [14], _03663_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [15], _02779_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _03695_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _03697_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _03699_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _03701_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _03703_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _03705_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _03707_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _03709_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _03711_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _03713_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _03715_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _03717_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _03719_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _03721_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _03723_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _02783_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [0], _05595_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [1], _05597_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [2], _05599_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [3], _05601_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [4], _05603_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [5], _05605_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [6], _05607_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [7], _05609_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [8], _05611_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [9], _05613_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [10], _05615_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [11], _05617_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [12], _05619_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [13], _05621_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [14], _05623_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [15], _05625_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [16], _05627_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [17], _05629_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [18], _05631_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [19], _05633_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [20], _05635_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [21], _05637_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [22], _05639_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [23], _05641_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [24], _05643_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [25], _05645_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [26], _05647_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [27], _05649_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [28], _05651_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [29], _05653_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [30], _05655_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [31], _03232_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _03161_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dack_ir , 1'b0);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [0], _05658_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [1], _05661_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [2], _05664_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [3], _05666_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [4], _03168_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [0], _05669_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [1], _05672_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [2], _05675_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [3], _05678_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [4], _05681_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [5], _05684_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [6], _05687_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [7], _03172_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [0], _05689_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [1], _05691_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [2], _05693_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [3], _05695_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [4], _05697_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [5], _05699_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [6], _05701_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [7], _03175_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [0], _05703_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [1], _05705_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [2], _05707_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [3], _05709_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [4], _05711_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [5], _05713_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [6], _05715_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [7], _03178_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _03181_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _03185_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], _05717_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _05719_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], _05721_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], _05723_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _05725_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], _05727_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], _05729_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [7], _03188_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [0], _05731_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [1], _05733_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _05735_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [3], _05737_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [4], _05739_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [5], _05741_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [6], _05743_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [7], _05745_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [8], _05747_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [9], _05749_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [10], _05751_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [11], _05753_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [12], _05755_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [13], _05757_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [14], _05759_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [15], _03191_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [0], _05761_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [1], _05763_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [2], _05765_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [3], _05767_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [4], _05769_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [5], _05771_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [6], _05773_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [7], _05775_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [8], _05777_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [9], _05779_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [10], _05781_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [11], _05783_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [12], _05785_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [13], _05787_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [14], _05789_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [15], _03194_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack , _03199_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_t , _03205_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_buff , _03202_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], _05791_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], _05793_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _05795_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], _05797_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _05799_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], _05801_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _05803_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _03208_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [0], _05805_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [1], _05807_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [2], _03210_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [0], _05809_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [1], _05811_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [2], _05813_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [3], _05815_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [4], _05817_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [5], _05819_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [6], _05821_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [7], _03212_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [0], _05823_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [1], _05825_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [2], _05827_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [3], _05829_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [4], _05831_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [5], _05833_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [6], _05835_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [7], _03215_);
  dff (\oc8051_top_1.oc8051_memory_interface1.reti , _03218_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [0], _05837_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [1], _05839_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [2], _05841_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [3], _05843_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [4], _05845_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [5], _05847_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [6], _05849_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [7], _03220_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdone , _03223_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst , _03226_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], _05851_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], _05853_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], _05855_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], _03229_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [0], _05857_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [1], _05859_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [2], _05861_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [3], _05863_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [4], _05865_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [5], _05867_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [6], _05869_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [7], _05871_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [8], _05873_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [9], _05875_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [10], _05877_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [11], _05879_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [12], _05881_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [13], _05883_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [14], _05885_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [15], _05887_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [16], _05889_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [17], _05891_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [18], _05893_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [19], _05895_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [20], _05897_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [21], _05899_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [22], _05901_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [23], _05903_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [24], _05905_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [25], _05907_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [26], _05909_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [27], _05911_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [28], _05913_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [29], _05915_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [30], _05917_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [31], _03234_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [0], _05919_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [1], _05921_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [2], _05923_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [3], _05925_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [4], _05927_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [5], _05929_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [6], _05931_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [7], _03236_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dwe_o , _03238_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dstb_o , _03240_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [0], _05933_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [1], _05935_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [2], _05937_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [3], _05939_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [4], _05941_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [5], _05943_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [6], _05945_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [7], _05947_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [8], _05949_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [9], _05951_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [10], _05953_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [11], _05955_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [12], _05957_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [13], _05959_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [14], _05961_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [15], _03242_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dmem_wait , _03244_);
  dff (\oc8051_top_1.oc8051_memory_interface1.istb_t , _03246_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imem_wait , _03248_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _05963_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _05965_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _05967_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _05969_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [4], _05971_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [5], _05973_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [6], _05975_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [7], _05977_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [8], _05979_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [9], _05981_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [10], _05983_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [11], _05985_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [12], _05987_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [13], _05989_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [14], _05991_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [15], _03250_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_ind , _03252_);
  dff (\oc8051_top_1.oc8051_ram_top1.rd_en_r , _08305_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _08467_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _08469_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _08471_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _08473_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _08475_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _08477_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _08479_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [7], _08308_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_addr_r , _08311_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [0], _08481_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [1], _08483_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [2], _08314_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0], _39004_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1], _39008_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2], _39013_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3], _39019_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4], _39025_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5], _39031_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6], _39037_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7], _39040_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0], _39083_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1], _39087_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2], _39091_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3], _39095_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4], _39099_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5], _39103_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6], _39107_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7], _39110_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0], _39281_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1], _39285_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2], _39289_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3], _39293_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4], _39297_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5], _39301_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6], _39305_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7], _39308_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0], _39246_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1], _39250_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2], _39254_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3], _39258_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4], _39262_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5], _39266_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6], _39270_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7], _39273_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0], _39215_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1], _39219_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2], _39222_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3], _39226_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4], _39230_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5], _39234_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6], _39238_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7], _39241_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0], _39183_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1], _39187_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2], _39191_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3], _39195_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4], _39199_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5], _39203_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6], _39207_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7], _39210_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0], _39151_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1], _39155_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2], _39159_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3], _39163_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4], _39167_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5], _39171_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6], _39175_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7], _39178_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0], _39116_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1], _39120_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2], _39124_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3], _39128_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4], _39132_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5], _39136_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6], _39140_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7], _39143_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0], _39048_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1], _39052_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2], _39056_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3], _39060_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4], _39064_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5], _39068_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6], _39072_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7], _39075_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0], _39313_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1], _39317_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2], _39321_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3], _39325_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4], _39329_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5], _39333_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6], _39337_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7], _39340_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0], _39474_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1], _39478_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2], _39482_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3], _39486_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4], _39490_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5], _39494_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6], _39498_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7], _39501_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0], _39442_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1], _39446_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2], _39450_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3], _39454_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4], _39458_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5], _39462_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6], _39466_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7], _39469_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0], _39410_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1], _39414_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2], _39418_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3], _39422_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4], _39426_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5], _39430_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6], _39434_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7], _39437_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0], _39377_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1], _39381_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2], _39385_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3], _39389_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4], _39393_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5], _39397_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6], _39401_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7], _39404_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0], _39345_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1], _39349_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2], _39353_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3], _39357_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4], _39361_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5], _39365_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6], _39369_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7], _39372_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0], _39506_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1], _39510_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2], _39514_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3], _39518_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4], _39522_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5], _39526_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6], _39530_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7], _38724_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0], _00042_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1], _00044_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2], _00046_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3], _00048_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4], _00050_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5], _00052_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6], _00054_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7], _38712_);
  dff (\oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  dff (\oc8051_top_1.oc8051_rom1.ea_int , 1'b1);
  dff (\oc8051_top_1.oc8051_sfr1.bit_out , _01521_);
  dff (\oc8051_top_1.oc8051_sfr1.wait_data , _01523_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [0], _02204_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [1], _02206_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [2], _02208_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [3], _02210_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [4], _02212_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [5], _02214_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [6], _02216_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [7], _01525_);
  dff (\oc8051_top_1.oc8051_sfr1.wr_bit_r , _01528_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], _08869_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], _08880_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], _08891_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3], _08902_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4], _08913_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], _08924_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], _08935_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], _07163_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0], _29076_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1], _29184_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2], _29294_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3], _29403_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4], _29511_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5], _29620_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6], _29730_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7], _05323_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], _39759_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], _39767_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], _39776_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], _39785_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], _39793_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], _39802_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], _39810_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7], _38754_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0], _39819_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1], _39827_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2], _39836_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3], _39844_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4], _39853_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5], _39861_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6], _39870_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7], _38774_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff , 1'b0);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff , 1'b0);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff , 1'b0);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie1_buff , _37580_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], _38571_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], _38573_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _38575_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3], _38577_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4], _38579_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], _38581_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _38583_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _37547_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], _38585_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _37582_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc , _37549_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _38587_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _38589_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], _37584_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _38591_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _38593_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], _37551_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], _38595_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [1], _37586_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _38597_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [1], _37588_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , _37571_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , _37573_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , _37575_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , _37576_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0], _38599_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1], _38601_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2], _38603_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], _37578_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0], _38605_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], _38607_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], _38609_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3], _38611_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4], _38613_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5], _38615_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6], _38617_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _37492_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0], _38619_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1], _38621_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2], _38623_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3], _38625_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4], _38626_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5], _38628_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6], _38630_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7], _37528_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0], _36859_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1], _36861_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2], _36863_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3], _36865_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4], _36867_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5], _36869_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6], _36871_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7], _19317_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0], _36873_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1], _36875_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2], _36877_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3], _36879_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4], _36881_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5], _36883_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6], _36885_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7], _19339_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0], _36887_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1], _36888_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2], _36890_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3], _36892_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4], _36894_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5], _36896_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6], _36898_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7], _19362_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0], _36900_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1], _36902_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2], _36904_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3], _36906_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4], _36908_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5], _36910_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6], _36912_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7], _19385_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1], _06388_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], _06399_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3], _06409_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4], _06420_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5], _06431_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6], _06442_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], _01571_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], _36625_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], _36633_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2], _36641_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3], _36649_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4], _36657_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5], _36665_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6], _36672_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7], _35441_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop , _35258_);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.bit_in , ABINPUT[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_in [0], ABINPUT[19]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_in [1], ABINPUT[20]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_in [2], ABINPUT[21]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_in [3], ABINPUT[22]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_in [4], ABINPUT[23]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_in [5], ABINPUT[24]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_in [6], ABINPUT[25]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_in [7], ABINPUT[26]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.data_in [0], ABINPUT[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.data_in [1], ABINPUT[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.data_in [2], ABINPUT[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.data_in [3], ABINPUT[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.data_in [4], ABINPUT[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.data_in [5], ABINPUT[8]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.data_in [6], ABINPUT[9]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.data_in [7], ABINPUT[10]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_in [0], ABINPUT[19]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_in [1], ABINPUT[20]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_in [2], ABINPUT[21]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_in [3], ABINPUT[22]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_in [4], ABINPUT[23]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_in [5], ABINPUT[24]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_in [6], ABINPUT[25]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_in [7], ABINPUT[26]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data2_in [0], ABINPUT[11]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data2_in [1], ABINPUT[12]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data2_in [2], ABINPUT[13]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data2_in [3], ABINPUT[14]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data2_in [4], ABINPUT[15]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data2_in [5], ABINPUT[16]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data2_in [6], ABINPUT[17]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data2_in [7], ABINPUT[18]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.cy_in , ABINPUT[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.ac_in , ABINPUT[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.ov_in , ABINPUT[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_in [0], ABINPUT[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_in [1], ABINPUT[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_in [2], ABINPUT[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_in [3], ABINPUT[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_in [4], ABINPUT[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_in [5], ABINPUT[8]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_in [6], ABINPUT[9]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_in [7], ABINPUT[10]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [0], psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [0], psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [1], \oc8051_top_1.oc8051_sfr1.psw_next [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [2], \oc8051_top_1.oc8051_sfr1.psw_next [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [3], \oc8051_top_1.oc8051_sfr1.psw_next [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [4], \oc8051_top_1.oc8051_sfr1.psw_next [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [5], \oc8051_top_1.oc8051_sfr1.psw_next [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [6], \oc8051_top_1.oc8051_sfr1.psw_next [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [7], \oc8051_top_1.oc8051_sfr1.psw_next [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [1], \oc8051_top_1.oc8051_sfr1.psw_next [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [2], \oc8051_top_1.oc8051_sfr1.psw_next [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [3], \oc8051_top_1.oc8051_sfr1.psw_next [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [4], \oc8051_top_1.oc8051_sfr1.psw_next [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [5], \oc8051_top_1.oc8051_sfr1.psw_next [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [6], \oc8051_top_1.oc8051_sfr1.psw_next [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [7], \oc8051_top_1.oc8051_sfr1.psw_next [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.bit_in , ABINPUT[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_in [0], ABINPUT[19]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_in [1], ABINPUT[20]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_in [2], ABINPUT[21]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_in [3], ABINPUT[22]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_in [4], ABINPUT[23]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_in [5], ABINPUT[24]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_in [6], ABINPUT[25]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_in [7], ABINPUT[26]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data2_in [0], ABINPUT[11]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data2_in [1], ABINPUT[12]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data2_in [2], ABINPUT[13]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data2_in [3], ABINPUT[14]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data2_in [4], ABINPUT[15]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data2_in [5], ABINPUT[16]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data2_in [6], ABINPUT[17]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data2_in [7], ABINPUT[18]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.p , psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.bit_in , ABINPUT[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.data_in [0], ABINPUT[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.data_in [1], ABINPUT[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.data_in [2], ABINPUT[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.data_in [3], ABINPUT[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.data_in [4], ABINPUT[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.data_in [5], ABINPUT[8]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.data_in [6], ABINPUT[9]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.data_in [7], ABINPUT[10]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.data_in [0], ABINPUT[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.data_in [1], ABINPUT[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.data_in [2], ABINPUT[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.data_in [3], ABINPUT[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.data_in [4], ABINPUT[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.data_in [5], ABINPUT[8]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.data_in [6], ABINPUT[9]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.data_in [7], ABINPUT[10]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.bit_in , ABINPUT[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [4], 1'b0);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [5], 1'b0);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell0.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell0.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell0.word [0], word_in[0]);
  buf(\oc8051_gm_cxrom_1.cell0.word [1], word_in[1]);
  buf(\oc8051_gm_cxrom_1.cell0.word [2], word_in[2]);
  buf(\oc8051_gm_cxrom_1.cell0.word [3], word_in[3]);
  buf(\oc8051_gm_cxrom_1.cell0.word [4], word_in[4]);
  buf(\oc8051_gm_cxrom_1.cell0.word [5], word_in[5]);
  buf(\oc8051_gm_cxrom_1.cell0.word [6], word_in[6]);
  buf(\oc8051_gm_cxrom_1.cell0.word [7], word_in[7]);
  buf(\oc8051_gm_cxrom_1.cell1.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell1.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell1.word [0], word_in[8]);
  buf(\oc8051_gm_cxrom_1.cell1.word [1], word_in[9]);
  buf(\oc8051_gm_cxrom_1.cell1.word [2], word_in[10]);
  buf(\oc8051_gm_cxrom_1.cell1.word [3], word_in[11]);
  buf(\oc8051_gm_cxrom_1.cell1.word [4], word_in[12]);
  buf(\oc8051_gm_cxrom_1.cell1.word [5], word_in[13]);
  buf(\oc8051_gm_cxrom_1.cell1.word [6], word_in[14]);
  buf(\oc8051_gm_cxrom_1.cell1.word [7], word_in[15]);
  buf(\oc8051_gm_cxrom_1.cell2.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell2.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell2.word [0], word_in[16]);
  buf(\oc8051_gm_cxrom_1.cell2.word [1], word_in[17]);
  buf(\oc8051_gm_cxrom_1.cell2.word [2], word_in[18]);
  buf(\oc8051_gm_cxrom_1.cell2.word [3], word_in[19]);
  buf(\oc8051_gm_cxrom_1.cell2.word [4], word_in[20]);
  buf(\oc8051_gm_cxrom_1.cell2.word [5], word_in[21]);
  buf(\oc8051_gm_cxrom_1.cell2.word [6], word_in[22]);
  buf(\oc8051_gm_cxrom_1.cell2.word [7], word_in[23]);
  buf(\oc8051_gm_cxrom_1.cell3.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell3.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell3.word [0], word_in[24]);
  buf(\oc8051_gm_cxrom_1.cell3.word [1], word_in[25]);
  buf(\oc8051_gm_cxrom_1.cell3.word [2], word_in[26]);
  buf(\oc8051_gm_cxrom_1.cell3.word [3], word_in[27]);
  buf(\oc8051_gm_cxrom_1.cell3.word [4], word_in[28]);
  buf(\oc8051_gm_cxrom_1.cell3.word [5], word_in[29]);
  buf(\oc8051_gm_cxrom_1.cell3.word [6], word_in[30]);
  buf(\oc8051_gm_cxrom_1.cell3.word [7], word_in[31]);
  buf(\oc8051_gm_cxrom_1.cell4.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell4.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell4.word [0], word_in[32]);
  buf(\oc8051_gm_cxrom_1.cell4.word [1], word_in[33]);
  buf(\oc8051_gm_cxrom_1.cell4.word [2], word_in[34]);
  buf(\oc8051_gm_cxrom_1.cell4.word [3], word_in[35]);
  buf(\oc8051_gm_cxrom_1.cell4.word [4], word_in[36]);
  buf(\oc8051_gm_cxrom_1.cell4.word [5], word_in[37]);
  buf(\oc8051_gm_cxrom_1.cell4.word [6], word_in[38]);
  buf(\oc8051_gm_cxrom_1.cell4.word [7], word_in[39]);
  buf(\oc8051_gm_cxrom_1.cell5.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell5.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell5.word [0], word_in[40]);
  buf(\oc8051_gm_cxrom_1.cell5.word [1], word_in[41]);
  buf(\oc8051_gm_cxrom_1.cell5.word [2], word_in[42]);
  buf(\oc8051_gm_cxrom_1.cell5.word [3], word_in[43]);
  buf(\oc8051_gm_cxrom_1.cell5.word [4], word_in[44]);
  buf(\oc8051_gm_cxrom_1.cell5.word [5], word_in[45]);
  buf(\oc8051_gm_cxrom_1.cell5.word [6], word_in[46]);
  buf(\oc8051_gm_cxrom_1.cell5.word [7], word_in[47]);
  buf(\oc8051_gm_cxrom_1.cell6.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell6.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell6.word [0], word_in[48]);
  buf(\oc8051_gm_cxrom_1.cell6.word [1], word_in[49]);
  buf(\oc8051_gm_cxrom_1.cell6.word [2], word_in[50]);
  buf(\oc8051_gm_cxrom_1.cell6.word [3], word_in[51]);
  buf(\oc8051_gm_cxrom_1.cell6.word [4], word_in[52]);
  buf(\oc8051_gm_cxrom_1.cell6.word [5], word_in[53]);
  buf(\oc8051_gm_cxrom_1.cell6.word [6], word_in[54]);
  buf(\oc8051_gm_cxrom_1.cell6.word [7], word_in[55]);
  buf(\oc8051_gm_cxrom_1.cell7.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell7.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell7.word [0], word_in[56]);
  buf(\oc8051_gm_cxrom_1.cell7.word [1], word_in[57]);
  buf(\oc8051_gm_cxrom_1.cell7.word [2], word_in[58]);
  buf(\oc8051_gm_cxrom_1.cell7.word [3], word_in[59]);
  buf(\oc8051_gm_cxrom_1.cell7.word [4], word_in[60]);
  buf(\oc8051_gm_cxrom_1.cell7.word [5], word_in[61]);
  buf(\oc8051_gm_cxrom_1.cell7.word [6], word_in[62]);
  buf(\oc8051_gm_cxrom_1.cell7.word [7], word_in[63]);
  buf(\oc8051_gm_cxrom_1.cell8.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell8.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell8.word [0], word_in[64]);
  buf(\oc8051_gm_cxrom_1.cell8.word [1], word_in[65]);
  buf(\oc8051_gm_cxrom_1.cell8.word [2], word_in[66]);
  buf(\oc8051_gm_cxrom_1.cell8.word [3], word_in[67]);
  buf(\oc8051_gm_cxrom_1.cell8.word [4], word_in[68]);
  buf(\oc8051_gm_cxrom_1.cell8.word [5], word_in[69]);
  buf(\oc8051_gm_cxrom_1.cell8.word [6], word_in[70]);
  buf(\oc8051_gm_cxrom_1.cell8.word [7], word_in[71]);
  buf(\oc8051_gm_cxrom_1.cell9.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell9.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell9.word [0], word_in[72]);
  buf(\oc8051_gm_cxrom_1.cell9.word [1], word_in[73]);
  buf(\oc8051_gm_cxrom_1.cell9.word [2], word_in[74]);
  buf(\oc8051_gm_cxrom_1.cell9.word [3], word_in[75]);
  buf(\oc8051_gm_cxrom_1.cell9.word [4], word_in[76]);
  buf(\oc8051_gm_cxrom_1.cell9.word [5], word_in[77]);
  buf(\oc8051_gm_cxrom_1.cell9.word [6], word_in[78]);
  buf(\oc8051_gm_cxrom_1.cell9.word [7], word_in[79]);
  buf(\oc8051_gm_cxrom_1.cell10.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell10.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell10.word [0], word_in[80]);
  buf(\oc8051_gm_cxrom_1.cell10.word [1], word_in[81]);
  buf(\oc8051_gm_cxrom_1.cell10.word [2], word_in[82]);
  buf(\oc8051_gm_cxrom_1.cell10.word [3], word_in[83]);
  buf(\oc8051_gm_cxrom_1.cell10.word [4], word_in[84]);
  buf(\oc8051_gm_cxrom_1.cell10.word [5], word_in[85]);
  buf(\oc8051_gm_cxrom_1.cell10.word [6], word_in[86]);
  buf(\oc8051_gm_cxrom_1.cell10.word [7], word_in[87]);
  buf(\oc8051_gm_cxrom_1.cell11.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell11.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell11.word [0], word_in[88]);
  buf(\oc8051_gm_cxrom_1.cell11.word [1], word_in[89]);
  buf(\oc8051_gm_cxrom_1.cell11.word [2], word_in[90]);
  buf(\oc8051_gm_cxrom_1.cell11.word [3], word_in[91]);
  buf(\oc8051_gm_cxrom_1.cell11.word [4], word_in[92]);
  buf(\oc8051_gm_cxrom_1.cell11.word [5], word_in[93]);
  buf(\oc8051_gm_cxrom_1.cell11.word [6], word_in[94]);
  buf(\oc8051_gm_cxrom_1.cell11.word [7], word_in[95]);
  buf(\oc8051_gm_cxrom_1.cell12.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell12.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell12.word [0], word_in[96]);
  buf(\oc8051_gm_cxrom_1.cell12.word [1], word_in[97]);
  buf(\oc8051_gm_cxrom_1.cell12.word [2], word_in[98]);
  buf(\oc8051_gm_cxrom_1.cell12.word [3], word_in[99]);
  buf(\oc8051_gm_cxrom_1.cell12.word [4], word_in[100]);
  buf(\oc8051_gm_cxrom_1.cell12.word [5], word_in[101]);
  buf(\oc8051_gm_cxrom_1.cell12.word [6], word_in[102]);
  buf(\oc8051_gm_cxrom_1.cell12.word [7], word_in[103]);
  buf(\oc8051_gm_cxrom_1.cell13.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell13.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell13.word [0], word_in[104]);
  buf(\oc8051_gm_cxrom_1.cell13.word [1], word_in[105]);
  buf(\oc8051_gm_cxrom_1.cell13.word [2], word_in[106]);
  buf(\oc8051_gm_cxrom_1.cell13.word [3], word_in[107]);
  buf(\oc8051_gm_cxrom_1.cell13.word [4], word_in[108]);
  buf(\oc8051_gm_cxrom_1.cell13.word [5], word_in[109]);
  buf(\oc8051_gm_cxrom_1.cell13.word [6], word_in[110]);
  buf(\oc8051_gm_cxrom_1.cell13.word [7], word_in[111]);
  buf(\oc8051_gm_cxrom_1.cell14.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell14.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell14.word [0], word_in[112]);
  buf(\oc8051_gm_cxrom_1.cell14.word [1], word_in[113]);
  buf(\oc8051_gm_cxrom_1.cell14.word [2], word_in[114]);
  buf(\oc8051_gm_cxrom_1.cell14.word [3], word_in[115]);
  buf(\oc8051_gm_cxrom_1.cell14.word [4], word_in[116]);
  buf(\oc8051_gm_cxrom_1.cell14.word [5], word_in[117]);
  buf(\oc8051_gm_cxrom_1.cell14.word [6], word_in[118]);
  buf(\oc8051_gm_cxrom_1.cell14.word [7], word_in[119]);
  buf(\oc8051_gm_cxrom_1.cell15.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell15.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell15.word [0], word_in[120]);
  buf(\oc8051_gm_cxrom_1.cell15.word [1], word_in[121]);
  buf(\oc8051_gm_cxrom_1.cell15.word [2], word_in[122]);
  buf(\oc8051_gm_cxrom_1.cell15.word [3], word_in[123]);
  buf(\oc8051_gm_cxrom_1.cell15.word [4], word_in[124]);
  buf(\oc8051_gm_cxrom_1.cell15.word [5], word_in[125]);
  buf(\oc8051_gm_cxrom_1.cell15.word [6], word_in[126]);
  buf(\oc8051_gm_cxrom_1.cell15.word [7], word_in[127]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_in , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.bit_in , ABINPUT[0]);
  buf(\oc8051_top_1.oc8051_sfr1.desAc , ABINPUT[1]);
  buf(\oc8051_top_1.oc8051_sfr1.desOv , ABINPUT[2]);
  buf(\oc8051_top_1.oc8051_sfr1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.des_acc [0], ABINPUT[19]);
  buf(\oc8051_top_1.oc8051_sfr1.des_acc [1], ABINPUT[20]);
  buf(\oc8051_top_1.oc8051_sfr1.des_acc [2], ABINPUT[21]);
  buf(\oc8051_top_1.oc8051_sfr1.des_acc [3], ABINPUT[22]);
  buf(\oc8051_top_1.oc8051_sfr1.des_acc [4], ABINPUT[23]);
  buf(\oc8051_top_1.oc8051_sfr1.des_acc [5], ABINPUT[24]);
  buf(\oc8051_top_1.oc8051_sfr1.des_acc [6], ABINPUT[25]);
  buf(\oc8051_top_1.oc8051_sfr1.des_acc [7], ABINPUT[26]);
  buf(\oc8051_top_1.oc8051_sfr1.dat1 [0], ABINPUT[3]);
  buf(\oc8051_top_1.oc8051_sfr1.dat1 [1], ABINPUT[4]);
  buf(\oc8051_top_1.oc8051_sfr1.dat1 [2], ABINPUT[5]);
  buf(\oc8051_top_1.oc8051_sfr1.dat1 [3], ABINPUT[6]);
  buf(\oc8051_top_1.oc8051_sfr1.dat1 [4], ABINPUT[7]);
  buf(\oc8051_top_1.oc8051_sfr1.dat1 [5], ABINPUT[8]);
  buf(\oc8051_top_1.oc8051_sfr1.dat1 [6], ABINPUT[9]);
  buf(\oc8051_top_1.oc8051_sfr1.dat1 [7], ABINPUT[10]);
  buf(\oc8051_top_1.oc8051_sfr1.dat2 [0], ABINPUT[11]);
  buf(\oc8051_top_1.oc8051_sfr1.dat2 [1], ABINPUT[12]);
  buf(\oc8051_top_1.oc8051_sfr1.dat2 [2], ABINPUT[13]);
  buf(\oc8051_top_1.oc8051_sfr1.dat2 [3], ABINPUT[14]);
  buf(\oc8051_top_1.oc8051_sfr1.dat2 [4], ABINPUT[15]);
  buf(\oc8051_top_1.oc8051_sfr1.dat2 [5], ABINPUT[16]);
  buf(\oc8051_top_1.oc8051_sfr1.dat2 [6], ABINPUT[17]);
  buf(\oc8051_top_1.oc8051_sfr1.dat2 [7], ABINPUT[18]);
  buf(\oc8051_top_1.oc8051_sfr1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [0], psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p , psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.ip [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_next [0], psw_impl[0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.rst , rst);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.wr_dat [0], ABINPUT[3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.wr_dat [1], ABINPUT[4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.wr_dat [2], ABINPUT[5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.wr_dat [3], ABINPUT[6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.wr_dat [4], ABINPUT[7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.wr_dat [5], ABINPUT[8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.wr_dat [6], ABINPUT[9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.wr_dat [7], ABINPUT[10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des_acc [0], ABINPUT[19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des_acc [1], ABINPUT[20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des_acc [2], ABINPUT[21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des_acc [3], ABINPUT[22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des_acc [4], ABINPUT[23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des_acc [5], ABINPUT[24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des_acc [6], ABINPUT[25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des_acc [7], ABINPUT[26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des1 [0], ABINPUT[3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des1 [1], ABINPUT[4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des1 [2], ABINPUT[5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des1 [3], ABINPUT[6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des1 [4], ABINPUT[7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des1 [5], ABINPUT[8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des1 [6], ABINPUT[9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des1 [7], ABINPUT[10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des2 [0], ABINPUT[11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des2 [1], ABINPUT[12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des2 [2], ABINPUT[13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des2 [3], ABINPUT[14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des2 [4], ABINPUT[15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des2 [5], ABINPUT[16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des2 [6], ABINPUT[17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des2 [7], ABINPUT[18]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [0], ABINPUT[19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [1], ABINPUT[20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [2], ABINPUT[21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [3], ABINPUT[22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [4], ABINPUT[23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [5], ABINPUT[24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [6], ABINPUT[25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [7], ABINPUT[26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [8], ABINPUT[11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [9], ABINPUT[12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [10], ABINPUT[13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [11], ABINPUT[14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [12], ABINPUT[15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [13], ABINPUT[16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [14], ABINPUT[17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [15], ABINPUT[18]);
  buf(\oc8051_top_1.oc8051_rom1.rst , rst);
  buf(\oc8051_top_1.oc8051_rom1.clk , clk);
  buf(\oc8051_top_1.oc8051_indi_addr1.clk , clk);
  buf(\oc8051_top_1.oc8051_indi_addr1.rst , rst);
  buf(\oc8051_top_1.oc8051_indi_addr1.data_in [0], ABINPUT[3]);
  buf(\oc8051_top_1.oc8051_indi_addr1.data_in [1], ABINPUT[4]);
  buf(\oc8051_top_1.oc8051_indi_addr1.data_in [2], ABINPUT[5]);
  buf(\oc8051_top_1.oc8051_indi_addr1.data_in [3], ABINPUT[6]);
  buf(\oc8051_top_1.oc8051_indi_addr1.data_in [4], ABINPUT[7]);
  buf(\oc8051_top_1.oc8051_indi_addr1.data_in [5], ABINPUT[8]);
  buf(\oc8051_top_1.oc8051_indi_addr1.data_in [6], ABINPUT[9]);
  buf(\oc8051_top_1.oc8051_indi_addr1.data_in [7], ABINPUT[10]);
  buf(\oc8051_top_1.oc8051_ram_top1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.bit_data_in , ABINPUT[0]);
  buf(\oc8051_top_1.oc8051_ram_top1.rst , rst);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_data [0], ABINPUT[3]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_data [1], ABINPUT[4]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_data [2], ABINPUT[5]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_data [3], ABINPUT[6]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_data [4], ABINPUT[7]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_data [5], ABINPUT[8]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_data [6], ABINPUT[9]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_data [7], ABINPUT[10]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  buf(\oc8051_top_1.oc8051_decoder1.clk , clk);
  buf(\oc8051_top_1.oc8051_decoder1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.oc8051_decoder1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.oc8051_comp1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_comp1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_comp1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_comp1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_comp1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_comp1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_comp1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_comp1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_comp1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_comp1.des [0], ABINPUT[27]);
  buf(\oc8051_top_1.oc8051_comp1.des [1], ABINPUT[28]);
  buf(\oc8051_top_1.oc8051_comp1.des [2], ABINPUT[29]);
  buf(\oc8051_top_1.oc8051_comp1.des [3], ABINPUT[30]);
  buf(\oc8051_top_1.oc8051_comp1.des [4], ABINPUT[31]);
  buf(\oc8051_top_1.oc8051_comp1.des [5], ABINPUT[32]);
  buf(\oc8051_top_1.oc8051_comp1.des [6], ABINPUT[33]);
  buf(\oc8051_top_1.oc8051_comp1.des [7], ABINPUT[34]);
  buf(\oc8051_gm_cxrom_1.clk , clk);
  buf(\oc8051_gm_cxrom_1.rst , rst);
  buf(\oc8051_gm_cxrom_1.word_in [0], word_in[0]);
  buf(\oc8051_gm_cxrom_1.word_in [1], word_in[1]);
  buf(\oc8051_gm_cxrom_1.word_in [2], word_in[2]);
  buf(\oc8051_gm_cxrom_1.word_in [3], word_in[3]);
  buf(\oc8051_gm_cxrom_1.word_in [4], word_in[4]);
  buf(\oc8051_gm_cxrom_1.word_in [5], word_in[5]);
  buf(\oc8051_gm_cxrom_1.word_in [6], word_in[6]);
  buf(\oc8051_gm_cxrom_1.word_in [7], word_in[7]);
  buf(\oc8051_gm_cxrom_1.word_in [8], word_in[8]);
  buf(\oc8051_gm_cxrom_1.word_in [9], word_in[9]);
  buf(\oc8051_gm_cxrom_1.word_in [10], word_in[10]);
  buf(\oc8051_gm_cxrom_1.word_in [11], word_in[11]);
  buf(\oc8051_gm_cxrom_1.word_in [12], word_in[12]);
  buf(\oc8051_gm_cxrom_1.word_in [13], word_in[13]);
  buf(\oc8051_gm_cxrom_1.word_in [14], word_in[14]);
  buf(\oc8051_gm_cxrom_1.word_in [15], word_in[15]);
  buf(\oc8051_gm_cxrom_1.word_in [16], word_in[16]);
  buf(\oc8051_gm_cxrom_1.word_in [17], word_in[17]);
  buf(\oc8051_gm_cxrom_1.word_in [18], word_in[18]);
  buf(\oc8051_gm_cxrom_1.word_in [19], word_in[19]);
  buf(\oc8051_gm_cxrom_1.word_in [20], word_in[20]);
  buf(\oc8051_gm_cxrom_1.word_in [21], word_in[21]);
  buf(\oc8051_gm_cxrom_1.word_in [22], word_in[22]);
  buf(\oc8051_gm_cxrom_1.word_in [23], word_in[23]);
  buf(\oc8051_gm_cxrom_1.word_in [24], word_in[24]);
  buf(\oc8051_gm_cxrom_1.word_in [25], word_in[25]);
  buf(\oc8051_gm_cxrom_1.word_in [26], word_in[26]);
  buf(\oc8051_gm_cxrom_1.word_in [27], word_in[27]);
  buf(\oc8051_gm_cxrom_1.word_in [28], word_in[28]);
  buf(\oc8051_gm_cxrom_1.word_in [29], word_in[29]);
  buf(\oc8051_gm_cxrom_1.word_in [30], word_in[30]);
  buf(\oc8051_gm_cxrom_1.word_in [31], word_in[31]);
  buf(\oc8051_gm_cxrom_1.word_in [32], word_in[32]);
  buf(\oc8051_gm_cxrom_1.word_in [33], word_in[33]);
  buf(\oc8051_gm_cxrom_1.word_in [34], word_in[34]);
  buf(\oc8051_gm_cxrom_1.word_in [35], word_in[35]);
  buf(\oc8051_gm_cxrom_1.word_in [36], word_in[36]);
  buf(\oc8051_gm_cxrom_1.word_in [37], word_in[37]);
  buf(\oc8051_gm_cxrom_1.word_in [38], word_in[38]);
  buf(\oc8051_gm_cxrom_1.word_in [39], word_in[39]);
  buf(\oc8051_gm_cxrom_1.word_in [40], word_in[40]);
  buf(\oc8051_gm_cxrom_1.word_in [41], word_in[41]);
  buf(\oc8051_gm_cxrom_1.word_in [42], word_in[42]);
  buf(\oc8051_gm_cxrom_1.word_in [43], word_in[43]);
  buf(\oc8051_gm_cxrom_1.word_in [44], word_in[44]);
  buf(\oc8051_gm_cxrom_1.word_in [45], word_in[45]);
  buf(\oc8051_gm_cxrom_1.word_in [46], word_in[46]);
  buf(\oc8051_gm_cxrom_1.word_in [47], word_in[47]);
  buf(\oc8051_gm_cxrom_1.word_in [48], word_in[48]);
  buf(\oc8051_gm_cxrom_1.word_in [49], word_in[49]);
  buf(\oc8051_gm_cxrom_1.word_in [50], word_in[50]);
  buf(\oc8051_gm_cxrom_1.word_in [51], word_in[51]);
  buf(\oc8051_gm_cxrom_1.word_in [52], word_in[52]);
  buf(\oc8051_gm_cxrom_1.word_in [53], word_in[53]);
  buf(\oc8051_gm_cxrom_1.word_in [54], word_in[54]);
  buf(\oc8051_gm_cxrom_1.word_in [55], word_in[55]);
  buf(\oc8051_gm_cxrom_1.word_in [56], word_in[56]);
  buf(\oc8051_gm_cxrom_1.word_in [57], word_in[57]);
  buf(\oc8051_gm_cxrom_1.word_in [58], word_in[58]);
  buf(\oc8051_gm_cxrom_1.word_in [59], word_in[59]);
  buf(\oc8051_gm_cxrom_1.word_in [60], word_in[60]);
  buf(\oc8051_gm_cxrom_1.word_in [61], word_in[61]);
  buf(\oc8051_gm_cxrom_1.word_in [62], word_in[62]);
  buf(\oc8051_gm_cxrom_1.word_in [63], word_in[63]);
  buf(\oc8051_gm_cxrom_1.word_in [64], word_in[64]);
  buf(\oc8051_gm_cxrom_1.word_in [65], word_in[65]);
  buf(\oc8051_gm_cxrom_1.word_in [66], word_in[66]);
  buf(\oc8051_gm_cxrom_1.word_in [67], word_in[67]);
  buf(\oc8051_gm_cxrom_1.word_in [68], word_in[68]);
  buf(\oc8051_gm_cxrom_1.word_in [69], word_in[69]);
  buf(\oc8051_gm_cxrom_1.word_in [70], word_in[70]);
  buf(\oc8051_gm_cxrom_1.word_in [71], word_in[71]);
  buf(\oc8051_gm_cxrom_1.word_in [72], word_in[72]);
  buf(\oc8051_gm_cxrom_1.word_in [73], word_in[73]);
  buf(\oc8051_gm_cxrom_1.word_in [74], word_in[74]);
  buf(\oc8051_gm_cxrom_1.word_in [75], word_in[75]);
  buf(\oc8051_gm_cxrom_1.word_in [76], word_in[76]);
  buf(\oc8051_gm_cxrom_1.word_in [77], word_in[77]);
  buf(\oc8051_gm_cxrom_1.word_in [78], word_in[78]);
  buf(\oc8051_gm_cxrom_1.word_in [79], word_in[79]);
  buf(\oc8051_gm_cxrom_1.word_in [80], word_in[80]);
  buf(\oc8051_gm_cxrom_1.word_in [81], word_in[81]);
  buf(\oc8051_gm_cxrom_1.word_in [82], word_in[82]);
  buf(\oc8051_gm_cxrom_1.word_in [83], word_in[83]);
  buf(\oc8051_gm_cxrom_1.word_in [84], word_in[84]);
  buf(\oc8051_gm_cxrom_1.word_in [85], word_in[85]);
  buf(\oc8051_gm_cxrom_1.word_in [86], word_in[86]);
  buf(\oc8051_gm_cxrom_1.word_in [87], word_in[87]);
  buf(\oc8051_gm_cxrom_1.word_in [88], word_in[88]);
  buf(\oc8051_gm_cxrom_1.word_in [89], word_in[89]);
  buf(\oc8051_gm_cxrom_1.word_in [90], word_in[90]);
  buf(\oc8051_gm_cxrom_1.word_in [91], word_in[91]);
  buf(\oc8051_gm_cxrom_1.word_in [92], word_in[92]);
  buf(\oc8051_gm_cxrom_1.word_in [93], word_in[93]);
  buf(\oc8051_gm_cxrom_1.word_in [94], word_in[94]);
  buf(\oc8051_gm_cxrom_1.word_in [95], word_in[95]);
  buf(\oc8051_gm_cxrom_1.word_in [96], word_in[96]);
  buf(\oc8051_gm_cxrom_1.word_in [97], word_in[97]);
  buf(\oc8051_gm_cxrom_1.word_in [98], word_in[98]);
  buf(\oc8051_gm_cxrom_1.word_in [99], word_in[99]);
  buf(\oc8051_gm_cxrom_1.word_in [100], word_in[100]);
  buf(\oc8051_gm_cxrom_1.word_in [101], word_in[101]);
  buf(\oc8051_gm_cxrom_1.word_in [102], word_in[102]);
  buf(\oc8051_gm_cxrom_1.word_in [103], word_in[103]);
  buf(\oc8051_gm_cxrom_1.word_in [104], word_in[104]);
  buf(\oc8051_gm_cxrom_1.word_in [105], word_in[105]);
  buf(\oc8051_gm_cxrom_1.word_in [106], word_in[106]);
  buf(\oc8051_gm_cxrom_1.word_in [107], word_in[107]);
  buf(\oc8051_gm_cxrom_1.word_in [108], word_in[108]);
  buf(\oc8051_gm_cxrom_1.word_in [109], word_in[109]);
  buf(\oc8051_gm_cxrom_1.word_in [110], word_in[110]);
  buf(\oc8051_gm_cxrom_1.word_in [111], word_in[111]);
  buf(\oc8051_gm_cxrom_1.word_in [112], word_in[112]);
  buf(\oc8051_gm_cxrom_1.word_in [113], word_in[113]);
  buf(\oc8051_gm_cxrom_1.word_in [114], word_in[114]);
  buf(\oc8051_gm_cxrom_1.word_in [115], word_in[115]);
  buf(\oc8051_gm_cxrom_1.word_in [116], word_in[116]);
  buf(\oc8051_gm_cxrom_1.word_in [117], word_in[117]);
  buf(\oc8051_gm_cxrom_1.word_in [118], word_in[118]);
  buf(\oc8051_gm_cxrom_1.word_in [119], word_in[119]);
  buf(\oc8051_gm_cxrom_1.word_in [120], word_in[120]);
  buf(\oc8051_gm_cxrom_1.word_in [121], word_in[121]);
  buf(\oc8051_gm_cxrom_1.word_in [122], word_in[122]);
  buf(\oc8051_gm_cxrom_1.word_in [123], word_in[123]);
  buf(\oc8051_gm_cxrom_1.word_in [124], word_in[124]);
  buf(\oc8051_gm_cxrom_1.word_in [125], word_in[125]);
  buf(\oc8051_gm_cxrom_1.word_in [126], word_in[126]);
  buf(\oc8051_gm_cxrom_1.word_in [127], word_in[127]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [0], \oc8051_golden_model_1.PC [0]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [1], \oc8051_golden_model_1.PC [1]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [2], \oc8051_golden_model_1.PC [2]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [3], \oc8051_golden_model_1.PC [3]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [4], \oc8051_golden_model_1.PC [4]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [5], \oc8051_golden_model_1.PC [5]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [6], \oc8051_golden_model_1.PC [6]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [7], \oc8051_golden_model_1.PC [7]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [8], \oc8051_golden_model_1.PC [8]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [9], \oc8051_golden_model_1.PC [9]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [10], \oc8051_golden_model_1.PC [10]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [11], \oc8051_golden_model_1.PC [11]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [12], \oc8051_golden_model_1.PC [12]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [13], \oc8051_golden_model_1.PC [13]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [14], \oc8051_golden_model_1.PC [14]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [15], \oc8051_golden_model_1.PC [15]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [0], \oc8051_golden_model_1.PC [0]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [1], \oc8051_golden_model_1.PC [1]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [2], \oc8051_golden_model_1.PC [2]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [3], \oc8051_golden_model_1.PC [3]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [4], \oc8051_golden_model_1.PC [4]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [5], \oc8051_golden_model_1.PC [5]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [6], \oc8051_golden_model_1.PC [6]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [7], \oc8051_golden_model_1.PC [7]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [8], \oc8051_golden_model_1.PC [8]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [9], \oc8051_golden_model_1.PC [9]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [10], \oc8051_golden_model_1.PC [10]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [11], \oc8051_golden_model_1.PC [11]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [12], \oc8051_golden_model_1.PC [12]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [13], \oc8051_golden_model_1.PC [13]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [14], \oc8051_golden_model_1.PC [14]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [15], \oc8051_golden_model_1.PC [15]);
  buf(\oc8051_golden_model_1.clk , clk);
  buf(\oc8051_golden_model_1.rst , rst);
  buf(\oc8051_golden_model_1.ACC_03 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_03 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_03 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_03 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_03 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_03 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_03 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_03 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_13 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_13 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_13 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_13 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_13 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_13 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_13 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_13 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.ACC_23 [0], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_23 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_23 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_23 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_23 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_23 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_23 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_23 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_33 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.ACC_33 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_33 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_33 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_33 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_33 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_33 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_33 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_c4 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_c4 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_c4 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_c4 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_c4 [4], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_c4 [5], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_c4 [6], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_c4 [7], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_d6 [0], \oc8051_golden_model_1.n2868 );
  buf(\oc8051_golden_model_1.ACC_d6 [1], \oc8051_golden_model_1.n2867 );
  buf(\oc8051_golden_model_1.ACC_d6 [2], \oc8051_golden_model_1.n2866 );
  buf(\oc8051_golden_model_1.ACC_d6 [3], \oc8051_golden_model_1.n2865 );
  buf(\oc8051_golden_model_1.ACC_d6 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_d6 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_d6 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_d6 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_d7 [0], \oc8051_golden_model_1.n2868 );
  buf(\oc8051_golden_model_1.ACC_d7 [1], \oc8051_golden_model_1.n2867 );
  buf(\oc8051_golden_model_1.ACC_d7 [2], \oc8051_golden_model_1.n2866 );
  buf(\oc8051_golden_model_1.ACC_d7 [3], \oc8051_golden_model_1.n2865 );
  buf(\oc8051_golden_model_1.ACC_d7 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_d7 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_d7 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_d7 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_e6 [0], \oc8051_golden_model_1.n2868 );
  buf(\oc8051_golden_model_1.ACC_e6 [1], \oc8051_golden_model_1.n2867 );
  buf(\oc8051_golden_model_1.ACC_e6 [2], \oc8051_golden_model_1.n2866 );
  buf(\oc8051_golden_model_1.ACC_e6 [3], \oc8051_golden_model_1.n2865 );
  buf(\oc8051_golden_model_1.ACC_e6 [4], \oc8051_golden_model_1.n2860 [4]);
  buf(\oc8051_golden_model_1.ACC_e6 [5], \oc8051_golden_model_1.n2860 [5]);
  buf(\oc8051_golden_model_1.ACC_e6 [6], \oc8051_golden_model_1.n2860 [6]);
  buf(\oc8051_golden_model_1.ACC_e6 [7], \oc8051_golden_model_1.n2860 [7]);
  buf(\oc8051_golden_model_1.ACC_e7 [0], \oc8051_golden_model_1.n2868 );
  buf(\oc8051_golden_model_1.ACC_e7 [1], \oc8051_golden_model_1.n2867 );
  buf(\oc8051_golden_model_1.ACC_e7 [2], \oc8051_golden_model_1.n2866 );
  buf(\oc8051_golden_model_1.ACC_e7 [3], \oc8051_golden_model_1.n2865 );
  buf(\oc8051_golden_model_1.ACC_e7 [4], \oc8051_golden_model_1.n2860 [4]);
  buf(\oc8051_golden_model_1.ACC_e7 [5], \oc8051_golden_model_1.n2860 [5]);
  buf(\oc8051_golden_model_1.ACC_e7 [6], \oc8051_golden_model_1.n2860 [6]);
  buf(\oc8051_golden_model_1.ACC_e7 [7], \oc8051_golden_model_1.n2860 [7]);
  buf(\oc8051_golden_model_1.PC_22 [0], \oc8051_golden_model_1.n2868 );
  buf(\oc8051_golden_model_1.PC_22 [1], \oc8051_golden_model_1.n2867 );
  buf(\oc8051_golden_model_1.PC_22 [2], \oc8051_golden_model_1.n2866 );
  buf(\oc8051_golden_model_1.PC_22 [3], \oc8051_golden_model_1.n2865 );
  buf(\oc8051_golden_model_1.PC_22 [4], \oc8051_golden_model_1.n2860 [4]);
  buf(\oc8051_golden_model_1.PC_22 [5], \oc8051_golden_model_1.n2860 [5]);
  buf(\oc8051_golden_model_1.PC_22 [6], \oc8051_golden_model_1.n2860 [6]);
  buf(\oc8051_golden_model_1.PC_22 [7], \oc8051_golden_model_1.n2860 [7]);
  buf(\oc8051_golden_model_1.PC_22 [8], \oc8051_golden_model_1.n2775 );
  buf(\oc8051_golden_model_1.PC_22 [9], \oc8051_golden_model_1.n2774 );
  buf(\oc8051_golden_model_1.PC_22 [10], \oc8051_golden_model_1.n2773 );
  buf(\oc8051_golden_model_1.PC_22 [11], \oc8051_golden_model_1.n2772 );
  buf(\oc8051_golden_model_1.PC_22 [12], \oc8051_golden_model_1.n2771 );
  buf(\oc8051_golden_model_1.PC_22 [13], \oc8051_golden_model_1.n2770 );
  buf(\oc8051_golden_model_1.PC_22 [14], \oc8051_golden_model_1.n2769 );
  buf(\oc8051_golden_model_1.PC_22 [15], \oc8051_golden_model_1.n2768 );
  buf(\oc8051_golden_model_1.PC_32 [0], \oc8051_golden_model_1.n2868 );
  buf(\oc8051_golden_model_1.PC_32 [1], \oc8051_golden_model_1.n2867 );
  buf(\oc8051_golden_model_1.PC_32 [2], \oc8051_golden_model_1.n2866 );
  buf(\oc8051_golden_model_1.PC_32 [3], \oc8051_golden_model_1.n2865 );
  buf(\oc8051_golden_model_1.PC_32 [4], \oc8051_golden_model_1.n2860 [4]);
  buf(\oc8051_golden_model_1.PC_32 [5], \oc8051_golden_model_1.n2860 [5]);
  buf(\oc8051_golden_model_1.PC_32 [6], \oc8051_golden_model_1.n2860 [6]);
  buf(\oc8051_golden_model_1.PC_32 [7], \oc8051_golden_model_1.n2860 [7]);
  buf(\oc8051_golden_model_1.PC_32 [8], \oc8051_golden_model_1.n2775 );
  buf(\oc8051_golden_model_1.PC_32 [9], \oc8051_golden_model_1.n2774 );
  buf(\oc8051_golden_model_1.PC_32 [10], \oc8051_golden_model_1.n2773 );
  buf(\oc8051_golden_model_1.PC_32 [11], \oc8051_golden_model_1.n2772 );
  buf(\oc8051_golden_model_1.PC_32 [12], \oc8051_golden_model_1.n2771 );
  buf(\oc8051_golden_model_1.PC_32 [13], \oc8051_golden_model_1.n2770 );
  buf(\oc8051_golden_model_1.PC_32 [14], \oc8051_golden_model_1.n2769 );
  buf(\oc8051_golden_model_1.PC_32 [15], \oc8051_golden_model_1.n2768 );
  buf(\oc8051_golden_model_1.PSW_00 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_00 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_00 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_00 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_00 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_00 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_00 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_00 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_01 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_01 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_01 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_01 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_01 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_01 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_01 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_01 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_02 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_02 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_02 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_02 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_02 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_02 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_02 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_02 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_03 [0], \oc8051_golden_model_1.n1047 [0]);
  buf(\oc8051_golden_model_1.PSW_03 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_03 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_03 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_03 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_03 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_03 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_03 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_04 [0], \oc8051_golden_model_1.n1064 [0]);
  buf(\oc8051_golden_model_1.PSW_04 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_04 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_04 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_04 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_04 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_04 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_04 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_06 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_06 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_06 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_06 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_06 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_06 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_06 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_06 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_07 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_07 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_07 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_07 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_07 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_07 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_07 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_07 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_08 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_08 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_08 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_08 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_08 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_08 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_08 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_08 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_09 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_09 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_09 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_09 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_09 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_09 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_09 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_09 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0a [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_0a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0b [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_0b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0c [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_0c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0d [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_0d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0e [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_0e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0f [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_0f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_11 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_11 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_11 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_11 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_11 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_11 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_11 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_11 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_12 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_12 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_12 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_12 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_12 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_12 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_12 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_12 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_13 [0], \oc8051_golden_model_1.n1284 [0]);
  buf(\oc8051_golden_model_1.PSW_13 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_13 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_13 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_13 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_13 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_13 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_13 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.PSW_14 [0], \oc8051_golden_model_1.n1301 [0]);
  buf(\oc8051_golden_model_1.PSW_14 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_14 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_14 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_14 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_14 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_14 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_14 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_16 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_16 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_16 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_16 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_16 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_16 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_16 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_16 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_17 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_17 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_17 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_17 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_17 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_17 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_17 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_17 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_18 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_18 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_18 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_18 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_18 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_18 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_18 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_18 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_19 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_19 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_19 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_19 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_19 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_19 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_19 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_19 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1a [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_1a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1b [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_1b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1c [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_1c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1d [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_1d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1e [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_1e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1f [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_1f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_20 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_20 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_20 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_20 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_20 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_20 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_20 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_20 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_21 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_21 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_21 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_21 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_21 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_21 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_21 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_21 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_22 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_22 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_22 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_22 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_22 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_22 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_22 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_22 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_23 [0], \oc8051_golden_model_1.n1361 [0]);
  buf(\oc8051_golden_model_1.PSW_23 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_23 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_23 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_23 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_23 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_23 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_23 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_24 [0], \oc8051_golden_model_1.n1402 [0]);
  buf(\oc8051_golden_model_1.PSW_24 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_24 [2], \oc8051_golden_model_1.n1402 [2]);
  buf(\oc8051_golden_model_1.PSW_24 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_24 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_24 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_24 [6], \oc8051_golden_model_1.n1402 [6]);
  buf(\oc8051_golden_model_1.PSW_24 [7], \oc8051_golden_model_1.n1402 [7]);
  buf(\oc8051_golden_model_1.PSW_25 [0], \oc8051_golden_model_1.n1457 [0]);
  buf(\oc8051_golden_model_1.PSW_25 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_25 [2], \oc8051_golden_model_1.n1457 [2]);
  buf(\oc8051_golden_model_1.PSW_25 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_25 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_25 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_25 [6], \oc8051_golden_model_1.n1457 [6]);
  buf(\oc8051_golden_model_1.PSW_25 [7], \oc8051_golden_model_1.n1457 [7]);
  buf(\oc8051_golden_model_1.PSW_26 [0], \oc8051_golden_model_1.n1507 [0]);
  buf(\oc8051_golden_model_1.PSW_26 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_26 [2], \oc8051_golden_model_1.n1493 [2]);
  buf(\oc8051_golden_model_1.PSW_26 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_26 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_26 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_26 [6], \oc8051_golden_model_1.n1507 [6]);
  buf(\oc8051_golden_model_1.PSW_26 [7], \oc8051_golden_model_1.n1493 [7]);
  buf(\oc8051_golden_model_1.PSW_27 [0], \oc8051_golden_model_1.n1507 [0]);
  buf(\oc8051_golden_model_1.PSW_27 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_27 [2], \oc8051_golden_model_1.n1507 [2]);
  buf(\oc8051_golden_model_1.PSW_27 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_27 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_27 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_27 [6], \oc8051_golden_model_1.n1507 [6]);
  buf(\oc8051_golden_model_1.PSW_27 [7], \oc8051_golden_model_1.n1507 [7]);
  buf(\oc8051_golden_model_1.PSW_28 [0], \oc8051_golden_model_1.n1564 [0]);
  buf(\oc8051_golden_model_1.PSW_28 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_28 [2], \oc8051_golden_model_1.n1548 [2]);
  buf(\oc8051_golden_model_1.PSW_28 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_28 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_28 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_28 [6], \oc8051_golden_model_1.n1564 [6]);
  buf(\oc8051_golden_model_1.PSW_28 [7], \oc8051_golden_model_1.n1548 [7]);
  buf(\oc8051_golden_model_1.PSW_29 [0], \oc8051_golden_model_1.n1564 [0]);
  buf(\oc8051_golden_model_1.PSW_29 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_29 [2], \oc8051_golden_model_1.n1548 [2]);
  buf(\oc8051_golden_model_1.PSW_29 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_29 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_29 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_29 [6], \oc8051_golden_model_1.n1564 [6]);
  buf(\oc8051_golden_model_1.PSW_29 [7], \oc8051_golden_model_1.n1548 [7]);
  buf(\oc8051_golden_model_1.PSW_2a [0], \oc8051_golden_model_1.n1564 [0]);
  buf(\oc8051_golden_model_1.PSW_2a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2a [2], \oc8051_golden_model_1.n1548 [2]);
  buf(\oc8051_golden_model_1.PSW_2a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2a [6], \oc8051_golden_model_1.n1561 [6]);
  buf(\oc8051_golden_model_1.PSW_2a [7], \oc8051_golden_model_1.n1548 [7]);
  buf(\oc8051_golden_model_1.PSW_2b [0], \oc8051_golden_model_1.n1564 [0]);
  buf(\oc8051_golden_model_1.PSW_2b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2b [2], \oc8051_golden_model_1.n1564 [2]);
  buf(\oc8051_golden_model_1.PSW_2b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2b [6], \oc8051_golden_model_1.n1561 [6]);
  buf(\oc8051_golden_model_1.PSW_2b [7], \oc8051_golden_model_1.n1564 [7]);
  buf(\oc8051_golden_model_1.PSW_2c [0], \oc8051_golden_model_1.n1564 [0]);
  buf(\oc8051_golden_model_1.PSW_2c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2c [2], \oc8051_golden_model_1.n1564 [2]);
  buf(\oc8051_golden_model_1.PSW_2c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2c [6], \oc8051_golden_model_1.n1561 [6]);
  buf(\oc8051_golden_model_1.PSW_2c [7], \oc8051_golden_model_1.n1564 [7]);
  buf(\oc8051_golden_model_1.PSW_2d [0], \oc8051_golden_model_1.n1564 [0]);
  buf(\oc8051_golden_model_1.PSW_2d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2d [2], \oc8051_golden_model_1.n1548 [2]);
  buf(\oc8051_golden_model_1.PSW_2d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2d [6], \oc8051_golden_model_1.n1564 [6]);
  buf(\oc8051_golden_model_1.PSW_2d [7], \oc8051_golden_model_1.n1548 [7]);
  buf(\oc8051_golden_model_1.PSW_2e [0], \oc8051_golden_model_1.n1564 [0]);
  buf(\oc8051_golden_model_1.PSW_2e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2e [2], \oc8051_golden_model_1.n1564 [2]);
  buf(\oc8051_golden_model_1.PSW_2e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2e [6], \oc8051_golden_model_1.n1564 [6]);
  buf(\oc8051_golden_model_1.PSW_2e [7], \oc8051_golden_model_1.n1564 [7]);
  buf(\oc8051_golden_model_1.PSW_2f [0], \oc8051_golden_model_1.n1564 [0]);
  buf(\oc8051_golden_model_1.PSW_2f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2f [2], \oc8051_golden_model_1.n1564 [2]);
  buf(\oc8051_golden_model_1.PSW_2f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2f [6], \oc8051_golden_model_1.n1564 [6]);
  buf(\oc8051_golden_model_1.PSW_2f [7], \oc8051_golden_model_1.n1564 [7]);
  buf(\oc8051_golden_model_1.PSW_30 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_30 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_30 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_30 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_30 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_30 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_30 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_30 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_31 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_31 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_31 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_31 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_31 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_31 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_31 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_31 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_32 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_32 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_32 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_32 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_32 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_32 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_32 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_32 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_33 [0], \oc8051_golden_model_1.n1587 [0]);
  buf(\oc8051_golden_model_1.PSW_33 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_33 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_33 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_33 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_33 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_33 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_33 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.PSW_34 [0], \oc8051_golden_model_1.n1623 [0]);
  buf(\oc8051_golden_model_1.PSW_34 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_34 [2], \oc8051_golden_model_1.n1623 [2]);
  buf(\oc8051_golden_model_1.PSW_34 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_34 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_34 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_34 [6], \oc8051_golden_model_1.n1623 [6]);
  buf(\oc8051_golden_model_1.PSW_34 [7], \oc8051_golden_model_1.n1623 [7]);
  buf(\oc8051_golden_model_1.PSW_35 [0], \oc8051_golden_model_1.n1656 [0]);
  buf(\oc8051_golden_model_1.PSW_35 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_35 [2], \oc8051_golden_model_1.n1656 [2]);
  buf(\oc8051_golden_model_1.PSW_35 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_35 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_35 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_35 [6], \oc8051_golden_model_1.n1656 [6]);
  buf(\oc8051_golden_model_1.PSW_35 [7], \oc8051_golden_model_1.n1656 [7]);
  buf(\oc8051_golden_model_1.PSW_36 [0], \oc8051_golden_model_1.n1689 [0]);
  buf(\oc8051_golden_model_1.PSW_36 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_36 [2], \oc8051_golden_model_1.n1689 [2]);
  buf(\oc8051_golden_model_1.PSW_36 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_36 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_36 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_36 [6], \oc8051_golden_model_1.n1689 [6]);
  buf(\oc8051_golden_model_1.PSW_36 [7], \oc8051_golden_model_1.n1689 [7]);
  buf(\oc8051_golden_model_1.PSW_37 [0], \oc8051_golden_model_1.n1689 [0]);
  buf(\oc8051_golden_model_1.PSW_37 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_37 [2], \oc8051_golden_model_1.n1689 [2]);
  buf(\oc8051_golden_model_1.PSW_37 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_37 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_37 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_37 [6], \oc8051_golden_model_1.n1689 [6]);
  buf(\oc8051_golden_model_1.PSW_37 [7], \oc8051_golden_model_1.n1689 [7]);
  buf(\oc8051_golden_model_1.PSW_38 [0], \oc8051_golden_model_1.n1722 [0]);
  buf(\oc8051_golden_model_1.PSW_38 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_38 [2], \oc8051_golden_model_1.n1722 [2]);
  buf(\oc8051_golden_model_1.PSW_38 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_38 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_38 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_38 [6], \oc8051_golden_model_1.n1722 [6]);
  buf(\oc8051_golden_model_1.PSW_38 [7], \oc8051_golden_model_1.n1722 [7]);
  buf(\oc8051_golden_model_1.PSW_39 [0], \oc8051_golden_model_1.n1722 [0]);
  buf(\oc8051_golden_model_1.PSW_39 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_39 [2], \oc8051_golden_model_1.n1722 [2]);
  buf(\oc8051_golden_model_1.PSW_39 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_39 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_39 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_39 [6], \oc8051_golden_model_1.n1722 [6]);
  buf(\oc8051_golden_model_1.PSW_39 [7], \oc8051_golden_model_1.n1722 [7]);
  buf(\oc8051_golden_model_1.PSW_3a [0], \oc8051_golden_model_1.n1722 [0]);
  buf(\oc8051_golden_model_1.PSW_3a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3a [2], \oc8051_golden_model_1.n1722 [2]);
  buf(\oc8051_golden_model_1.PSW_3a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3a [6], \oc8051_golden_model_1.n1722 [6]);
  buf(\oc8051_golden_model_1.PSW_3a [7], \oc8051_golden_model_1.n1722 [7]);
  buf(\oc8051_golden_model_1.PSW_3b [0], \oc8051_golden_model_1.n1722 [0]);
  buf(\oc8051_golden_model_1.PSW_3b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3b [2], \oc8051_golden_model_1.n1722 [2]);
  buf(\oc8051_golden_model_1.PSW_3b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3b [6], \oc8051_golden_model_1.n1722 [6]);
  buf(\oc8051_golden_model_1.PSW_3b [7], \oc8051_golden_model_1.n1722 [7]);
  buf(\oc8051_golden_model_1.PSW_3c [0], \oc8051_golden_model_1.n1722 [0]);
  buf(\oc8051_golden_model_1.PSW_3c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3c [2], \oc8051_golden_model_1.n1722 [2]);
  buf(\oc8051_golden_model_1.PSW_3c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3c [6], \oc8051_golden_model_1.n1722 [6]);
  buf(\oc8051_golden_model_1.PSW_3c [7], \oc8051_golden_model_1.n1722 [7]);
  buf(\oc8051_golden_model_1.PSW_3d [0], \oc8051_golden_model_1.n1722 [0]);
  buf(\oc8051_golden_model_1.PSW_3d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3d [2], \oc8051_golden_model_1.n1722 [2]);
  buf(\oc8051_golden_model_1.PSW_3d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3d [6], \oc8051_golden_model_1.n1722 [6]);
  buf(\oc8051_golden_model_1.PSW_3d [7], \oc8051_golden_model_1.n1722 [7]);
  buf(\oc8051_golden_model_1.PSW_3e [0], \oc8051_golden_model_1.n1722 [0]);
  buf(\oc8051_golden_model_1.PSW_3e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3e [2], \oc8051_golden_model_1.n1722 [2]);
  buf(\oc8051_golden_model_1.PSW_3e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3e [6], \oc8051_golden_model_1.n1722 [6]);
  buf(\oc8051_golden_model_1.PSW_3e [7], \oc8051_golden_model_1.n1722 [7]);
  buf(\oc8051_golden_model_1.PSW_3f [0], \oc8051_golden_model_1.n1722 [0]);
  buf(\oc8051_golden_model_1.PSW_3f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3f [2], \oc8051_golden_model_1.n1722 [2]);
  buf(\oc8051_golden_model_1.PSW_3f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3f [6], \oc8051_golden_model_1.n1722 [6]);
  buf(\oc8051_golden_model_1.PSW_3f [7], \oc8051_golden_model_1.n1722 [7]);
  buf(\oc8051_golden_model_1.PSW_40 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_40 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_40 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_40 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_40 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_40 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_40 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_40 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_41 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_41 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_41 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_41 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_41 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_41 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_41 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_41 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_42 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_42 [1], \oc8051_golden_model_1.n1749 [1]);
  buf(\oc8051_golden_model_1.PSW_42 [2], \oc8051_golden_model_1.n1749 [2]);
  buf(\oc8051_golden_model_1.PSW_42 [3], \oc8051_golden_model_1.n1749 [3]);
  buf(\oc8051_golden_model_1.PSW_42 [4], \oc8051_golden_model_1.n1749 [4]);
  buf(\oc8051_golden_model_1.PSW_42 [5], \oc8051_golden_model_1.n1749 [5]);
  buf(\oc8051_golden_model_1.PSW_42 [6], \oc8051_golden_model_1.n1749 [6]);
  buf(\oc8051_golden_model_1.PSW_42 [7], \oc8051_golden_model_1.n1749 [7]);
  buf(\oc8051_golden_model_1.PSW_44 [0], \oc8051_golden_model_1.n1805 [0]);
  buf(\oc8051_golden_model_1.PSW_44 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_44 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_44 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_44 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_44 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_44 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_44 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_45 [0], \oc8051_golden_model_1.n1822 [0]);
  buf(\oc8051_golden_model_1.PSW_45 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_45 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_45 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_45 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_45 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_45 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_45 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_46 [0], \oc8051_golden_model_1.n1839 [0]);
  buf(\oc8051_golden_model_1.PSW_46 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_46 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_46 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_46 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_46 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_46 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_46 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_47 [0], \oc8051_golden_model_1.n1839 [0]);
  buf(\oc8051_golden_model_1.PSW_47 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_47 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_47 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_47 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_47 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_47 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_47 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_48 [0], \oc8051_golden_model_1.n1856 [0]);
  buf(\oc8051_golden_model_1.PSW_48 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_48 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_48 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_48 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_48 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_48 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_48 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_49 [0], \oc8051_golden_model_1.n1856 [0]);
  buf(\oc8051_golden_model_1.PSW_49 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_49 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_49 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_49 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_49 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_49 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_49 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4a [0], \oc8051_golden_model_1.n1856 [0]);
  buf(\oc8051_golden_model_1.PSW_4a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4b [0], \oc8051_golden_model_1.n1856 [0]);
  buf(\oc8051_golden_model_1.PSW_4b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4c [0], \oc8051_golden_model_1.n1856 [0]);
  buf(\oc8051_golden_model_1.PSW_4c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4d [0], \oc8051_golden_model_1.n1856 [0]);
  buf(\oc8051_golden_model_1.PSW_4d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4e [0], \oc8051_golden_model_1.n1856 [0]);
  buf(\oc8051_golden_model_1.PSW_4e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4f [0], \oc8051_golden_model_1.n1856 [0]);
  buf(\oc8051_golden_model_1.PSW_4f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_50 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_50 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_50 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_50 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_50 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_50 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_50 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_50 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_51 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_51 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_51 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_51 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_51 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_51 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_51 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_51 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_52 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_52 [1], \oc8051_golden_model_1.n1881 [1]);
  buf(\oc8051_golden_model_1.PSW_52 [2], \oc8051_golden_model_1.n1881 [2]);
  buf(\oc8051_golden_model_1.PSW_52 [3], \oc8051_golden_model_1.n1881 [3]);
  buf(\oc8051_golden_model_1.PSW_52 [4], \oc8051_golden_model_1.n1881 [4]);
  buf(\oc8051_golden_model_1.PSW_52 [5], \oc8051_golden_model_1.n1881 [5]);
  buf(\oc8051_golden_model_1.PSW_52 [6], \oc8051_golden_model_1.n1881 [6]);
  buf(\oc8051_golden_model_1.PSW_52 [7], \oc8051_golden_model_1.n1881 [7]);
  buf(\oc8051_golden_model_1.PSW_54 [0], \oc8051_golden_model_1.n1937 [0]);
  buf(\oc8051_golden_model_1.PSW_54 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_54 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_54 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_54 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_54 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_54 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_54 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_55 [0], \oc8051_golden_model_1.n1954 [0]);
  buf(\oc8051_golden_model_1.PSW_55 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_55 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_55 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_55 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_55 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_55 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_55 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_56 [0], \oc8051_golden_model_1.n1971 [0]);
  buf(\oc8051_golden_model_1.PSW_56 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_56 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_56 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_56 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_56 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_56 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_56 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_57 [0], \oc8051_golden_model_1.n1971 [0]);
  buf(\oc8051_golden_model_1.PSW_57 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_57 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_57 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_57 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_57 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_57 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_57 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_58 [0], \oc8051_golden_model_1.n1988 [0]);
  buf(\oc8051_golden_model_1.PSW_58 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_58 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_58 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_58 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_58 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_58 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_58 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_59 [0], \oc8051_golden_model_1.n1988 [0]);
  buf(\oc8051_golden_model_1.PSW_59 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_59 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_59 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_59 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_59 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_59 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_59 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5a [0], \oc8051_golden_model_1.n1988 [0]);
  buf(\oc8051_golden_model_1.PSW_5a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5b [0], \oc8051_golden_model_1.n1988 [0]);
  buf(\oc8051_golden_model_1.PSW_5b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5c [0], \oc8051_golden_model_1.n1988 [0]);
  buf(\oc8051_golden_model_1.PSW_5c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5d [0], \oc8051_golden_model_1.n1988 [0]);
  buf(\oc8051_golden_model_1.PSW_5d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5e [0], \oc8051_golden_model_1.n1988 [0]);
  buf(\oc8051_golden_model_1.PSW_5e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5f [0], \oc8051_golden_model_1.n1988 [0]);
  buf(\oc8051_golden_model_1.PSW_5f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_60 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_60 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_60 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_60 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_60 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_60 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_60 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_60 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_61 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_61 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_61 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_61 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_61 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_61 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_61 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_61 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_64 [0], \oc8051_golden_model_1.n2086 [0]);
  buf(\oc8051_golden_model_1.PSW_64 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_64 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_64 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_64 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_64 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_64 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_64 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_65 [0], \oc8051_golden_model_1.n2103 [0]);
  buf(\oc8051_golden_model_1.PSW_65 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_65 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_65 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_65 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_65 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_65 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_65 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_66 [0], \oc8051_golden_model_1.n2120 [0]);
  buf(\oc8051_golden_model_1.PSW_66 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_66 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_66 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_66 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_66 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_66 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_66 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_67 [0], \oc8051_golden_model_1.n2120 [0]);
  buf(\oc8051_golden_model_1.PSW_67 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_67 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_67 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_67 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_67 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_67 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_67 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_68 [0], \oc8051_golden_model_1.n2137 [0]);
  buf(\oc8051_golden_model_1.PSW_68 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_68 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_68 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_68 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_68 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_68 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_68 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_69 [0], \oc8051_golden_model_1.n2137 [0]);
  buf(\oc8051_golden_model_1.PSW_69 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_69 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_69 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_69 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_69 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_69 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_69 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6a [0], \oc8051_golden_model_1.n2137 [0]);
  buf(\oc8051_golden_model_1.PSW_6a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6b [0], \oc8051_golden_model_1.n2137 [0]);
  buf(\oc8051_golden_model_1.PSW_6b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6c [0], \oc8051_golden_model_1.n2137 [0]);
  buf(\oc8051_golden_model_1.PSW_6c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6d [0], \oc8051_golden_model_1.n2137 [0]);
  buf(\oc8051_golden_model_1.PSW_6d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6e [0], \oc8051_golden_model_1.n2137 [0]);
  buf(\oc8051_golden_model_1.PSW_6e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6f [0], \oc8051_golden_model_1.n2137 [0]);
  buf(\oc8051_golden_model_1.PSW_6f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_70 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_70 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_70 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_70 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_70 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_70 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_70 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_70 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_71 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_71 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_71 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_71 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_71 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_71 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_71 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_71 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_72 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_72 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_72 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_72 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_72 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_72 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_72 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_72 [7], \oc8051_golden_model_1.n2145 [7]);
  buf(\oc8051_golden_model_1.PSW_73 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_73 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_73 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_73 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_73 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_73 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_73 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_73 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_74 [0], \oc8051_golden_model_1.n2161 [0]);
  buf(\oc8051_golden_model_1.PSW_74 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_74 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_74 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_74 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_74 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_74 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_74 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_76 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_76 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_76 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_76 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_76 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_76 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_76 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_76 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_77 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_77 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_77 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_77 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_77 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_77 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_77 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_77 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_78 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_78 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_78 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_78 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_78 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_78 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_78 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_78 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_79 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_79 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_79 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_79 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_79 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_79 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_79 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_79 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7a [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_7a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7b [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_7b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7c [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_7c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7d [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_7d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7e [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_7e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7f [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_7f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_80 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_80 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_80 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_80 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_80 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_80 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_80 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_80 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_81 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_81 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_81 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_81 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_81 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_81 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_81 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_81 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_82 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_82 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_82 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_82 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_82 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_82 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_82 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_82 [7], \oc8051_golden_model_1.n2203 [7]);
  buf(\oc8051_golden_model_1.PSW_83 [0], \oc8051_golden_model_1.n2161 [0]);
  buf(\oc8051_golden_model_1.PSW_83 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_83 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_83 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_83 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_83 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_83 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_83 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_84 [0], \oc8051_golden_model_1.n2229 [0]);
  buf(\oc8051_golden_model_1.PSW_84 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_84 [2], \oc8051_golden_model_1.n2229 [2]);
  buf(\oc8051_golden_model_1.PSW_84 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_84 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_84 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_84 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_84 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_90 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_90 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_90 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_90 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_90 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_90 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_90 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_90 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_91 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_91 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_91 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_91 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_91 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_91 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_91 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_91 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_93 [0], \oc8051_golden_model_1.n2161 [0]);
  buf(\oc8051_golden_model_1.PSW_93 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_93 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_93 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_93 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_93 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_93 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_93 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_94 [0], \oc8051_golden_model_1.n2470 [0]);
  buf(\oc8051_golden_model_1.PSW_94 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_94 [2], \oc8051_golden_model_1.n2470 [2]);
  buf(\oc8051_golden_model_1.PSW_94 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_94 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_94 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_94 [6], \oc8051_golden_model_1.n2470 [6]);
  buf(\oc8051_golden_model_1.PSW_94 [7], \oc8051_golden_model_1.n2470 [7]);
  buf(\oc8051_golden_model_1.PSW_95 [0], \oc8051_golden_model_1.n2500 [0]);
  buf(\oc8051_golden_model_1.PSW_95 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_95 [2], \oc8051_golden_model_1.n2500 [2]);
  buf(\oc8051_golden_model_1.PSW_95 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_95 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_95 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_95 [6], \oc8051_golden_model_1.n2500 [6]);
  buf(\oc8051_golden_model_1.PSW_95 [7], \oc8051_golden_model_1.n2500 [7]);
  buf(\oc8051_golden_model_1.PSW_96 [0], \oc8051_golden_model_1.n2530 [0]);
  buf(\oc8051_golden_model_1.PSW_96 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_96 [2], \oc8051_golden_model_1.n2530 [2]);
  buf(\oc8051_golden_model_1.PSW_96 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_96 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_96 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_96 [6], \oc8051_golden_model_1.n2530 [6]);
  buf(\oc8051_golden_model_1.PSW_96 [7], \oc8051_golden_model_1.n2530 [7]);
  buf(\oc8051_golden_model_1.PSW_97 [0], \oc8051_golden_model_1.n2530 [0]);
  buf(\oc8051_golden_model_1.PSW_97 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_97 [2], \oc8051_golden_model_1.n2530 [2]);
  buf(\oc8051_golden_model_1.PSW_97 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_97 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_97 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_97 [6], \oc8051_golden_model_1.n2530 [6]);
  buf(\oc8051_golden_model_1.PSW_97 [7], \oc8051_golden_model_1.n2530 [7]);
  buf(\oc8051_golden_model_1.PSW_98 [0], \oc8051_golden_model_1.n2560 [0]);
  buf(\oc8051_golden_model_1.PSW_98 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_98 [2], \oc8051_golden_model_1.n2560 [2]);
  buf(\oc8051_golden_model_1.PSW_98 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_98 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_98 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_98 [6], \oc8051_golden_model_1.n2560 [6]);
  buf(\oc8051_golden_model_1.PSW_98 [7], \oc8051_golden_model_1.n2560 [7]);
  buf(\oc8051_golden_model_1.PSW_99 [0], \oc8051_golden_model_1.n2560 [0]);
  buf(\oc8051_golden_model_1.PSW_99 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_99 [2], \oc8051_golden_model_1.n2560 [2]);
  buf(\oc8051_golden_model_1.PSW_99 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_99 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_99 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_99 [6], \oc8051_golden_model_1.n2560 [6]);
  buf(\oc8051_golden_model_1.PSW_99 [7], \oc8051_golden_model_1.n2560 [7]);
  buf(\oc8051_golden_model_1.PSW_9a [0], \oc8051_golden_model_1.n2560 [0]);
  buf(\oc8051_golden_model_1.PSW_9a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9a [2], \oc8051_golden_model_1.n2560 [2]);
  buf(\oc8051_golden_model_1.PSW_9a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9a [6], \oc8051_golden_model_1.n2560 [6]);
  buf(\oc8051_golden_model_1.PSW_9a [7], \oc8051_golden_model_1.n2560 [7]);
  buf(\oc8051_golden_model_1.PSW_9b [0], \oc8051_golden_model_1.n2560 [0]);
  buf(\oc8051_golden_model_1.PSW_9b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9b [2], \oc8051_golden_model_1.n2560 [2]);
  buf(\oc8051_golden_model_1.PSW_9b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9b [6], \oc8051_golden_model_1.n2560 [6]);
  buf(\oc8051_golden_model_1.PSW_9b [7], \oc8051_golden_model_1.n2560 [7]);
  buf(\oc8051_golden_model_1.PSW_9c [0], \oc8051_golden_model_1.n2560 [0]);
  buf(\oc8051_golden_model_1.PSW_9c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9c [2], \oc8051_golden_model_1.n2560 [2]);
  buf(\oc8051_golden_model_1.PSW_9c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9c [6], \oc8051_golden_model_1.n2560 [6]);
  buf(\oc8051_golden_model_1.PSW_9c [7], \oc8051_golden_model_1.n2560 [7]);
  buf(\oc8051_golden_model_1.PSW_9d [0], \oc8051_golden_model_1.n2560 [0]);
  buf(\oc8051_golden_model_1.PSW_9d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9d [2], \oc8051_golden_model_1.n2560 [2]);
  buf(\oc8051_golden_model_1.PSW_9d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9d [6], \oc8051_golden_model_1.n2560 [6]);
  buf(\oc8051_golden_model_1.PSW_9d [7], \oc8051_golden_model_1.n2560 [7]);
  buf(\oc8051_golden_model_1.PSW_9e [0], \oc8051_golden_model_1.n2560 [0]);
  buf(\oc8051_golden_model_1.PSW_9e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9e [2], \oc8051_golden_model_1.n2560 [2]);
  buf(\oc8051_golden_model_1.PSW_9e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9e [6], \oc8051_golden_model_1.n2560 [6]);
  buf(\oc8051_golden_model_1.PSW_9e [7], \oc8051_golden_model_1.n2560 [7]);
  buf(\oc8051_golden_model_1.PSW_9f [0], \oc8051_golden_model_1.n2560 [0]);
  buf(\oc8051_golden_model_1.PSW_9f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9f [2], \oc8051_golden_model_1.n2560 [2]);
  buf(\oc8051_golden_model_1.PSW_9f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9f [6], \oc8051_golden_model_1.n2560 [6]);
  buf(\oc8051_golden_model_1.PSW_9f [7], \oc8051_golden_model_1.n2560 [7]);
  buf(\oc8051_golden_model_1.PSW_a0 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_a0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a0 [7], \oc8051_golden_model_1.n2565 [7]);
  buf(\oc8051_golden_model_1.PSW_a1 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_a1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a2 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_a2 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a2 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a2 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a2 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a2 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a2 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a2 [7], \oc8051_golden_model_1.n2568 [7]);
  buf(\oc8051_golden_model_1.PSW_a3 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_a3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a3 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a4 [0], \oc8051_golden_model_1.n2596 [0]);
  buf(\oc8051_golden_model_1.PSW_a4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a4 [2], \oc8051_golden_model_1.n2596 [2]);
  buf(\oc8051_golden_model_1.PSW_a4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a4 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_a5 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_a5 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a5 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a5 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a5 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a5 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a5 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a5 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a6 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_a6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a7 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_a7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a8 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_a8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a9 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_a9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_aa [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_aa [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_aa [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_aa [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_aa [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_aa [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_aa [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_aa [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ab [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_ab [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ab [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ab [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ab [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ab [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ab [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ab [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ac [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_ac [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ac [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ac [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ac [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ac [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ac [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ac [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ad [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_ad [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ad [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ad [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ad [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ad [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ad [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ad [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ae [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_ae [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ae [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ae [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ae [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ae [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ae [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ae [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_af [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_af [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_af [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_af [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_af [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_af [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_af [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_af [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_b0 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_b0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b0 [7], \oc8051_golden_model_1.n2602 [7]);
  buf(\oc8051_golden_model_1.PSW_b1 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_b1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_b3 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_b3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b3 [7], \oc8051_golden_model_1.n2637 [7]);
  buf(\oc8051_golden_model_1.PSW_b4 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_b4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b4 [7], \oc8051_golden_model_1.n2645 [7]);
  buf(\oc8051_golden_model_1.PSW_b5 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_b5 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b5 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b5 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b5 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b5 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b5 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b5 [7], \oc8051_golden_model_1.n2653 [7]);
  buf(\oc8051_golden_model_1.PSW_b6 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_b6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b6 [7], \oc8051_golden_model_1.n2661 [7]);
  buf(\oc8051_golden_model_1.PSW_b7 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_b7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b7 [7], \oc8051_golden_model_1.n2661 [7]);
  buf(\oc8051_golden_model_1.PSW_b8 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_b8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b8 [7], \oc8051_golden_model_1.n2669 [7]);
  buf(\oc8051_golden_model_1.PSW_b9 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_b9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b9 [7], \oc8051_golden_model_1.n2669 [7]);
  buf(\oc8051_golden_model_1.PSW_ba [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_ba [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ba [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ba [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ba [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ba [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ba [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ba [7], \oc8051_golden_model_1.n2669 [7]);
  buf(\oc8051_golden_model_1.PSW_bb [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_bb [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bb [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bb [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bb [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bb [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bb [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bb [7], \oc8051_golden_model_1.n2669 [7]);
  buf(\oc8051_golden_model_1.PSW_bc [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_bc [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bc [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bc [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bc [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bc [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bc [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bc [7], \oc8051_golden_model_1.n2669 [7]);
  buf(\oc8051_golden_model_1.PSW_bd [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_bd [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bd [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bd [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bd [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bd [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bd [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bd [7], \oc8051_golden_model_1.n2669 [7]);
  buf(\oc8051_golden_model_1.PSW_be [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_be [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_be [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_be [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_be [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_be [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_be [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_be [7], \oc8051_golden_model_1.n2669 [7]);
  buf(\oc8051_golden_model_1.PSW_bf [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_bf [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bf [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bf [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bf [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bf [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bf [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bf [7], \oc8051_golden_model_1.n2669 [7]);
  buf(\oc8051_golden_model_1.PSW_c0 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_c0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c0 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c1 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_c1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c3 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_c3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c3 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_c4 [0], \oc8051_golden_model_1.n2714 [0]);
  buf(\oc8051_golden_model_1.PSW_c4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c4 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c6 [0], \oc8051_golden_model_1.n2767 [0]);
  buf(\oc8051_golden_model_1.PSW_c6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c7 [0], \oc8051_golden_model_1.n2767 [0]);
  buf(\oc8051_golden_model_1.PSW_c7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c8 [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_c8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c9 [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_c9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ca [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_ca [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ca [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ca [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ca [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ca [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ca [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ca [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_cb [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_cb [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_cb [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_cb [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_cb [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_cb [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_cb [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_cb [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_cc [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_cc [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_cc [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_cc [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_cc [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_cc [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_cc [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_cc [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_cd [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_cd [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_cd [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_cd [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_cd [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_cd [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_cd [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_cd [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ce [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_ce [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ce [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ce [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ce [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ce [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ce [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ce [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_cf [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_cf [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_cf [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_cf [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_cf [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_cf [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_cf [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_cf [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d1 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_d1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d3 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_d3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d3 [7], 1'b1);
  buf(\oc8051_golden_model_1.PSW_d4 [0], \oc8051_golden_model_1.n2854 [0]);
  buf(\oc8051_golden_model_1.PSW_d4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d4 [7], \oc8051_golden_model_1.n2854 [7]);
  buf(\oc8051_golden_model_1.PSW_d6 [0], \oc8051_golden_model_1.n2876 [0]);
  buf(\oc8051_golden_model_1.PSW_d6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d7 [0], \oc8051_golden_model_1.n2876 [0]);
  buf(\oc8051_golden_model_1.PSW_d7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d8 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_d8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d9 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_d9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_da [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_da [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_da [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_da [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_da [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_da [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_da [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_da [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_db [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_db [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_db [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_db [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_db [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_db [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_db [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_db [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_dc [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_dc [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_dc [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_dc [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_dc [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_dc [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_dc [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_dc [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_dd [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_dd [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_dd [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_dd [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_dd [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_dd [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_dd [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_dd [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_de [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_de [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_de [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_de [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_de [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_de [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_de [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_de [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_df [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_df [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_df [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_df [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_df [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_df [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_df [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_df [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e1 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_e1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e4 [0], \oc8051_golden_model_1.n2895 [0]);
  buf(\oc8051_golden_model_1.PSW_e4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e4 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e5 [0], \oc8051_golden_model_1.n2896 [0]);
  buf(\oc8051_golden_model_1.PSW_e5 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e5 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e5 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e5 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e5 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e5 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e5 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e6 [0], \oc8051_golden_model_1.n2767 [0]);
  buf(\oc8051_golden_model_1.PSW_e6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e7 [0], \oc8051_golden_model_1.n2767 [0]);
  buf(\oc8051_golden_model_1.PSW_e7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e8 [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_e8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e9 [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_e9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ea [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_ea [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ea [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ea [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ea [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ea [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ea [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ea [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_eb [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_eb [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_eb [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_eb [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_eb [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_eb [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_eb [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_eb [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ec [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_ec [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ec [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ec [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ec [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ec [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ec [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ec [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ed [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_ed [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ed [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ed [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ed [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ed [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ed [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ed [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ee [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_ee [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ee [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ee [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ee [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ee [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ee [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ee [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ef [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_ef [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ef [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ef [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ef [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ef [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ef [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ef [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f1 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_f1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f4 [0], \oc8051_golden_model_1.n2913 [0]);
  buf(\oc8051_golden_model_1.PSW_f4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f4 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f5 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_f5 [1], \oc8051_golden_model_1.n2914 [1]);
  buf(\oc8051_golden_model_1.PSW_f5 [2], \oc8051_golden_model_1.n2914 [2]);
  buf(\oc8051_golden_model_1.PSW_f5 [3], \oc8051_golden_model_1.n2914 [3]);
  buf(\oc8051_golden_model_1.PSW_f5 [4], \oc8051_golden_model_1.n2914 [4]);
  buf(\oc8051_golden_model_1.PSW_f5 [5], \oc8051_golden_model_1.n2914 [5]);
  buf(\oc8051_golden_model_1.PSW_f5 [6], \oc8051_golden_model_1.n2914 [6]);
  buf(\oc8051_golden_model_1.PSW_f5 [7], \oc8051_golden_model_1.n2914 [7]);
  buf(\oc8051_golden_model_1.PSW_f6 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_f6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f7 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_f7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f8 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_f8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f9 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_f9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_fa [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_fa [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_fa [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_fa [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_fa [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_fa [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_fa [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_fa [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_fb [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_fb [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_fb [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_fb [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_fb [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_fb [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_fb [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_fb [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_fc [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_fc [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_fc [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_fc [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_fc [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_fc [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_fc [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_fc [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_fd [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_fd [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_fd [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_fd [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_fd [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_fd [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_fd [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_fd [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_fe [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_fe [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_fe [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_fe [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_fe [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_fe [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_fe [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_fe [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ff [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_ff [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ff [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ff [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ff [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ff [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ff [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ff [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [0], \oc8051_golden_model_1.n2775 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [1], \oc8051_golden_model_1.n2774 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [2], \oc8051_golden_model_1.n2773 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [3], \oc8051_golden_model_1.n2772 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [4], \oc8051_golden_model_1.n2771 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [5], \oc8051_golden_model_1.n2770 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [6], \oc8051_golden_model_1.n2769 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [7], \oc8051_golden_model_1.n2768 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [0], \oc8051_golden_model_1.n2868 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [1], \oc8051_golden_model_1.n2867 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [2], \oc8051_golden_model_1.n2866 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [3], \oc8051_golden_model_1.n2865 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [4], \oc8051_golden_model_1.n2860 [4]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [5], \oc8051_golden_model_1.n2860 [5]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [6], \oc8051_golden_model_1.n2860 [6]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [7], \oc8051_golden_model_1.n2860 [7]);
  buf(\oc8051_golden_model_1.n0006 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0006 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0007 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0007 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0007 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0011 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0011 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0011 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0019 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0019 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0019 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0023 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0023 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0023 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0023 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0027 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0027 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0027 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0031 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0031 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0031 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0031 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0035 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0035 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0035 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0035 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0039 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0039 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0573 [0], \oc8051_golden_model_1.n2775 );
  buf(\oc8051_golden_model_1.n0573 [1], \oc8051_golden_model_1.n2774 );
  buf(\oc8051_golden_model_1.n0573 [2], \oc8051_golden_model_1.n2773 );
  buf(\oc8051_golden_model_1.n0573 [3], \oc8051_golden_model_1.n2772 );
  buf(\oc8051_golden_model_1.n0573 [4], \oc8051_golden_model_1.n2771 );
  buf(\oc8051_golden_model_1.n0573 [5], \oc8051_golden_model_1.n2770 );
  buf(\oc8051_golden_model_1.n0573 [6], \oc8051_golden_model_1.n2769 );
  buf(\oc8051_golden_model_1.n0573 [7], \oc8051_golden_model_1.n2768 );
  buf(\oc8051_golden_model_1.n0606 [0], \oc8051_golden_model_1.n2868 );
  buf(\oc8051_golden_model_1.n0606 [1], \oc8051_golden_model_1.n2867 );
  buf(\oc8051_golden_model_1.n0606 [2], \oc8051_golden_model_1.n2866 );
  buf(\oc8051_golden_model_1.n0606 [3], \oc8051_golden_model_1.n2865 );
  buf(\oc8051_golden_model_1.n0606 [4], \oc8051_golden_model_1.n2860 [4]);
  buf(\oc8051_golden_model_1.n0606 [5], \oc8051_golden_model_1.n2860 [5]);
  buf(\oc8051_golden_model_1.n0606 [6], \oc8051_golden_model_1.n2860 [6]);
  buf(\oc8051_golden_model_1.n0606 [7], \oc8051_golden_model_1.n2860 [7]);
  buf(\oc8051_golden_model_1.n0713 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n0713 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n0713 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n0713 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n0713 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n0713 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n0713 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n0713 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n0713 [8], 1'b0);
  buf(\oc8051_golden_model_1.n0713 [9], 1'b0);
  buf(\oc8051_golden_model_1.n0713 [10], 1'b0);
  buf(\oc8051_golden_model_1.n0713 [11], 1'b0);
  buf(\oc8051_golden_model_1.n0713 [12], 1'b0);
  buf(\oc8051_golden_model_1.n0713 [13], 1'b0);
  buf(\oc8051_golden_model_1.n0713 [14], 1'b0);
  buf(\oc8051_golden_model_1.n0713 [15], 1'b0);
  buf(\oc8051_golden_model_1.n0745 [0], \oc8051_golden_model_1.DPL [0]);
  buf(\oc8051_golden_model_1.n0745 [1], \oc8051_golden_model_1.DPL [1]);
  buf(\oc8051_golden_model_1.n0745 [2], \oc8051_golden_model_1.DPL [2]);
  buf(\oc8051_golden_model_1.n0745 [3], \oc8051_golden_model_1.DPL [3]);
  buf(\oc8051_golden_model_1.n0745 [4], \oc8051_golden_model_1.DPL [4]);
  buf(\oc8051_golden_model_1.n0745 [5], \oc8051_golden_model_1.DPL [5]);
  buf(\oc8051_golden_model_1.n0745 [6], \oc8051_golden_model_1.DPL [6]);
  buf(\oc8051_golden_model_1.n0745 [7], \oc8051_golden_model_1.DPL [7]);
  buf(\oc8051_golden_model_1.n0745 [8], \oc8051_golden_model_1.DPH [0]);
  buf(\oc8051_golden_model_1.n0745 [9], \oc8051_golden_model_1.DPH [1]);
  buf(\oc8051_golden_model_1.n0745 [10], \oc8051_golden_model_1.DPH [2]);
  buf(\oc8051_golden_model_1.n0745 [11], \oc8051_golden_model_1.DPH [3]);
  buf(\oc8051_golden_model_1.n0745 [12], \oc8051_golden_model_1.DPH [4]);
  buf(\oc8051_golden_model_1.n0745 [13], \oc8051_golden_model_1.DPH [5]);
  buf(\oc8051_golden_model_1.n0745 [14], \oc8051_golden_model_1.DPH [6]);
  buf(\oc8051_golden_model_1.n0745 [15], \oc8051_golden_model_1.DPH [7]);
  buf(\oc8051_golden_model_1.n1004 [0], \oc8051_golden_model_1.n2775 );
  buf(\oc8051_golden_model_1.n1004 [1], \oc8051_golden_model_1.n2774 );
  buf(\oc8051_golden_model_1.n1004 [2], \oc8051_golden_model_1.n2773 );
  buf(\oc8051_golden_model_1.n1004 [3], \oc8051_golden_model_1.n2772 );
  buf(\oc8051_golden_model_1.n1004 [4], \oc8051_golden_model_1.n2771 );
  buf(\oc8051_golden_model_1.n1004 [5], \oc8051_golden_model_1.n2770 );
  buf(\oc8051_golden_model_1.n1004 [6], \oc8051_golden_model_1.n2769 );
  buf(\oc8051_golden_model_1.n1004 [7], \oc8051_golden_model_1.n2768 );
  buf(\oc8051_golden_model_1.n1004 [8], \oc8051_golden_model_1.P2 [0]);
  buf(\oc8051_golden_model_1.n1004 [9], \oc8051_golden_model_1.P2 [1]);
  buf(\oc8051_golden_model_1.n1004 [10], \oc8051_golden_model_1.P2 [2]);
  buf(\oc8051_golden_model_1.n1004 [11], \oc8051_golden_model_1.P2 [3]);
  buf(\oc8051_golden_model_1.n1004 [12], \oc8051_golden_model_1.P2 [4]);
  buf(\oc8051_golden_model_1.n1004 [13], \oc8051_golden_model_1.P2 [5]);
  buf(\oc8051_golden_model_1.n1004 [14], \oc8051_golden_model_1.P2 [6]);
  buf(\oc8051_golden_model_1.n1004 [15], \oc8051_golden_model_1.P2 [7]);
  buf(\oc8051_golden_model_1.n1008 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1008 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1008 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1008 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1008 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1008 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1008 [6], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1009 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1010 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1011 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1012 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1013 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1014 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1015 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1016 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1023 , \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.n1024 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.n1024 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1024 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1024 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1024 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1024 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1024 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1024 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1031 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1031 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1031 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1031 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1031 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1031 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1031 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1031 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1032 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1033 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1034 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1035 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1036 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1037 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1038 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1039 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1046 , \oc8051_golden_model_1.n1047 [0]);
  buf(\oc8051_golden_model_1.n1047 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1047 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1047 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1047 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1047 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1047 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1047 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1063 , \oc8051_golden_model_1.n1064 [0]);
  buf(\oc8051_golden_model_1.n1064 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1064 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1064 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1064 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1064 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1064 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1064 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1157 [0], \oc8051_golden_model_1.n2775 );
  buf(\oc8051_golden_model_1.n1157 [1], \oc8051_golden_model_1.n2774 );
  buf(\oc8051_golden_model_1.n1157 [2], \oc8051_golden_model_1.n2773 );
  buf(\oc8051_golden_model_1.n1157 [3], \oc8051_golden_model_1.n2772 );
  buf(\oc8051_golden_model_1.n1159 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1159 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1159 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1159 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1161 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1161 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1161 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1161 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1162 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1162 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1162 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1162 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1163 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1163 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1163 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1163 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1164 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1164 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1164 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1164 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1165 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1165 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1165 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1165 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1166 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1166 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1166 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1166 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1167 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1167 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1167 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1167 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1214 , \oc8051_golden_model_1.n2568 [7]);
  buf(\oc8051_golden_model_1.n1259 , \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1260 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1260 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1260 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1260 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1260 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1260 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1260 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1260 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1260 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1261 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1261 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1261 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1261 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1261 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1261 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1261 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1261 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1261 [8], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1262 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1262 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1262 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1262 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1262 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1262 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1262 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1262 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1263 , \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1264 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1264 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1264 [2], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1265 , \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1266 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1266 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1267 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1267 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1267 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1267 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1267 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1267 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1267 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1267 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1268 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1268 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1268 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1268 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1268 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1268 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1268 [6], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1269 , \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1270 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1271 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1272 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1273 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1274 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1275 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1276 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1283 , \oc8051_golden_model_1.n1284 [0]);
  buf(\oc8051_golden_model_1.n1284 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1284 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1284 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1284 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1284 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1284 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1284 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1300 , \oc8051_golden_model_1.n1301 [0]);
  buf(\oc8051_golden_model_1.n1301 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1301 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1301 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1301 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1301 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1301 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1301 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1343 [0], \oc8051_golden_model_1.n2868 );
  buf(\oc8051_golden_model_1.n1343 [1], \oc8051_golden_model_1.n2867 );
  buf(\oc8051_golden_model_1.n1343 [2], \oc8051_golden_model_1.n2866 );
  buf(\oc8051_golden_model_1.n1343 [3], \oc8051_golden_model_1.n2865 );
  buf(\oc8051_golden_model_1.n1343 [4], \oc8051_golden_model_1.n2860 [4]);
  buf(\oc8051_golden_model_1.n1343 [5], \oc8051_golden_model_1.n2860 [5]);
  buf(\oc8051_golden_model_1.n1343 [6], \oc8051_golden_model_1.n2860 [6]);
  buf(\oc8051_golden_model_1.n1343 [7], \oc8051_golden_model_1.n2860 [7]);
  buf(\oc8051_golden_model_1.n1343 [8], \oc8051_golden_model_1.n2775 );
  buf(\oc8051_golden_model_1.n1343 [9], \oc8051_golden_model_1.n2774 );
  buf(\oc8051_golden_model_1.n1343 [10], \oc8051_golden_model_1.n2773 );
  buf(\oc8051_golden_model_1.n1343 [11], \oc8051_golden_model_1.n2772 );
  buf(\oc8051_golden_model_1.n1343 [12], \oc8051_golden_model_1.n2771 );
  buf(\oc8051_golden_model_1.n1343 [13], \oc8051_golden_model_1.n2770 );
  buf(\oc8051_golden_model_1.n1343 [14], \oc8051_golden_model_1.n2769 );
  buf(\oc8051_golden_model_1.n1343 [15], \oc8051_golden_model_1.n2768 );
  buf(\oc8051_golden_model_1.n1345 [0], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1345 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1345 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1345 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1345 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1345 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1345 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1345 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1346 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1347 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1348 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1349 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1350 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1351 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1352 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1353 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1360 , \oc8051_golden_model_1.n1361 [0]);
  buf(\oc8051_golden_model_1.n1361 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1361 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1361 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1361 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1361 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1361 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1361 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1363 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1363 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1363 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1363 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1363 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1363 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1363 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1363 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1363 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1367 [8], \oc8051_golden_model_1.n1402 [7]);
  buf(\oc8051_golden_model_1.n1368 , \oc8051_golden_model_1.n1402 [7]);
  buf(\oc8051_golden_model_1.n1369 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1369 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1369 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1369 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1370 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1370 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1370 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1370 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1370 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1374 [4], \oc8051_golden_model_1.n1402 [6]);
  buf(\oc8051_golden_model_1.n1375 , \oc8051_golden_model_1.n1402 [6]);
  buf(\oc8051_golden_model_1.n1376 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1376 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1376 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1376 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1376 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1376 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1376 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1376 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1376 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1384 , \oc8051_golden_model_1.n1402 [2]);
  buf(\oc8051_golden_model_1.n1385 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1385 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1385 [2], \oc8051_golden_model_1.n1402 [2]);
  buf(\oc8051_golden_model_1.n1385 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1385 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1385 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1385 [6], \oc8051_golden_model_1.n1402 [6]);
  buf(\oc8051_golden_model_1.n1385 [7], \oc8051_golden_model_1.n1402 [7]);
  buf(\oc8051_golden_model_1.n1386 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1386 [1], \oc8051_golden_model_1.n1402 [2]);
  buf(\oc8051_golden_model_1.n1386 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1386 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1386 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1386 [5], \oc8051_golden_model_1.n1402 [6]);
  buf(\oc8051_golden_model_1.n1386 [6], \oc8051_golden_model_1.n1402 [7]);
  buf(\oc8051_golden_model_1.n1401 , \oc8051_golden_model_1.n1402 [0]);
  buf(\oc8051_golden_model_1.n1402 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1402 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1402 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1402 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1424 [8], \oc8051_golden_model_1.n1457 [7]);
  buf(\oc8051_golden_model_1.n1425 , \oc8051_golden_model_1.n1457 [7]);
  buf(\oc8051_golden_model_1.n1430 [4], \oc8051_golden_model_1.n1457 [6]);
  buf(\oc8051_golden_model_1.n1431 , \oc8051_golden_model_1.n1457 [6]);
  buf(\oc8051_golden_model_1.n1439 , \oc8051_golden_model_1.n1457 [2]);
  buf(\oc8051_golden_model_1.n1440 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1440 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1440 [2], \oc8051_golden_model_1.n1457 [2]);
  buf(\oc8051_golden_model_1.n1440 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1440 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1440 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1440 [6], \oc8051_golden_model_1.n1457 [6]);
  buf(\oc8051_golden_model_1.n1440 [7], \oc8051_golden_model_1.n1457 [7]);
  buf(\oc8051_golden_model_1.n1441 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1441 [1], \oc8051_golden_model_1.n1457 [2]);
  buf(\oc8051_golden_model_1.n1441 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1441 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1441 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1441 [5], \oc8051_golden_model_1.n1457 [6]);
  buf(\oc8051_golden_model_1.n1441 [6], \oc8051_golden_model_1.n1457 [7]);
  buf(\oc8051_golden_model_1.n1456 , \oc8051_golden_model_1.n1457 [0]);
  buf(\oc8051_golden_model_1.n1457 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1457 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1457 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1457 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1459 [0], \oc8051_golden_model_1.n2868 );
  buf(\oc8051_golden_model_1.n1459 [1], \oc8051_golden_model_1.n2867 );
  buf(\oc8051_golden_model_1.n1459 [2], \oc8051_golden_model_1.n2866 );
  buf(\oc8051_golden_model_1.n1459 [3], \oc8051_golden_model_1.n2865 );
  buf(\oc8051_golden_model_1.n1459 [4], \oc8051_golden_model_1.n2860 [4]);
  buf(\oc8051_golden_model_1.n1459 [5], \oc8051_golden_model_1.n2860 [5]);
  buf(\oc8051_golden_model_1.n1459 [6], \oc8051_golden_model_1.n2860 [6]);
  buf(\oc8051_golden_model_1.n1459 [7], \oc8051_golden_model_1.n2860 [7]);
  buf(\oc8051_golden_model_1.n1459 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1461 [8], \oc8051_golden_model_1.n1493 [7]);
  buf(\oc8051_golden_model_1.n1462 , \oc8051_golden_model_1.n1493 [7]);
  buf(\oc8051_golden_model_1.n1463 [0], \oc8051_golden_model_1.n2868 );
  buf(\oc8051_golden_model_1.n1463 [1], \oc8051_golden_model_1.n2867 );
  buf(\oc8051_golden_model_1.n1463 [2], \oc8051_golden_model_1.n2866 );
  buf(\oc8051_golden_model_1.n1463 [3], \oc8051_golden_model_1.n2865 );
  buf(\oc8051_golden_model_1.n1464 [0], \oc8051_golden_model_1.n2868 );
  buf(\oc8051_golden_model_1.n1464 [1], \oc8051_golden_model_1.n2867 );
  buf(\oc8051_golden_model_1.n1464 [2], \oc8051_golden_model_1.n2866 );
  buf(\oc8051_golden_model_1.n1464 [3], \oc8051_golden_model_1.n2865 );
  buf(\oc8051_golden_model_1.n1464 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1466 [4], \oc8051_golden_model_1.n1507 [6]);
  buf(\oc8051_golden_model_1.n1467 , \oc8051_golden_model_1.n1507 [6]);
  buf(\oc8051_golden_model_1.n1468 [0], \oc8051_golden_model_1.n2868 );
  buf(\oc8051_golden_model_1.n1468 [1], \oc8051_golden_model_1.n2867 );
  buf(\oc8051_golden_model_1.n1468 [2], \oc8051_golden_model_1.n2866 );
  buf(\oc8051_golden_model_1.n1468 [3], \oc8051_golden_model_1.n2865 );
  buf(\oc8051_golden_model_1.n1468 [4], \oc8051_golden_model_1.n2860 [4]);
  buf(\oc8051_golden_model_1.n1468 [5], \oc8051_golden_model_1.n2860 [5]);
  buf(\oc8051_golden_model_1.n1468 [6], \oc8051_golden_model_1.n2860 [6]);
  buf(\oc8051_golden_model_1.n1468 [7], \oc8051_golden_model_1.n2860 [7]);
  buf(\oc8051_golden_model_1.n1468 [8], \oc8051_golden_model_1.n2860 [7]);
  buf(\oc8051_golden_model_1.n1475 , \oc8051_golden_model_1.n1493 [2]);
  buf(\oc8051_golden_model_1.n1476 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1476 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1476 [2], \oc8051_golden_model_1.n1493 [2]);
  buf(\oc8051_golden_model_1.n1476 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1476 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1476 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1476 [6], \oc8051_golden_model_1.n1507 [6]);
  buf(\oc8051_golden_model_1.n1476 [7], \oc8051_golden_model_1.n1493 [7]);
  buf(\oc8051_golden_model_1.n1477 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1477 [1], \oc8051_golden_model_1.n1493 [2]);
  buf(\oc8051_golden_model_1.n1477 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1477 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1477 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1477 [5], \oc8051_golden_model_1.n1507 [6]);
  buf(\oc8051_golden_model_1.n1477 [6], \oc8051_golden_model_1.n1493 [7]);
  buf(\oc8051_golden_model_1.n1492 , \oc8051_golden_model_1.n1507 [0]);
  buf(\oc8051_golden_model_1.n1493 [0], \oc8051_golden_model_1.n1507 [0]);
  buf(\oc8051_golden_model_1.n1493 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1493 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1493 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1493 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1493 [6], \oc8051_golden_model_1.n1507 [6]);
  buf(\oc8051_golden_model_1.n1496 [8], \oc8051_golden_model_1.n1507 [7]);
  buf(\oc8051_golden_model_1.n1497 , \oc8051_golden_model_1.n1507 [7]);
  buf(\oc8051_golden_model_1.n1504 , \oc8051_golden_model_1.n1507 [2]);
  buf(\oc8051_golden_model_1.n1505 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1505 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1505 [2], \oc8051_golden_model_1.n1507 [2]);
  buf(\oc8051_golden_model_1.n1505 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1505 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1505 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1505 [6], \oc8051_golden_model_1.n1507 [6]);
  buf(\oc8051_golden_model_1.n1505 [7], \oc8051_golden_model_1.n1507 [7]);
  buf(\oc8051_golden_model_1.n1506 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1506 [1], \oc8051_golden_model_1.n1507 [2]);
  buf(\oc8051_golden_model_1.n1506 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1506 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1506 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1506 [5], \oc8051_golden_model_1.n1507 [6]);
  buf(\oc8051_golden_model_1.n1506 [6], \oc8051_golden_model_1.n1507 [7]);
  buf(\oc8051_golden_model_1.n1507 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1507 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1507 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1507 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1509 [0], \oc8051_golden_model_1.n2775 );
  buf(\oc8051_golden_model_1.n1509 [1], \oc8051_golden_model_1.n2774 );
  buf(\oc8051_golden_model_1.n1509 [2], \oc8051_golden_model_1.n2773 );
  buf(\oc8051_golden_model_1.n1509 [3], \oc8051_golden_model_1.n2772 );
  buf(\oc8051_golden_model_1.n1509 [4], \oc8051_golden_model_1.n2771 );
  buf(\oc8051_golden_model_1.n1509 [5], \oc8051_golden_model_1.n2770 );
  buf(\oc8051_golden_model_1.n1509 [6], \oc8051_golden_model_1.n2769 );
  buf(\oc8051_golden_model_1.n1509 [7], \oc8051_golden_model_1.n2768 );
  buf(\oc8051_golden_model_1.n1509 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1511 [8], \oc8051_golden_model_1.n1548 [7]);
  buf(\oc8051_golden_model_1.n1512 , \oc8051_golden_model_1.n1548 [7]);
  buf(\oc8051_golden_model_1.n1513 [0], \oc8051_golden_model_1.n2775 );
  buf(\oc8051_golden_model_1.n1513 [1], \oc8051_golden_model_1.n2774 );
  buf(\oc8051_golden_model_1.n1513 [2], \oc8051_golden_model_1.n2773 );
  buf(\oc8051_golden_model_1.n1513 [3], \oc8051_golden_model_1.n2772 );
  buf(\oc8051_golden_model_1.n1513 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1515 [4], \oc8051_golden_model_1.n1564 [6]);
  buf(\oc8051_golden_model_1.n1516 , \oc8051_golden_model_1.n1564 [6]);
  buf(\oc8051_golden_model_1.n1517 [0], \oc8051_golden_model_1.n2775 );
  buf(\oc8051_golden_model_1.n1517 [1], \oc8051_golden_model_1.n2774 );
  buf(\oc8051_golden_model_1.n1517 [2], \oc8051_golden_model_1.n2773 );
  buf(\oc8051_golden_model_1.n1517 [3], \oc8051_golden_model_1.n2772 );
  buf(\oc8051_golden_model_1.n1517 [4], \oc8051_golden_model_1.n2771 );
  buf(\oc8051_golden_model_1.n1517 [5], \oc8051_golden_model_1.n2770 );
  buf(\oc8051_golden_model_1.n1517 [6], \oc8051_golden_model_1.n2769 );
  buf(\oc8051_golden_model_1.n1517 [7], \oc8051_golden_model_1.n2768 );
  buf(\oc8051_golden_model_1.n1517 [8], \oc8051_golden_model_1.n2768 );
  buf(\oc8051_golden_model_1.n1524 , \oc8051_golden_model_1.n1548 [2]);
  buf(\oc8051_golden_model_1.n1525 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1525 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1525 [2], \oc8051_golden_model_1.n1548 [2]);
  buf(\oc8051_golden_model_1.n1525 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1525 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1525 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1525 [6], \oc8051_golden_model_1.n1564 [6]);
  buf(\oc8051_golden_model_1.n1525 [7], \oc8051_golden_model_1.n1548 [7]);
  buf(\oc8051_golden_model_1.n1526 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1526 [1], \oc8051_golden_model_1.n1548 [2]);
  buf(\oc8051_golden_model_1.n1526 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1526 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1526 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1526 [5], \oc8051_golden_model_1.n1564 [6]);
  buf(\oc8051_golden_model_1.n1526 [6], \oc8051_golden_model_1.n1548 [7]);
  buf(\oc8051_golden_model_1.n1541 , \oc8051_golden_model_1.n1564 [0]);
  buf(\oc8051_golden_model_1.n1542 [0], \oc8051_golden_model_1.n1564 [0]);
  buf(\oc8051_golden_model_1.n1542 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1542 [2], \oc8051_golden_model_1.n1548 [2]);
  buf(\oc8051_golden_model_1.n1542 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1542 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1542 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1542 [6], \oc8051_golden_model_1.n1564 [6]);
  buf(\oc8051_golden_model_1.n1542 [7], \oc8051_golden_model_1.n1548 [7]);
  buf(\oc8051_golden_model_1.n1544 [4], \oc8051_golden_model_1.n1561 [6]);
  buf(\oc8051_golden_model_1.n1545 , \oc8051_golden_model_1.n1561 [6]);
  buf(\oc8051_golden_model_1.n1546 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1546 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1546 [2], \oc8051_golden_model_1.n1548 [2]);
  buf(\oc8051_golden_model_1.n1546 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1546 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1546 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1546 [6], \oc8051_golden_model_1.n1561 [6]);
  buf(\oc8051_golden_model_1.n1546 [7], \oc8051_golden_model_1.n1548 [7]);
  buf(\oc8051_golden_model_1.n1547 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1547 [1], \oc8051_golden_model_1.n1548 [2]);
  buf(\oc8051_golden_model_1.n1547 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1547 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1547 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1547 [5], \oc8051_golden_model_1.n1561 [6]);
  buf(\oc8051_golden_model_1.n1547 [6], \oc8051_golden_model_1.n1548 [7]);
  buf(\oc8051_golden_model_1.n1548 [0], \oc8051_golden_model_1.n1564 [0]);
  buf(\oc8051_golden_model_1.n1548 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1548 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1548 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1548 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1548 [6], \oc8051_golden_model_1.n1561 [6]);
  buf(\oc8051_golden_model_1.n1550 [8], \oc8051_golden_model_1.n1564 [7]);
  buf(\oc8051_golden_model_1.n1551 , \oc8051_golden_model_1.n1564 [7]);
  buf(\oc8051_golden_model_1.n1558 , \oc8051_golden_model_1.n1564 [2]);
  buf(\oc8051_golden_model_1.n1559 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1559 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1559 [2], \oc8051_golden_model_1.n1564 [2]);
  buf(\oc8051_golden_model_1.n1559 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1559 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1559 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1559 [6], \oc8051_golden_model_1.n1561 [6]);
  buf(\oc8051_golden_model_1.n1559 [7], \oc8051_golden_model_1.n1564 [7]);
  buf(\oc8051_golden_model_1.n1560 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1560 [1], \oc8051_golden_model_1.n1564 [2]);
  buf(\oc8051_golden_model_1.n1560 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1560 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1560 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1560 [5], \oc8051_golden_model_1.n1561 [6]);
  buf(\oc8051_golden_model_1.n1560 [6], \oc8051_golden_model_1.n1564 [7]);
  buf(\oc8051_golden_model_1.n1561 [0], \oc8051_golden_model_1.n1564 [0]);
  buf(\oc8051_golden_model_1.n1561 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1561 [2], \oc8051_golden_model_1.n1564 [2]);
  buf(\oc8051_golden_model_1.n1561 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1561 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1561 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1561 [7], \oc8051_golden_model_1.n1564 [7]);
  buf(\oc8051_golden_model_1.n1562 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1562 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1562 [2], \oc8051_golden_model_1.n1564 [2]);
  buf(\oc8051_golden_model_1.n1562 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1562 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1562 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1562 [6], \oc8051_golden_model_1.n1564 [6]);
  buf(\oc8051_golden_model_1.n1562 [7], \oc8051_golden_model_1.n1564 [7]);
  buf(\oc8051_golden_model_1.n1563 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1563 [1], \oc8051_golden_model_1.n1564 [2]);
  buf(\oc8051_golden_model_1.n1563 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1563 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1563 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1563 [5], \oc8051_golden_model_1.n1564 [6]);
  buf(\oc8051_golden_model_1.n1563 [6], \oc8051_golden_model_1.n1564 [7]);
  buf(\oc8051_golden_model_1.n1564 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1564 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1564 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1564 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1567 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1567 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1567 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1567 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1567 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1567 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1567 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1567 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1567 [8], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1568 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1568 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1568 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1568 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1568 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1568 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1568 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1568 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1568 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1569 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1569 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1569 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1569 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1569 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1569 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1569 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1569 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1570 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1570 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1570 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1570 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1570 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1570 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1570 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1570 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1571 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1571 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1571 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1571 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1571 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1571 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1571 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1572 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1573 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1574 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1575 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1576 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1577 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1578 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1579 , \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1586 , \oc8051_golden_model_1.n1587 [0]);
  buf(\oc8051_golden_model_1.n1587 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1587 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1587 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1587 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1587 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1587 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1587 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1588 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1588 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1588 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1588 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1588 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1588 [5], 1'b0);
  buf(\oc8051_golden_model_1.n1588 [6], 1'b0);
  buf(\oc8051_golden_model_1.n1588 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1591 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1591 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1591 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1591 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1591 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1591 [5], 1'b0);
  buf(\oc8051_golden_model_1.n1591 [6], 1'b0);
  buf(\oc8051_golden_model_1.n1591 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1591 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1593 [8], \oc8051_golden_model_1.n1623 [7]);
  buf(\oc8051_golden_model_1.n1594 , \oc8051_golden_model_1.n1623 [7]);
  buf(\oc8051_golden_model_1.n1595 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1595 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1595 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1595 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1595 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1597 [4], \oc8051_golden_model_1.n1623 [6]);
  buf(\oc8051_golden_model_1.n1598 , \oc8051_golden_model_1.n1623 [6]);
  buf(\oc8051_golden_model_1.n1605 , \oc8051_golden_model_1.n1623 [2]);
  buf(\oc8051_golden_model_1.n1606 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1606 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1606 [2], \oc8051_golden_model_1.n1623 [2]);
  buf(\oc8051_golden_model_1.n1606 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1606 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1606 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1606 [6], \oc8051_golden_model_1.n1623 [6]);
  buf(\oc8051_golden_model_1.n1606 [7], \oc8051_golden_model_1.n1623 [7]);
  buf(\oc8051_golden_model_1.n1607 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1607 [1], \oc8051_golden_model_1.n1623 [2]);
  buf(\oc8051_golden_model_1.n1607 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1607 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1607 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1607 [5], \oc8051_golden_model_1.n1623 [6]);
  buf(\oc8051_golden_model_1.n1607 [6], \oc8051_golden_model_1.n1623 [7]);
  buf(\oc8051_golden_model_1.n1622 , \oc8051_golden_model_1.n1623 [0]);
  buf(\oc8051_golden_model_1.n1623 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1623 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1623 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1623 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1627 [8], \oc8051_golden_model_1.n1656 [7]);
  buf(\oc8051_golden_model_1.n1628 , \oc8051_golden_model_1.n1656 [7]);
  buf(\oc8051_golden_model_1.n1630 [4], \oc8051_golden_model_1.n1656 [6]);
  buf(\oc8051_golden_model_1.n1631 , \oc8051_golden_model_1.n1656 [6]);
  buf(\oc8051_golden_model_1.n1638 , \oc8051_golden_model_1.n1656 [2]);
  buf(\oc8051_golden_model_1.n1639 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1639 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1639 [2], \oc8051_golden_model_1.n1656 [2]);
  buf(\oc8051_golden_model_1.n1639 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1639 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1639 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1639 [6], \oc8051_golden_model_1.n1656 [6]);
  buf(\oc8051_golden_model_1.n1639 [7], \oc8051_golden_model_1.n1656 [7]);
  buf(\oc8051_golden_model_1.n1640 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1640 [1], \oc8051_golden_model_1.n1656 [2]);
  buf(\oc8051_golden_model_1.n1640 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1640 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1640 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1640 [5], \oc8051_golden_model_1.n1656 [6]);
  buf(\oc8051_golden_model_1.n1640 [6], \oc8051_golden_model_1.n1656 [7]);
  buf(\oc8051_golden_model_1.n1655 , \oc8051_golden_model_1.n1656 [0]);
  buf(\oc8051_golden_model_1.n1656 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1656 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1656 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1656 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1660 [8], \oc8051_golden_model_1.n1689 [7]);
  buf(\oc8051_golden_model_1.n1661 , \oc8051_golden_model_1.n1689 [7]);
  buf(\oc8051_golden_model_1.n1663 [4], \oc8051_golden_model_1.n1689 [6]);
  buf(\oc8051_golden_model_1.n1664 , \oc8051_golden_model_1.n1689 [6]);
  buf(\oc8051_golden_model_1.n1671 , \oc8051_golden_model_1.n1689 [2]);
  buf(\oc8051_golden_model_1.n1672 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1672 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1672 [2], \oc8051_golden_model_1.n1689 [2]);
  buf(\oc8051_golden_model_1.n1672 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1672 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1672 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1672 [6], \oc8051_golden_model_1.n1689 [6]);
  buf(\oc8051_golden_model_1.n1672 [7], \oc8051_golden_model_1.n1689 [7]);
  buf(\oc8051_golden_model_1.n1673 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1673 [1], \oc8051_golden_model_1.n1689 [2]);
  buf(\oc8051_golden_model_1.n1673 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1673 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1673 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1673 [5], \oc8051_golden_model_1.n1689 [6]);
  buf(\oc8051_golden_model_1.n1673 [6], \oc8051_golden_model_1.n1689 [7]);
  buf(\oc8051_golden_model_1.n1688 , \oc8051_golden_model_1.n1689 [0]);
  buf(\oc8051_golden_model_1.n1689 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1689 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1689 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1689 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1693 [8], \oc8051_golden_model_1.n1722 [7]);
  buf(\oc8051_golden_model_1.n1694 , \oc8051_golden_model_1.n1722 [7]);
  buf(\oc8051_golden_model_1.n1696 [4], \oc8051_golden_model_1.n1722 [6]);
  buf(\oc8051_golden_model_1.n1697 , \oc8051_golden_model_1.n1722 [6]);
  buf(\oc8051_golden_model_1.n1704 , \oc8051_golden_model_1.n1722 [2]);
  buf(\oc8051_golden_model_1.n1705 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1705 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1705 [2], \oc8051_golden_model_1.n1722 [2]);
  buf(\oc8051_golden_model_1.n1705 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1705 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1705 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1705 [6], \oc8051_golden_model_1.n1722 [6]);
  buf(\oc8051_golden_model_1.n1705 [7], \oc8051_golden_model_1.n1722 [7]);
  buf(\oc8051_golden_model_1.n1706 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1706 [1], \oc8051_golden_model_1.n1722 [2]);
  buf(\oc8051_golden_model_1.n1706 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1706 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1706 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1706 [5], \oc8051_golden_model_1.n1722 [6]);
  buf(\oc8051_golden_model_1.n1706 [6], \oc8051_golden_model_1.n1722 [7]);
  buf(\oc8051_golden_model_1.n1721 , \oc8051_golden_model_1.n1722 [0]);
  buf(\oc8051_golden_model_1.n1722 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1722 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1722 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1722 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1747 [1], \oc8051_golden_model_1.n1749 [1]);
  buf(\oc8051_golden_model_1.n1747 [2], \oc8051_golden_model_1.n1749 [2]);
  buf(\oc8051_golden_model_1.n1747 [3], \oc8051_golden_model_1.n1749 [3]);
  buf(\oc8051_golden_model_1.n1747 [4], \oc8051_golden_model_1.n1749 [4]);
  buf(\oc8051_golden_model_1.n1747 [5], \oc8051_golden_model_1.n1749 [5]);
  buf(\oc8051_golden_model_1.n1747 [6], \oc8051_golden_model_1.n1749 [6]);
  buf(\oc8051_golden_model_1.n1747 [7], \oc8051_golden_model_1.n1749 [7]);
  buf(\oc8051_golden_model_1.n1748 [0], \oc8051_golden_model_1.n1749 [1]);
  buf(\oc8051_golden_model_1.n1748 [1], \oc8051_golden_model_1.n1749 [2]);
  buf(\oc8051_golden_model_1.n1748 [2], \oc8051_golden_model_1.n1749 [3]);
  buf(\oc8051_golden_model_1.n1748 [3], \oc8051_golden_model_1.n1749 [4]);
  buf(\oc8051_golden_model_1.n1748 [4], \oc8051_golden_model_1.n1749 [5]);
  buf(\oc8051_golden_model_1.n1748 [5], \oc8051_golden_model_1.n1749 [6]);
  buf(\oc8051_golden_model_1.n1748 [6], \oc8051_golden_model_1.n1749 [7]);
  buf(\oc8051_golden_model_1.n1749 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.n1804 , \oc8051_golden_model_1.n1805 [0]);
  buf(\oc8051_golden_model_1.n1805 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1805 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1805 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1805 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1805 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1805 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1805 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1821 , \oc8051_golden_model_1.n1822 [0]);
  buf(\oc8051_golden_model_1.n1822 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1822 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1822 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1822 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1822 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1822 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1822 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1838 , \oc8051_golden_model_1.n1839 [0]);
  buf(\oc8051_golden_model_1.n1839 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1839 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1839 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1839 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1839 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1839 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1839 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1855 , \oc8051_golden_model_1.n1856 [0]);
  buf(\oc8051_golden_model_1.n1856 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1856 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1856 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1856 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1856 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1856 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1856 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1879 [1], \oc8051_golden_model_1.n1881 [1]);
  buf(\oc8051_golden_model_1.n1879 [2], \oc8051_golden_model_1.n1881 [2]);
  buf(\oc8051_golden_model_1.n1879 [3], \oc8051_golden_model_1.n1881 [3]);
  buf(\oc8051_golden_model_1.n1879 [4], \oc8051_golden_model_1.n1881 [4]);
  buf(\oc8051_golden_model_1.n1879 [5], \oc8051_golden_model_1.n1881 [5]);
  buf(\oc8051_golden_model_1.n1879 [6], \oc8051_golden_model_1.n1881 [6]);
  buf(\oc8051_golden_model_1.n1879 [7], \oc8051_golden_model_1.n1881 [7]);
  buf(\oc8051_golden_model_1.n1880 [0], \oc8051_golden_model_1.n1881 [1]);
  buf(\oc8051_golden_model_1.n1880 [1], \oc8051_golden_model_1.n1881 [2]);
  buf(\oc8051_golden_model_1.n1880 [2], \oc8051_golden_model_1.n1881 [3]);
  buf(\oc8051_golden_model_1.n1880 [3], \oc8051_golden_model_1.n1881 [4]);
  buf(\oc8051_golden_model_1.n1880 [4], \oc8051_golden_model_1.n1881 [5]);
  buf(\oc8051_golden_model_1.n1880 [5], \oc8051_golden_model_1.n1881 [6]);
  buf(\oc8051_golden_model_1.n1880 [6], \oc8051_golden_model_1.n1881 [7]);
  buf(\oc8051_golden_model_1.n1881 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.n1936 , \oc8051_golden_model_1.n1937 [0]);
  buf(\oc8051_golden_model_1.n1937 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1937 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1937 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1937 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1937 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1937 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1937 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1953 , \oc8051_golden_model_1.n1954 [0]);
  buf(\oc8051_golden_model_1.n1954 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1954 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1954 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1954 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1954 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1954 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1954 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1970 , \oc8051_golden_model_1.n1971 [0]);
  buf(\oc8051_golden_model_1.n1971 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1971 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1971 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1971 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1971 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1971 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1971 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1987 , \oc8051_golden_model_1.n1988 [0]);
  buf(\oc8051_golden_model_1.n1988 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1988 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1988 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1988 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1988 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1988 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1988 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2085 , \oc8051_golden_model_1.n2086 [0]);
  buf(\oc8051_golden_model_1.n2086 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2086 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2086 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2086 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2086 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2086 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2086 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2102 , \oc8051_golden_model_1.n2103 [0]);
  buf(\oc8051_golden_model_1.n2103 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2103 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2103 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2103 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2103 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2103 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2103 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2119 , \oc8051_golden_model_1.n2120 [0]);
  buf(\oc8051_golden_model_1.n2120 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2120 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2120 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2120 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2120 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2120 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2120 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2136 , \oc8051_golden_model_1.n2137 [0]);
  buf(\oc8051_golden_model_1.n2137 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2137 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2137 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2137 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2137 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2137 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2137 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2141 , \oc8051_golden_model_1.n2145 [7]);
  buf(\oc8051_golden_model_1.n2142 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2142 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2142 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2142 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2142 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2142 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2142 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2143 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2143 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2143 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2143 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2143 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2143 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2143 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2143 [7], \oc8051_golden_model_1.n2145 [7]);
  buf(\oc8051_golden_model_1.n2144 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2144 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2144 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2144 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2144 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2144 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2144 [6], \oc8051_golden_model_1.n2145 [7]);
  buf(\oc8051_golden_model_1.n2145 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.n2145 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2145 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2145 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2145 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2145 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2145 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2160 , \oc8051_golden_model_1.n2161 [0]);
  buf(\oc8051_golden_model_1.n2161 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2161 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2161 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2161 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2161 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2161 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2161 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2200 , \oc8051_golden_model_1.n2203 [7]);
  buf(\oc8051_golden_model_1.n2201 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2201 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2201 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2201 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2201 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2201 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2201 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2201 [7], \oc8051_golden_model_1.n2203 [7]);
  buf(\oc8051_golden_model_1.n2202 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2202 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2202 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2202 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2202 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2202 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2202 [6], \oc8051_golden_model_1.n2203 [7]);
  buf(\oc8051_golden_model_1.n2203 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.n2203 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2203 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2203 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2203 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2203 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2203 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2210 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2210 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2210 [2], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2210 [3], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2211 , \oc8051_golden_model_1.n2229 [2]);
  buf(\oc8051_golden_model_1.n2212 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2212 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2212 [2], \oc8051_golden_model_1.n2229 [2]);
  buf(\oc8051_golden_model_1.n2212 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2212 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2212 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2212 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2212 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2213 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2213 [1], \oc8051_golden_model_1.n2229 [2]);
  buf(\oc8051_golden_model_1.n2213 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2213 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2213 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2213 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2213 [6], 1'b0);
  buf(\oc8051_golden_model_1.n2228 , \oc8051_golden_model_1.n2229 [0]);
  buf(\oc8051_golden_model_1.n2229 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2229 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2229 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2229 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2229 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2229 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2441 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2441 [1], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2441 [2], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2441 [3], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2441 [4], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2441 [5], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2441 [6], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2441 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2444 , \oc8051_golden_model_1.n2470 [7]);
  buf(\oc8051_golden_model_1.n2446 , \oc8051_golden_model_1.n2470 [6]);
  buf(\oc8051_golden_model_1.n2452 , \oc8051_golden_model_1.n2470 [2]);
  buf(\oc8051_golden_model_1.n2453 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2453 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2453 [2], \oc8051_golden_model_1.n2470 [2]);
  buf(\oc8051_golden_model_1.n2453 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2453 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2453 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2453 [6], \oc8051_golden_model_1.n2470 [6]);
  buf(\oc8051_golden_model_1.n2453 [7], \oc8051_golden_model_1.n2470 [7]);
  buf(\oc8051_golden_model_1.n2454 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2454 [1], \oc8051_golden_model_1.n2470 [2]);
  buf(\oc8051_golden_model_1.n2454 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2454 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2454 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2454 [5], \oc8051_golden_model_1.n2470 [6]);
  buf(\oc8051_golden_model_1.n2454 [6], \oc8051_golden_model_1.n2470 [7]);
  buf(\oc8051_golden_model_1.n2469 , \oc8051_golden_model_1.n2470 [0]);
  buf(\oc8051_golden_model_1.n2470 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2470 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2470 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2470 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2474 , \oc8051_golden_model_1.n2500 [7]);
  buf(\oc8051_golden_model_1.n2476 , \oc8051_golden_model_1.n2500 [6]);
  buf(\oc8051_golden_model_1.n2482 , \oc8051_golden_model_1.n2500 [2]);
  buf(\oc8051_golden_model_1.n2483 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2483 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2483 [2], \oc8051_golden_model_1.n2500 [2]);
  buf(\oc8051_golden_model_1.n2483 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2483 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2483 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2483 [6], \oc8051_golden_model_1.n2500 [6]);
  buf(\oc8051_golden_model_1.n2483 [7], \oc8051_golden_model_1.n2500 [7]);
  buf(\oc8051_golden_model_1.n2484 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2484 [1], \oc8051_golden_model_1.n2500 [2]);
  buf(\oc8051_golden_model_1.n2484 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2484 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2484 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2484 [5], \oc8051_golden_model_1.n2500 [6]);
  buf(\oc8051_golden_model_1.n2484 [6], \oc8051_golden_model_1.n2500 [7]);
  buf(\oc8051_golden_model_1.n2499 , \oc8051_golden_model_1.n2500 [0]);
  buf(\oc8051_golden_model_1.n2500 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2500 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2500 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2500 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2504 , \oc8051_golden_model_1.n2530 [7]);
  buf(\oc8051_golden_model_1.n2506 , \oc8051_golden_model_1.n2530 [6]);
  buf(\oc8051_golden_model_1.n2512 , \oc8051_golden_model_1.n2530 [2]);
  buf(\oc8051_golden_model_1.n2513 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2513 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2513 [2], \oc8051_golden_model_1.n2530 [2]);
  buf(\oc8051_golden_model_1.n2513 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2513 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2513 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2513 [6], \oc8051_golden_model_1.n2530 [6]);
  buf(\oc8051_golden_model_1.n2513 [7], \oc8051_golden_model_1.n2530 [7]);
  buf(\oc8051_golden_model_1.n2514 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2514 [1], \oc8051_golden_model_1.n2530 [2]);
  buf(\oc8051_golden_model_1.n2514 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2514 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2514 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2514 [5], \oc8051_golden_model_1.n2530 [6]);
  buf(\oc8051_golden_model_1.n2514 [6], \oc8051_golden_model_1.n2530 [7]);
  buf(\oc8051_golden_model_1.n2529 , \oc8051_golden_model_1.n2530 [0]);
  buf(\oc8051_golden_model_1.n2530 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2530 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2530 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2530 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2534 , \oc8051_golden_model_1.n2560 [7]);
  buf(\oc8051_golden_model_1.n2536 , \oc8051_golden_model_1.n2560 [6]);
  buf(\oc8051_golden_model_1.n2542 , \oc8051_golden_model_1.n2560 [2]);
  buf(\oc8051_golden_model_1.n2543 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2543 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2543 [2], \oc8051_golden_model_1.n2560 [2]);
  buf(\oc8051_golden_model_1.n2543 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2543 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2543 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2543 [6], \oc8051_golden_model_1.n2560 [6]);
  buf(\oc8051_golden_model_1.n2543 [7], \oc8051_golden_model_1.n2560 [7]);
  buf(\oc8051_golden_model_1.n2544 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2544 [1], \oc8051_golden_model_1.n2560 [2]);
  buf(\oc8051_golden_model_1.n2544 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2544 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2544 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2544 [5], \oc8051_golden_model_1.n2560 [6]);
  buf(\oc8051_golden_model_1.n2544 [6], \oc8051_golden_model_1.n2560 [7]);
  buf(\oc8051_golden_model_1.n2559 , \oc8051_golden_model_1.n2560 [0]);
  buf(\oc8051_golden_model_1.n2560 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2560 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2560 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2560 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2562 , \oc8051_golden_model_1.n2565 [7]);
  buf(\oc8051_golden_model_1.n2563 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2563 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2563 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2563 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2563 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2563 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2563 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2563 [7], \oc8051_golden_model_1.n2565 [7]);
  buf(\oc8051_golden_model_1.n2564 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2564 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2564 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2564 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2564 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2564 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2564 [6], \oc8051_golden_model_1.n2565 [7]);
  buf(\oc8051_golden_model_1.n2565 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.n2565 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2565 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2565 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2565 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2565 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2565 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2566 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2566 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2566 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2566 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2566 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2566 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2566 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2566 [7], \oc8051_golden_model_1.n2568 [7]);
  buf(\oc8051_golden_model_1.n2567 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2567 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2567 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2567 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2567 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2567 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2567 [6], \oc8051_golden_model_1.n2568 [7]);
  buf(\oc8051_golden_model_1.n2568 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.n2568 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2568 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2568 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2568 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2568 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2568 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2572 [0], \oc8051_golden_model_1.B [0]);
  buf(\oc8051_golden_model_1.n2572 [1], \oc8051_golden_model_1.B [1]);
  buf(\oc8051_golden_model_1.n2572 [2], \oc8051_golden_model_1.B [2]);
  buf(\oc8051_golden_model_1.n2572 [3], \oc8051_golden_model_1.B [3]);
  buf(\oc8051_golden_model_1.n2572 [4], \oc8051_golden_model_1.B [4]);
  buf(\oc8051_golden_model_1.n2572 [5], \oc8051_golden_model_1.B [5]);
  buf(\oc8051_golden_model_1.n2572 [6], \oc8051_golden_model_1.B [6]);
  buf(\oc8051_golden_model_1.n2572 [7], \oc8051_golden_model_1.B [7]);
  buf(\oc8051_golden_model_1.n2572 [8], 1'b0);
  buf(\oc8051_golden_model_1.n2572 [9], 1'b0);
  buf(\oc8051_golden_model_1.n2572 [10], 1'b0);
  buf(\oc8051_golden_model_1.n2572 [11], 1'b0);
  buf(\oc8051_golden_model_1.n2572 [12], 1'b0);
  buf(\oc8051_golden_model_1.n2572 [13], 1'b0);
  buf(\oc8051_golden_model_1.n2572 [14], 1'b0);
  buf(\oc8051_golden_model_1.n2572 [15], 1'b0);
  buf(\oc8051_golden_model_1.n2578 , \oc8051_golden_model_1.n2596 [2]);
  buf(\oc8051_golden_model_1.n2579 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2579 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2579 [2], \oc8051_golden_model_1.n2596 [2]);
  buf(\oc8051_golden_model_1.n2579 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2579 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2579 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2579 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2579 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2580 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2580 [1], \oc8051_golden_model_1.n2596 [2]);
  buf(\oc8051_golden_model_1.n2580 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2580 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2580 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2580 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2580 [6], 1'b0);
  buf(\oc8051_golden_model_1.n2595 , \oc8051_golden_model_1.n2596 [0]);
  buf(\oc8051_golden_model_1.n2596 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2596 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2596 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2596 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2596 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2596 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2599 , \oc8051_golden_model_1.n2602 [7]);
  buf(\oc8051_golden_model_1.n2600 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2600 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2600 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2600 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2600 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2600 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2600 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2600 [7], \oc8051_golden_model_1.n2602 [7]);
  buf(\oc8051_golden_model_1.n2601 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2601 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2601 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2601 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2601 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2601 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2601 [6], \oc8051_golden_model_1.n2602 [7]);
  buf(\oc8051_golden_model_1.n2602 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.n2602 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2602 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2602 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2602 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2602 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2602 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2634 , \oc8051_golden_model_1.n2637 [7]);
  buf(\oc8051_golden_model_1.n2635 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2635 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2635 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2635 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2635 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2635 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2635 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2635 [7], \oc8051_golden_model_1.n2637 [7]);
  buf(\oc8051_golden_model_1.n2636 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2636 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2636 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2636 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2636 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2636 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2636 [6], \oc8051_golden_model_1.n2637 [7]);
  buf(\oc8051_golden_model_1.n2637 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.n2637 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2637 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2637 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2637 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2637 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2637 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2642 , \oc8051_golden_model_1.n2645 [7]);
  buf(\oc8051_golden_model_1.n2643 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2643 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2643 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2643 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2643 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2643 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2643 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2643 [7], \oc8051_golden_model_1.n2645 [7]);
  buf(\oc8051_golden_model_1.n2644 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2644 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2644 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2644 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2644 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2644 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2644 [6], \oc8051_golden_model_1.n2645 [7]);
  buf(\oc8051_golden_model_1.n2645 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.n2645 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2645 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2645 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2645 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2645 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2645 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2650 , \oc8051_golden_model_1.n2653 [7]);
  buf(\oc8051_golden_model_1.n2651 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2651 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2651 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2651 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2651 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2651 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2651 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2651 [7], \oc8051_golden_model_1.n2653 [7]);
  buf(\oc8051_golden_model_1.n2652 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2652 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2652 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2652 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2652 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2652 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2652 [6], \oc8051_golden_model_1.n2653 [7]);
  buf(\oc8051_golden_model_1.n2653 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.n2653 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2653 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2653 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2653 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2653 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2653 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2658 , \oc8051_golden_model_1.n2661 [7]);
  buf(\oc8051_golden_model_1.n2659 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2659 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2659 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2659 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2659 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2659 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2659 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2659 [7], \oc8051_golden_model_1.n2661 [7]);
  buf(\oc8051_golden_model_1.n2660 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2660 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2660 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2660 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2660 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2660 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2660 [6], \oc8051_golden_model_1.n2661 [7]);
  buf(\oc8051_golden_model_1.n2661 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.n2661 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2661 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2661 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2661 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2661 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2661 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2666 , \oc8051_golden_model_1.n2669 [7]);
  buf(\oc8051_golden_model_1.n2667 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2667 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2667 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2667 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2667 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2667 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2667 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2667 [7], \oc8051_golden_model_1.n2669 [7]);
  buf(\oc8051_golden_model_1.n2668 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2668 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2668 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2668 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2668 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2668 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2668 [6], \oc8051_golden_model_1.n2669 [7]);
  buf(\oc8051_golden_model_1.n2669 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.n2669 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2669 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2669 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2669 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2669 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2669 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2694 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2694 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2694 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2694 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2694 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2694 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2694 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2694 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2695 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2695 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2695 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2695 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2695 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2695 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2695 [6], 1'b0);
  buf(\oc8051_golden_model_1.n2696 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.n2696 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2696 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2696 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2696 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2696 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2696 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2696 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2697 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2697 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2697 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2697 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2698 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2698 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2698 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2698 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2698 [4], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n2698 [5], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n2698 [6], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n2698 [7], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n2699 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n2700 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n2701 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n2702 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n2703 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2704 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2705 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2706 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2713 , \oc8051_golden_model_1.n2714 [0]);
  buf(\oc8051_golden_model_1.n2714 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2714 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2714 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2714 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2714 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2714 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2714 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2734 [1], \oc8051_golden_model_1.n2914 [1]);
  buf(\oc8051_golden_model_1.n2734 [2], \oc8051_golden_model_1.n2914 [2]);
  buf(\oc8051_golden_model_1.n2734 [3], \oc8051_golden_model_1.n2914 [3]);
  buf(\oc8051_golden_model_1.n2734 [4], \oc8051_golden_model_1.n2914 [4]);
  buf(\oc8051_golden_model_1.n2734 [5], \oc8051_golden_model_1.n2914 [5]);
  buf(\oc8051_golden_model_1.n2734 [6], \oc8051_golden_model_1.n2914 [6]);
  buf(\oc8051_golden_model_1.n2734 [7], \oc8051_golden_model_1.n2914 [7]);
  buf(\oc8051_golden_model_1.n2735 [0], \oc8051_golden_model_1.n2914 [1]);
  buf(\oc8051_golden_model_1.n2735 [1], \oc8051_golden_model_1.n2914 [2]);
  buf(\oc8051_golden_model_1.n2735 [2], \oc8051_golden_model_1.n2914 [3]);
  buf(\oc8051_golden_model_1.n2735 [3], \oc8051_golden_model_1.n2914 [4]);
  buf(\oc8051_golden_model_1.n2735 [4], \oc8051_golden_model_1.n2914 [5]);
  buf(\oc8051_golden_model_1.n2735 [5], \oc8051_golden_model_1.n2914 [6]);
  buf(\oc8051_golden_model_1.n2735 [6], \oc8051_golden_model_1.n2914 [7]);
  buf(\oc8051_golden_model_1.n2750 , \oc8051_golden_model_1.n2896 [0]);
  buf(\oc8051_golden_model_1.n2751 [0], \oc8051_golden_model_1.n2896 [0]);
  buf(\oc8051_golden_model_1.n2751 [1], \oc8051_golden_model_1.n2914 [1]);
  buf(\oc8051_golden_model_1.n2751 [2], \oc8051_golden_model_1.n2914 [2]);
  buf(\oc8051_golden_model_1.n2751 [3], \oc8051_golden_model_1.n2914 [3]);
  buf(\oc8051_golden_model_1.n2751 [4], \oc8051_golden_model_1.n2914 [4]);
  buf(\oc8051_golden_model_1.n2751 [5], \oc8051_golden_model_1.n2914 [5]);
  buf(\oc8051_golden_model_1.n2751 [6], \oc8051_golden_model_1.n2914 [6]);
  buf(\oc8051_golden_model_1.n2751 [7], \oc8051_golden_model_1.n2914 [7]);
  buf(\oc8051_golden_model_1.n2752 , \oc8051_golden_model_1.n2860 [7]);
  buf(\oc8051_golden_model_1.n2753 , \oc8051_golden_model_1.n2860 [6]);
  buf(\oc8051_golden_model_1.n2754 , \oc8051_golden_model_1.n2860 [5]);
  buf(\oc8051_golden_model_1.n2755 , \oc8051_golden_model_1.n2860 [4]);
  buf(\oc8051_golden_model_1.n2756 , \oc8051_golden_model_1.n2865 );
  buf(\oc8051_golden_model_1.n2757 , \oc8051_golden_model_1.n2866 );
  buf(\oc8051_golden_model_1.n2758 , \oc8051_golden_model_1.n2867 );
  buf(\oc8051_golden_model_1.n2759 , \oc8051_golden_model_1.n2868 );
  buf(\oc8051_golden_model_1.n2766 , \oc8051_golden_model_1.n2767 [0]);
  buf(\oc8051_golden_model_1.n2767 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2767 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2767 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2767 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2767 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2767 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2767 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2782 , \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.n2783 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2783 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2783 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2783 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2783 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2783 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2783 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2815 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2815 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2815 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2815 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2815 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2815 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2815 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2815 [7], 1'b1);
  buf(\oc8051_golden_model_1.n2816 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2816 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2816 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2816 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2816 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2816 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2816 [6], 1'b1);
  buf(\oc8051_golden_model_1.n2817 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.n2817 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2817 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2817 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2817 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2817 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2817 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2817 [7], 1'b1);
  buf(\oc8051_golden_model_1.n2836 , \oc8051_golden_model_1.n2854 [7]);
  buf(\oc8051_golden_model_1.n2837 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2837 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2837 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2837 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2837 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2837 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2837 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2837 [7], \oc8051_golden_model_1.n2854 [7]);
  buf(\oc8051_golden_model_1.n2838 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2838 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2838 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2838 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2838 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2838 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2838 [6], \oc8051_golden_model_1.n2854 [7]);
  buf(\oc8051_golden_model_1.n2853 , \oc8051_golden_model_1.n2854 [0]);
  buf(\oc8051_golden_model_1.n2854 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2854 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2854 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2854 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2854 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2854 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2858 [0], \oc8051_golden_model_1.n2868 );
  buf(\oc8051_golden_model_1.n2858 [1], \oc8051_golden_model_1.n2867 );
  buf(\oc8051_golden_model_1.n2858 [2], \oc8051_golden_model_1.n2866 );
  buf(\oc8051_golden_model_1.n2858 [3], \oc8051_golden_model_1.n2865 );
  buf(\oc8051_golden_model_1.n2858 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2858 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2858 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2858 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2859 [0], \oc8051_golden_model_1.n2860 [4]);
  buf(\oc8051_golden_model_1.n2859 [1], \oc8051_golden_model_1.n2860 [5]);
  buf(\oc8051_golden_model_1.n2859 [2], \oc8051_golden_model_1.n2860 [6]);
  buf(\oc8051_golden_model_1.n2859 [3], \oc8051_golden_model_1.n2860 [7]);
  buf(\oc8051_golden_model_1.n2860 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n2860 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n2860 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n2860 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n2861 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2862 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2863 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2864 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2875 , \oc8051_golden_model_1.n2876 [0]);
  buf(\oc8051_golden_model_1.n2876 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2876 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2876 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2876 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2876 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2876 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2876 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2894 , \oc8051_golden_model_1.n2895 [0]);
  buf(\oc8051_golden_model_1.n2895 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2895 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2895 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2895 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2895 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2895 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2895 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2896 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2896 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2896 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2896 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2896 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2896 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2896 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2912 , \oc8051_golden_model_1.n2913 [0]);
  buf(\oc8051_golden_model_1.n2913 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2913 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2913 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2913 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2913 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2913 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2913 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_top_1.sub_result [0], ABINPUT[27]);
  buf(\oc8051_top_1.sub_result [1], ABINPUT[28]);
  buf(\oc8051_top_1.sub_result [2], ABINPUT[29]);
  buf(\oc8051_top_1.sub_result [3], ABINPUT[30]);
  buf(\oc8051_top_1.sub_result [4], ABINPUT[31]);
  buf(\oc8051_top_1.sub_result [5], ABINPUT[32]);
  buf(\oc8051_top_1.sub_result [6], ABINPUT[33]);
  buf(\oc8051_top_1.sub_result [7], ABINPUT[34]);
  buf(\oc8051_top_1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.rd_ind , \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  buf(\oc8051_top_1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.ABINPUT [0], ABINPUT[0]);
  buf(\oc8051_top_1.ABINPUT [1], ABINPUT[1]);
  buf(\oc8051_top_1.ABINPUT [2], ABINPUT[2]);
  buf(\oc8051_top_1.ABINPUT [3], ABINPUT[3]);
  buf(\oc8051_top_1.ABINPUT [4], ABINPUT[4]);
  buf(\oc8051_top_1.ABINPUT [5], ABINPUT[5]);
  buf(\oc8051_top_1.ABINPUT [6], ABINPUT[6]);
  buf(\oc8051_top_1.ABINPUT [7], ABINPUT[7]);
  buf(\oc8051_top_1.ABINPUT [8], ABINPUT[8]);
  buf(\oc8051_top_1.ABINPUT [9], ABINPUT[9]);
  buf(\oc8051_top_1.ABINPUT [10], ABINPUT[10]);
  buf(\oc8051_top_1.ABINPUT [11], ABINPUT[11]);
  buf(\oc8051_top_1.ABINPUT [12], ABINPUT[12]);
  buf(\oc8051_top_1.ABINPUT [13], ABINPUT[13]);
  buf(\oc8051_top_1.ABINPUT [14], ABINPUT[14]);
  buf(\oc8051_top_1.ABINPUT [15], ABINPUT[15]);
  buf(\oc8051_top_1.ABINPUT [16], ABINPUT[16]);
  buf(\oc8051_top_1.ABINPUT [17], ABINPUT[17]);
  buf(\oc8051_top_1.ABINPUT [18], ABINPUT[18]);
  buf(\oc8051_top_1.ABINPUT [19], ABINPUT[19]);
  buf(\oc8051_top_1.ABINPUT [20], ABINPUT[20]);
  buf(\oc8051_top_1.ABINPUT [21], ABINPUT[21]);
  buf(\oc8051_top_1.ABINPUT [22], ABINPUT[22]);
  buf(\oc8051_top_1.ABINPUT [23], ABINPUT[23]);
  buf(\oc8051_top_1.ABINPUT [24], ABINPUT[24]);
  buf(\oc8051_top_1.ABINPUT [25], ABINPUT[25]);
  buf(\oc8051_top_1.ABINPUT [26], ABINPUT[26]);
  buf(\oc8051_top_1.ABINPUT [27], ABINPUT[27]);
  buf(\oc8051_top_1.ABINPUT [28], ABINPUT[28]);
  buf(\oc8051_top_1.ABINPUT [29], ABINPUT[29]);
  buf(\oc8051_top_1.ABINPUT [30], ABINPUT[30]);
  buf(\oc8051_top_1.ABINPUT [31], ABINPUT[31]);
  buf(\oc8051_top_1.ABINPUT [32], ABINPUT[32]);
  buf(\oc8051_top_1.ABINPUT [33], ABINPUT[33]);
  buf(\oc8051_top_1.ABINPUT [34], ABINPUT[34]);
  buf(\oc8051_top_1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.desOv , ABINPUT[2]);
  buf(\oc8051_top_1.desAc , ABINPUT[1]);
  buf(\oc8051_top_1.desCy , ABINPUT[0]);
  buf(\oc8051_top_1.des2 [0], ABINPUT[11]);
  buf(\oc8051_top_1.des2 [1], ABINPUT[12]);
  buf(\oc8051_top_1.des2 [2], ABINPUT[13]);
  buf(\oc8051_top_1.des2 [3], ABINPUT[14]);
  buf(\oc8051_top_1.des2 [4], ABINPUT[15]);
  buf(\oc8051_top_1.des2 [5], ABINPUT[16]);
  buf(\oc8051_top_1.des2 [6], ABINPUT[17]);
  buf(\oc8051_top_1.des2 [7], ABINPUT[18]);
  buf(\oc8051_top_1.des1 [0], ABINPUT[3]);
  buf(\oc8051_top_1.des1 [1], ABINPUT[4]);
  buf(\oc8051_top_1.des1 [2], ABINPUT[5]);
  buf(\oc8051_top_1.des1 [3], ABINPUT[6]);
  buf(\oc8051_top_1.des1 [4], ABINPUT[7]);
  buf(\oc8051_top_1.des1 [5], ABINPUT[8]);
  buf(\oc8051_top_1.des1 [6], ABINPUT[9]);
  buf(\oc8051_top_1.des1 [7], ABINPUT[10]);
  buf(\oc8051_top_1.des_acc [0], ABINPUT[19]);
  buf(\oc8051_top_1.des_acc [1], ABINPUT[20]);
  buf(\oc8051_top_1.des_acc [2], ABINPUT[21]);
  buf(\oc8051_top_1.des_acc [3], ABINPUT[22]);
  buf(\oc8051_top_1.des_acc [4], ABINPUT[23]);
  buf(\oc8051_top_1.des_acc [5], ABINPUT[24]);
  buf(\oc8051_top_1.des_acc [6], ABINPUT[25]);
  buf(\oc8051_top_1.des_acc [7], ABINPUT[26]);
  buf(\oc8051_top_1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.wb_rst_i , rst);
  buf(\oc8051_top_1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.wr_dat [0], ABINPUT[3]);
  buf(\oc8051_top_1.wr_dat [1], ABINPUT[4]);
  buf(\oc8051_top_1.wr_dat [2], ABINPUT[5]);
  buf(\oc8051_top_1.wr_dat [3], ABINPUT[6]);
  buf(\oc8051_top_1.wr_dat [4], ABINPUT[7]);
  buf(\oc8051_top_1.wr_dat [5], ABINPUT[8]);
  buf(\oc8051_top_1.wr_dat [6], ABINPUT[9]);
  buf(\oc8051_top_1.wr_dat [7], ABINPUT[10]);
  buf(\oc8051_top_1.sfr_out [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.sfr_out [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.sfr_out [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.sfr_out [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.sfr_out [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.sfr_out [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.sfr_out [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.sfr_out [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.src_sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.src_sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.wb_clk_i , clk);
  buf(\oc8051_top_1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.p3_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.p3_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.p3_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.p3_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.p3_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.p3_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.p3_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.p3_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.p2_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.p2_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.p2_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.p2_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.p2_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.p2_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.p2_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.p2_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.p1_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.p1_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.p1_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.p1_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.p1_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.p1_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.p1_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.p1_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.p0_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.p0_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.p0_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.p0_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.p0_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.p0_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.p0_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.p0_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.cxrom_data_out [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.cxrom_data_out [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.cxrom_data_out [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.cxrom_data_out [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.cxrom_data_out [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.cxrom_data_out [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.cxrom_data_out [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.cxrom_data_out [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.cxrom_data_out [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.cxrom_data_out [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.cxrom_data_out [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.cxrom_data_out [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.cxrom_data_out [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.cxrom_data_out [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.cxrom_data_out [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.cxrom_data_out [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.cxrom_data_out [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.cxrom_data_out [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.cxrom_data_out [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.cxrom_data_out [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.cxrom_data_out [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.cxrom_data_out [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.cxrom_data_out [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.cxrom_data_out [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.cxrom_data_out [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.cxrom_data_out [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.cxrom_data_out [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.cxrom_data_out [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.cxrom_data_out [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.cxrom_data_out [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.cxrom_data_out [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.cxrom_data_out [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.wbd_adr_o [0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(\oc8051_top_1.wbd_adr_o [1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(\oc8051_top_1.wbd_adr_o [2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(\oc8051_top_1.wbd_adr_o [3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(\oc8051_top_1.wbd_adr_o [4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(\oc8051_top_1.wbd_adr_o [5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(\oc8051_top_1.wbd_adr_o [6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(\oc8051_top_1.wbd_adr_o [7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(\oc8051_top_1.wbd_adr_o [8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(\oc8051_top_1.wbd_adr_o [9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(\oc8051_top_1.wbd_adr_o [10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(\oc8051_top_1.wbd_adr_o [11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(\oc8051_top_1.wbd_adr_o [12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(\oc8051_top_1.wbd_adr_o [13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(\oc8051_top_1.wbd_adr_o [14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(\oc8051_top_1.wbd_adr_o [15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(\oc8051_top_1.wbd_dat_o [0], \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  buf(\oc8051_top_1.wbd_dat_o [1], \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  buf(\oc8051_top_1.wbd_dat_o [2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  buf(\oc8051_top_1.wbd_dat_o [3], \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  buf(\oc8051_top_1.wbd_dat_o [4], \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  buf(\oc8051_top_1.wbd_dat_o [5], \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  buf(\oc8051_top_1.wbd_dat_o [6], \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  buf(\oc8051_top_1.wbd_dat_o [7], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  buf(\oc8051_top_1.wbd_cyc_o , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.wbd_stb_o , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.wbd_we_o , \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  buf(\oc8051_top_1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(\oc8051_top_1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(\oc8051_top_1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(\oc8051_top_1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(\oc8051_top_1.ie [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(\oc8051_top_1.ie [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(\oc8051_top_1.ie [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(\oc8051_top_1.ie [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(\oc8051_top_1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.psw [0], psw_impl[0]);
  buf(\oc8051_top_1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_top_1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_top_1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_top_1.pc_log_prev [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_top_1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_top_1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_top_1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_top_1.pc_log_prev [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_top_1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_top_1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_top_1.pc_log_prev [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_top_1.pc_log_prev [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_top_1.pc_log_prev [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_top_1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_top_1.pc_log_prev [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_top_1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_top_1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_top_1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_top_1.pc_log [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_top_1.pc_log [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_top_1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_top_1.pc_log [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_top_1.pc_log [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_top_1.pc_log [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_top_1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_top_1.pc_log [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_top_1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_top_1.pc_log [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_top_1.pc_log [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_top_1.pc_log [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_top_1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_top_1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(rd_rom_0_addr[0], \oc8051_golden_model_1.PC [0]);
  buf(rd_rom_0_addr[1], \oc8051_golden_model_1.PC [1]);
  buf(rd_rom_0_addr[2], \oc8051_golden_model_1.PC [2]);
  buf(rd_rom_0_addr[3], \oc8051_golden_model_1.PC [3]);
  buf(rd_rom_0_addr[4], \oc8051_golden_model_1.PC [4]);
  buf(rd_rom_0_addr[5], \oc8051_golden_model_1.PC [5]);
  buf(rd_rom_0_addr[6], \oc8051_golden_model_1.PC [6]);
  buf(rd_rom_0_addr[7], \oc8051_golden_model_1.PC [7]);
  buf(rd_rom_0_addr[8], \oc8051_golden_model_1.PC [8]);
  buf(rd_rom_0_addr[9], \oc8051_golden_model_1.PC [9]);
  buf(rd_rom_0_addr[10], \oc8051_golden_model_1.PC [10]);
  buf(rd_rom_0_addr[11], \oc8051_golden_model_1.PC [11]);
  buf(rd_rom_0_addr[12], \oc8051_golden_model_1.PC [12]);
  buf(rd_rom_0_addr[13], \oc8051_golden_model_1.PC [13]);
  buf(rd_rom_0_addr[14], \oc8051_golden_model_1.PC [14]);
  buf(rd_rom_0_addr[15], \oc8051_golden_model_1.PC [15]);
  buf(TMOD_gm[0], \oc8051_golden_model_1.TMOD [0]);
  buf(TMOD_gm[1], \oc8051_golden_model_1.TMOD [1]);
  buf(TMOD_gm[2], \oc8051_golden_model_1.TMOD [2]);
  buf(TMOD_gm[3], \oc8051_golden_model_1.TMOD [3]);
  buf(TMOD_gm[4], \oc8051_golden_model_1.TMOD [4]);
  buf(TMOD_gm[5], \oc8051_golden_model_1.TMOD [5]);
  buf(TMOD_gm[6], \oc8051_golden_model_1.TMOD [6]);
  buf(TMOD_gm[7], \oc8051_golden_model_1.TMOD [7]);
  buf(TL1_gm[0], \oc8051_golden_model_1.TL1 [0]);
  buf(TL1_gm[1], \oc8051_golden_model_1.TL1 [1]);
  buf(TL1_gm[2], \oc8051_golden_model_1.TL1 [2]);
  buf(TL1_gm[3], \oc8051_golden_model_1.TL1 [3]);
  buf(TL1_gm[4], \oc8051_golden_model_1.TL1 [4]);
  buf(TL1_gm[5], \oc8051_golden_model_1.TL1 [5]);
  buf(TL1_gm[6], \oc8051_golden_model_1.TL1 [6]);
  buf(TL1_gm[7], \oc8051_golden_model_1.TL1 [7]);
  buf(TL0_gm[0], \oc8051_golden_model_1.TL0 [0]);
  buf(TL0_gm[1], \oc8051_golden_model_1.TL0 [1]);
  buf(TL0_gm[2], \oc8051_golden_model_1.TL0 [2]);
  buf(TL0_gm[3], \oc8051_golden_model_1.TL0 [3]);
  buf(TL0_gm[4], \oc8051_golden_model_1.TL0 [4]);
  buf(TL0_gm[5], \oc8051_golden_model_1.TL0 [5]);
  buf(TL0_gm[6], \oc8051_golden_model_1.TL0 [6]);
  buf(TL0_gm[7], \oc8051_golden_model_1.TL0 [7]);
  buf(TH1_gm[0], \oc8051_golden_model_1.TH1 [0]);
  buf(TH1_gm[1], \oc8051_golden_model_1.TH1 [1]);
  buf(TH1_gm[2], \oc8051_golden_model_1.TH1 [2]);
  buf(TH1_gm[3], \oc8051_golden_model_1.TH1 [3]);
  buf(TH1_gm[4], \oc8051_golden_model_1.TH1 [4]);
  buf(TH1_gm[5], \oc8051_golden_model_1.TH1 [5]);
  buf(TH1_gm[6], \oc8051_golden_model_1.TH1 [6]);
  buf(TH1_gm[7], \oc8051_golden_model_1.TH1 [7]);
  buf(TH0_gm[0], \oc8051_golden_model_1.TH0 [0]);
  buf(TH0_gm[1], \oc8051_golden_model_1.TH0 [1]);
  buf(TH0_gm[2], \oc8051_golden_model_1.TH0 [2]);
  buf(TH0_gm[3], \oc8051_golden_model_1.TH0 [3]);
  buf(TH0_gm[4], \oc8051_golden_model_1.TH0 [4]);
  buf(TH0_gm[5], \oc8051_golden_model_1.TH0 [5]);
  buf(TH0_gm[6], \oc8051_golden_model_1.TH0 [6]);
  buf(TH0_gm[7], \oc8051_golden_model_1.TH0 [7]);
  buf(TCON_gm[0], \oc8051_golden_model_1.TCON [0]);
  buf(TCON_gm[1], \oc8051_golden_model_1.TCON [1]);
  buf(TCON_gm[2], \oc8051_golden_model_1.TCON [2]);
  buf(TCON_gm[3], \oc8051_golden_model_1.TCON [3]);
  buf(TCON_gm[4], \oc8051_golden_model_1.TCON [4]);
  buf(TCON_gm[5], \oc8051_golden_model_1.TCON [5]);
  buf(TCON_gm[6], \oc8051_golden_model_1.TCON [6]);
  buf(TCON_gm[7], \oc8051_golden_model_1.TCON [7]);
  buf(SP_gm[0], \oc8051_golden_model_1.SP [0]);
  buf(SP_gm[1], \oc8051_golden_model_1.SP [1]);
  buf(SP_gm[2], \oc8051_golden_model_1.SP [2]);
  buf(SP_gm[3], \oc8051_golden_model_1.SP [3]);
  buf(SP_gm[4], \oc8051_golden_model_1.SP [4]);
  buf(SP_gm[5], \oc8051_golden_model_1.SP [5]);
  buf(SP_gm[6], \oc8051_golden_model_1.SP [6]);
  buf(SP_gm[7], \oc8051_golden_model_1.SP [7]);
  buf(SCON_gm[0], \oc8051_golden_model_1.SCON [0]);
  buf(SCON_gm[1], \oc8051_golden_model_1.SCON [1]);
  buf(SCON_gm[2], \oc8051_golden_model_1.SCON [2]);
  buf(SCON_gm[3], \oc8051_golden_model_1.SCON [3]);
  buf(SCON_gm[4], \oc8051_golden_model_1.SCON [4]);
  buf(SCON_gm[5], \oc8051_golden_model_1.SCON [5]);
  buf(SCON_gm[6], \oc8051_golden_model_1.SCON [6]);
  buf(SCON_gm[7], \oc8051_golden_model_1.SCON [7]);
  buf(SBUF_gm[0], \oc8051_golden_model_1.SBUF [0]);
  buf(SBUF_gm[1], \oc8051_golden_model_1.SBUF [1]);
  buf(SBUF_gm[2], \oc8051_golden_model_1.SBUF [2]);
  buf(SBUF_gm[3], \oc8051_golden_model_1.SBUF [3]);
  buf(SBUF_gm[4], \oc8051_golden_model_1.SBUF [4]);
  buf(SBUF_gm[5], \oc8051_golden_model_1.SBUF [5]);
  buf(SBUF_gm[6], \oc8051_golden_model_1.SBUF [6]);
  buf(SBUF_gm[7], \oc8051_golden_model_1.SBUF [7]);
  buf(PSW_gm[0], \oc8051_golden_model_1.PSW [0]);
  buf(PSW_gm[1], \oc8051_golden_model_1.PSW [1]);
  buf(PSW_gm[2], \oc8051_golden_model_1.PSW [2]);
  buf(PSW_gm[3], \oc8051_golden_model_1.PSW [3]);
  buf(PSW_gm[4], \oc8051_golden_model_1.PSW [4]);
  buf(PSW_gm[5], \oc8051_golden_model_1.PSW [5]);
  buf(PSW_gm[6], \oc8051_golden_model_1.PSW [6]);
  buf(PSW_gm[7], \oc8051_golden_model_1.PSW [7]);
  buf(PCON_gm[0], \oc8051_golden_model_1.PCON [0]);
  buf(PCON_gm[1], \oc8051_golden_model_1.PCON [1]);
  buf(PCON_gm[2], \oc8051_golden_model_1.PCON [2]);
  buf(PCON_gm[3], \oc8051_golden_model_1.PCON [3]);
  buf(PCON_gm[4], \oc8051_golden_model_1.PCON [4]);
  buf(PCON_gm[5], \oc8051_golden_model_1.PCON [5]);
  buf(PCON_gm[6], \oc8051_golden_model_1.PCON [6]);
  buf(PCON_gm[7], \oc8051_golden_model_1.PCON [7]);
  buf(P3_gm[0], \oc8051_golden_model_1.P3 [0]);
  buf(P3_gm[1], \oc8051_golden_model_1.P3 [1]);
  buf(P3_gm[2], \oc8051_golden_model_1.P3 [2]);
  buf(P3_gm[3], \oc8051_golden_model_1.P3 [3]);
  buf(P3_gm[4], \oc8051_golden_model_1.P3 [4]);
  buf(P3_gm[5], \oc8051_golden_model_1.P3 [5]);
  buf(P3_gm[6], \oc8051_golden_model_1.P3 [6]);
  buf(P3_gm[7], \oc8051_golden_model_1.P3 [7]);
  buf(P2_gm[0], \oc8051_golden_model_1.P2 [0]);
  buf(P2_gm[1], \oc8051_golden_model_1.P2 [1]);
  buf(P2_gm[2], \oc8051_golden_model_1.P2 [2]);
  buf(P2_gm[3], \oc8051_golden_model_1.P2 [3]);
  buf(P2_gm[4], \oc8051_golden_model_1.P2 [4]);
  buf(P2_gm[5], \oc8051_golden_model_1.P2 [5]);
  buf(P2_gm[6], \oc8051_golden_model_1.P2 [6]);
  buf(P2_gm[7], \oc8051_golden_model_1.P2 [7]);
  buf(P1_gm[0], \oc8051_golden_model_1.P1 [0]);
  buf(P1_gm[1], \oc8051_golden_model_1.P1 [1]);
  buf(P1_gm[2], \oc8051_golden_model_1.P1 [2]);
  buf(P1_gm[3], \oc8051_golden_model_1.P1 [3]);
  buf(P1_gm[4], \oc8051_golden_model_1.P1 [4]);
  buf(P1_gm[5], \oc8051_golden_model_1.P1 [5]);
  buf(P1_gm[6], \oc8051_golden_model_1.P1 [6]);
  buf(P1_gm[7], \oc8051_golden_model_1.P1 [7]);
  buf(P0_gm[0], \oc8051_golden_model_1.P0 [0]);
  buf(P0_gm[1], \oc8051_golden_model_1.P0 [1]);
  buf(P0_gm[2], \oc8051_golden_model_1.P0 [2]);
  buf(P0_gm[3], \oc8051_golden_model_1.P0 [3]);
  buf(P0_gm[4], \oc8051_golden_model_1.P0 [4]);
  buf(P0_gm[5], \oc8051_golden_model_1.P0 [5]);
  buf(P0_gm[6], \oc8051_golden_model_1.P0 [6]);
  buf(P0_gm[7], \oc8051_golden_model_1.P0 [7]);
  buf(IP_gm[0], \oc8051_golden_model_1.IP [0]);
  buf(IP_gm[1], \oc8051_golden_model_1.IP [1]);
  buf(IP_gm[2], \oc8051_golden_model_1.IP [2]);
  buf(IP_gm[3], \oc8051_golden_model_1.IP [3]);
  buf(IP_gm[4], \oc8051_golden_model_1.IP [4]);
  buf(IP_gm[5], \oc8051_golden_model_1.IP [5]);
  buf(IP_gm[6], \oc8051_golden_model_1.IP [6]);
  buf(IP_gm[7], \oc8051_golden_model_1.IP [7]);
  buf(IE_gm[0], \oc8051_golden_model_1.IE [0]);
  buf(IE_gm[1], \oc8051_golden_model_1.IE [1]);
  buf(IE_gm[2], \oc8051_golden_model_1.IE [2]);
  buf(IE_gm[3], \oc8051_golden_model_1.IE [3]);
  buf(IE_gm[4], \oc8051_golden_model_1.IE [4]);
  buf(IE_gm[5], \oc8051_golden_model_1.IE [5]);
  buf(IE_gm[6], \oc8051_golden_model_1.IE [6]);
  buf(IE_gm[7], \oc8051_golden_model_1.IE [7]);
  buf(DPH_gm[0], \oc8051_golden_model_1.DPH [0]);
  buf(DPH_gm[1], \oc8051_golden_model_1.DPH [1]);
  buf(DPH_gm[2], \oc8051_golden_model_1.DPH [2]);
  buf(DPH_gm[3], \oc8051_golden_model_1.DPH [3]);
  buf(DPH_gm[4], \oc8051_golden_model_1.DPH [4]);
  buf(DPH_gm[5], \oc8051_golden_model_1.DPH [5]);
  buf(DPH_gm[6], \oc8051_golden_model_1.DPH [6]);
  buf(DPH_gm[7], \oc8051_golden_model_1.DPH [7]);
  buf(DPL_gm[0], \oc8051_golden_model_1.DPL [0]);
  buf(DPL_gm[1], \oc8051_golden_model_1.DPL [1]);
  buf(DPL_gm[2], \oc8051_golden_model_1.DPL [2]);
  buf(DPL_gm[3], \oc8051_golden_model_1.DPL [3]);
  buf(DPL_gm[4], \oc8051_golden_model_1.DPL [4]);
  buf(DPL_gm[5], \oc8051_golden_model_1.DPL [5]);
  buf(DPL_gm[6], \oc8051_golden_model_1.DPL [6]);
  buf(DPL_gm[7], \oc8051_golden_model_1.DPL [7]);
  buf(B_gm[0], \oc8051_golden_model_1.B [0]);
  buf(B_gm[1], \oc8051_golden_model_1.B [1]);
  buf(B_gm[2], \oc8051_golden_model_1.B [2]);
  buf(B_gm[3], \oc8051_golden_model_1.B [3]);
  buf(B_gm[4], \oc8051_golden_model_1.B [4]);
  buf(B_gm[5], \oc8051_golden_model_1.B [5]);
  buf(B_gm[6], \oc8051_golden_model_1.B [6]);
  buf(B_gm[7], \oc8051_golden_model_1.B [7]);
  buf(ACC_gm[0], \oc8051_golden_model_1.ACC [0]);
  buf(ACC_gm[1], \oc8051_golden_model_1.ACC [1]);
  buf(ACC_gm[2], \oc8051_golden_model_1.ACC [2]);
  buf(ACC_gm[3], \oc8051_golden_model_1.ACC [3]);
  buf(ACC_gm[4], \oc8051_golden_model_1.ACC [4]);
  buf(ACC_gm[5], \oc8051_golden_model_1.ACC [5]);
  buf(ACC_gm[6], \oc8051_golden_model_1.ACC [6]);
  buf(ACC_gm[7], \oc8051_golden_model_1.ACC [7]);
  buf(dptr_impl[0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(dptr_impl[1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(dptr_impl[2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(dptr_impl[3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(dptr_impl[4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(dptr_impl[5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(dptr_impl[6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(dptr_impl[7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(dptr_impl[8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(dptr_impl[9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(dptr_impl[10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(dptr_impl[11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(dptr_impl[12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(dptr_impl[13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(dptr_impl[14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(dptr_impl[15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(b_reg_impl[0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(b_reg_impl[1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(b_reg_impl[2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(b_reg_impl[3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(b_reg_impl[4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(b_reg_impl[5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(b_reg_impl[6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(b_reg_impl[7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(acc_impl[0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(acc_impl[1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(acc_impl[2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(acc_impl[3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(acc_impl[4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(acc_impl[5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(acc_impl[6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(acc_impl[7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(psw_impl[1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(psw_impl[2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(psw_impl[3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(psw_impl[4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(psw_impl[5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(psw_impl[6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(psw_impl[7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(pc_impl[0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(pc_impl[1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(pc_impl[2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(pc_impl[3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(pc_impl[4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(pc_impl[5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(pc_impl[6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(pc_impl[7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(pc_impl[8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(pc_impl[9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(pc_impl[10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(pc_impl[11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(pc_impl[12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(pc_impl[13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(pc_impl[14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(pc_impl[15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(cxrom_data_out[0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(cxrom_data_out[1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(cxrom_data_out[2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(cxrom_data_out[3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(cxrom_data_out[4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(cxrom_data_out[5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(cxrom_data_out[6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(cxrom_data_out[7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(cxrom_data_out[8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(cxrom_data_out[9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(cxrom_data_out[10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(cxrom_data_out[11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(cxrom_data_out[12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(cxrom_data_out[13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(cxrom_data_out[14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(cxrom_data_out[15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(cxrom_data_out[16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(cxrom_data_out[17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(cxrom_data_out[18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(cxrom_data_out[19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(cxrom_data_out[20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(cxrom_data_out[21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(cxrom_data_out[22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(cxrom_data_out[23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(cxrom_data_out[24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(cxrom_data_out[25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(cxrom_data_out[26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(cxrom_data_out[27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(cxrom_data_out[28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(cxrom_data_out[29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(cxrom_data_out[30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(cxrom_data_out[31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(wbd_adr_o[0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(wbd_adr_o[1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(wbd_adr_o[2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(wbd_adr_o[3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(wbd_adr_o[4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(wbd_adr_o[5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(wbd_adr_o[6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(wbd_adr_o[7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(wbd_adr_o[8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(wbd_adr_o[9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(wbd_adr_o[10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(wbd_adr_o[11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(wbd_adr_o[12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(wbd_adr_o[13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(wbd_adr_o[14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(wbd_adr_o[15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(wbd_dat_o[0], \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  buf(wbd_dat_o[1], \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  buf(wbd_dat_o[2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  buf(wbd_dat_o[3], \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  buf(wbd_dat_o[4], \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  buf(wbd_dat_o[5], \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  buf(wbd_dat_o[6], \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  buf(wbd_dat_o[7], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  buf(wbd_cyc_o, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_stb_o, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_we_o, \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  buf(p3_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(p3_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(p3_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(p3_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(p3_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(p3_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(p3_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(p3_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(p2_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(p2_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(p2_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(p2_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(p2_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(p2_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(p2_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(p2_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(p1_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(p1_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(p1_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(p1_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(p1_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(p1_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(p1_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(p1_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(p0_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(p0_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(p0_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(p0_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(p0_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(p0_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(p0_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(p0_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
endmodule
