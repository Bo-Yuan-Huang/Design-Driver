
module oc8051_fv_top(clk, rst, word_in, p0_in, p1_in, p2_in, p3_in, rxd_i, t0_i, t1_i, t2_i, t2ex_i, property_invalid_jc, ABINPUT);
  wire _00000_;
  wire _00001_;
  wire _00002_;
  wire _00003_;
  wire _00004_;
  wire _00005_;
  wire _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  wire _08001_;
  wire _08002_;
  wire _08003_;
  wire _08004_;
  wire _08005_;
  wire _08006_;
  wire _08007_;
  wire _08008_;
  wire _08009_;
  wire _08010_;
  wire _08011_;
  wire _08012_;
  wire _08013_;
  wire _08014_;
  wire _08015_;
  wire _08016_;
  wire _08017_;
  wire _08018_;
  wire _08019_;
  wire _08020_;
  wire _08021_;
  wire _08022_;
  wire _08023_;
  wire _08024_;
  wire _08025_;
  wire _08026_;
  wire _08027_;
  wire _08028_;
  wire _08029_;
  wire _08030_;
  wire _08031_;
  wire _08032_;
  wire _08033_;
  wire _08034_;
  wire _08035_;
  wire _08036_;
  wire _08037_;
  wire _08038_;
  wire _08039_;
  wire _08040_;
  wire _08041_;
  wire _08042_;
  wire _08043_;
  wire _08044_;
  wire _08045_;
  wire _08046_;
  wire _08047_;
  wire _08048_;
  wire _08049_;
  wire _08050_;
  wire _08051_;
  wire _08052_;
  wire _08053_;
  wire _08054_;
  wire _08055_;
  wire _08056_;
  wire _08057_;
  wire _08058_;
  wire _08059_;
  wire _08060_;
  wire _08061_;
  wire _08062_;
  wire _08063_;
  wire _08064_;
  wire _08065_;
  wire _08066_;
  wire _08067_;
  wire _08068_;
  wire _08069_;
  wire _08070_;
  wire _08071_;
  wire _08072_;
  wire _08073_;
  wire _08074_;
  wire _08075_;
  wire _08076_;
  wire _08077_;
  wire _08078_;
  wire _08079_;
  wire _08080_;
  wire _08081_;
  wire _08082_;
  wire _08083_;
  wire _08084_;
  wire _08085_;
  wire _08086_;
  wire _08087_;
  wire _08088_;
  wire _08089_;
  wire _08090_;
  wire _08091_;
  wire _08092_;
  wire _08093_;
  wire _08094_;
  wire _08095_;
  wire _08096_;
  wire _08097_;
  wire _08098_;
  wire _08099_;
  wire _08100_;
  wire _08101_;
  wire _08102_;
  wire _08103_;
  wire _08104_;
  wire _08105_;
  wire _08106_;
  wire _08107_;
  wire _08108_;
  wire _08109_;
  wire _08110_;
  wire _08111_;
  wire _08112_;
  wire _08113_;
  wire _08114_;
  wire _08115_;
  wire _08116_;
  wire _08117_;
  wire _08118_;
  wire _08119_;
  wire _08120_;
  wire _08121_;
  wire _08122_;
  wire _08123_;
  wire _08124_;
  wire _08125_;
  wire _08126_;
  wire _08127_;
  wire _08128_;
  wire _08129_;
  wire _08130_;
  wire _08131_;
  wire _08132_;
  wire _08133_;
  wire _08134_;
  wire _08135_;
  wire _08136_;
  wire _08137_;
  wire _08138_;
  wire _08139_;
  wire _08140_;
  wire _08141_;
  wire _08142_;
  wire _08143_;
  wire _08144_;
  wire _08145_;
  wire _08146_;
  wire _08147_;
  wire _08148_;
  wire _08149_;
  wire _08150_;
  wire _08151_;
  wire _08152_;
  wire _08153_;
  wire _08154_;
  wire _08155_;
  wire _08156_;
  wire _08157_;
  wire _08158_;
  wire _08159_;
  wire _08160_;
  wire _08161_;
  wire _08162_;
  wire _08163_;
  wire _08164_;
  wire _08165_;
  wire _08166_;
  wire _08167_;
  wire _08168_;
  wire _08169_;
  wire _08170_;
  wire _08171_;
  wire _08172_;
  wire _08173_;
  wire _08174_;
  wire _08175_;
  wire _08176_;
  wire _08177_;
  wire _08178_;
  wire _08179_;
  wire _08180_;
  wire _08181_;
  wire _08182_;
  wire _08183_;
  wire _08184_;
  wire _08185_;
  wire _08186_;
  wire _08187_;
  wire _08188_;
  wire _08189_;
  wire _08190_;
  wire _08191_;
  wire _08192_;
  wire _08193_;
  wire _08194_;
  wire _08195_;
  wire _08196_;
  wire _08197_;
  wire _08198_;
  wire _08199_;
  wire _08200_;
  wire _08201_;
  wire _08202_;
  wire _08203_;
  wire _08204_;
  wire _08205_;
  wire _08206_;
  wire _08207_;
  wire _08208_;
  wire _08209_;
  wire _08210_;
  wire _08211_;
  wire _08212_;
  wire _08213_;
  wire _08214_;
  wire _08215_;
  wire _08216_;
  wire _08217_;
  wire _08218_;
  wire _08219_;
  wire _08220_;
  wire _08221_;
  wire _08222_;
  wire _08223_;
  wire _08224_;
  wire _08225_;
  wire _08226_;
  wire _08227_;
  wire _08228_;
  wire _08229_;
  wire _08230_;
  wire _08231_;
  wire _08232_;
  wire _08233_;
  wire _08234_;
  wire _08235_;
  wire _08236_;
  wire _08237_;
  wire _08238_;
  wire _08239_;
  wire _08240_;
  wire _08241_;
  wire _08242_;
  wire _08243_;
  wire _08244_;
  wire _08245_;
  wire _08246_;
  wire _08247_;
  wire _08248_;
  wire _08249_;
  wire _08250_;
  wire _08251_;
  wire _08252_;
  wire _08253_;
  wire _08254_;
  wire _08255_;
  wire _08256_;
  wire _08257_;
  wire _08258_;
  wire _08259_;
  wire _08260_;
  wire _08261_;
  wire _08262_;
  wire _08263_;
  wire _08264_;
  wire _08265_;
  wire _08266_;
  wire _08267_;
  wire _08268_;
  wire _08269_;
  wire _08270_;
  wire _08271_;
  wire _08272_;
  wire _08273_;
  wire _08274_;
  wire _08275_;
  wire _08276_;
  wire _08277_;
  wire _08278_;
  wire _08279_;
  wire _08280_;
  wire _08281_;
  wire _08282_;
  wire _08283_;
  wire _08284_;
  wire _08285_;
  wire _08286_;
  wire _08287_;
  wire _08288_;
  wire _08289_;
  wire _08290_;
  wire _08291_;
  wire _08292_;
  wire _08293_;
  wire _08294_;
  wire _08295_;
  wire _08296_;
  wire _08297_;
  wire _08298_;
  wire _08299_;
  wire _08300_;
  wire _08301_;
  wire _08302_;
  wire _08303_;
  wire _08304_;
  wire _08305_;
  wire _08306_;
  wire _08307_;
  wire _08308_;
  wire _08309_;
  wire _08310_;
  wire _08311_;
  wire _08312_;
  wire _08313_;
  wire _08314_;
  wire _08315_;
  wire _08316_;
  wire _08317_;
  wire _08318_;
  wire _08319_;
  wire _08320_;
  wire _08321_;
  wire _08322_;
  wire _08323_;
  wire _08324_;
  wire _08325_;
  wire _08326_;
  wire _08327_;
  wire _08328_;
  wire _08329_;
  wire _08330_;
  wire _08331_;
  wire _08332_;
  wire _08333_;
  wire _08334_;
  wire _08335_;
  wire _08336_;
  wire _08337_;
  wire _08338_;
  wire _08339_;
  wire _08340_;
  wire _08341_;
  wire _08342_;
  wire _08343_;
  wire _08344_;
  wire _08345_;
  wire _08346_;
  wire _08347_;
  wire _08348_;
  wire _08349_;
  wire _08350_;
  wire _08351_;
  wire _08352_;
  wire _08353_;
  wire _08354_;
  wire _08355_;
  wire _08356_;
  wire _08357_;
  wire _08358_;
  wire _08359_;
  wire _08360_;
  wire _08361_;
  wire _08362_;
  wire _08363_;
  wire _08364_;
  wire _08365_;
  wire _08366_;
  wire _08367_;
  wire _08368_;
  wire _08369_;
  wire _08370_;
  wire _08371_;
  wire _08372_;
  wire _08373_;
  wire _08374_;
  wire _08375_;
  wire _08376_;
  wire _08377_;
  wire _08378_;
  wire _08379_;
  wire _08380_;
  wire _08381_;
  wire _08382_;
  wire _08383_;
  wire _08384_;
  wire _08385_;
  wire _08386_;
  wire _08387_;
  wire _08388_;
  wire _08389_;
  wire _08390_;
  wire _08391_;
  wire _08392_;
  wire _08393_;
  wire _08394_;
  wire _08395_;
  wire _08396_;
  wire _08397_;
  wire _08398_;
  wire _08399_;
  wire _08400_;
  wire _08401_;
  wire _08402_;
  wire _08403_;
  wire _08404_;
  wire _08405_;
  wire _08406_;
  wire _08407_;
  wire _08408_;
  wire _08409_;
  wire _08410_;
  wire _08411_;
  wire _08412_;
  wire _08413_;
  wire _08414_;
  wire _08415_;
  wire _08416_;
  wire _08417_;
  wire _08418_;
  wire _08419_;
  wire _08420_;
  wire _08421_;
  wire _08422_;
  wire _08423_;
  wire _08424_;
  wire _08425_;
  wire _08426_;
  wire _08427_;
  wire _08428_;
  wire _08429_;
  wire _08430_;
  wire _08431_;
  wire _08432_;
  wire _08433_;
  wire _08434_;
  wire _08435_;
  wire _08436_;
  wire _08437_;
  wire _08438_;
  wire _08439_;
  wire _08440_;
  wire _08441_;
  wire _08442_;
  wire _08443_;
  wire _08444_;
  wire _08445_;
  wire _08446_;
  wire _08447_;
  wire _08448_;
  wire _08449_;
  wire _08450_;
  wire _08451_;
  wire _08452_;
  wire _08453_;
  wire _08454_;
  wire _08455_;
  wire _08456_;
  wire _08457_;
  wire _08458_;
  wire _08459_;
  wire _08460_;
  wire _08461_;
  wire _08462_;
  wire _08463_;
  wire _08464_;
  wire _08465_;
  wire _08466_;
  wire _08467_;
  wire _08468_;
  wire _08469_;
  wire _08470_;
  wire _08471_;
  wire _08472_;
  wire _08473_;
  wire _08474_;
  wire _08475_;
  wire _08476_;
  wire _08477_;
  wire _08478_;
  wire _08479_;
  wire _08480_;
  wire _08481_;
  wire _08482_;
  wire _08483_;
  wire _08484_;
  wire _08485_;
  wire _08486_;
  wire _08487_;
  wire _08488_;
  wire _08489_;
  wire _08490_;
  wire _08491_;
  wire _08492_;
  wire _08493_;
  wire _08494_;
  wire _08495_;
  wire _08496_;
  wire _08497_;
  wire _08498_;
  wire _08499_;
  wire _08500_;
  wire _08501_;
  wire _08502_;
  wire _08503_;
  wire _08504_;
  wire _08505_;
  wire _08506_;
  wire _08507_;
  wire _08508_;
  wire _08509_;
  wire _08510_;
  wire _08511_;
  wire _08512_;
  wire _08513_;
  wire _08514_;
  wire _08515_;
  wire _08516_;
  wire _08517_;
  wire _08518_;
  wire _08519_;
  wire _08520_;
  wire _08521_;
  wire _08522_;
  wire _08523_;
  wire _08524_;
  wire _08525_;
  wire _08526_;
  wire _08527_;
  wire _08528_;
  wire _08529_;
  wire _08530_;
  wire _08531_;
  wire _08532_;
  wire _08533_;
  wire _08534_;
  wire _08535_;
  wire _08536_;
  wire _08537_;
  wire _08538_;
  wire _08539_;
  wire _08540_;
  wire _08541_;
  wire _08542_;
  wire _08543_;
  wire _08544_;
  wire _08545_;
  wire _08546_;
  wire _08547_;
  wire _08548_;
  wire _08549_;
  wire _08550_;
  wire _08551_;
  wire _08552_;
  wire _08553_;
  wire _08554_;
  wire _08555_;
  wire _08556_;
  wire _08557_;
  wire _08558_;
  wire _08559_;
  wire _08560_;
  wire _08561_;
  wire _08562_;
  wire _08563_;
  wire _08564_;
  wire _08565_;
  wire _08566_;
  wire _08567_;
  wire _08568_;
  wire _08569_;
  wire _08570_;
  wire _08571_;
  wire _08572_;
  wire _08573_;
  wire _08574_;
  wire _08575_;
  wire _08576_;
  wire _08577_;
  wire _08578_;
  wire _08579_;
  wire _08580_;
  wire _08581_;
  wire _08582_;
  wire _08583_;
  wire _08584_;
  wire _08585_;
  wire _08586_;
  wire _08587_;
  wire _08588_;
  wire _08589_;
  wire _08590_;
  wire _08591_;
  wire _08592_;
  wire _08593_;
  wire _08594_;
  wire _08595_;
  wire _08596_;
  wire _08597_;
  wire _08598_;
  wire _08599_;
  wire _08600_;
  wire _08601_;
  wire _08602_;
  wire _08603_;
  wire _08604_;
  wire _08605_;
  wire _08606_;
  wire _08607_;
  wire _08608_;
  wire _08609_;
  wire _08610_;
  wire _08611_;
  wire _08612_;
  wire _08613_;
  wire _08614_;
  wire _08615_;
  wire _08616_;
  wire _08617_;
  wire _08618_;
  wire _08619_;
  wire _08620_;
  wire _08621_;
  wire _08622_;
  wire _08623_;
  wire _08624_;
  wire _08625_;
  wire _08626_;
  wire _08627_;
  wire _08628_;
  wire _08629_;
  wire _08630_;
  wire _08631_;
  wire _08632_;
  wire _08633_;
  wire _08634_;
  wire _08635_;
  wire _08636_;
  wire _08637_;
  wire _08638_;
  wire _08639_;
  wire _08640_;
  wire _08641_;
  wire _08642_;
  wire _08643_;
  wire _08644_;
  wire _08645_;
  wire _08646_;
  wire _08647_;
  wire _08648_;
  wire _08649_;
  wire _08650_;
  wire _08651_;
  wire _08652_;
  wire _08653_;
  wire _08654_;
  wire _08655_;
  wire _08656_;
  wire _08657_;
  wire _08658_;
  wire _08659_;
  wire _08660_;
  wire _08661_;
  wire _08662_;
  wire _08663_;
  wire _08664_;
  wire _08665_;
  wire _08666_;
  wire _08667_;
  wire _08668_;
  wire _08669_;
  wire _08670_;
  wire _08671_;
  wire _08672_;
  wire _08673_;
  wire _08674_;
  wire _08675_;
  wire _08676_;
  wire _08677_;
  wire _08678_;
  wire _08679_;
  wire _08680_;
  wire _08681_;
  wire _08682_;
  wire _08683_;
  wire _08684_;
  wire _08685_;
  wire _08686_;
  wire _08687_;
  wire _08688_;
  wire _08689_;
  wire _08690_;
  wire _08691_;
  wire _08692_;
  wire _08693_;
  wire _08694_;
  wire _08695_;
  wire _08696_;
  wire _08697_;
  wire _08698_;
  wire _08699_;
  wire _08700_;
  wire _08701_;
  wire _08702_;
  wire _08703_;
  wire _08704_;
  wire _08705_;
  wire _08706_;
  wire _08707_;
  wire _08708_;
  wire _08709_;
  wire _08710_;
  wire _08711_;
  wire _08712_;
  wire _08713_;
  wire _08714_;
  wire _08715_;
  wire _08716_;
  wire _08717_;
  wire _08718_;
  wire _08719_;
  wire _08720_;
  wire _08721_;
  wire _08722_;
  wire _08723_;
  wire _08724_;
  wire _08725_;
  wire _08726_;
  wire _08727_;
  wire _08728_;
  wire _08729_;
  wire _08730_;
  wire _08731_;
  wire _08732_;
  wire _08733_;
  wire _08734_;
  wire _08735_;
  wire _08736_;
  wire _08737_;
  wire _08738_;
  wire _08739_;
  wire _08740_;
  wire _08741_;
  wire _08742_;
  wire _08743_;
  wire _08744_;
  wire _08745_;
  wire _08746_;
  wire _08747_;
  wire _08748_;
  wire _08749_;
  wire _08750_;
  wire _08751_;
  wire _08752_;
  wire _08753_;
  wire _08754_;
  wire _08755_;
  wire _08756_;
  wire _08757_;
  wire _08758_;
  wire _08759_;
  wire _08760_;
  wire _08761_;
  wire _08762_;
  wire _08763_;
  wire _08764_;
  wire _08765_;
  wire _08766_;
  wire _08767_;
  wire _08768_;
  wire _08769_;
  wire _08770_;
  wire _08771_;
  wire _08772_;
  wire _08773_;
  wire _08774_;
  wire _08775_;
  wire _08776_;
  wire _08777_;
  wire _08778_;
  wire _08779_;
  wire _08780_;
  wire _08781_;
  wire _08782_;
  wire _08783_;
  wire _08784_;
  wire _08785_;
  wire _08786_;
  wire _08787_;
  wire _08788_;
  wire _08789_;
  wire _08790_;
  wire _08791_;
  wire _08792_;
  wire _08793_;
  wire _08794_;
  wire _08795_;
  wire _08796_;
  wire _08797_;
  wire _08798_;
  wire _08799_;
  wire _08800_;
  wire _08801_;
  wire _08802_;
  wire _08803_;
  wire _08804_;
  wire _08805_;
  wire _08806_;
  wire _08807_;
  wire _08808_;
  wire _08809_;
  wire _08810_;
  wire _08811_;
  wire _08812_;
  wire _08813_;
  wire _08814_;
  wire _08815_;
  wire _08816_;
  wire _08817_;
  wire _08818_;
  wire _08819_;
  wire _08820_;
  wire _08821_;
  wire _08822_;
  wire _08823_;
  wire _08824_;
  wire _08825_;
  wire _08826_;
  wire _08827_;
  wire _08828_;
  wire _08829_;
  wire _08830_;
  wire _08831_;
  wire _08832_;
  wire _08833_;
  wire _08834_;
  wire _08835_;
  wire _08836_;
  wire _08837_;
  wire _08838_;
  wire _08839_;
  wire _08840_;
  wire _08841_;
  wire _08842_;
  wire _08843_;
  wire _08844_;
  wire _08845_;
  wire _08846_;
  wire _08847_;
  wire _08848_;
  wire _08849_;
  wire _08850_;
  wire _08851_;
  wire _08852_;
  wire _08853_;
  wire _08854_;
  wire _08855_;
  wire _08856_;
  wire _08857_;
  wire _08858_;
  wire _08859_;
  wire _08860_;
  wire _08861_;
  wire _08862_;
  wire _08863_;
  wire _08864_;
  wire _08865_;
  wire _08866_;
  wire _08867_;
  wire _08868_;
  wire _08869_;
  wire _08870_;
  wire _08871_;
  wire _08872_;
  wire _08873_;
  wire _08874_;
  wire _08875_;
  wire _08876_;
  wire _08877_;
  wire _08878_;
  wire _08879_;
  wire _08880_;
  wire _08881_;
  wire _08882_;
  wire _08883_;
  wire _08884_;
  wire _08885_;
  wire _08886_;
  wire _08887_;
  wire _08888_;
  wire _08889_;
  wire _08890_;
  wire _08891_;
  wire _08892_;
  wire _08893_;
  wire _08894_;
  wire _08895_;
  wire _08896_;
  wire _08897_;
  wire _08898_;
  wire _08899_;
  wire _08900_;
  wire _08901_;
  wire _08902_;
  wire _08903_;
  wire _08904_;
  wire _08905_;
  wire _08906_;
  wire _08907_;
  wire _08908_;
  wire _08909_;
  wire _08910_;
  wire _08911_;
  wire _08912_;
  wire _08913_;
  wire _08914_;
  wire _08915_;
  wire _08916_;
  wire _08917_;
  wire _08918_;
  wire _08919_;
  wire _08920_;
  wire _08921_;
  wire _08922_;
  wire _08923_;
  wire _08924_;
  wire _08925_;
  wire _08926_;
  wire _08927_;
  wire _08928_;
  wire _08929_;
  wire _08930_;
  wire _08931_;
  wire _08932_;
  wire _08933_;
  wire _08934_;
  wire _08935_;
  wire _08936_;
  wire _08937_;
  wire _08938_;
  wire _08939_;
  wire _08940_;
  wire _08941_;
  wire _08942_;
  wire _08943_;
  wire _08944_;
  wire _08945_;
  wire _08946_;
  wire _08947_;
  wire _08948_;
  wire _08949_;
  wire _08950_;
  wire _08951_;
  wire _08952_;
  wire _08953_;
  wire _08954_;
  wire _08955_;
  wire _08956_;
  wire _08957_;
  wire _08958_;
  wire _08959_;
  wire _08960_;
  wire _08961_;
  wire _08962_;
  wire _08963_;
  wire _08964_;
  wire _08965_;
  wire _08966_;
  wire _08967_;
  wire _08968_;
  wire _08969_;
  wire _08970_;
  wire _08971_;
  wire _08972_;
  wire _08973_;
  wire _08974_;
  wire _08975_;
  wire _08976_;
  wire _08977_;
  wire _08978_;
  wire _08979_;
  wire _08980_;
  wire _08981_;
  wire _08982_;
  wire _08983_;
  wire _08984_;
  wire _08985_;
  wire _08986_;
  wire _08987_;
  wire _08988_;
  wire _08989_;
  wire _08990_;
  wire _08991_;
  wire _08992_;
  wire _08993_;
  wire _08994_;
  wire _08995_;
  wire _08996_;
  wire _08997_;
  wire _08998_;
  wire _08999_;
  wire _09000_;
  wire _09001_;
  wire _09002_;
  wire _09003_;
  wire _09004_;
  wire _09005_;
  wire _09006_;
  wire _09007_;
  wire _09008_;
  wire _09009_;
  wire _09010_;
  wire _09011_;
  wire _09012_;
  wire _09013_;
  wire _09014_;
  wire _09015_;
  wire _09016_;
  wire _09017_;
  wire _09018_;
  wire _09019_;
  wire _09020_;
  wire _09021_;
  wire _09022_;
  wire _09023_;
  wire _09024_;
  wire _09025_;
  wire _09026_;
  wire _09027_;
  wire _09028_;
  wire _09029_;
  wire _09030_;
  wire _09031_;
  wire _09032_;
  wire _09033_;
  wire _09034_;
  wire _09035_;
  wire _09036_;
  wire _09037_;
  wire _09038_;
  wire _09039_;
  wire _09040_;
  wire _09041_;
  wire _09042_;
  wire _09043_;
  wire _09044_;
  wire _09045_;
  wire _09046_;
  wire _09047_;
  wire _09048_;
  wire _09049_;
  wire _09050_;
  wire _09051_;
  wire _09052_;
  wire _09053_;
  wire _09054_;
  wire _09055_;
  wire _09056_;
  wire _09057_;
  wire _09058_;
  wire _09059_;
  wire _09060_;
  wire _09061_;
  wire _09062_;
  wire _09063_;
  wire _09064_;
  wire _09065_;
  wire _09066_;
  wire _09067_;
  wire _09068_;
  wire _09069_;
  wire _09070_;
  wire _09071_;
  wire _09072_;
  wire _09073_;
  wire _09074_;
  wire _09075_;
  wire _09076_;
  wire _09077_;
  wire _09078_;
  wire _09079_;
  wire _09080_;
  wire _09081_;
  wire _09082_;
  wire _09083_;
  wire _09084_;
  wire _09085_;
  wire _09086_;
  wire _09087_;
  wire _09088_;
  wire _09089_;
  wire _09090_;
  wire _09091_;
  wire _09092_;
  wire _09093_;
  wire _09094_;
  wire _09095_;
  wire _09096_;
  wire _09097_;
  wire _09098_;
  wire _09099_;
  wire _09100_;
  wire _09101_;
  wire _09102_;
  wire _09103_;
  wire _09104_;
  wire _09105_;
  wire _09106_;
  wire _09107_;
  wire _09108_;
  wire _09109_;
  wire _09110_;
  wire _09111_;
  wire _09112_;
  wire _09113_;
  wire _09114_;
  wire _09115_;
  wire _09116_;
  wire _09117_;
  wire _09118_;
  wire _09119_;
  wire _09120_;
  wire _09121_;
  wire _09122_;
  wire _09123_;
  wire _09124_;
  wire _09125_;
  wire _09126_;
  wire _09127_;
  wire _09128_;
  wire _09129_;
  wire _09130_;
  wire _09131_;
  wire _09132_;
  wire _09133_;
  wire _09134_;
  wire _09135_;
  wire _09136_;
  wire _09137_;
  wire _09138_;
  wire _09139_;
  wire _09140_;
  wire _09141_;
  wire _09142_;
  wire _09143_;
  wire _09144_;
  wire _09145_;
  wire _09146_;
  wire _09147_;
  wire _09148_;
  wire _09149_;
  wire _09150_;
  wire _09151_;
  wire _09152_;
  wire _09153_;
  wire _09154_;
  wire _09155_;
  wire _09156_;
  wire _09157_;
  wire _09158_;
  wire _09159_;
  wire _09160_;
  wire _09161_;
  wire _09162_;
  wire _09163_;
  wire _09164_;
  wire _09165_;
  wire _09166_;
  wire _09167_;
  wire _09168_;
  wire _09169_;
  wire _09170_;
  wire _09171_;
  wire _09172_;
  wire _09173_;
  wire _09174_;
  wire _09175_;
  wire _09176_;
  wire _09177_;
  wire _09178_;
  wire _09179_;
  wire _09180_;
  wire _09181_;
  wire _09182_;
  wire _09183_;
  wire _09184_;
  wire _09185_;
  wire _09186_;
  wire _09187_;
  wire _09188_;
  wire _09189_;
  wire _09190_;
  wire _09191_;
  wire _09192_;
  wire _09193_;
  wire _09194_;
  wire _09195_;
  wire _09196_;
  wire _09197_;
  wire _09198_;
  wire _09199_;
  wire _09200_;
  wire _09201_;
  wire _09202_;
  wire _09203_;
  wire _09204_;
  wire _09205_;
  wire _09206_;
  wire _09207_;
  wire _09208_;
  wire _09209_;
  wire _09210_;
  wire _09211_;
  wire _09212_;
  wire _09213_;
  wire _09214_;
  wire _09215_;
  wire _09216_;
  wire _09217_;
  wire _09218_;
  wire _09219_;
  wire _09220_;
  wire _09221_;
  wire _09222_;
  wire _09223_;
  wire _09224_;
  wire _09225_;
  wire _09226_;
  wire _09227_;
  wire _09228_;
  wire _09229_;
  wire _09230_;
  wire _09231_;
  wire _09232_;
  wire _09233_;
  wire _09234_;
  wire _09235_;
  wire _09236_;
  wire _09237_;
  wire _09238_;
  wire _09239_;
  wire _09240_;
  wire _09241_;
  wire _09242_;
  wire _09243_;
  wire _09244_;
  wire _09245_;
  wire _09246_;
  wire _09247_;
  wire _09248_;
  wire _09249_;
  wire _09250_;
  wire _09251_;
  wire _09252_;
  wire _09253_;
  wire _09254_;
  wire _09255_;
  wire _09256_;
  wire _09257_;
  wire _09258_;
  wire _09259_;
  wire _09260_;
  wire _09261_;
  wire _09262_;
  wire _09263_;
  wire _09264_;
  wire _09265_;
  wire _09266_;
  wire _09267_;
  wire _09268_;
  wire _09269_;
  wire _09270_;
  wire _09271_;
  wire _09272_;
  wire _09273_;
  wire _09274_;
  wire _09275_;
  wire _09276_;
  wire _09277_;
  wire _09278_;
  wire _09279_;
  wire _09280_;
  wire _09281_;
  wire _09282_;
  wire _09283_;
  wire _09284_;
  wire _09285_;
  wire _09286_;
  wire _09287_;
  wire _09288_;
  wire _09289_;
  wire _09290_;
  wire _09291_;
  wire _09292_;
  wire _09293_;
  wire _09294_;
  wire _09295_;
  wire _09296_;
  wire _09297_;
  wire _09298_;
  wire _09299_;
  wire _09300_;
  wire _09301_;
  wire _09302_;
  wire _09303_;
  wire _09304_;
  wire _09305_;
  wire _09306_;
  wire _09307_;
  wire _09308_;
  wire _09309_;
  wire _09310_;
  wire _09311_;
  wire _09312_;
  wire _09313_;
  wire _09314_;
  wire _09315_;
  wire _09316_;
  wire _09317_;
  wire _09318_;
  wire _09319_;
  wire _09320_;
  wire _09321_;
  wire _09322_;
  wire _09323_;
  wire _09324_;
  wire _09325_;
  wire _09326_;
  wire _09327_;
  wire _09328_;
  wire _09329_;
  wire _09330_;
  wire _09331_;
  wire _09332_;
  wire _09333_;
  wire _09334_;
  wire _09335_;
  wire _09336_;
  wire _09337_;
  wire _09338_;
  wire _09339_;
  wire _09340_;
  wire _09341_;
  wire _09342_;
  wire _09343_;
  wire _09344_;
  wire _09345_;
  wire _09346_;
  wire _09347_;
  wire _09348_;
  wire _09349_;
  wire _09350_;
  wire _09351_;
  wire _09352_;
  wire _09353_;
  wire _09354_;
  wire _09355_;
  wire _09356_;
  wire _09357_;
  wire _09358_;
  wire _09359_;
  wire _09360_;
  wire _09361_;
  wire _09362_;
  wire _09363_;
  wire _09364_;
  wire _09365_;
  wire _09366_;
  wire _09367_;
  wire _09368_;
  wire _09369_;
  wire _09370_;
  wire _09371_;
  wire _09372_;
  wire _09373_;
  wire _09374_;
  wire _09375_;
  wire _09376_;
  wire _09377_;
  wire _09378_;
  wire _09379_;
  wire _09380_;
  wire _09381_;
  wire _09382_;
  wire _09383_;
  wire _09384_;
  wire _09385_;
  wire _09386_;
  wire _09387_;
  wire _09388_;
  wire _09389_;
  wire _09390_;
  wire _09391_;
  wire _09392_;
  wire _09393_;
  wire _09394_;
  wire _09395_;
  wire _09396_;
  wire _09397_;
  wire _09398_;
  wire _09399_;
  wire _09400_;
  wire _09401_;
  wire _09402_;
  wire _09403_;
  wire _09404_;
  wire _09405_;
  wire _09406_;
  wire _09407_;
  wire _09408_;
  wire _09409_;
  wire _09410_;
  wire _09411_;
  wire _09412_;
  wire _09413_;
  wire _09414_;
  wire _09415_;
  wire _09416_;
  wire _09417_;
  wire _09418_;
  wire _09419_;
  wire _09420_;
  wire _09421_;
  wire _09422_;
  wire _09423_;
  wire _09424_;
  wire _09425_;
  wire _09426_;
  wire _09427_;
  wire _09428_;
  wire _09429_;
  wire _09430_;
  wire _09431_;
  wire _09432_;
  wire _09433_;
  wire _09434_;
  wire _09435_;
  wire _09436_;
  wire _09437_;
  wire _09438_;
  wire _09439_;
  wire _09440_;
  wire _09441_;
  wire _09442_;
  wire _09443_;
  wire _09444_;
  wire _09445_;
  wire _09446_;
  wire _09447_;
  wire _09448_;
  wire _09449_;
  wire _09450_;
  wire _09451_;
  wire _09452_;
  wire _09453_;
  wire _09454_;
  wire _09455_;
  wire _09456_;
  wire _09457_;
  wire _09458_;
  wire _09459_;
  wire _09460_;
  wire _09461_;
  wire _09462_;
  wire _09463_;
  wire _09464_;
  wire _09465_;
  wire _09466_;
  wire _09467_;
  wire _09468_;
  wire _09469_;
  wire _09470_;
  wire _09471_;
  wire _09472_;
  wire _09473_;
  wire _09474_;
  wire _09475_;
  wire _09476_;
  wire _09477_;
  wire _09478_;
  wire _09479_;
  wire _09480_;
  wire _09481_;
  wire _09482_;
  wire _09483_;
  wire _09484_;
  wire _09485_;
  wire _09486_;
  wire _09487_;
  wire _09488_;
  wire _09489_;
  wire _09490_;
  wire _09491_;
  wire _09492_;
  wire _09493_;
  wire _09494_;
  wire _09495_;
  wire _09496_;
  wire _09497_;
  wire _09498_;
  wire _09499_;
  wire _09500_;
  wire _09501_;
  wire _09502_;
  wire _09503_;
  wire _09504_;
  wire _09505_;
  wire _09506_;
  wire _09507_;
  wire _09508_;
  wire _09509_;
  wire _09510_;
  wire _09511_;
  wire _09512_;
  wire _09513_;
  wire _09514_;
  wire _09515_;
  wire _09516_;
  wire _09517_;
  wire _09518_;
  wire _09519_;
  wire _09520_;
  wire _09521_;
  wire _09522_;
  wire _09523_;
  wire _09524_;
  wire _09525_;
  wire _09526_;
  wire _09527_;
  wire _09528_;
  wire _09529_;
  wire _09530_;
  wire _09531_;
  wire _09532_;
  wire _09533_;
  wire _09534_;
  wire _09535_;
  wire _09536_;
  wire _09537_;
  wire _09538_;
  wire _09539_;
  wire _09540_;
  wire _09541_;
  wire _09542_;
  wire _09543_;
  wire _09544_;
  wire _09545_;
  wire _09546_;
  wire _09547_;
  wire _09548_;
  wire _09549_;
  wire _09550_;
  wire _09551_;
  wire _09552_;
  wire _09553_;
  wire _09554_;
  wire _09555_;
  wire _09556_;
  wire _09557_;
  wire _09558_;
  wire _09559_;
  wire _09560_;
  wire _09561_;
  wire _09562_;
  wire _09563_;
  wire _09564_;
  wire _09565_;
  wire _09566_;
  wire _09567_;
  wire _09568_;
  wire _09569_;
  wire _09570_;
  wire _09571_;
  wire _09572_;
  wire _09573_;
  wire _09574_;
  wire _09575_;
  wire _09576_;
  wire _09577_;
  wire _09578_;
  wire _09579_;
  wire _09580_;
  wire _09581_;
  wire _09582_;
  wire _09583_;
  wire _09584_;
  wire _09585_;
  wire _09586_;
  wire _09587_;
  wire _09588_;
  wire _09589_;
  wire _09590_;
  wire _09591_;
  wire _09592_;
  wire _09593_;
  wire _09594_;
  wire _09595_;
  wire _09596_;
  wire _09597_;
  wire _09598_;
  wire _09599_;
  wire _09600_;
  wire _09601_;
  wire _09602_;
  wire _09603_;
  wire _09604_;
  wire _09605_;
  wire _09606_;
  wire _09607_;
  wire _09608_;
  wire _09609_;
  wire _09610_;
  wire _09611_;
  wire _09612_;
  wire _09613_;
  wire _09614_;
  wire _09615_;
  wire _09616_;
  wire _09617_;
  wire _09618_;
  wire _09619_;
  wire _09620_;
  wire _09621_;
  wire _09622_;
  wire _09623_;
  wire _09624_;
  wire _09625_;
  wire _09626_;
  wire _09627_;
  wire _09628_;
  wire _09629_;
  wire _09630_;
  wire _09631_;
  wire _09632_;
  wire _09633_;
  wire _09634_;
  wire _09635_;
  wire _09636_;
  wire _09637_;
  wire _09638_;
  wire _09639_;
  wire _09640_;
  wire _09641_;
  wire _09642_;
  wire _09643_;
  wire _09644_;
  wire _09645_;
  wire _09646_;
  wire _09647_;
  wire _09648_;
  wire _09649_;
  wire _09650_;
  wire _09651_;
  wire _09652_;
  wire _09653_;
  wire _09654_;
  wire _09655_;
  wire _09656_;
  wire _09657_;
  wire _09658_;
  wire _09659_;
  wire _09660_;
  wire _09661_;
  wire _09662_;
  wire _09663_;
  wire _09664_;
  wire _09665_;
  wire _09666_;
  wire _09667_;
  wire _09668_;
  wire _09669_;
  wire _09670_;
  wire _09671_;
  wire _09672_;
  wire _09673_;
  wire _09674_;
  wire _09675_;
  wire _09676_;
  wire _09677_;
  wire _09678_;
  wire _09679_;
  wire _09680_;
  wire _09681_;
  wire _09682_;
  wire _09683_;
  wire _09684_;
  wire _09685_;
  wire _09686_;
  wire _09687_;
  wire _09688_;
  wire _09689_;
  wire _09690_;
  wire _09691_;
  wire _09692_;
  wire _09693_;
  wire _09694_;
  wire _09695_;
  wire _09696_;
  wire _09697_;
  wire _09698_;
  wire _09699_;
  wire _09700_;
  wire _09701_;
  wire _09702_;
  wire _09703_;
  wire _09704_;
  wire _09705_;
  wire _09706_;
  wire _09707_;
  wire _09708_;
  wire _09709_;
  wire _09710_;
  wire _09711_;
  wire _09712_;
  wire _09713_;
  wire _09714_;
  wire _09715_;
  wire _09716_;
  wire _09717_;
  wire _09718_;
  wire _09719_;
  wire _09720_;
  wire _09721_;
  wire _09722_;
  wire _09723_;
  wire _09724_;
  wire _09725_;
  wire _09726_;
  wire _09727_;
  wire _09728_;
  wire _09729_;
  wire _09730_;
  wire _09731_;
  wire _09732_;
  wire _09733_;
  wire _09734_;
  wire _09735_;
  wire _09736_;
  wire _09737_;
  wire _09738_;
  wire _09739_;
  wire _09740_;
  wire _09741_;
  wire _09742_;
  wire _09743_;
  wire _09744_;
  wire _09745_;
  wire _09746_;
  wire _09747_;
  wire _09748_;
  wire _09749_;
  wire _09750_;
  wire _09751_;
  wire _09752_;
  wire _09753_;
  wire _09754_;
  wire _09755_;
  wire _09756_;
  wire _09757_;
  wire _09758_;
  wire _09759_;
  wire _09760_;
  wire _09761_;
  wire _09762_;
  wire _09763_;
  wire _09764_;
  wire _09765_;
  wire _09766_;
  wire _09767_;
  wire _09768_;
  wire _09769_;
  wire _09770_;
  wire _09771_;
  wire _09772_;
  wire _09773_;
  wire _09774_;
  wire _09775_;
  wire _09776_;
  wire _09777_;
  wire _09778_;
  wire _09779_;
  wire _09780_;
  wire _09781_;
  wire _09782_;
  wire _09783_;
  wire _09784_;
  wire _09785_;
  wire _09786_;
  wire _09787_;
  wire _09788_;
  wire _09789_;
  wire _09790_;
  wire _09791_;
  wire _09792_;
  wire _09793_;
  wire _09794_;
  wire _09795_;
  wire _09796_;
  wire _09797_;
  wire _09798_;
  wire _09799_;
  wire _09800_;
  wire _09801_;
  wire _09802_;
  wire _09803_;
  wire _09804_;
  wire _09805_;
  wire _09806_;
  wire _09807_;
  wire _09808_;
  wire _09809_;
  wire _09810_;
  wire _09811_;
  wire _09812_;
  wire _09813_;
  wire _09814_;
  wire _09815_;
  wire _09816_;
  wire _09817_;
  wire _09818_;
  wire _09819_;
  wire _09820_;
  wire _09821_;
  wire _09822_;
  wire _09823_;
  wire _09824_;
  wire _09825_;
  wire _09826_;
  wire _09827_;
  wire _09828_;
  wire _09829_;
  wire _09830_;
  wire _09831_;
  wire _09832_;
  wire _09833_;
  wire _09834_;
  wire _09835_;
  wire _09836_;
  wire _09837_;
  wire _09838_;
  wire _09839_;
  wire _09840_;
  wire _09841_;
  wire _09842_;
  wire _09843_;
  wire _09844_;
  wire _09845_;
  wire _09846_;
  wire _09847_;
  wire _09848_;
  wire _09849_;
  wire _09850_;
  wire _09851_;
  wire _09852_;
  wire _09853_;
  wire _09854_;
  wire _09855_;
  wire _09856_;
  wire _09857_;
  wire _09858_;
  wire _09859_;
  wire _09860_;
  wire _09861_;
  wire _09862_;
  wire _09863_;
  wire _09864_;
  wire _09865_;
  wire _09866_;
  wire _09867_;
  wire _09868_;
  wire _09869_;
  wire _09870_;
  wire _09871_;
  wire _09872_;
  wire _09873_;
  wire _09874_;
  wire _09875_;
  wire _09876_;
  wire _09877_;
  wire _09878_;
  wire _09879_;
  wire _09880_;
  wire _09881_;
  wire _09882_;
  wire _09883_;
  wire _09884_;
  wire _09885_;
  wire _09886_;
  wire _09887_;
  wire _09888_;
  wire _09889_;
  wire _09890_;
  wire _09891_;
  wire _09892_;
  wire _09893_;
  wire _09894_;
  wire _09895_;
  wire _09896_;
  wire _09897_;
  wire _09898_;
  wire _09899_;
  wire _09900_;
  wire _09901_;
  wire _09902_;
  wire _09903_;
  wire _09904_;
  wire _09905_;
  wire _09906_;
  wire _09907_;
  wire _09908_;
  wire _09909_;
  wire _09910_;
  wire _09911_;
  wire _09912_;
  wire _09913_;
  wire _09914_;
  wire _09915_;
  wire _09916_;
  wire _09917_;
  wire _09918_;
  wire _09919_;
  wire _09920_;
  wire _09921_;
  wire _09922_;
  wire _09923_;
  wire _09924_;
  wire _09925_;
  wire _09926_;
  wire _09927_;
  wire _09928_;
  wire _09929_;
  wire _09930_;
  wire _09931_;
  wire _09932_;
  wire _09933_;
  wire _09934_;
  wire _09935_;
  wire _09936_;
  wire _09937_;
  wire _09938_;
  wire _09939_;
  wire _09940_;
  wire _09941_;
  wire _09942_;
  wire _09943_;
  wire _09944_;
  wire _09945_;
  wire _09946_;
  wire _09947_;
  wire _09948_;
  wire _09949_;
  wire _09950_;
  wire _09951_;
  wire _09952_;
  wire _09953_;
  wire _09954_;
  wire _09955_;
  wire _09956_;
  wire _09957_;
  wire _09958_;
  wire _09959_;
  wire _09960_;
  wire _09961_;
  wire _09962_;
  wire _09963_;
  wire _09964_;
  wire _09965_;
  wire _09966_;
  wire _09967_;
  wire _09968_;
  wire _09969_;
  wire _09970_;
  wire _09971_;
  wire _09972_;
  wire _09973_;
  wire _09974_;
  wire _09975_;
  wire _09976_;
  wire _09977_;
  wire _09978_;
  wire _09979_;
  wire _09980_;
  wire _09981_;
  wire _09982_;
  wire _09983_;
  wire _09984_;
  wire _09985_;
  wire _09986_;
  wire _09987_;
  wire _09988_;
  wire _09989_;
  wire _09990_;
  wire _09991_;
  wire _09992_;
  wire _09993_;
  wire _09994_;
  wire _09995_;
  wire _09996_;
  wire _09997_;
  wire _09998_;
  wire _09999_;
  wire _10000_;
  wire _10001_;
  wire _10002_;
  wire _10003_;
  wire _10004_;
  wire _10005_;
  wire _10006_;
  wire _10007_;
  wire _10008_;
  wire _10009_;
  wire _10010_;
  wire _10011_;
  wire _10012_;
  wire _10013_;
  wire _10014_;
  wire _10015_;
  wire _10016_;
  wire _10017_;
  wire _10018_;
  wire _10019_;
  wire _10020_;
  wire _10021_;
  wire _10022_;
  wire _10023_;
  wire _10024_;
  wire _10025_;
  wire _10026_;
  wire _10027_;
  wire _10028_;
  wire _10029_;
  wire _10030_;
  wire _10031_;
  wire _10032_;
  wire _10033_;
  wire _10034_;
  wire _10035_;
  wire _10036_;
  wire _10037_;
  wire _10038_;
  wire _10039_;
  wire _10040_;
  wire _10041_;
  wire _10042_;
  wire _10043_;
  wire _10044_;
  wire _10045_;
  wire _10046_;
  wire _10047_;
  wire _10048_;
  wire _10049_;
  wire _10050_;
  wire _10051_;
  wire _10052_;
  wire _10053_;
  wire _10054_;
  wire _10055_;
  wire _10056_;
  wire _10057_;
  wire _10058_;
  wire _10059_;
  wire _10060_;
  wire _10061_;
  wire _10062_;
  wire _10063_;
  wire _10064_;
  wire _10065_;
  wire _10066_;
  wire _10067_;
  wire _10068_;
  wire _10069_;
  wire _10070_;
  wire _10071_;
  wire _10072_;
  wire _10073_;
  wire _10074_;
  wire _10075_;
  wire _10076_;
  wire _10077_;
  wire _10078_;
  wire _10079_;
  wire _10080_;
  wire _10081_;
  wire _10082_;
  wire _10083_;
  wire _10084_;
  wire _10085_;
  wire _10086_;
  wire _10087_;
  wire _10088_;
  wire _10089_;
  wire _10090_;
  wire _10091_;
  wire _10092_;
  wire _10093_;
  wire _10094_;
  wire _10095_;
  wire _10096_;
  wire _10097_;
  wire _10098_;
  wire _10099_;
  wire _10100_;
  wire _10101_;
  wire _10102_;
  wire _10103_;
  wire _10104_;
  wire _10105_;
  wire _10106_;
  wire _10107_;
  wire _10108_;
  wire _10109_;
  wire _10110_;
  wire _10111_;
  wire _10112_;
  wire _10113_;
  wire _10114_;
  wire _10115_;
  wire _10116_;
  wire _10117_;
  wire _10118_;
  wire _10119_;
  wire _10120_;
  wire _10121_;
  wire _10122_;
  wire _10123_;
  wire _10124_;
  wire _10125_;
  wire _10126_;
  wire _10127_;
  wire _10128_;
  wire _10129_;
  wire _10130_;
  wire _10131_;
  wire _10132_;
  wire _10133_;
  wire _10134_;
  wire _10135_;
  wire _10136_;
  wire _10137_;
  wire _10138_;
  wire _10139_;
  wire _10140_;
  wire _10141_;
  wire _10142_;
  wire _10143_;
  wire _10144_;
  wire _10145_;
  wire _10146_;
  wire _10147_;
  wire _10148_;
  wire _10149_;
  wire _10150_;
  wire _10151_;
  wire _10152_;
  wire _10153_;
  wire _10154_;
  wire _10155_;
  wire _10156_;
  wire _10157_;
  wire _10158_;
  wire _10159_;
  wire _10160_;
  wire _10161_;
  wire _10162_;
  wire _10163_;
  wire _10164_;
  wire _10165_;
  wire _10166_;
  wire _10167_;
  wire _10168_;
  wire _10169_;
  wire _10170_;
  wire _10171_;
  wire _10172_;
  wire _10173_;
  wire _10174_;
  wire _10175_;
  wire _10176_;
  wire _10177_;
  wire _10178_;
  wire _10179_;
  wire _10180_;
  wire _10181_;
  wire _10182_;
  wire _10183_;
  wire _10184_;
  wire _10185_;
  wire _10186_;
  wire _10187_;
  wire _10188_;
  wire _10189_;
  wire _10190_;
  wire _10191_;
  wire _10192_;
  wire _10193_;
  wire _10194_;
  wire _10195_;
  wire _10196_;
  wire _10197_;
  wire _10198_;
  wire _10199_;
  wire _10200_;
  wire _10201_;
  wire _10202_;
  wire _10203_;
  wire _10204_;
  wire _10205_;
  wire _10206_;
  wire _10207_;
  wire _10208_;
  wire _10209_;
  wire _10210_;
  wire _10211_;
  wire _10212_;
  wire _10213_;
  wire _10214_;
  wire _10215_;
  wire _10216_;
  wire _10217_;
  wire _10218_;
  wire _10219_;
  wire _10220_;
  wire _10221_;
  wire _10222_;
  wire _10223_;
  wire _10224_;
  wire _10225_;
  wire _10226_;
  wire _10227_;
  wire _10228_;
  wire _10229_;
  wire _10230_;
  wire _10231_;
  wire _10232_;
  wire _10233_;
  wire _10234_;
  wire _10235_;
  wire _10236_;
  wire _10237_;
  wire _10238_;
  wire _10239_;
  wire _10240_;
  wire _10241_;
  wire _10242_;
  wire _10243_;
  wire _10244_;
  wire _10245_;
  wire _10246_;
  wire _10247_;
  wire _10248_;
  wire _10249_;
  wire _10250_;
  wire _10251_;
  wire _10252_;
  wire _10253_;
  wire _10254_;
  wire _10255_;
  wire _10256_;
  wire _10257_;
  wire _10258_;
  wire _10259_;
  wire _10260_;
  wire _10261_;
  wire _10262_;
  wire _10263_;
  wire _10264_;
  wire _10265_;
  wire _10266_;
  wire _10267_;
  wire _10268_;
  wire _10269_;
  wire _10270_;
  wire _10271_;
  wire _10272_;
  wire _10273_;
  wire _10274_;
  wire _10275_;
  wire _10276_;
  wire _10277_;
  wire _10278_;
  wire _10279_;
  wire _10280_;
  wire _10281_;
  wire _10282_;
  wire _10283_;
  wire _10284_;
  wire _10285_;
  wire _10286_;
  wire _10287_;
  wire _10288_;
  wire _10289_;
  wire _10290_;
  wire _10291_;
  wire _10292_;
  wire _10293_;
  wire _10294_;
  wire _10295_;
  wire _10296_;
  wire _10297_;
  wire _10298_;
  wire _10299_;
  wire _10300_;
  wire _10301_;
  wire _10302_;
  wire _10303_;
  wire _10304_;
  wire _10305_;
  wire _10306_;
  wire _10307_;
  wire _10308_;
  wire _10309_;
  wire _10310_;
  wire _10311_;
  wire _10312_;
  wire _10313_;
  wire _10314_;
  wire _10315_;
  wire _10316_;
  wire _10317_;
  wire _10318_;
  wire _10319_;
  wire _10320_;
  wire _10321_;
  wire _10322_;
  wire _10323_;
  wire _10324_;
  wire _10325_;
  wire _10326_;
  wire _10327_;
  wire _10328_;
  wire _10329_;
  wire _10330_;
  wire _10331_;
  wire _10332_;
  wire _10333_;
  wire _10334_;
  wire _10335_;
  wire _10336_;
  wire _10337_;
  wire _10338_;
  wire _10339_;
  wire _10340_;
  wire _10341_;
  wire _10342_;
  wire _10343_;
  wire _10344_;
  wire _10345_;
  wire _10346_;
  wire _10347_;
  wire _10348_;
  wire _10349_;
  wire _10350_;
  wire _10351_;
  wire _10352_;
  wire _10353_;
  wire _10354_;
  wire _10355_;
  wire _10356_;
  wire _10357_;
  wire _10358_;
  wire _10359_;
  wire _10360_;
  wire _10361_;
  wire _10362_;
  wire _10363_;
  wire _10364_;
  wire _10365_;
  wire _10366_;
  wire _10367_;
  wire _10368_;
  wire _10369_;
  wire _10370_;
  wire _10371_;
  wire _10372_;
  wire _10373_;
  wire _10374_;
  wire _10375_;
  wire _10376_;
  wire _10377_;
  wire _10378_;
  wire _10379_;
  wire _10380_;
  wire _10381_;
  wire _10382_;
  wire _10383_;
  wire _10384_;
  wire _10385_;
  wire _10386_;
  wire _10387_;
  wire _10388_;
  wire _10389_;
  wire _10390_;
  wire _10391_;
  wire _10392_;
  wire _10393_;
  wire _10394_;
  wire _10395_;
  wire _10396_;
  wire _10397_;
  wire _10398_;
  wire _10399_;
  wire _10400_;
  wire _10401_;
  wire _10402_;
  wire _10403_;
  wire _10404_;
  wire _10405_;
  wire _10406_;
  wire _10407_;
  wire _10408_;
  wire _10409_;
  wire _10410_;
  wire _10411_;
  wire _10412_;
  wire _10413_;
  wire _10414_;
  wire _10415_;
  wire _10416_;
  wire _10417_;
  wire _10418_;
  wire _10419_;
  wire _10420_;
  wire _10421_;
  wire _10422_;
  wire _10423_;
  wire _10424_;
  wire _10425_;
  wire _10426_;
  wire _10427_;
  wire _10428_;
  wire _10429_;
  wire _10430_;
  wire _10431_;
  wire _10432_;
  wire _10433_;
  wire _10434_;
  wire _10435_;
  wire _10436_;
  wire _10437_;
  wire _10438_;
  wire _10439_;
  wire _10440_;
  wire _10441_;
  wire _10442_;
  wire _10443_;
  wire _10444_;
  wire _10445_;
  wire _10446_;
  wire _10447_;
  wire _10448_;
  wire _10449_;
  wire _10450_;
  wire _10451_;
  wire _10452_;
  wire _10453_;
  wire _10454_;
  wire _10455_;
  wire _10456_;
  wire _10457_;
  wire _10458_;
  wire _10459_;
  wire _10460_;
  wire _10461_;
  wire _10462_;
  wire _10463_;
  wire _10464_;
  wire _10465_;
  wire _10466_;
  wire _10467_;
  wire _10468_;
  wire _10469_;
  wire _10470_;
  wire _10471_;
  wire _10472_;
  wire _10473_;
  wire _10474_;
  wire _10475_;
  wire _10476_;
  wire _10477_;
  wire _10478_;
  wire _10479_;
  wire _10480_;
  wire _10481_;
  wire _10482_;
  wire _10483_;
  wire _10484_;
  wire _10485_;
  wire _10486_;
  wire _10487_;
  wire _10488_;
  wire _10489_;
  wire _10490_;
  wire _10491_;
  wire _10492_;
  wire _10493_;
  wire _10494_;
  wire _10495_;
  wire _10496_;
  wire _10497_;
  wire _10498_;
  wire _10499_;
  wire _10500_;
  wire _10501_;
  wire _10502_;
  wire _10503_;
  wire _10504_;
  wire _10505_;
  wire _10506_;
  wire _10507_;
  wire _10508_;
  wire _10509_;
  wire _10510_;
  wire _10511_;
  wire _10512_;
  wire _10513_;
  wire _10514_;
  wire _10515_;
  wire _10516_;
  wire _10517_;
  wire _10518_;
  wire _10519_;
  wire _10520_;
  wire _10521_;
  wire _10522_;
  wire _10523_;
  wire _10524_;
  wire _10525_;
  wire _10526_;
  wire _10527_;
  wire _10528_;
  wire _10529_;
  wire _10530_;
  wire _10531_;
  wire _10532_;
  wire _10533_;
  wire _10534_;
  wire _10535_;
  wire _10536_;
  wire _10537_;
  wire _10538_;
  wire _10539_;
  wire _10540_;
  wire _10541_;
  wire _10542_;
  wire _10543_;
  wire _10544_;
  wire _10545_;
  wire _10546_;
  wire _10547_;
  wire _10548_;
  wire _10549_;
  wire _10550_;
  wire _10551_;
  wire _10552_;
  wire _10553_;
  wire _10554_;
  wire _10555_;
  wire _10556_;
  wire _10557_;
  wire _10558_;
  wire _10559_;
  wire _10560_;
  wire _10561_;
  wire _10562_;
  wire _10563_;
  wire _10564_;
  wire _10565_;
  wire _10566_;
  wire _10567_;
  wire _10568_;
  wire _10569_;
  wire _10570_;
  wire _10571_;
  wire _10572_;
  wire _10573_;
  wire _10574_;
  wire _10575_;
  wire _10576_;
  wire _10577_;
  wire _10578_;
  wire _10579_;
  wire _10580_;
  wire _10581_;
  wire _10582_;
  wire _10583_;
  wire _10584_;
  wire _10585_;
  wire _10586_;
  wire _10587_;
  wire _10588_;
  wire _10589_;
  wire _10590_;
  wire _10591_;
  wire _10592_;
  wire _10593_;
  wire _10594_;
  wire _10595_;
  wire _10596_;
  wire _10597_;
  wire _10598_;
  wire _10599_;
  wire _10600_;
  wire _10601_;
  wire _10602_;
  wire _10603_;
  wire _10604_;
  wire _10605_;
  wire _10606_;
  wire _10607_;
  wire _10608_;
  wire _10609_;
  wire _10610_;
  wire _10611_;
  wire _10612_;
  wire _10613_;
  wire _10614_;
  wire _10615_;
  wire _10616_;
  wire _10617_;
  wire _10618_;
  wire _10619_;
  wire _10620_;
  wire _10621_;
  wire _10622_;
  wire _10623_;
  wire _10624_;
  wire _10625_;
  wire _10626_;
  wire _10627_;
  wire _10628_;
  wire _10629_;
  wire _10630_;
  wire _10631_;
  wire _10632_;
  wire _10633_;
  wire _10634_;
  wire _10635_;
  wire _10636_;
  wire _10637_;
  wire _10638_;
  wire _10639_;
  wire _10640_;
  wire _10641_;
  wire _10642_;
  wire _10643_;
  wire _10644_;
  wire _10645_;
  wire _10646_;
  wire _10647_;
  wire _10648_;
  wire _10649_;
  wire _10650_;
  wire _10651_;
  wire _10652_;
  wire _10653_;
  wire _10654_;
  wire _10655_;
  wire _10656_;
  wire _10657_;
  wire _10658_;
  wire _10659_;
  wire _10660_;
  wire _10661_;
  wire _10662_;
  wire _10663_;
  wire _10664_;
  wire _10665_;
  wire _10666_;
  wire _10667_;
  wire _10668_;
  wire _10669_;
  wire _10670_;
  wire _10671_;
  wire _10672_;
  wire _10673_;
  wire _10674_;
  wire _10675_;
  wire _10676_;
  wire _10677_;
  wire _10678_;
  wire _10679_;
  wire _10680_;
  wire _10681_;
  wire _10682_;
  wire _10683_;
  wire _10684_;
  wire _10685_;
  wire _10686_;
  wire _10687_;
  wire _10688_;
  wire _10689_;
  wire _10690_;
  wire _10691_;
  wire _10692_;
  wire _10693_;
  wire _10694_;
  wire _10695_;
  wire _10696_;
  wire _10697_;
  wire _10698_;
  wire _10699_;
  wire _10700_;
  wire _10701_;
  wire _10702_;
  wire _10703_;
  wire _10704_;
  wire _10705_;
  wire _10706_;
  wire _10707_;
  wire _10708_;
  wire _10709_;
  wire _10710_;
  wire _10711_;
  wire _10712_;
  wire _10713_;
  wire _10714_;
  wire _10715_;
  wire _10716_;
  wire _10717_;
  wire _10718_;
  wire _10719_;
  wire _10720_;
  wire _10721_;
  wire _10722_;
  wire _10723_;
  wire _10724_;
  wire _10725_;
  wire _10726_;
  wire _10727_;
  wire _10728_;
  wire _10729_;
  wire _10730_;
  wire _10731_;
  wire _10732_;
  wire _10733_;
  wire _10734_;
  wire _10735_;
  wire _10736_;
  wire _10737_;
  wire _10738_;
  wire _10739_;
  wire _10740_;
  wire _10741_;
  wire _10742_;
  wire _10743_;
  wire _10744_;
  wire _10745_;
  wire _10746_;
  wire _10747_;
  wire _10748_;
  wire _10749_;
  wire _10750_;
  wire _10751_;
  wire _10752_;
  wire _10753_;
  wire _10754_;
  wire _10755_;
  wire _10756_;
  wire _10757_;
  wire _10758_;
  wire _10759_;
  wire _10760_;
  wire _10761_;
  wire _10762_;
  wire _10763_;
  wire _10764_;
  wire _10765_;
  wire _10766_;
  wire _10767_;
  wire _10768_;
  wire _10769_;
  wire _10770_;
  wire _10771_;
  wire _10772_;
  wire _10773_;
  wire _10774_;
  wire _10775_;
  wire _10776_;
  wire _10777_;
  wire _10778_;
  wire _10779_;
  wire _10780_;
  wire _10781_;
  wire _10782_;
  wire _10783_;
  wire _10784_;
  wire _10785_;
  wire _10786_;
  wire _10787_;
  wire _10788_;
  wire _10789_;
  wire _10790_;
  wire _10791_;
  wire _10792_;
  wire _10793_;
  wire _10794_;
  wire _10795_;
  wire _10796_;
  wire _10797_;
  wire _10798_;
  wire _10799_;
  wire _10800_;
  wire _10801_;
  wire _10802_;
  wire _10803_;
  wire _10804_;
  wire _10805_;
  wire _10806_;
  wire _10807_;
  wire _10808_;
  wire _10809_;
  wire _10810_;
  wire _10811_;
  wire _10812_;
  wire _10813_;
  wire _10814_;
  wire _10815_;
  wire _10816_;
  wire _10817_;
  wire _10818_;
  wire _10819_;
  wire _10820_;
  wire _10821_;
  wire _10822_;
  wire _10823_;
  wire _10824_;
  wire _10825_;
  wire _10826_;
  wire _10827_;
  wire _10828_;
  wire _10829_;
  wire _10830_;
  wire _10831_;
  wire _10832_;
  wire _10833_;
  wire _10834_;
  wire _10835_;
  wire _10836_;
  wire _10837_;
  wire _10838_;
  wire _10839_;
  wire _10840_;
  wire _10841_;
  wire _10842_;
  wire _10843_;
  wire _10844_;
  wire _10845_;
  wire _10846_;
  wire _10847_;
  wire _10848_;
  wire _10849_;
  wire _10850_;
  wire _10851_;
  wire _10852_;
  wire _10853_;
  wire _10854_;
  wire _10855_;
  wire _10856_;
  wire _10857_;
  wire _10858_;
  wire _10859_;
  wire _10860_;
  wire _10861_;
  wire _10862_;
  wire _10863_;
  wire _10864_;
  wire _10865_;
  wire _10866_;
  wire _10867_;
  wire _10868_;
  wire _10869_;
  wire _10870_;
  wire _10871_;
  wire _10872_;
  wire _10873_;
  wire _10874_;
  wire _10875_;
  wire _10876_;
  wire _10877_;
  wire _10878_;
  wire _10879_;
  wire _10880_;
  wire _10881_;
  wire _10882_;
  wire _10883_;
  wire _10884_;
  wire _10885_;
  wire _10886_;
  wire _10887_;
  wire _10888_;
  wire _10889_;
  wire _10890_;
  wire _10891_;
  wire _10892_;
  wire _10893_;
  wire _10894_;
  wire _10895_;
  wire _10896_;
  wire _10897_;
  wire _10898_;
  wire _10899_;
  wire _10900_;
  wire _10901_;
  wire _10902_;
  wire _10903_;
  wire _10904_;
  wire _10905_;
  wire _10906_;
  wire _10907_;
  wire _10908_;
  wire _10909_;
  wire _10910_;
  wire _10911_;
  wire _10912_;
  wire _10913_;
  wire _10914_;
  wire _10915_;
  wire _10916_;
  wire _10917_;
  wire _10918_;
  wire _10919_;
  wire _10920_;
  wire _10921_;
  wire _10922_;
  wire _10923_;
  wire _10924_;
  wire _10925_;
  wire _10926_;
  wire _10927_;
  wire _10928_;
  wire _10929_;
  wire _10930_;
  wire _10931_;
  wire _10932_;
  wire _10933_;
  wire _10934_;
  wire _10935_;
  wire _10936_;
  wire _10937_;
  wire _10938_;
  wire _10939_;
  wire _10940_;
  wire _10941_;
  wire _10942_;
  wire _10943_;
  wire _10944_;
  wire _10945_;
  wire _10946_;
  wire _10947_;
  wire _10948_;
  wire _10949_;
  wire _10950_;
  wire _10951_;
  wire _10952_;
  wire _10953_;
  wire _10954_;
  wire _10955_;
  wire _10956_;
  wire _10957_;
  wire _10958_;
  wire _10959_;
  wire _10960_;
  wire _10961_;
  wire _10962_;
  wire _10963_;
  wire _10964_;
  wire _10965_;
  wire _10966_;
  wire _10967_;
  wire _10968_;
  wire _10969_;
  wire _10970_;
  wire _10971_;
  wire _10972_;
  wire _10973_;
  wire _10974_;
  wire _10975_;
  wire _10976_;
  wire _10977_;
  wire _10978_;
  wire _10979_;
  wire _10980_;
  wire _10981_;
  wire _10982_;
  wire _10983_;
  wire _10984_;
  wire _10985_;
  wire _10986_;
  wire _10987_;
  wire _10988_;
  wire _10989_;
  wire _10990_;
  wire _10991_;
  wire _10992_;
  wire _10993_;
  wire _10994_;
  wire _10995_;
  wire _10996_;
  wire _10997_;
  wire _10998_;
  wire _10999_;
  wire _11000_;
  wire _11001_;
  wire _11002_;
  wire _11003_;
  wire _11004_;
  wire _11005_;
  wire _11006_;
  wire _11007_;
  wire _11008_;
  wire _11009_;
  wire _11010_;
  wire _11011_;
  wire _11012_;
  wire _11013_;
  wire _11014_;
  wire _11015_;
  wire _11016_;
  wire _11017_;
  wire _11018_;
  wire _11019_;
  wire _11020_;
  wire _11021_;
  wire _11022_;
  wire _11023_;
  wire _11024_;
  wire _11025_;
  wire _11026_;
  wire _11027_;
  wire _11028_;
  wire _11029_;
  wire _11030_;
  wire _11031_;
  wire _11032_;
  wire _11033_;
  wire _11034_;
  wire _11035_;
  wire _11036_;
  wire _11037_;
  wire _11038_;
  wire _11039_;
  wire _11040_;
  wire _11041_;
  wire _11042_;
  wire _11043_;
  wire _11044_;
  wire _11045_;
  wire _11046_;
  wire _11047_;
  wire _11048_;
  wire _11049_;
  wire _11050_;
  wire _11051_;
  wire _11052_;
  wire _11053_;
  wire _11054_;
  wire _11055_;
  wire _11056_;
  wire _11057_;
  wire _11058_;
  wire _11059_;
  wire _11060_;
  wire _11061_;
  wire _11062_;
  wire _11063_;
  wire _11064_;
  wire _11065_;
  wire _11066_;
  wire _11067_;
  wire _11068_;
  wire _11069_;
  wire _11070_;
  wire _11071_;
  wire _11072_;
  wire _11073_;
  wire _11074_;
  wire _11075_;
  wire _11076_;
  wire _11077_;
  wire _11078_;
  wire _11079_;
  wire _11080_;
  wire _11081_;
  wire _11082_;
  wire _11083_;
  wire _11084_;
  wire _11085_;
  wire _11086_;
  wire _11087_;
  wire _11088_;
  wire _11089_;
  wire _11090_;
  wire _11091_;
  wire _11092_;
  wire _11093_;
  wire _11094_;
  wire _11095_;
  wire _11096_;
  wire _11097_;
  wire _11098_;
  wire _11099_;
  wire _11100_;
  wire _11101_;
  wire _11102_;
  wire _11103_;
  wire _11104_;
  wire _11105_;
  wire _11106_;
  wire _11107_;
  wire _11108_;
  wire _11109_;
  wire _11110_;
  wire _11111_;
  wire _11112_;
  wire _11113_;
  wire _11114_;
  wire _11115_;
  wire _11116_;
  wire _11117_;
  wire _11118_;
  wire _11119_;
  wire _11120_;
  wire _11121_;
  wire _11122_;
  wire _11123_;
  wire _11124_;
  wire _11125_;
  wire _11126_;
  wire _11127_;
  wire _11128_;
  wire _11129_;
  wire _11130_;
  wire _11131_;
  wire _11132_;
  wire _11133_;
  wire _11134_;
  wire _11135_;
  wire _11136_;
  wire _11137_;
  wire _11138_;
  wire _11139_;
  wire _11140_;
  wire _11141_;
  wire _11142_;
  wire _11143_;
  wire _11144_;
  wire _11145_;
  wire _11146_;
  wire _11147_;
  wire _11148_;
  wire _11149_;
  wire _11150_;
  wire _11151_;
  wire _11152_;
  wire _11153_;
  wire _11154_;
  wire _11155_;
  wire _11156_;
  wire _11157_;
  wire _11158_;
  wire _11159_;
  wire _11160_;
  wire _11161_;
  wire _11162_;
  wire _11163_;
  wire _11164_;
  wire _11165_;
  wire _11166_;
  wire _11167_;
  wire _11168_;
  wire _11169_;
  wire _11170_;
  wire _11171_;
  wire _11172_;
  wire _11173_;
  wire _11174_;
  wire _11175_;
  wire _11176_;
  wire _11177_;
  wire _11178_;
  wire _11179_;
  wire _11180_;
  wire _11181_;
  wire _11182_;
  wire _11183_;
  wire _11184_;
  wire _11185_;
  wire _11186_;
  wire _11187_;
  wire _11188_;
  wire _11189_;
  wire _11190_;
  wire _11191_;
  wire _11192_;
  wire _11193_;
  wire _11194_;
  wire _11195_;
  wire _11196_;
  wire _11197_;
  wire _11198_;
  wire _11199_;
  wire _11200_;
  wire _11201_;
  wire _11202_;
  wire _11203_;
  wire _11204_;
  wire _11205_;
  wire _11206_;
  wire _11207_;
  wire _11208_;
  wire _11209_;
  wire _11210_;
  wire _11211_;
  wire _11212_;
  wire _11213_;
  wire _11214_;
  wire _11215_;
  wire _11216_;
  wire _11217_;
  wire _11218_;
  wire _11219_;
  wire _11220_;
  wire _11221_;
  wire _11222_;
  wire _11223_;
  wire _11224_;
  wire _11225_;
  wire _11226_;
  wire _11227_;
  wire _11228_;
  wire _11229_;
  wire _11230_;
  wire _11231_;
  wire _11232_;
  wire _11233_;
  wire _11234_;
  wire _11235_;
  wire _11236_;
  wire _11237_;
  wire _11238_;
  wire _11239_;
  wire _11240_;
  wire _11241_;
  wire _11242_;
  wire _11243_;
  wire _11244_;
  wire _11245_;
  wire _11246_;
  wire _11247_;
  wire _11248_;
  wire _11249_;
  wire _11250_;
  wire _11251_;
  wire _11252_;
  wire _11253_;
  wire _11254_;
  wire _11255_;
  wire _11256_;
  wire _11257_;
  wire _11258_;
  wire _11259_;
  wire _11260_;
  wire _11261_;
  wire _11262_;
  wire _11263_;
  wire _11264_;
  wire _11265_;
  wire _11266_;
  wire _11267_;
  wire _11268_;
  wire _11269_;
  wire _11270_;
  wire _11271_;
  wire _11272_;
  wire _11273_;
  wire _11274_;
  wire _11275_;
  wire _11276_;
  wire _11277_;
  wire _11278_;
  wire _11279_;
  wire _11280_;
  wire _11281_;
  wire _11282_;
  wire _11283_;
  wire _11284_;
  wire _11285_;
  wire _11286_;
  wire _11287_;
  wire _11288_;
  wire _11289_;
  wire _11290_;
  wire _11291_;
  wire _11292_;
  wire _11293_;
  wire _11294_;
  wire _11295_;
  wire _11296_;
  wire _11297_;
  wire _11298_;
  wire _11299_;
  wire _11300_;
  wire _11301_;
  wire _11302_;
  wire _11303_;
  wire _11304_;
  wire _11305_;
  wire _11306_;
  wire _11307_;
  wire _11308_;
  wire _11309_;
  wire _11310_;
  wire _11311_;
  wire _11312_;
  wire _11313_;
  wire _11314_;
  wire _11315_;
  wire _11316_;
  wire _11317_;
  wire _11318_;
  wire _11319_;
  wire _11320_;
  wire _11321_;
  wire _11322_;
  wire _11323_;
  wire _11324_;
  wire _11325_;
  wire _11326_;
  wire _11327_;
  wire _11328_;
  wire _11329_;
  wire _11330_;
  wire _11331_;
  wire _11332_;
  wire _11333_;
  wire _11334_;
  wire _11335_;
  wire _11336_;
  wire _11337_;
  wire _11338_;
  wire _11339_;
  wire _11340_;
  wire _11341_;
  wire _11342_;
  wire _11343_;
  wire _11344_;
  wire _11345_;
  wire _11346_;
  wire _11347_;
  wire _11348_;
  wire _11349_;
  wire _11350_;
  wire _11351_;
  wire _11352_;
  wire _11353_;
  wire _11354_;
  wire _11355_;
  wire _11356_;
  wire _11357_;
  wire _11358_;
  wire _11359_;
  wire _11360_;
  wire _11361_;
  wire _11362_;
  wire _11363_;
  wire _11364_;
  wire _11365_;
  wire _11366_;
  wire _11367_;
  wire _11368_;
  wire _11369_;
  wire _11370_;
  wire _11371_;
  wire _11372_;
  wire _11373_;
  wire _11374_;
  wire _11375_;
  wire _11376_;
  wire _11377_;
  wire _11378_;
  wire _11379_;
  wire _11380_;
  wire _11381_;
  wire _11382_;
  wire _11383_;
  wire _11384_;
  wire _11385_;
  wire _11386_;
  wire _11387_;
  wire _11388_;
  wire _11389_;
  wire _11390_;
  wire _11391_;
  wire _11392_;
  wire _11393_;
  wire _11394_;
  wire _11395_;
  wire _11396_;
  wire _11397_;
  wire _11398_;
  wire _11399_;
  wire _11400_;
  wire _11401_;
  wire _11402_;
  wire _11403_;
  wire _11404_;
  wire _11405_;
  wire _11406_;
  wire _11407_;
  wire _11408_;
  wire _11409_;
  wire _11410_;
  wire _11411_;
  wire _11412_;
  wire _11413_;
  wire _11414_;
  wire _11415_;
  wire _11416_;
  wire _11417_;
  wire _11418_;
  wire _11419_;
  wire _11420_;
  wire _11421_;
  wire _11422_;
  wire _11423_;
  wire _11424_;
  wire _11425_;
  wire _11426_;
  wire _11427_;
  wire _11428_;
  wire _11429_;
  wire _11430_;
  wire _11431_;
  wire _11432_;
  wire _11433_;
  wire _11434_;
  wire _11435_;
  wire _11436_;
  wire _11437_;
  wire _11438_;
  wire _11439_;
  wire _11440_;
  wire _11441_;
  wire _11442_;
  wire _11443_;
  wire _11444_;
  wire _11445_;
  wire _11446_;
  wire _11447_;
  wire _11448_;
  wire _11449_;
  wire _11450_;
  wire _11451_;
  wire _11452_;
  wire _11453_;
  wire _11454_;
  wire _11455_;
  wire _11456_;
  wire _11457_;
  wire _11458_;
  wire _11459_;
  wire _11460_;
  wire _11461_;
  wire _11462_;
  wire _11463_;
  wire _11464_;
  wire _11465_;
  wire _11466_;
  wire _11467_;
  wire _11468_;
  wire _11469_;
  wire _11470_;
  wire _11471_;
  wire _11472_;
  wire _11473_;
  wire _11474_;
  wire _11475_;
  wire _11476_;
  wire _11477_;
  wire _11478_;
  wire _11479_;
  wire _11480_;
  wire _11481_;
  wire _11482_;
  wire _11483_;
  wire _11484_;
  wire _11485_;
  wire _11486_;
  wire _11487_;
  wire _11488_;
  wire _11489_;
  wire _11490_;
  wire _11491_;
  wire _11492_;
  wire _11493_;
  wire _11494_;
  wire _11495_;
  wire _11496_;
  wire _11497_;
  wire _11498_;
  wire _11499_;
  wire _11500_;
  wire _11501_;
  wire _11502_;
  wire _11503_;
  wire _11504_;
  wire _11505_;
  wire _11506_;
  wire _11507_;
  wire _11508_;
  wire _11509_;
  wire _11510_;
  wire _11511_;
  wire _11512_;
  wire _11513_;
  wire _11514_;
  wire _11515_;
  wire _11516_;
  wire _11517_;
  wire _11518_;
  wire _11519_;
  wire _11520_;
  wire _11521_;
  wire _11522_;
  wire _11523_;
  wire _11524_;
  wire _11525_;
  wire _11526_;
  wire _11527_;
  wire _11528_;
  wire _11529_;
  wire _11530_;
  wire _11531_;
  wire _11532_;
  wire _11533_;
  wire _11534_;
  wire _11535_;
  wire _11536_;
  wire _11537_;
  wire _11538_;
  wire _11539_;
  wire _11540_;
  wire _11541_;
  wire _11542_;
  wire _11543_;
  wire _11544_;
  wire _11545_;
  wire _11546_;
  wire _11547_;
  wire _11548_;
  wire _11549_;
  wire _11550_;
  wire _11551_;
  wire _11552_;
  wire _11553_;
  wire _11554_;
  wire _11555_;
  wire _11556_;
  wire _11557_;
  wire _11558_;
  wire _11559_;
  wire _11560_;
  wire _11561_;
  wire _11562_;
  wire _11563_;
  wire _11564_;
  wire _11565_;
  wire _11566_;
  wire _11567_;
  wire _11568_;
  wire _11569_;
  wire _11570_;
  wire _11571_;
  wire _11572_;
  wire _11573_;
  wire _11574_;
  wire _11575_;
  wire _11576_;
  wire _11577_;
  wire _11578_;
  wire _11579_;
  wire _11580_;
  wire _11581_;
  wire _11582_;
  wire _11583_;
  wire _11584_;
  wire _11585_;
  wire _11586_;
  wire _11587_;
  wire _11588_;
  wire _11589_;
  wire _11590_;
  wire _11591_;
  wire _11592_;
  wire _11593_;
  wire _11594_;
  wire _11595_;
  wire _11596_;
  wire _11597_;
  wire _11598_;
  wire _11599_;
  wire _11600_;
  wire _11601_;
  wire _11602_;
  wire _11603_;
  wire _11604_;
  wire _11605_;
  wire _11606_;
  wire _11607_;
  wire _11608_;
  wire _11609_;
  wire _11610_;
  wire _11611_;
  wire _11612_;
  wire _11613_;
  wire _11614_;
  wire _11615_;
  wire _11616_;
  wire _11617_;
  wire _11618_;
  wire _11619_;
  wire _11620_;
  wire _11621_;
  wire _11622_;
  wire _11623_;
  wire _11624_;
  wire _11625_;
  wire _11626_;
  wire _11627_;
  wire _11628_;
  wire _11629_;
  wire _11630_;
  wire _11631_;
  wire _11632_;
  wire _11633_;
  wire _11634_;
  wire _11635_;
  wire _11636_;
  wire _11637_;
  wire _11638_;
  wire _11639_;
  wire _11640_;
  wire _11641_;
  wire _11642_;
  wire _11643_;
  wire _11644_;
  wire _11645_;
  wire _11646_;
  wire _11647_;
  wire _11648_;
  wire _11649_;
  wire _11650_;
  wire _11651_;
  wire _11652_;
  wire _11653_;
  wire _11654_;
  wire _11655_;
  wire _11656_;
  wire _11657_;
  wire _11658_;
  wire _11659_;
  wire _11660_;
  wire _11661_;
  wire _11662_;
  wire _11663_;
  wire _11664_;
  wire _11665_;
  wire _11666_;
  wire _11667_;
  wire _11668_;
  wire _11669_;
  wire _11670_;
  wire _11671_;
  wire _11672_;
  wire _11673_;
  wire _11674_;
  wire _11675_;
  wire _11676_;
  wire _11677_;
  wire _11678_;
  wire _11679_;
  wire _11680_;
  wire _11681_;
  wire _11682_;
  wire _11683_;
  wire _11684_;
  wire _11685_;
  wire _11686_;
  wire _11687_;
  wire _11688_;
  wire _11689_;
  wire _11690_;
  wire _11691_;
  wire _11692_;
  wire _11693_;
  wire _11694_;
  wire _11695_;
  wire _11696_;
  wire _11697_;
  wire _11698_;
  wire _11699_;
  wire _11700_;
  wire _11701_;
  wire _11702_;
  wire _11703_;
  wire _11704_;
  wire _11705_;
  wire _11706_;
  wire _11707_;
  wire _11708_;
  wire _11709_;
  wire _11710_;
  wire _11711_;
  wire _11712_;
  wire _11713_;
  wire _11714_;
  wire _11715_;
  wire _11716_;
  wire _11717_;
  wire _11718_;
  wire _11719_;
  wire _11720_;
  wire _11721_;
  wire _11722_;
  wire _11723_;
  wire _11724_;
  wire _11725_;
  wire _11726_;
  wire _11727_;
  wire _11728_;
  wire _11729_;
  wire _11730_;
  wire _11731_;
  wire _11732_;
  wire _11733_;
  wire _11734_;
  wire _11735_;
  wire _11736_;
  wire _11737_;
  wire _11738_;
  wire _11739_;
  wire _11740_;
  wire _11741_;
  wire _11742_;
  wire _11743_;
  wire _11744_;
  wire _11745_;
  wire _11746_;
  wire _11747_;
  wire _11748_;
  wire _11749_;
  wire _11750_;
  wire _11751_;
  wire _11752_;
  wire _11753_;
  wire _11754_;
  wire _11755_;
  wire _11756_;
  wire _11757_;
  wire _11758_;
  wire _11759_;
  wire _11760_;
  wire _11761_;
  wire _11762_;
  wire _11763_;
  wire _11764_;
  wire _11765_;
  wire _11766_;
  wire _11767_;
  wire _11768_;
  wire _11769_;
  wire _11770_;
  wire _11771_;
  wire _11772_;
  wire _11773_;
  wire _11774_;
  wire _11775_;
  wire _11776_;
  wire _11777_;
  wire _11778_;
  wire _11779_;
  wire _11780_;
  wire _11781_;
  wire _11782_;
  wire _11783_;
  wire _11784_;
  wire _11785_;
  wire _11786_;
  wire _11787_;
  wire _11788_;
  wire _11789_;
  wire _11790_;
  wire _11791_;
  wire _11792_;
  wire _11793_;
  wire _11794_;
  wire _11795_;
  wire _11796_;
  wire _11797_;
  wire _11798_;
  wire _11799_;
  wire _11800_;
  wire _11801_;
  wire _11802_;
  wire _11803_;
  wire _11804_;
  wire _11805_;
  wire _11806_;
  wire _11807_;
  wire _11808_;
  wire _11809_;
  wire _11810_;
  wire _11811_;
  wire _11812_;
  wire _11813_;
  wire _11814_;
  wire _11815_;
  wire _11816_;
  wire _11817_;
  wire _11818_;
  wire _11819_;
  wire _11820_;
  wire _11821_;
  wire _11822_;
  wire _11823_;
  wire _11824_;
  wire _11825_;
  wire _11826_;
  wire _11827_;
  wire _11828_;
  wire _11829_;
  wire _11830_;
  wire _11831_;
  wire _11832_;
  wire _11833_;
  wire _11834_;
  wire _11835_;
  wire _11836_;
  wire _11837_;
  wire _11838_;
  wire _11839_;
  wire _11840_;
  wire _11841_;
  wire _11842_;
  wire _11843_;
  wire _11844_;
  wire _11845_;
  wire _11846_;
  wire _11847_;
  wire _11848_;
  wire _11849_;
  wire _11850_;
  wire _11851_;
  wire _11852_;
  wire _11853_;
  wire _11854_;
  wire _11855_;
  wire _11856_;
  wire _11857_;
  wire _11858_;
  wire _11859_;
  wire _11860_;
  wire _11861_;
  wire _11862_;
  wire _11863_;
  wire _11864_;
  wire _11865_;
  wire _11866_;
  wire _11867_;
  wire _11868_;
  wire _11869_;
  wire _11870_;
  wire _11871_;
  wire _11872_;
  wire _11873_;
  wire _11874_;
  wire _11875_;
  wire _11876_;
  wire _11877_;
  wire _11878_;
  wire _11879_;
  wire _11880_;
  wire _11881_;
  wire _11882_;
  wire _11883_;
  wire _11884_;
  wire _11885_;
  wire _11886_;
  wire _11887_;
  wire _11888_;
  wire _11889_;
  wire _11890_;
  wire _11891_;
  wire _11892_;
  wire _11893_;
  wire _11894_;
  wire _11895_;
  wire _11896_;
  wire _11897_;
  wire _11898_;
  wire _11899_;
  wire _11900_;
  wire _11901_;
  wire _11902_;
  wire _11903_;
  wire _11904_;
  wire _11905_;
  wire _11906_;
  wire _11907_;
  wire _11908_;
  wire _11909_;
  wire _11910_;
  wire _11911_;
  wire _11912_;
  wire _11913_;
  wire _11914_;
  wire _11915_;
  wire _11916_;
  wire _11917_;
  wire _11918_;
  wire _11919_;
  wire _11920_;
  wire _11921_;
  wire _11922_;
  wire _11923_;
  wire _11924_;
  wire _11925_;
  wire _11926_;
  wire _11927_;
  wire _11928_;
  wire _11929_;
  wire _11930_;
  wire _11931_;
  wire _11932_;
  wire _11933_;
  wire _11934_;
  wire _11935_;
  wire _11936_;
  wire _11937_;
  wire _11938_;
  wire _11939_;
  wire _11940_;
  wire _11941_;
  wire _11942_;
  wire _11943_;
  wire _11944_;
  wire _11945_;
  wire _11946_;
  wire _11947_;
  wire _11948_;
  wire _11949_;
  wire _11950_;
  wire _11951_;
  wire _11952_;
  wire _11953_;
  wire _11954_;
  wire _11955_;
  wire _11956_;
  wire _11957_;
  wire _11958_;
  wire _11959_;
  wire _11960_;
  wire _11961_;
  wire _11962_;
  wire _11963_;
  wire _11964_;
  wire _11965_;
  wire _11966_;
  wire _11967_;
  wire _11968_;
  wire _11969_;
  wire _11970_;
  wire _11971_;
  wire _11972_;
  wire _11973_;
  wire _11974_;
  wire _11975_;
  wire _11976_;
  wire _11977_;
  wire _11978_;
  wire _11979_;
  wire _11980_;
  wire _11981_;
  wire _11982_;
  wire _11983_;
  wire _11984_;
  wire _11985_;
  wire _11986_;
  wire _11987_;
  wire _11988_;
  wire _11989_;
  wire _11990_;
  wire _11991_;
  wire _11992_;
  wire _11993_;
  wire _11994_;
  wire _11995_;
  wire _11996_;
  wire _11997_;
  wire _11998_;
  wire _11999_;
  wire _12000_;
  wire _12001_;
  wire _12002_;
  wire _12003_;
  wire _12004_;
  wire _12005_;
  wire _12006_;
  wire _12007_;
  wire _12008_;
  wire _12009_;
  wire _12010_;
  wire _12011_;
  wire _12012_;
  wire _12013_;
  wire _12014_;
  wire _12015_;
  wire _12016_;
  wire _12017_;
  wire _12018_;
  wire _12019_;
  wire _12020_;
  wire _12021_;
  wire _12022_;
  wire _12023_;
  wire _12024_;
  wire _12025_;
  wire _12026_;
  wire _12027_;
  wire _12028_;
  wire _12029_;
  wire _12030_;
  wire _12031_;
  wire _12032_;
  wire _12033_;
  wire _12034_;
  wire _12035_;
  wire _12036_;
  wire _12037_;
  wire _12038_;
  wire _12039_;
  wire _12040_;
  wire _12041_;
  wire _12042_;
  wire _12043_;
  wire _12044_;
  wire _12045_;
  wire _12046_;
  wire _12047_;
  wire _12048_;
  wire _12049_;
  wire _12050_;
  wire _12051_;
  wire _12052_;
  wire _12053_;
  wire _12054_;
  wire _12055_;
  wire _12056_;
  wire _12057_;
  wire _12058_;
  wire _12059_;
  wire _12060_;
  wire _12061_;
  wire _12062_;
  wire _12063_;
  wire _12064_;
  wire _12065_;
  wire _12066_;
  wire _12067_;
  wire _12068_;
  wire _12069_;
  wire _12070_;
  wire _12071_;
  wire _12072_;
  wire _12073_;
  wire _12074_;
  wire _12075_;
  wire _12076_;
  wire _12077_;
  wire _12078_;
  wire _12079_;
  wire _12080_;
  wire _12081_;
  wire _12082_;
  wire _12083_;
  wire _12084_;
  wire _12085_;
  wire _12086_;
  wire _12087_;
  wire _12088_;
  wire _12089_;
  wire _12090_;
  wire _12091_;
  wire _12092_;
  wire _12093_;
  wire _12094_;
  wire _12095_;
  wire _12096_;
  wire _12097_;
  wire _12098_;
  wire _12099_;
  wire _12100_;
  wire _12101_;
  wire _12102_;
  wire _12103_;
  wire _12104_;
  wire _12105_;
  wire _12106_;
  wire _12107_;
  wire _12108_;
  wire _12109_;
  wire _12110_;
  wire _12111_;
  wire _12112_;
  wire _12113_;
  wire _12114_;
  wire _12115_;
  wire _12116_;
  wire _12117_;
  wire _12118_;
  wire _12119_;
  wire _12120_;
  wire _12121_;
  wire _12122_;
  wire _12123_;
  wire _12124_;
  wire _12125_;
  wire _12126_;
  wire _12127_;
  wire _12128_;
  wire _12129_;
  wire _12130_;
  wire _12131_;
  wire _12132_;
  wire _12133_;
  wire _12134_;
  wire _12135_;
  wire _12136_;
  wire _12137_;
  wire _12138_;
  wire _12139_;
  wire _12140_;
  wire _12141_;
  wire _12142_;
  wire _12143_;
  wire _12144_;
  wire _12145_;
  wire _12146_;
  wire _12147_;
  wire _12148_;
  wire _12149_;
  wire _12150_;
  wire _12151_;
  wire _12152_;
  wire _12153_;
  wire _12154_;
  wire _12155_;
  wire _12156_;
  wire _12157_;
  wire _12158_;
  wire _12159_;
  wire _12160_;
  wire _12161_;
  wire _12162_;
  wire _12163_;
  wire _12164_;
  wire _12165_;
  wire _12166_;
  wire _12167_;
  wire _12168_;
  wire _12169_;
  wire _12170_;
  wire _12171_;
  wire _12172_;
  wire _12173_;
  wire _12174_;
  wire _12175_;
  wire _12176_;
  wire _12177_;
  wire _12178_;
  wire _12179_;
  wire _12180_;
  wire _12181_;
  wire _12182_;
  wire _12183_;
  wire _12184_;
  wire _12185_;
  wire _12186_;
  wire _12187_;
  wire _12188_;
  wire _12189_;
  wire _12190_;
  wire _12191_;
  wire _12192_;
  wire _12193_;
  wire _12194_;
  wire _12195_;
  wire _12196_;
  wire _12197_;
  wire _12198_;
  wire _12199_;
  wire _12200_;
  wire _12201_;
  wire _12202_;
  wire _12203_;
  wire _12204_;
  wire _12205_;
  wire _12206_;
  wire _12207_;
  wire _12208_;
  wire _12209_;
  wire _12210_;
  wire _12211_;
  wire _12212_;
  wire _12213_;
  wire _12214_;
  wire _12215_;
  wire _12216_;
  wire _12217_;
  wire _12218_;
  wire _12219_;
  wire _12220_;
  wire _12221_;
  wire _12222_;
  wire _12223_;
  wire _12224_;
  wire _12225_;
  wire _12226_;
  wire _12227_;
  wire _12228_;
  wire _12229_;
  wire _12230_;
  wire _12231_;
  wire _12232_;
  wire _12233_;
  wire _12234_;
  wire _12235_;
  wire _12236_;
  wire _12237_;
  wire _12238_;
  wire _12239_;
  wire _12240_;
  wire _12241_;
  wire _12242_;
  wire _12243_;
  wire _12244_;
  wire _12245_;
  wire _12246_;
  wire _12247_;
  wire _12248_;
  wire _12249_;
  wire _12250_;
  wire _12251_;
  wire _12252_;
  wire _12253_;
  wire _12254_;
  wire _12255_;
  wire _12256_;
  wire _12257_;
  wire _12258_;
  wire _12259_;
  wire _12260_;
  wire _12261_;
  wire _12262_;
  wire _12263_;
  wire _12264_;
  wire _12265_;
  wire _12266_;
  wire _12267_;
  wire _12268_;
  wire _12269_;
  wire _12270_;
  wire _12271_;
  wire _12272_;
  wire _12273_;
  wire _12274_;
  wire _12275_;
  wire _12276_;
  wire _12277_;
  wire _12278_;
  wire _12279_;
  wire _12280_;
  wire _12281_;
  wire _12282_;
  wire _12283_;
  wire _12284_;
  wire _12285_;
  wire _12286_;
  wire _12287_;
  wire _12288_;
  wire _12289_;
  wire _12290_;
  wire _12291_;
  wire _12292_;
  wire _12293_;
  wire _12294_;
  wire _12295_;
  wire _12296_;
  wire _12297_;
  wire _12298_;
  wire _12299_;
  wire _12300_;
  wire _12301_;
  wire _12302_;
  wire _12303_;
  wire _12304_;
  wire _12305_;
  wire _12306_;
  wire _12307_;
  wire _12308_;
  wire _12309_;
  wire _12310_;
  wire _12311_;
  wire _12312_;
  wire _12313_;
  wire _12314_;
  wire _12315_;
  wire _12316_;
  wire _12317_;
  wire _12318_;
  wire _12319_;
  wire _12320_;
  wire _12321_;
  wire _12322_;
  wire _12323_;
  wire _12324_;
  wire _12325_;
  wire _12326_;
  wire _12327_;
  wire _12328_;
  wire _12329_;
  wire _12330_;
  wire _12331_;
  wire _12332_;
  wire _12333_;
  wire _12334_;
  wire _12335_;
  wire _12336_;
  wire _12337_;
  wire _12338_;
  wire _12339_;
  wire _12340_;
  wire _12341_;
  wire _12342_;
  wire _12343_;
  wire _12344_;
  wire _12345_;
  wire _12346_;
  wire _12347_;
  wire _12348_;
  wire _12349_;
  wire _12350_;
  wire _12351_;
  wire _12352_;
  wire _12353_;
  wire _12354_;
  wire _12355_;
  wire _12356_;
  wire _12357_;
  wire _12358_;
  wire _12359_;
  wire _12360_;
  wire _12361_;
  wire _12362_;
  wire _12363_;
  wire _12364_;
  wire _12365_;
  wire _12366_;
  wire _12367_;
  wire _12368_;
  wire _12369_;
  wire _12370_;
  wire _12371_;
  wire _12372_;
  wire _12373_;
  wire _12374_;
  wire _12375_;
  wire _12376_;
  wire _12377_;
  wire _12378_;
  wire _12379_;
  wire _12380_;
  wire _12381_;
  wire _12382_;
  wire _12383_;
  wire _12384_;
  wire _12385_;
  wire _12386_;
  wire _12387_;
  wire _12388_;
  wire _12389_;
  wire _12390_;
  wire _12391_;
  wire _12392_;
  wire _12393_;
  wire _12394_;
  wire _12395_;
  wire _12396_;
  wire _12397_;
  wire _12398_;
  wire _12399_;
  wire _12400_;
  wire _12401_;
  wire _12402_;
  wire _12403_;
  wire _12404_;
  wire _12405_;
  wire _12406_;
  wire _12407_;
  wire _12408_;
  wire _12409_;
  wire _12410_;
  wire _12411_;
  wire _12412_;
  wire _12413_;
  wire _12414_;
  wire _12415_;
  wire _12416_;
  wire _12417_;
  wire _12418_;
  wire _12419_;
  wire _12420_;
  wire _12421_;
  wire _12422_;
  wire _12423_;
  wire _12424_;
  wire _12425_;
  wire _12426_;
  wire _12427_;
  wire _12428_;
  wire _12429_;
  wire _12430_;
  wire _12431_;
  wire _12432_;
  wire _12433_;
  wire _12434_;
  wire _12435_;
  wire _12436_;
  wire _12437_;
  wire _12438_;
  wire _12439_;
  wire _12440_;
  wire _12441_;
  wire _12442_;
  wire _12443_;
  wire _12444_;
  wire _12445_;
  wire _12446_;
  wire _12447_;
  wire _12448_;
  wire _12449_;
  wire _12450_;
  wire _12451_;
  wire _12452_;
  wire _12453_;
  wire _12454_;
  wire _12455_;
  wire _12456_;
  wire _12457_;
  wire _12458_;
  wire _12459_;
  wire _12460_;
  wire _12461_;
  wire _12462_;
  wire _12463_;
  wire _12464_;
  wire _12465_;
  wire _12466_;
  wire _12467_;
  wire _12468_;
  wire _12469_;
  wire _12470_;
  wire _12471_;
  wire _12472_;
  wire _12473_;
  wire _12474_;
  wire _12475_;
  wire _12476_;
  wire _12477_;
  wire _12478_;
  wire _12479_;
  wire _12480_;
  wire _12481_;
  wire _12482_;
  wire _12483_;
  wire _12484_;
  wire _12485_;
  wire _12486_;
  wire _12487_;
  wire _12488_;
  wire _12489_;
  wire _12490_;
  wire _12491_;
  wire _12492_;
  wire _12493_;
  wire _12494_;
  wire _12495_;
  wire _12496_;
  wire _12497_;
  wire _12498_;
  wire _12499_;
  wire _12500_;
  wire _12501_;
  wire _12502_;
  wire _12503_;
  wire _12504_;
  wire _12505_;
  wire _12506_;
  wire _12507_;
  wire _12508_;
  wire _12509_;
  wire _12510_;
  wire _12511_;
  wire _12512_;
  wire _12513_;
  wire _12514_;
  wire _12515_;
  wire _12516_;
  wire _12517_;
  wire _12518_;
  wire _12519_;
  wire _12520_;
  wire _12521_;
  wire _12522_;
  wire _12523_;
  wire _12524_;
  wire _12525_;
  wire _12526_;
  wire _12527_;
  wire _12528_;
  wire _12529_;
  wire _12530_;
  wire _12531_;
  wire _12532_;
  wire _12533_;
  wire _12534_;
  wire _12535_;
  wire _12536_;
  wire _12537_;
  wire _12538_;
  wire _12539_;
  wire _12540_;
  wire _12541_;
  wire _12542_;
  wire _12543_;
  wire _12544_;
  wire _12545_;
  wire _12546_;
  wire _12547_;
  wire _12548_;
  wire _12549_;
  wire _12550_;
  wire _12551_;
  wire _12552_;
  wire _12553_;
  wire _12554_;
  wire _12555_;
  wire _12556_;
  wire _12557_;
  wire _12558_;
  wire _12559_;
  wire _12560_;
  wire _12561_;
  wire _12562_;
  wire _12563_;
  wire _12564_;
  wire _12565_;
  wire _12566_;
  wire _12567_;
  wire _12568_;
  wire _12569_;
  wire _12570_;
  wire _12571_;
  wire _12572_;
  wire _12573_;
  wire _12574_;
  wire _12575_;
  wire _12576_;
  wire _12577_;
  wire _12578_;
  wire _12579_;
  wire _12580_;
  wire _12581_;
  wire _12582_;
  wire _12583_;
  wire _12584_;
  wire _12585_;
  wire _12586_;
  wire _12587_;
  wire _12588_;
  wire _12589_;
  wire _12590_;
  wire _12591_;
  wire _12592_;
  wire _12593_;
  wire _12594_;
  wire _12595_;
  wire _12596_;
  wire _12597_;
  wire _12598_;
  wire _12599_;
  wire _12600_;
  wire _12601_;
  wire _12602_;
  wire _12603_;
  wire _12604_;
  wire _12605_;
  wire _12606_;
  wire _12607_;
  wire _12608_;
  wire _12609_;
  wire _12610_;
  wire _12611_;
  wire _12612_;
  wire _12613_;
  wire _12614_;
  wire _12615_;
  wire _12616_;
  wire _12617_;
  wire _12618_;
  wire _12619_;
  wire _12620_;
  wire _12621_;
  wire _12622_;
  wire _12623_;
  wire _12624_;
  wire _12625_;
  wire _12626_;
  wire _12627_;
  wire _12628_;
  wire _12629_;
  wire _12630_;
  wire _12631_;
  wire _12632_;
  wire _12633_;
  wire _12634_;
  wire _12635_;
  wire _12636_;
  wire _12637_;
  wire _12638_;
  wire _12639_;
  wire _12640_;
  wire _12641_;
  wire _12642_;
  wire _12643_;
  wire _12644_;
  wire _12645_;
  wire _12646_;
  wire _12647_;
  wire _12648_;
  wire _12649_;
  wire _12650_;
  wire _12651_;
  wire _12652_;
  wire _12653_;
  wire _12654_;
  wire _12655_;
  wire _12656_;
  wire _12657_;
  wire _12658_;
  wire _12659_;
  wire _12660_;
  wire _12661_;
  wire _12662_;
  wire _12663_;
  wire _12664_;
  wire _12665_;
  wire _12666_;
  wire _12667_;
  wire _12668_;
  wire _12669_;
  wire _12670_;
  wire _12671_;
  wire _12672_;
  wire _12673_;
  wire _12674_;
  wire _12675_;
  wire _12676_;
  wire _12677_;
  wire _12678_;
  wire _12679_;
  wire _12680_;
  wire _12681_;
  wire _12682_;
  wire _12683_;
  wire _12684_;
  wire _12685_;
  wire _12686_;
  wire _12687_;
  wire _12688_;
  wire _12689_;
  wire _12690_;
  wire _12691_;
  wire _12692_;
  wire _12693_;
  wire _12694_;
  wire _12695_;
  wire _12696_;
  wire _12697_;
  wire _12698_;
  wire _12699_;
  wire _12700_;
  wire _12701_;
  wire _12702_;
  wire _12703_;
  wire _12704_;
  wire _12705_;
  wire _12706_;
  wire _12707_;
  wire _12708_;
  wire _12709_;
  wire _12710_;
  wire _12711_;
  wire _12712_;
  wire _12713_;
  wire _12714_;
  wire _12715_;
  wire _12716_;
  wire _12717_;
  wire _12718_;
  wire _12719_;
  wire _12720_;
  wire _12721_;
  wire _12722_;
  wire _12723_;
  wire _12724_;
  wire _12725_;
  wire _12726_;
  wire _12727_;
  wire _12728_;
  wire _12729_;
  wire _12730_;
  wire _12731_;
  wire _12732_;
  wire _12733_;
  wire _12734_;
  wire _12735_;
  wire _12736_;
  wire _12737_;
  wire _12738_;
  wire _12739_;
  wire _12740_;
  wire _12741_;
  wire _12742_;
  wire _12743_;
  wire _12744_;
  wire _12745_;
  wire _12746_;
  wire _12747_;
  wire _12748_;
  wire _12749_;
  wire _12750_;
  wire _12751_;
  wire _12752_;
  wire _12753_;
  wire _12754_;
  wire _12755_;
  wire _12756_;
  wire _12757_;
  wire _12758_;
  wire _12759_;
  wire _12760_;
  wire _12761_;
  wire _12762_;
  wire _12763_;
  wire _12764_;
  wire _12765_;
  wire _12766_;
  wire _12767_;
  wire _12768_;
  wire _12769_;
  wire _12770_;
  wire _12771_;
  wire _12772_;
  wire _12773_;
  wire _12774_;
  wire _12775_;
  wire _12776_;
  wire _12777_;
  wire _12778_;
  wire _12779_;
  wire _12780_;
  wire _12781_;
  wire _12782_;
  wire _12783_;
  wire _12784_;
  wire _12785_;
  wire _12786_;
  wire _12787_;
  wire _12788_;
  wire _12789_;
  wire _12790_;
  wire _12791_;
  wire _12792_;
  wire _12793_;
  wire _12794_;
  wire _12795_;
  wire _12796_;
  wire _12797_;
  wire _12798_;
  wire _12799_;
  wire _12800_;
  wire _12801_;
  wire _12802_;
  wire _12803_;
  wire _12804_;
  wire _12805_;
  wire _12806_;
  wire _12807_;
  wire _12808_;
  wire _12809_;
  wire _12810_;
  wire _12811_;
  wire _12812_;
  wire _12813_;
  wire _12814_;
  wire _12815_;
  wire _12816_;
  wire _12817_;
  wire _12818_;
  wire _12819_;
  wire _12820_;
  wire _12821_;
  wire _12822_;
  wire _12823_;
  wire _12824_;
  wire _12825_;
  wire _12826_;
  wire _12827_;
  wire _12828_;
  wire _12829_;
  wire _12830_;
  wire _12831_;
  wire _12832_;
  wire _12833_;
  wire _12834_;
  wire _12835_;
  wire _12836_;
  wire _12837_;
  wire _12838_;
  wire _12839_;
  wire _12840_;
  wire _12841_;
  wire _12842_;
  wire _12843_;
  wire _12844_;
  wire _12845_;
  wire _12846_;
  wire _12847_;
  wire _12848_;
  wire _12849_;
  wire _12850_;
  wire _12851_;
  wire _12852_;
  wire _12853_;
  wire _12854_;
  wire _12855_;
  wire _12856_;
  wire _12857_;
  wire _12858_;
  wire _12859_;
  wire _12860_;
  wire _12861_;
  wire _12862_;
  wire _12863_;
  wire _12864_;
  wire _12865_;
  wire _12866_;
  wire _12867_;
  wire _12868_;
  wire _12869_;
  wire _12870_;
  wire _12871_;
  wire _12872_;
  wire _12873_;
  wire _12874_;
  wire _12875_;
  wire _12876_;
  wire _12877_;
  wire _12878_;
  wire _12879_;
  wire _12880_;
  wire _12881_;
  wire _12882_;
  wire _12883_;
  wire _12884_;
  wire _12885_;
  wire _12886_;
  wire _12887_;
  wire _12888_;
  wire _12889_;
  wire _12890_;
  wire _12891_;
  wire _12892_;
  wire _12893_;
  wire _12894_;
  wire _12895_;
  wire _12896_;
  wire _12897_;
  wire _12898_;
  wire _12899_;
  wire _12900_;
  wire _12901_;
  wire _12902_;
  wire _12903_;
  wire _12904_;
  wire _12905_;
  wire _12906_;
  wire _12907_;
  wire _12908_;
  wire _12909_;
  wire _12910_;
  wire _12911_;
  wire _12912_;
  wire _12913_;
  wire _12914_;
  wire _12915_;
  wire _12916_;
  wire _12917_;
  wire _12918_;
  wire _12919_;
  wire _12920_;
  wire _12921_;
  wire _12922_;
  wire _12923_;
  wire _12924_;
  wire _12925_;
  wire _12926_;
  wire _12927_;
  wire _12928_;
  wire _12929_;
  wire _12930_;
  wire _12931_;
  wire _12932_;
  wire _12933_;
  wire _12934_;
  wire _12935_;
  wire _12936_;
  wire _12937_;
  wire _12938_;
  wire _12939_;
  wire _12940_;
  wire _12941_;
  wire _12942_;
  wire _12943_;
  wire _12944_;
  wire _12945_;
  wire _12946_;
  wire _12947_;
  wire _12948_;
  wire _12949_;
  wire _12950_;
  wire _12951_;
  wire _12952_;
  wire _12953_;
  wire _12954_;
  wire _12955_;
  wire _12956_;
  wire _12957_;
  wire _12958_;
  wire _12959_;
  wire _12960_;
  wire _12961_;
  wire _12962_;
  wire _12963_;
  wire _12964_;
  wire _12965_;
  wire _12966_;
  wire _12967_;
  wire _12968_;
  wire _12969_;
  wire _12970_;
  wire _12971_;
  wire _12972_;
  wire _12973_;
  wire _12974_;
  wire _12975_;
  wire _12976_;
  wire _12977_;
  wire _12978_;
  wire _12979_;
  wire _12980_;
  wire _12981_;
  wire _12982_;
  wire _12983_;
  wire _12984_;
  wire _12985_;
  wire _12986_;
  wire _12987_;
  wire _12988_;
  wire _12989_;
  wire _12990_;
  wire _12991_;
  wire _12992_;
  wire _12993_;
  wire _12994_;
  wire _12995_;
  wire _12996_;
  wire _12997_;
  wire _12998_;
  wire _12999_;
  wire _13000_;
  wire _13001_;
  wire _13002_;
  wire _13003_;
  wire _13004_;
  wire _13005_;
  wire _13006_;
  wire _13007_;
  wire _13008_;
  wire _13009_;
  wire _13010_;
  wire _13011_;
  wire _13012_;
  wire _13013_;
  wire _13014_;
  wire _13015_;
  wire _13016_;
  wire _13017_;
  wire _13018_;
  wire _13019_;
  wire _13020_;
  wire _13021_;
  wire _13022_;
  wire _13023_;
  wire _13024_;
  wire _13025_;
  wire _13026_;
  wire _13027_;
  wire _13028_;
  wire _13029_;
  wire _13030_;
  wire _13031_;
  wire _13032_;
  wire _13033_;
  wire _13034_;
  wire _13035_;
  wire _13036_;
  wire _13037_;
  wire _13038_;
  wire _13039_;
  wire _13040_;
  wire _13041_;
  wire _13042_;
  wire _13043_;
  wire _13044_;
  wire _13045_;
  wire _13046_;
  wire _13047_;
  wire _13048_;
  wire _13049_;
  wire _13050_;
  wire _13051_;
  wire _13052_;
  wire _13053_;
  wire _13054_;
  wire _13055_;
  wire _13056_;
  wire _13057_;
  wire _13058_;
  wire _13059_;
  wire _13060_;
  wire _13061_;
  wire _13062_;
  wire _13063_;
  wire _13064_;
  wire _13065_;
  wire _13066_;
  wire _13067_;
  wire _13068_;
  wire _13069_;
  wire _13070_;
  wire _13071_;
  wire _13072_;
  wire _13073_;
  wire _13074_;
  wire _13075_;
  wire _13076_;
  wire _13077_;
  wire _13078_;
  wire _13079_;
  wire _13080_;
  wire _13081_;
  wire _13082_;
  wire _13083_;
  wire _13084_;
  wire _13085_;
  wire _13086_;
  wire _13087_;
  wire _13088_;
  wire _13089_;
  wire _13090_;
  wire _13091_;
  wire _13092_;
  wire _13093_;
  wire _13094_;
  wire _13095_;
  wire _13096_;
  wire _13097_;
  wire _13098_;
  wire _13099_;
  wire _13100_;
  wire _13101_;
  wire _13102_;
  wire _13103_;
  wire _13104_;
  wire _13105_;
  wire _13106_;
  wire _13107_;
  wire _13108_;
  wire _13109_;
  wire _13110_;
  wire _13111_;
  wire _13112_;
  wire _13113_;
  wire _13114_;
  wire _13115_;
  wire _13116_;
  wire _13117_;
  wire _13118_;
  wire _13119_;
  wire _13120_;
  wire _13121_;
  wire _13122_;
  wire _13123_;
  wire _13124_;
  wire _13125_;
  wire _13126_;
  wire _13127_;
  wire _13128_;
  wire _13129_;
  wire _13130_;
  wire _13131_;
  wire _13132_;
  wire _13133_;
  wire _13134_;
  wire _13135_;
  wire _13136_;
  wire _13137_;
  wire _13138_;
  wire _13139_;
  wire _13140_;
  wire _13141_;
  wire _13142_;
  wire _13143_;
  wire _13144_;
  wire _13145_;
  wire _13146_;
  wire _13147_;
  wire _13148_;
  wire _13149_;
  wire _13150_;
  wire _13151_;
  wire _13152_;
  wire _13153_;
  wire _13154_;
  wire _13155_;
  wire _13156_;
  wire _13157_;
  wire _13158_;
  wire _13159_;
  wire _13160_;
  wire _13161_;
  wire _13162_;
  wire _13163_;
  wire _13164_;
  wire _13165_;
  wire _13166_;
  wire _13167_;
  wire _13168_;
  wire _13169_;
  wire _13170_;
  wire _13171_;
  wire _13172_;
  wire _13173_;
  wire _13174_;
  wire _13175_;
  wire _13176_;
  wire _13177_;
  wire _13178_;
  wire _13179_;
  wire _13180_;
  wire _13181_;
  wire _13182_;
  wire _13183_;
  wire _13184_;
  wire _13185_;
  wire _13186_;
  wire _13187_;
  wire _13188_;
  wire _13189_;
  wire _13190_;
  wire _13191_;
  wire _13192_;
  wire _13193_;
  wire _13194_;
  wire _13195_;
  wire _13196_;
  wire _13197_;
  wire _13198_;
  wire _13199_;
  wire _13200_;
  wire _13201_;
  wire _13202_;
  wire _13203_;
  wire _13204_;
  wire _13205_;
  wire _13206_;
  wire _13207_;
  wire _13208_;
  wire _13209_;
  wire _13210_;
  wire _13211_;
  wire _13212_;
  wire _13213_;
  wire _13214_;
  wire _13215_;
  wire _13216_;
  wire _13217_;
  wire _13218_;
  wire _13219_;
  wire _13220_;
  wire _13221_;
  wire _13222_;
  wire _13223_;
  wire _13224_;
  wire _13225_;
  wire _13226_;
  wire _13227_;
  wire _13228_;
  wire _13229_;
  wire _13230_;
  wire _13231_;
  wire _13232_;
  wire _13233_;
  wire _13234_;
  wire _13235_;
  wire _13236_;
  wire _13237_;
  wire _13238_;
  wire _13239_;
  wire _13240_;
  wire _13241_;
  wire _13242_;
  wire _13243_;
  wire _13244_;
  wire _13245_;
  wire _13246_;
  wire _13247_;
  wire _13248_;
  wire _13249_;
  wire _13250_;
  wire _13251_;
  wire _13252_;
  wire _13253_;
  wire _13254_;
  wire _13255_;
  wire _13256_;
  wire _13257_;
  wire _13258_;
  wire _13259_;
  wire _13260_;
  wire _13261_;
  wire _13262_;
  wire _13263_;
  wire _13264_;
  wire _13265_;
  wire _13266_;
  wire _13267_;
  wire _13268_;
  wire _13269_;
  wire _13270_;
  wire _13271_;
  wire _13272_;
  wire _13273_;
  wire _13274_;
  wire _13275_;
  wire _13276_;
  wire _13277_;
  wire _13278_;
  wire _13279_;
  wire _13280_;
  wire _13281_;
  wire _13282_;
  wire _13283_;
  wire _13284_;
  wire _13285_;
  wire _13286_;
  wire _13287_;
  wire _13288_;
  wire _13289_;
  wire _13290_;
  wire _13291_;
  wire _13292_;
  wire _13293_;
  wire _13294_;
  wire _13295_;
  wire _13296_;
  wire _13297_;
  wire _13298_;
  wire _13299_;
  wire _13300_;
  wire _13301_;
  wire _13302_;
  wire _13303_;
  wire _13304_;
  wire _13305_;
  wire _13306_;
  wire _13307_;
  wire _13308_;
  wire _13309_;
  wire _13310_;
  wire _13311_;
  wire _13312_;
  wire _13313_;
  wire _13314_;
  wire _13315_;
  wire _13316_;
  wire _13317_;
  wire _13318_;
  wire _13319_;
  wire _13320_;
  wire _13321_;
  wire _13322_;
  wire _13323_;
  wire _13324_;
  wire _13325_;
  wire _13326_;
  wire _13327_;
  wire _13328_;
  wire _13329_;
  wire _13330_;
  wire _13331_;
  wire _13332_;
  wire _13333_;
  wire _13334_;
  wire _13335_;
  wire _13336_;
  wire _13337_;
  wire _13338_;
  wire _13339_;
  wire _13340_;
  wire _13341_;
  wire _13342_;
  wire _13343_;
  wire _13344_;
  wire _13345_;
  wire _13346_;
  wire _13347_;
  wire _13348_;
  wire _13349_;
  wire _13350_;
  wire _13351_;
  wire _13352_;
  wire _13353_;
  wire _13354_;
  wire _13355_;
  wire _13356_;
  wire _13357_;
  wire _13358_;
  wire _13359_;
  wire _13360_;
  wire _13361_;
  wire _13362_;
  wire _13363_;
  wire _13364_;
  wire _13365_;
  wire _13366_;
  wire _13367_;
  wire _13368_;
  wire _13369_;
  wire _13370_;
  wire _13371_;
  wire _13372_;
  wire _13373_;
  wire _13374_;
  wire _13375_;
  wire _13376_;
  wire _13377_;
  wire _13378_;
  wire _13379_;
  wire _13380_;
  wire _13381_;
  wire _13382_;
  wire _13383_;
  wire _13384_;
  wire _13385_;
  wire _13386_;
  wire _13387_;
  wire _13388_;
  wire _13389_;
  wire _13390_;
  wire _13391_;
  wire _13392_;
  wire _13393_;
  wire _13394_;
  wire _13395_;
  wire _13396_;
  wire _13397_;
  wire _13398_;
  wire _13399_;
  wire _13400_;
  wire _13401_;
  wire _13402_;
  wire _13403_;
  wire _13404_;
  wire _13405_;
  wire _13406_;
  wire _13407_;
  wire _13408_;
  wire _13409_;
  wire _13410_;
  wire _13411_;
  wire _13412_;
  wire _13413_;
  wire _13414_;
  wire _13415_;
  wire _13416_;
  wire _13417_;
  wire _13418_;
  wire _13419_;
  wire _13420_;
  wire _13421_;
  wire _13422_;
  wire _13423_;
  wire _13424_;
  wire _13425_;
  wire _13426_;
  wire _13427_;
  wire _13428_;
  wire _13429_;
  wire _13430_;
  wire _13431_;
  wire _13432_;
  wire _13433_;
  wire _13434_;
  wire _13435_;
  wire _13436_;
  wire _13437_;
  wire _13438_;
  wire _13439_;
  wire _13440_;
  wire _13441_;
  wire _13442_;
  wire _13443_;
  wire _13444_;
  wire _13445_;
  wire _13446_;
  wire _13447_;
  wire _13448_;
  wire _13449_;
  wire _13450_;
  wire _13451_;
  wire _13452_;
  wire _13453_;
  wire _13454_;
  wire _13455_;
  wire _13456_;
  wire _13457_;
  wire _13458_;
  wire _13459_;
  wire _13460_;
  wire _13461_;
  wire _13462_;
  wire _13463_;
  wire _13464_;
  wire _13465_;
  wire _13466_;
  wire _13467_;
  wire _13468_;
  wire _13469_;
  wire _13470_;
  wire _13471_;
  wire _13472_;
  wire _13473_;
  wire _13474_;
  wire _13475_;
  wire _13476_;
  wire _13477_;
  wire _13478_;
  wire _13479_;
  wire _13480_;
  wire _13481_;
  wire _13482_;
  wire _13483_;
  wire _13484_;
  wire _13485_;
  wire _13486_;
  wire _13487_;
  wire _13488_;
  wire _13489_;
  wire _13490_;
  wire _13491_;
  wire _13492_;
  wire _13493_;
  wire _13494_;
  wire _13495_;
  wire _13496_;
  wire _13497_;
  wire _13498_;
  wire _13499_;
  wire _13500_;
  wire _13501_;
  wire _13502_;
  wire _13503_;
  wire _13504_;
  wire _13505_;
  wire _13506_;
  wire _13507_;
  wire _13508_;
  wire _13509_;
  wire _13510_;
  wire _13511_;
  wire _13512_;
  wire _13513_;
  wire _13514_;
  wire _13515_;
  wire _13516_;
  wire _13517_;
  wire _13518_;
  wire _13519_;
  wire _13520_;
  wire _13521_;
  wire _13522_;
  wire _13523_;
  wire _13524_;
  wire _13525_;
  wire _13526_;
  wire _13527_;
  wire _13528_;
  wire _13529_;
  wire _13530_;
  wire _13531_;
  wire _13532_;
  wire _13533_;
  wire _13534_;
  wire _13535_;
  wire _13536_;
  wire _13537_;
  wire _13538_;
  wire _13539_;
  wire _13540_;
  wire _13541_;
  wire _13542_;
  wire _13543_;
  wire _13544_;
  wire _13545_;
  wire _13546_;
  wire _13547_;
  wire _13548_;
  wire _13549_;
  wire _13550_;
  wire _13551_;
  wire _13552_;
  wire _13553_;
  wire _13554_;
  wire _13555_;
  wire _13556_;
  wire _13557_;
  wire _13558_;
  wire _13559_;
  wire _13560_;
  wire _13561_;
  wire _13562_;
  wire _13563_;
  wire _13564_;
  wire _13565_;
  wire _13566_;
  wire _13567_;
  wire _13568_;
  wire _13569_;
  wire _13570_;
  wire _13571_;
  wire _13572_;
  wire _13573_;
  wire _13574_;
  wire _13575_;
  wire _13576_;
  wire _13577_;
  wire _13578_;
  wire _13579_;
  wire _13580_;
  wire _13581_;
  wire _13582_;
  wire _13583_;
  wire _13584_;
  wire _13585_;
  wire _13586_;
  wire _13587_;
  wire _13588_;
  wire _13589_;
  wire _13590_;
  wire _13591_;
  wire _13592_;
  wire _13593_;
  wire _13594_;
  wire _13595_;
  wire _13596_;
  wire _13597_;
  wire _13598_;
  wire _13599_;
  wire _13600_;
  wire _13601_;
  wire _13602_;
  wire _13603_;
  wire _13604_;
  wire _13605_;
  wire _13606_;
  wire _13607_;
  wire _13608_;
  wire _13609_;
  wire _13610_;
  wire _13611_;
  wire _13612_;
  wire _13613_;
  wire _13614_;
  wire _13615_;
  wire _13616_;
  wire _13617_;
  wire _13618_;
  wire _13619_;
  wire _13620_;
  wire _13621_;
  wire _13622_;
  wire _13623_;
  wire _13624_;
  wire _13625_;
  wire _13626_;
  wire _13627_;
  wire _13628_;
  wire _13629_;
  wire _13630_;
  wire _13631_;
  wire _13632_;
  wire _13633_;
  wire _13634_;
  wire _13635_;
  wire _13636_;
  wire _13637_;
  wire _13638_;
  wire _13639_;
  wire _13640_;
  wire _13641_;
  wire _13642_;
  wire _13643_;
  wire _13644_;
  wire _13645_;
  wire _13646_;
  wire _13647_;
  wire _13648_;
  wire _13649_;
  wire _13650_;
  wire _13651_;
  wire _13652_;
  wire _13653_;
  wire _13654_;
  wire _13655_;
  wire _13656_;
  wire _13657_;
  wire _13658_;
  wire _13659_;
  wire _13660_;
  wire _13661_;
  wire _13662_;
  wire _13663_;
  wire _13664_;
  wire _13665_;
  wire _13666_;
  wire _13667_;
  wire _13668_;
  wire _13669_;
  wire _13670_;
  wire _13671_;
  wire _13672_;
  wire _13673_;
  wire _13674_;
  wire _13675_;
  wire _13676_;
  wire _13677_;
  wire _13678_;
  wire _13679_;
  wire _13680_;
  wire _13681_;
  wire _13682_;
  wire _13683_;
  wire _13684_;
  wire _13685_;
  wire _13686_;
  wire _13687_;
  wire _13688_;
  wire _13689_;
  wire _13690_;
  wire _13691_;
  wire _13692_;
  wire _13693_;
  wire _13694_;
  wire _13695_;
  wire _13696_;
  wire _13697_;
  wire _13698_;
  wire _13699_;
  wire _13700_;
  wire _13701_;
  wire _13702_;
  wire _13703_;
  wire _13704_;
  wire _13705_;
  wire _13706_;
  wire _13707_;
  wire _13708_;
  wire _13709_;
  wire _13710_;
  wire _13711_;
  wire _13712_;
  wire _13713_;
  wire _13714_;
  wire _13715_;
  wire _13716_;
  wire _13717_;
  wire _13718_;
  wire _13719_;
  wire _13720_;
  wire _13721_;
  wire _13722_;
  wire _13723_;
  wire _13724_;
  wire _13725_;
  wire _13726_;
  wire _13727_;
  wire _13728_;
  wire _13729_;
  wire _13730_;
  wire _13731_;
  wire _13732_;
  wire _13733_;
  wire _13734_;
  wire _13735_;
  wire _13736_;
  wire _13737_;
  wire _13738_;
  wire _13739_;
  wire _13740_;
  wire _13741_;
  wire _13742_;
  wire _13743_;
  wire _13744_;
  wire _13745_;
  wire _13746_;
  wire _13747_;
  wire _13748_;
  wire _13749_;
  wire _13750_;
  wire _13751_;
  wire _13752_;
  wire _13753_;
  wire _13754_;
  wire _13755_;
  wire _13756_;
  wire _13757_;
  wire _13758_;
  wire _13759_;
  wire _13760_;
  wire _13761_;
  wire _13762_;
  wire _13763_;
  wire _13764_;
  wire _13765_;
  wire _13766_;
  wire _13767_;
  wire _13768_;
  wire _13769_;
  wire _13770_;
  wire _13771_;
  wire _13772_;
  wire _13773_;
  wire _13774_;
  wire _13775_;
  wire _13776_;
  wire _13777_;
  wire _13778_;
  wire _13779_;
  wire _13780_;
  wire _13781_;
  wire _13782_;
  wire _13783_;
  wire _13784_;
  wire _13785_;
  wire _13786_;
  wire _13787_;
  wire _13788_;
  wire _13789_;
  wire _13790_;
  wire _13791_;
  wire _13792_;
  wire _13793_;
  wire _13794_;
  wire _13795_;
  wire _13796_;
  wire _13797_;
  wire _13798_;
  wire _13799_;
  wire _13800_;
  wire _13801_;
  wire _13802_;
  wire _13803_;
  wire _13804_;
  wire _13805_;
  wire _13806_;
  wire _13807_;
  wire _13808_;
  wire _13809_;
  wire _13810_;
  wire _13811_;
  wire _13812_;
  wire _13813_;
  wire _13814_;
  wire _13815_;
  wire _13816_;
  wire _13817_;
  wire _13818_;
  wire _13819_;
  wire _13820_;
  wire _13821_;
  wire _13822_;
  wire _13823_;
  wire _13824_;
  wire _13825_;
  wire _13826_;
  wire _13827_;
  wire _13828_;
  wire _13829_;
  wire _13830_;
  wire _13831_;
  wire _13832_;
  wire _13833_;
  wire _13834_;
  wire _13835_;
  wire _13836_;
  wire _13837_;
  wire _13838_;
  wire _13839_;
  wire _13840_;
  wire _13841_;
  wire _13842_;
  wire _13843_;
  wire _13844_;
  wire _13845_;
  wire _13846_;
  wire _13847_;
  wire _13848_;
  wire _13849_;
  wire _13850_;
  wire _13851_;
  wire _13852_;
  wire _13853_;
  wire _13854_;
  wire _13855_;
  wire _13856_;
  wire _13857_;
  wire _13858_;
  wire _13859_;
  wire _13860_;
  wire _13861_;
  wire _13862_;
  wire _13863_;
  wire _13864_;
  wire _13865_;
  wire _13866_;
  wire _13867_;
  wire _13868_;
  wire _13869_;
  wire _13870_;
  wire _13871_;
  wire _13872_;
  wire _13873_;
  wire _13874_;
  wire _13875_;
  wire _13876_;
  wire _13877_;
  wire _13878_;
  wire _13879_;
  wire _13880_;
  wire _13881_;
  wire _13882_;
  wire _13883_;
  wire _13884_;
  wire _13885_;
  wire _13886_;
  wire _13887_;
  wire _13888_;
  wire _13889_;
  wire _13890_;
  wire _13891_;
  wire _13892_;
  wire _13893_;
  wire _13894_;
  wire _13895_;
  wire _13896_;
  wire _13897_;
  wire _13898_;
  wire _13899_;
  wire _13900_;
  wire _13901_;
  wire _13902_;
  wire _13903_;
  wire _13904_;
  wire _13905_;
  input [8:0] ABINPUT;
  input clk;
  wire [31:0] cxrom_data_out;
  wire cy;
  wire cy_reg;
  wire first_instr;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein0 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein1 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein2 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein3 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout0 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout1 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout2 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout3 ;
  wire \oc8051_symbolic_cxrom1.clk ;
  wire [31:0] \oc8051_symbolic_cxrom1.cxrom_data_out ;
  wire [15:0] \oc8051_symbolic_cxrom1.pc1 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc10 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc12 ;
  wire [15:0] \oc8051_symbolic_cxrom1.pc2 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc20 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc22 ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[0] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[10] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[11] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[12] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[13] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[14] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[15] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[1] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[2] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[3] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[4] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[5] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[6] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[7] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[8] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[9] ;
  wire [15:0] \oc8051_symbolic_cxrom1.regvalid ;
  wire \oc8051_symbolic_cxrom1.rst ;
  wire [31:0] \oc8051_symbolic_cxrom1.word_in ;
  wire [8:0] \oc8051_top_1.ABINPUT ;
  wire [7:0] \oc8051_top_1.acc ;
  wire \oc8051_top_1.bit_data ;
  wire [31:0] \oc8051_top_1.cxrom_data_out ;
  wire \oc8051_top_1.cy ;
  wire [1:0] \oc8051_top_1.cy_sel ;
  wire \oc8051_top_1.decoder_new_valid_pc ;
  wire [7:0] \oc8051_top_1.dptr_hi ;
  wire [7:0] \oc8051_top_1.dptr_lo ;
  wire [31:0] \oc8051_top_1.idat_onchip ;
  wire \oc8051_top_1.int_ack ;
  wire [7:0] \oc8051_top_1.int_src ;
  wire \oc8051_top_1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.mem_act ;
  wire \oc8051_top_1.oc8051_alu1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.divsrc2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.des2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div0 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.div_out ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.rst ;
  wire [5:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.rst ;
  wire [15:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul ;
  wire \oc8051_top_1.oc8051_alu1.rst ;
  wire \oc8051_top_1.oc8051_alu1.srcAc ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.acc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.clk ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.dptr ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op1_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op2_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op3_r ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.pc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_alu_src_sel1.sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_alu_src_sel1.sel2 ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.sel3 ;
  wire [7:0] \oc8051_top_1.oc8051_comp1.acc ;
  wire \oc8051_top_1.oc8051_comp1.cy ;
  wire \oc8051_top_1.oc8051_cy_select1.cy_in ;
  wire [1:0] \oc8051_top_1.oc8051_cy_select1.cy_sel ;
  wire [3:0] \oc8051_top_1.oc8051_decoder1.alu_op ;
  wire \oc8051_top_1.oc8051_decoder1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.cy_sel ;
  wire \oc8051_top_1.oc8051_decoder1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.mem_act ;
  wire \oc8051_top_1.oc8051_decoder1.new_valid_pc ;
  wire [7:0] \oc8051_top_1.oc8051_decoder1.op ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.psw_set ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_wr_sel ;
  wire \oc8051_top_1.oc8051_decoder1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.src_sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.src_sel2 ;
  wire \oc8051_top_1.oc8051_decoder1.src_sel3 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.state ;
  wire \oc8051_top_1.oc8051_decoder1.wait_data ;
  wire \oc8051_top_1.oc8051_decoder1.wr ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.wr_sfr ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[7] ;
  wire \oc8051_top_1.oc8051_indi_addr1.clk ;
  wire \oc8051_top_1.oc8051_indi_addr1.rst ;
  wire \oc8051_top_1.oc8051_indi_addr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.acc ;
  wire \oc8051_top_1.oc8051_memory_interface1.bit_in ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.cdata ;
  wire \oc8051_top_1.oc8051_memory_interface1.cdone ;
  wire \oc8051_top_1.oc8051_memory_interface1.clk ;
  wire \oc8051_top_1.oc8051_memory_interface1.decoder_new_valid_pc ;
  wire \oc8051_top_1.oc8051_memory_interface1.dmem_wait ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dptr ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.iadr_t ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_cur ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_old ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_onchip ;
  wire \oc8051_top_1.oc8051_memory_interface1.imem_wait ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm2_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.in_ram ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_t ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_v ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_vec_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.istb_t ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op2_buff ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op3_buff ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.op_pos ;
  wire \oc8051_top_1.oc8051_memory_interface1.out_of_rst ;
  wire [3:0] \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_buf ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_for_ajmp ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log_prev ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_out ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_addr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_ind ;
  wire \oc8051_top_1.oc8051_memory_interface1.reti ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ri_r ;
  wire [4:0] \oc8051_top_1.oc8051_memory_interface1.rn_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.sfr ;
  wire \oc8051_top_1.oc8051_memory_interface1.sfr_bit ;
  wire \oc8051_top_1.oc8051_rom1.clk ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.cxrom_data_out ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.data_o ;
  wire \oc8051_top_1.oc8051_rom1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.b_reg ;
  wire \oc8051_top_1.oc8051_sfr1.bit_out ;
  wire \oc8051_top_1.oc8051_sfr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.cy ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_lo ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.int_ack ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ip ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ack ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.t2_int ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.uart_int ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.p ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.set ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd ;
  wire [11:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp ;
  wire [10:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.pres_ow ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.prescaler ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.psw_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.rxd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.srcAc ;
  wire \oc8051_top_1.oc8051_sfr1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.t2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.tc2_int ;
  wire \oc8051_top_1.oc8051_sfr1.tclk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.tf0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.uart_int ;
  wire \oc8051_top_1.oc8051_sfr1.wait_data ;
  wire \oc8051_top_1.oc8051_sfr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.p0_i ;
  wire [7:0] \oc8051_top_1.p0_o ;
  wire [7:0] \oc8051_top_1.p1_i ;
  wire [7:0] \oc8051_top_1.p1_o ;
  wire [7:0] \oc8051_top_1.p2_i ;
  wire [7:0] \oc8051_top_1.p2_o ;
  wire [7:0] \oc8051_top_1.p3_i ;
  wire [7:0] \oc8051_top_1.p3_o ;
  wire [15:0] \oc8051_top_1.pc ;
  wire [15:0] \oc8051_top_1.pc_log ;
  wire \oc8051_top_1.pc_log_change ;
  wire [15:0] \oc8051_top_1.pc_log_prev ;
  wire [1:0] \oc8051_top_1.psw_set ;
  wire [7:0] \oc8051_top_1.ram_data ;
  wire \oc8051_top_1.rd_ind ;
  wire \oc8051_top_1.reti ;
  wire \oc8051_top_1.rxd_i ;
  wire \oc8051_top_1.sfr_bit ;
  wire [7:0] \oc8051_top_1.sfr_out ;
  wire \oc8051_top_1.srcAc ;
  wire [2:0] \oc8051_top_1.src_sel1 ;
  wire [1:0] \oc8051_top_1.src_sel2 ;
  wire \oc8051_top_1.src_sel3 ;
  wire \oc8051_top_1.t0_i ;
  wire \oc8051_top_1.t1_i ;
  wire \oc8051_top_1.t2_i ;
  wire \oc8051_top_1.t2ex_i ;
  wire \oc8051_top_1.wait_data ;
  wire \oc8051_top_1.wb_clk_i ;
  wire \oc8051_top_1.wb_rst_i ;
  input [7:0] p0_in;
  wire [7:0] p0_out;
  input [7:0] p1_in;
  wire [7:0] p1_out;
  input [7:0] p2_in;
  wire [7:0] p2_out;
  input [7:0] p3_in;
  wire [7:0] p3_out;
  wire [15:0] pc1;
  wire [15:0] pc1_plus_2;
  wire [15:0] pc2;
  wire pc_log_change;
  wire pc_log_change_r;
  output property_invalid_jc;
  input rst;
  input rxd_i;
  input t0_i;
  input t1_i;
  input t2_i;
  input t2ex_i;
  input [31:0] word_in;
  not _13906_ (_05542_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nand _13907_ (_05543_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _13908_ (_05544_, _05543_, _05542_);
  not _13909_ (_05545_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _13910_ (_05546_, \oc8051_top_1.oc8051_decoder1.state [1], \oc8051_top_1.oc8051_decoder1.state [0]);
  and _13911_ (_05547_, _05546_, _05545_);
  not _13912_ (_05548_, _05547_);
  nor _13913_ (_05549_, _05548_, _05544_);
  nor _13914_ (_05550_, _05549_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _13915_ (_05551_, _05550_, \oc8051_top_1.oc8051_rom1.data_o [17]);
  not _13916_ (_05552_, rst);
  not _13917_ (_05553_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  nand _13918_ (_05554_, _05550_, _05553_);
  and _13919_ (_05555_, _05554_, _05552_);
  and _13920_ (_00395_, _05555_, _05551_);
  not _13921_ (_05556_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and _13922_ (_05557_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _05556_);
  and _13923_ (_05558_, _05557_, _05552_);
  not _13924_ (_05559_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  nor _13925_ (_05560_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  nor _13926_ (_05561_, _05560_, _05559_);
  and _13927_ (_05562_, _05561_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re );
  not _13928_ (_05563_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  nor _13929_ (_05564_, _05563_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  not _13930_ (_05565_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  nor _13931_ (_05566_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], _05565_);
  and _13932_ (_05567_, _05566_, _05564_);
  and _13933_ (_05568_, _05567_, _05562_);
  and _13934_ (_05569_, _05559_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  not _13935_ (_05570_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  and _13936_ (_05571_, _05560_, _05570_);
  and _13937_ (_05572_, _05571_, _05569_);
  not _13938_ (_05573_, _05560_);
  and _13939_ (_05574_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and _13940_ (_05575_, _05574_, _05573_);
  nor _13941_ (_05576_, _05575_, _05572_);
  nor _13942_ (_05577_, _05576_, _05562_);
  or _13943_ (_05579_, _05577_, _05568_);
  and _13944_ (_05580_, _05560_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  and _13945_ (_05582_, _05580_, \oc8051_top_1.oc8051_sfr1.pres_ow );
  or _13946_ (_05583_, _05582_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  or _13947_ (_05584_, _05583_, _05579_);
  and _13948_ (_05585_, _05552_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor _13949_ (_05586_, _05582_, _05568_);
  or _13950_ (_05587_, _05586_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  and _13951_ (_05588_, _05587_, _05585_);
  and _13952_ (_05589_, _05588_, _05584_);
  or _13953_ (_01099_, _05589_, _05558_);
  nor _13954_ (_05590_, rst, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and _13955_ (_05591_, _05590_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  or _13956_ (_05592_, _05575_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  not _13957_ (_05593_, _05562_);
  nor _13958_ (_05594_, _05567_, _05593_);
  and _13959_ (_05595_, _05594_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  nor _13960_ (_05596_, _05562_, _05572_);
  or _13961_ (_05597_, _05596_, _05595_);
  and _13962_ (_05598_, _05597_, _05592_);
  not _13963_ (_05599_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  nor _13964_ (_05600_, _05586_, _05599_);
  or _13965_ (_05601_, _05600_, _05598_);
  nand _13966_ (_05602_, _05582_, _05599_);
  and _13967_ (_05603_, _05602_, _05585_);
  and _13968_ (_05604_, _05603_, _05601_);
  or _13969_ (_03276_, _05604_, _05591_);
  not _13970_ (_05605_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  nor _13971_ (_05606_, \oc8051_top_1.oc8051_memory_interface1.imem_wait , \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and _13972_ (_05607_, _05606_, _05605_);
  and _13973_ (_05608_, _05607_, _05547_);
  not _13974_ (_05609_, _05608_);
  not _13975_ (_05611_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  or _13976_ (_05612_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  or _13977_ (_05613_, _05612_, _05542_);
  or _13978_ (_05614_, _05613_, _05611_);
  not _13979_ (_05615_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  or _13980_ (_05616_, _05543_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  or _13981_ (_05617_, _05616_, _05615_);
  and _13982_ (_05618_, _05617_, _05614_);
  and _13983_ (_05619_, _05612_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nand _13984_ (_05620_, _05619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nand _13985_ (_05621_, _05620_, _05618_);
  not _13986_ (_05622_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and _13987_ (_05623_, _05622_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nand _13988_ (_05624_, _05623_, _05542_);
  not _13989_ (_05625_, _05624_);
  nand _13990_ (_05626_, _05625_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor _13991_ (_05627_, _05612_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nand _13992_ (_05628_, _05627_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  nand _13993_ (_05629_, _05628_, _05626_);
  nor _13994_ (_05630_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nand _13995_ (_05631_, _05630_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  not _13996_ (_05632_, _05631_);
  and _13997_ (_05633_, _05632_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  or _13998_ (_05634_, _05633_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  or _13999_ (_05635_, _05634_, _05629_);
  or _14000_ (_05636_, _05635_, _05621_);
  or _14001_ (_05637_, _05636_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  not _14002_ (_05638_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor _14003_ (_05639_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], _05638_);
  not _14004_ (_05640_, _05639_);
  and _14005_ (_05641_, _05640_, _05637_);
  or _14006_ (_05642_, _05641_, _05609_);
  not _14007_ (_05643_, _05607_);
  nor _14008_ (_05644_, _05547_, \oc8051_top_1.oc8051_decoder1.op [1]);
  nor _14009_ (_05645_, _05644_, _05643_);
  nand _14010_ (_05646_, _05645_, _05642_);
  nand _14011_ (_05647_, _05619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nand _14012_ (_05648_, _05625_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  and _14013_ (_05649_, _05648_, _05647_);
  not _14014_ (_05650_, _05616_);
  nand _14015_ (_05651_, _05650_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  not _14016_ (_05652_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  or _14017_ (_05653_, _05631_, _05652_);
  and _14018_ (_05654_, _05653_, _05651_);
  nand _14019_ (_05655_, _05627_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  not _14020_ (_05656_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  or _14021_ (_05657_, _05613_, _05656_);
  and _14022_ (_05658_, _05657_, _05655_);
  and _14023_ (_05659_, _05658_, _05654_);
  and _14024_ (_05660_, _05659_, _05649_);
  or _14025_ (_05661_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  or _14026_ (_05662_, _05661_, _05660_);
  and _14027_ (_05663_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], \oc8051_top_1.oc8051_memory_interface1.cdone );
  not _14028_ (_05664_, _05663_);
  and _14029_ (_05665_, _05664_, _05662_);
  nand _14030_ (_05666_, _05665_, _05608_);
  nor _14031_ (_05667_, _05547_, \oc8051_top_1.oc8051_decoder1.op [0]);
  nor _14032_ (_05668_, _05667_, _05643_);
  and _14033_ (_05669_, _05668_, _05666_);
  and _14034_ (_05670_, _05669_, _05646_);
  not _14035_ (_05671_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nand _14036_ (_05673_, _05632_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nand _14037_ (_05674_, _05625_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  and _14038_ (_05675_, _05674_, _05673_);
  nand _14039_ (_05676_, _05619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  not _14040_ (_05677_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  or _14041_ (_05678_, _05613_, _05677_);
  and _14042_ (_05679_, _05678_, _05676_);
  nand _14043_ (_05680_, _05627_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  nand _14044_ (_05681_, _05650_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  and _14045_ (_05682_, _05681_, _05680_);
  and _14046_ (_05683_, _05682_, _05679_);
  nand _14047_ (_05684_, _05683_, _05675_);
  nand _14048_ (_05685_, _05684_, _05671_);
  nand _14049_ (_05686_, _05685_, _05638_);
  nor _14050_ (_05687_, _05638_, \oc8051_top_1.oc8051_memory_interface1.cdata [2]);
  not _14051_ (_05688_, _05687_);
  and _14052_ (_05689_, _05688_, _05686_);
  or _14053_ (_05690_, _05689_, _05609_);
  nor _14054_ (_05691_, _05547_, \oc8051_top_1.oc8051_decoder1.op [2]);
  nor _14055_ (_05692_, _05691_, _05643_);
  and _14056_ (_05693_, _05692_, _05690_);
  nand _14057_ (_05694_, _05627_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  not _14058_ (_05695_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  or _14059_ (_05696_, _05631_, _05695_);
  and _14060_ (_05697_, _05696_, _05694_);
  nand _14061_ (_05698_, _05619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  not _14062_ (_05699_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  or _14063_ (_05700_, _05613_, _05699_);
  and _14064_ (_05701_, _05700_, _05698_);
  nand _14065_ (_05702_, _05650_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nand _14066_ (_05703_, _05625_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  and _14067_ (_05704_, _05703_, _05702_);
  and _14068_ (_05705_, _05704_, _05701_);
  and _14069_ (_05706_, _05705_, _05697_);
  or _14070_ (_05707_, _05706_, _05661_);
  and _14071_ (_05708_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], \oc8051_top_1.oc8051_memory_interface1.cdone );
  not _14072_ (_05709_, _05708_);
  nand _14073_ (_05710_, _05709_, _05707_);
  or _14074_ (_05711_, _05710_, _05609_);
  nor _14075_ (_05712_, _05547_, \oc8051_top_1.oc8051_decoder1.op [3]);
  nor _14076_ (_05713_, _05712_, _05643_);
  nand _14077_ (_05714_, _05713_, _05711_);
  and _14078_ (_05715_, _05714_, _05693_);
  and _14079_ (_05716_, _05715_, _05670_);
  and _14080_ (_05717_, _05627_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  and _14081_ (_05718_, _05650_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  and _14082_ (_05719_, _05632_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  or _14083_ (_05720_, _05719_, _05718_);
  or _14084_ (_05721_, _05720_, _05717_);
  and _14085_ (_05722_, _05625_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  or _14086_ (_05723_, _05722_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and _14087_ (_05724_, _05619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  not _14088_ (_05725_, _05613_);
  and _14089_ (_05726_, _05725_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  or _14090_ (_05727_, _05726_, _05724_);
  or _14091_ (_05728_, _05727_, _05723_);
  or _14092_ (_05729_, _05728_, _05721_);
  or _14093_ (_05730_, _05729_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor _14094_ (_05731_, _05638_, \oc8051_top_1.oc8051_memory_interface1.cdata [4]);
  not _14095_ (_05732_, _05731_);
  and _14096_ (_05733_, _05732_, _05730_);
  or _14097_ (_05734_, _05733_, _05609_);
  nor _14098_ (_05735_, _05547_, \oc8051_top_1.oc8051_decoder1.op [4]);
  nor _14099_ (_05736_, _05735_, _05643_);
  and _14100_ (_05737_, _05736_, _05734_);
  not _14101_ (_05738_, _05737_);
  nor _14102_ (_05739_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nand _14103_ (_05740_, _05619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  nand _14104_ (_05741_, _05625_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  and _14105_ (_05742_, _05741_, _05740_);
  not _14106_ (_05743_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  or _14107_ (_05744_, _05616_, _05743_);
  nand _14108_ (_05745_, _05632_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  and _14109_ (_05746_, _05745_, _05744_);
  nand _14110_ (_05747_, _05627_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  not _14111_ (_05748_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  or _14112_ (_05749_, _05613_, _05748_);
  and _14113_ (_05750_, _05749_, _05747_);
  and _14114_ (_05751_, _05750_, _05746_);
  nand _14115_ (_05752_, _05751_, _05742_);
  nand _14116_ (_05753_, _05752_, _05739_);
  and _14117_ (_05754_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.cdata [5]);
  not _14118_ (_05755_, _05754_);
  and _14119_ (_05756_, _05755_, _05753_);
  nand _14120_ (_05757_, _05756_, _05608_);
  nor _14121_ (_05758_, _05547_, \oc8051_top_1.oc8051_decoder1.op [5]);
  nor _14122_ (_05759_, _05758_, _05643_);
  and _14123_ (_05760_, _05759_, _05757_);
  not _14124_ (_05761_, _05760_);
  not _14125_ (_05762_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  or _14126_ (_05763_, _05613_, _05762_);
  not _14127_ (_05765_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  or _14128_ (_05766_, _05624_, _05765_);
  and _14129_ (_05767_, _05766_, _05763_);
  not _14130_ (_05768_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  or _14131_ (_05769_, _05616_, _05768_);
  not _14132_ (_05770_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  or _14133_ (_05771_, _05631_, _05770_);
  and _14134_ (_05772_, _05771_, _05769_);
  and _14135_ (_05773_, _05772_, _05767_);
  nand _14136_ (_05774_, _05619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nand _14137_ (_05775_, _05627_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  and _14138_ (_05776_, _05775_, _05774_);
  and _14139_ (_05777_, _05776_, _05773_);
  or _14140_ (_05778_, _05777_, _05661_);
  and _14141_ (_05779_, \oc8051_top_1.oc8051_memory_interface1.cdata [7], \oc8051_top_1.oc8051_memory_interface1.cdone );
  not _14142_ (_05780_, _05779_);
  nand _14143_ (_05781_, _05780_, _05778_);
  or _14144_ (_05782_, _05781_, _05609_);
  nor _14145_ (_05783_, _05547_, \oc8051_top_1.oc8051_decoder1.op [7]);
  nor _14146_ (_05784_, _05783_, _05643_);
  nand _14147_ (_05785_, _05784_, _05782_);
  not _14148_ (_05786_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  or _14149_ (_05787_, _05613_, _05786_);
  not _14150_ (_05788_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  or _14151_ (_05789_, _05624_, _05788_);
  and _14152_ (_05790_, _05789_, _05787_);
  not _14153_ (_05791_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  or _14154_ (_05792_, _05616_, _05791_);
  nand _14155_ (_05793_, _05632_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  and _14156_ (_05794_, _05793_, _05792_);
  and _14157_ (_05795_, _05794_, _05790_);
  nand _14158_ (_05796_, _05619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nand _14159_ (_05797_, _05627_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  and _14160_ (_05798_, _05797_, _05796_);
  and _14161_ (_05799_, _05798_, _05795_);
  or _14162_ (_05800_, _05799_, _05661_);
  and _14163_ (_05801_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], \oc8051_top_1.oc8051_memory_interface1.cdone );
  not _14164_ (_05802_, _05801_);
  nand _14165_ (_05803_, _05802_, _05800_);
  or _14166_ (_05804_, _05803_, _05609_);
  nor _14167_ (_05805_, _05547_, \oc8051_top_1.oc8051_decoder1.op [6]);
  nor _14168_ (_05806_, _05805_, _05643_);
  nand _14169_ (_05807_, _05806_, _05804_);
  and _14170_ (_05808_, _05807_, _05785_);
  and _14171_ (_05809_, _05808_, _05761_);
  and _14172_ (_05810_, _05809_, _05738_);
  and _14173_ (_05811_, _05810_, _05716_);
  and _14174_ (_05812_, _05784_, _05782_);
  nor _14175_ (_05813_, _05807_, _05760_);
  and _14176_ (_05814_, _05813_, _05812_);
  and _14177_ (_05815_, _05737_, _05716_);
  and _14178_ (_05816_, _05815_, _05814_);
  or _14179_ (_05817_, _05816_, _05811_);
  not _14180_ (_05818_, _05669_);
  not _14181_ (_05819_, _05646_);
  not _14182_ (_05820_, _05714_);
  nor _14183_ (_05821_, _05820_, _05693_);
  and _14184_ (_05822_, _05821_, _05819_);
  and _14185_ (_05823_, _05822_, _05818_);
  and _14186_ (_05824_, _05809_, _05737_);
  and _14187_ (_05825_, _05824_, _05823_);
  and _14188_ (_05826_, _05807_, _05812_);
  and _14189_ (_05827_, _05826_, _05760_);
  and _14190_ (_05828_, _05827_, _05737_);
  and _14191_ (_05829_, _05828_, _05823_);
  and _14192_ (_05830_, _05814_, _05738_);
  and _14193_ (_05831_, _05830_, _05823_);
  nor _14194_ (_05832_, _05831_, _05829_);
  not _14195_ (_05833_, _05832_);
  or _14196_ (_05834_, _05833_, _05825_);
  or _14197_ (_05835_, _05834_, _05817_);
  not _14198_ (_05836_, _05807_);
  and _14199_ (_05837_, _05836_, _05760_);
  and _14200_ (_05838_, _05837_, _05815_);
  and _14201_ (_05839_, _05826_, _05761_);
  and _14202_ (_05840_, _05839_, _05737_);
  and _14203_ (_05841_, _05840_, _05823_);
  and _14204_ (_05842_, _05815_, _05809_);
  or _14205_ (_05843_, _05842_, _05841_);
  or _14206_ (_05844_, _05843_, _05838_);
  and _14207_ (_05845_, _05830_, _05716_);
  and _14208_ (_05846_, _05814_, _05737_);
  and _14209_ (_05847_, _05846_, _05823_);
  or _14210_ (_05848_, _05847_, _05845_);
  and _14211_ (_05849_, _05818_, _05646_);
  and _14212_ (_05850_, _05849_, _05821_);
  and _14213_ (_05851_, _05850_, _05814_);
  nor _14214_ (_05852_, _05807_, _05812_);
  and _14215_ (_05853_, _05852_, _05760_);
  and _14216_ (_05854_, _05853_, _05738_);
  and _14217_ (_05855_, _05854_, _05822_);
  nor _14218_ (_05856_, _05855_, _05851_);
  and _14219_ (_05857_, _05839_, _05738_);
  and _14220_ (_05858_, _05857_, _05716_);
  and _14221_ (_05859_, _05852_, _05761_);
  and _14222_ (_05860_, _05859_, _05738_);
  and _14223_ (_05861_, _05860_, _05822_);
  nor _14224_ (_05862_, _05861_, _05858_);
  nand _14225_ (_05864_, _05862_, _05856_);
  or _14226_ (_05865_, _05864_, _05848_);
  or _14227_ (_05867_, _05865_, _05844_);
  or _14228_ (_05868_, _05867_, _05835_);
  and _14229_ (_05869_, _05821_, _05670_);
  and _14230_ (_05870_, _05869_, _05737_);
  and _14231_ (_05872_, _05857_, _05820_);
  or _14232_ (_05873_, _05872_, _05870_);
  nor _14233_ (_05874_, _05737_, _05646_);
  and _14234_ (_05875_, _05874_, _05715_);
  and _14235_ (_05876_, _05875_, _05839_);
  and _14236_ (_05877_, _05859_, _05737_);
  and _14237_ (_05878_, _05877_, _05822_);
  or _14238_ (_05879_, _05878_, _05876_);
  or _14239_ (_05880_, _05879_, _05873_);
  or _14240_ (_05881_, _05880_, _05868_);
  and _14241_ (_05882_, _05881_, _05547_);
  and _14242_ (_05883_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  not _14243_ (_05884_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and _14244_ (_05885_, \oc8051_top_1.oc8051_decoder1.state [1], _05545_);
  and _14245_ (_05886_, _05885_, _05884_);
  and _14246_ (_05887_, _05850_, _05824_);
  and _14247_ (_05888_, _05887_, _05886_);
  or _14248_ (_05889_, _05870_, _05825_);
  and _14249_ (_05890_, _05889_, _05886_);
  not _14250_ (_05891_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and _14251_ (_05892_, \oc8051_top_1.oc8051_decoder1.state [0], _05545_);
  and _14252_ (_05893_, _05892_, _05891_);
  and _14253_ (_05894_, _05849_, _05715_);
  and _14254_ (_05895_, _05827_, _05738_);
  and _14255_ (_05896_, _05895_, _05894_);
  and _14256_ (_05897_, _05894_, _05857_);
  nor _14257_ (_05898_, _05897_, _05896_);
  not _14258_ (_05900_, _05898_);
  and _14259_ (_05901_, _05900_, _05893_);
  or _14260_ (_05902_, _05901_, _05890_);
  or _14261_ (_05903_, _05902_, _05888_);
  or _14262_ (_05904_, _05903_, _05883_);
  or _14263_ (_05905_, _05904_, _05882_);
  and _14264_ (_04490_, _05905_, _05552_);
  or _14265_ (_05906_, _05550_, \oc8051_top_1.oc8051_rom1.data_o [22]);
  not _14266_ (_05907_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  nand _14267_ (_05908_, _05550_, _05907_);
  and _14268_ (_05909_, _05908_, _05552_);
  and _14269_ (_05764_, _05909_, _05906_);
  not _14270_ (_05910_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  nor _14271_ (_05911_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  nor _14272_ (_05912_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and _14273_ (_05913_, _05912_, _05911_);
  or _14274_ (_05914_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  nor _14275_ (_05915_, _05914_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  and _14276_ (_05916_, _05915_, _05913_);
  and _14277_ (_05917_, _05916_, _05910_);
  and _14278_ (_05918_, _05917_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  or _14279_ (_05919_, _05918_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and _14280_ (_07307_, _05919_, _05552_);
  or _14281_ (_05920_, _05550_, \oc8051_top_1.oc8051_rom1.data_o [27]);
  not _14282_ (_05921_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  nand _14283_ (_05922_, _05550_, _05921_);
  and _14284_ (_05923_, _05922_, _05552_);
  and _14285_ (_08287_, _05923_, _05920_);
  and _14286_ (_05924_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  and _14287_ (_05925_, _05924_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  and _14288_ (_05926_, _05925_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  and _14289_ (_05927_, _05926_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  and _14290_ (_05928_, _05927_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  and _14291_ (_05930_, _05928_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  not _14292_ (_05931_, _05930_);
  not _14293_ (_05933_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and _14294_ (_05934_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _05545_);
  and _14295_ (_05935_, _05934_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  and _14296_ (_05936_, _05935_, _05933_);
  not _14297_ (_05937_, _05936_);
  nor _14298_ (_05938_, _05928_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor _14299_ (_05939_, _05938_, _05937_);
  and _14300_ (_05940_, _05939_, _05931_);
  not _14301_ (_05941_, _05940_);
  not _14302_ (_05942_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  and _14303_ (_05943_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _05545_);
  and _14304_ (_05944_, _05943_, _05942_);
  and _14305_ (_05945_, _05944_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and _14306_ (_05946_, _05945_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [6]);
  not _14307_ (_05947_, _05946_);
  and _14308_ (_05948_, _05944_, _05933_);
  and _14309_ (_05949_, _05948_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [6]);
  not _14310_ (_05950_, _05949_);
  nor _14311_ (_05951_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  and _14312_ (_05952_, _05951_, _05934_);
  and _14313_ (_05953_, _05952_, \oc8051_top_1.oc8051_memory_interface1.ri_r [6]);
  and _14314_ (_05954_, _05935_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  nor _14315_ (_05955_, _05954_, _05953_);
  and _14316_ (_05956_, _05955_, _05950_);
  and _14317_ (_05957_, _05956_, _05947_);
  and _14318_ (_05958_, _05957_, _05941_);
  not _14319_ (_05959_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  nor _14320_ (_05960_, _05930_, _05959_);
  and _14321_ (_05961_, _05930_, _05959_);
  nor _14322_ (_05962_, _05961_, _05960_);
  nor _14323_ (_05963_, _05962_, _05937_);
  not _14324_ (_05964_, _05963_);
  and _14325_ (_05965_, _05952_, \oc8051_top_1.oc8051_memory_interface1.ri_r [7]);
  and _14326_ (_05966_, _05945_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [7]);
  and _14327_ (_05967_, _05948_, \oc8051_top_1.oc8051_memory_interface1.imm_r [7]);
  or _14328_ (_05968_, _05967_, _05966_);
  or _14329_ (_05969_, _05968_, _05954_);
  nor _14330_ (_05970_, _05969_, _05965_);
  and _14331_ (_05971_, _05970_, _05964_);
  and _14332_ (_05972_, _05971_, _05958_);
  not _14333_ (_05973_, _05927_);
  nor _14334_ (_05974_, _05926_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  nor _14335_ (_05975_, _05974_, _05937_);
  and _14336_ (_05976_, _05975_, _05973_);
  not _14337_ (_05977_, _05976_);
  and _14338_ (_05978_, _05948_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [4]);
  not _14339_ (_05979_, _05978_);
  and _14340_ (_05980_, _05952_, \oc8051_top_1.oc8051_memory_interface1.ri_r [4]);
  nor _14341_ (_05981_, _05980_, _05954_);
  and _14342_ (_05982_, _05981_, _05979_);
  and _14343_ (_05983_, _05945_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [4]);
  and _14344_ (_05984_, _05951_, _05942_);
  or _14345_ (_05985_, _05984_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and _14346_ (_05986_, _05985_, \oc8051_top_1.oc8051_memory_interface1.rn_r [4]);
  nor _14347_ (_05987_, _05986_, _05983_);
  and _14348_ (_05988_, _05987_, _05982_);
  and _14349_ (_05989_, _05988_, _05977_);
  not _14350_ (_05990_, _05928_);
  nor _14351_ (_05991_, _05927_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor _14352_ (_05992_, _05991_, _05937_);
  and _14353_ (_05993_, _05992_, _05990_);
  not _14354_ (_05994_, _05993_);
  and _14355_ (_05995_, _05952_, \oc8051_top_1.oc8051_memory_interface1.ri_r [5]);
  and _14356_ (_05996_, _05945_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  and _14357_ (_05997_, _05948_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [5]);
  or _14358_ (_05998_, _05997_, _05996_);
  or _14359_ (_05999_, _05998_, _05954_);
  nor _14360_ (_06000_, _05999_, _05995_);
  and _14361_ (_06001_, _06000_, _05994_);
  and _14362_ (_06002_, _06001_, _05989_);
  and _14363_ (_06003_, _06002_, _05972_);
  and _14364_ (_06004_, _05945_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [3]);
  and _14365_ (_06006_, _05948_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [3]);
  nor _14366_ (_06008_, _06006_, _06004_);
  not _14367_ (_06009_, _05926_);
  nor _14368_ (_06010_, _05925_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor _14369_ (_06011_, _06010_, _05937_);
  and _14370_ (_06012_, _06011_, _06009_);
  and _14371_ (_06014_, _05952_, \oc8051_top_1.oc8051_memory_interface1.ri_r [3]);
  and _14372_ (_06015_, _05985_, \oc8051_top_1.oc8051_memory_interface1.rn_r [3]);
  nor _14373_ (_06016_, _06015_, _06014_);
  not _14374_ (_06018_, _06016_);
  nor _14375_ (_06019_, _06018_, _06012_);
  and _14376_ (_06020_, _06019_, _06008_);
  and _14377_ (_06021_, _05985_, \oc8051_top_1.oc8051_memory_interface1.rn_r [0]);
  and _14378_ (_06022_, _05952_, \oc8051_top_1.oc8051_memory_interface1.ri_r [0]);
  nor _14379_ (_06023_, _06022_, _06021_);
  and _14380_ (_06024_, _05945_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [0]);
  not _14381_ (_06025_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and _14382_ (_06026_, _05936_, _06025_);
  and _14383_ (_06027_, _05948_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [0]);
  or _14384_ (_06028_, _06027_, _06026_);
  nor _14385_ (_06029_, _06028_, _06024_);
  and _14386_ (_06030_, _06029_, _06023_);
  not _14387_ (_06031_, _06030_);
  nor _14388_ (_06032_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  nor _14389_ (_06033_, _06032_, _05924_);
  and _14390_ (_06034_, _06033_, _05936_);
  and _14391_ (_06035_, _05952_, \oc8051_top_1.oc8051_memory_interface1.ri_r [1]);
  nor _14392_ (_06037_, _06035_, _06034_);
  and _14393_ (_06038_, _05945_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [1]);
  and _14394_ (_06039_, _05948_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [1]);
  and _14395_ (_06040_, _05985_, \oc8051_top_1.oc8051_memory_interface1.rn_r [1]);
  or _14396_ (_06041_, _06040_, _06039_);
  nor _14397_ (_06042_, _06041_, _06038_);
  and _14398_ (_06043_, _06042_, _06037_);
  nor _14399_ (_06044_, _05924_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor _14400_ (_06045_, _06044_, _05925_);
  and _14401_ (_06046_, _06045_, _05936_);
  and _14402_ (_06047_, _05952_, \oc8051_top_1.oc8051_memory_interface1.ri_r [2]);
  nor _14403_ (_06048_, _06047_, _06046_);
  and _14404_ (_06049_, _05945_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [2]);
  and _14405_ (_06050_, _05948_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [2]);
  and _14406_ (_06051_, _05985_, \oc8051_top_1.oc8051_memory_interface1.rn_r [2]);
  or _14407_ (_06052_, _06051_, _06050_);
  nor _14408_ (_06053_, _06052_, _06049_);
  and _14409_ (_06054_, _06053_, _06048_);
  and _14410_ (_06055_, _06054_, _06043_);
  and _14411_ (_06056_, _06055_, _06031_);
  and _14412_ (_06057_, _06056_, _06020_);
  and _14413_ (_06058_, _06057_, _06003_);
  and _14414_ (_06059_, _06043_, _06030_);
  and _14415_ (_06060_, _06059_, _06054_);
  and _14416_ (_06061_, _06060_, _06020_);
  and _14417_ (_06062_, _06061_, _06003_);
  or _14418_ (_06063_, _06062_, _06058_);
  not _14419_ (_06064_, _06020_);
  and _14420_ (_06065_, _06060_, _06064_);
  not _14421_ (_06066_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and _14422_ (_06067_, \oc8051_top_1.oc8051_decoder1.wr , _05545_);
  and _14423_ (_06068_, _06067_, _06066_);
  and _14424_ (_06069_, _06055_, _06003_);
  nand _14425_ (_06070_, _06069_, _06068_);
  or _14426_ (_06071_, _06070_, _06065_);
  or _14427_ (_06072_, _06071_, _06063_);
  and _14428_ (_06073_, _06072_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  not _14429_ (_06074_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [5]);
  not _14430_ (_06075_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  or _14431_ (_06076_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], _06075_);
  or _14432_ (_06077_, _06076_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  or _14433_ (_06078_, _06077_, _06074_);
  not _14434_ (_06079_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  not _14435_ (_06080_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and _14436_ (_06081_, _06080_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  nand _14437_ (_06082_, _06081_, _06075_);
  or _14438_ (_06083_, _06082_, _06079_);
  and _14439_ (_06084_, _06083_, _06078_);
  not _14440_ (_06085_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  or _14441_ (_06086_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  or _14442_ (_06087_, _06086_, _06080_);
  or _14443_ (_06088_, _06087_, _06085_);
  or _14444_ (_06089_, _06076_, _06080_);
  not _14445_ (_06090_, _06089_);
  nand _14446_ (_06091_, _06090_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and _14447_ (_06092_, _06091_, _06088_);
  and _14448_ (_06093_, _06092_, _06084_);
  nor _14449_ (_06094_, _06086_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  not _14450_ (_06095_, _06094_);
  not _14451_ (_06096_, \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  and _14452_ (_06097_, _06096_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r );
  or _14453_ (_06098_, _06097_, ABINPUT[6]);
  nand _14454_ (_06099_, _06096_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r );
  or _14455_ (_06100_, _06099_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  nand _14456_ (_06101_, _06100_, _06098_);
  or _14457_ (_06102_, _06101_, _06095_);
  not _14458_ (_06103_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and _14459_ (_06104_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  nand _14460_ (_06105_, _06104_, _06080_);
  or _14461_ (_06106_, _06105_, _06103_);
  and _14462_ (_06107_, _06104_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  nand _14463_ (_06108_, _06107_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [5]);
  and _14464_ (_06109_, _06108_, _06106_);
  and _14465_ (_06110_, _06109_, _06102_);
  nand _14466_ (_06111_, _06110_, _06093_);
  and _14467_ (_06112_, \oc8051_top_1.oc8051_decoder1.alu_op [3], _05545_);
  and _14468_ (_06113_, \oc8051_top_1.oc8051_decoder1.alu_op [2], _05545_);
  nor _14469_ (_06114_, _06113_, _06112_);
  and _14470_ (_06115_, \oc8051_top_1.oc8051_decoder1.alu_op [0], _05545_);
  and _14471_ (_06116_, \oc8051_top_1.oc8051_decoder1.alu_op [1], _05545_);
  nor _14472_ (_06117_, _06116_, _06115_);
  and _14473_ (_06118_, _06117_, _06114_);
  not _14474_ (_06119_, _06118_);
  and _14475_ (_06120_, _06115_, _06114_);
  not _14476_ (_06121_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  not _14477_ (_06122_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and _14478_ (_06123_, _06113_, _06122_);
  and _14479_ (_06124_, _06123_, _06121_);
  nor _14480_ (_06125_, _06124_, _06120_);
  and _14481_ (_06126_, _06125_, _06119_);
  and _14482_ (_06127_, _06112_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and _14483_ (_06128_, _06127_, _06121_);
  not _14484_ (_06129_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and _14485_ (_06130_, _06112_, _06129_);
  and _14486_ (_06131_, _06130_, _06116_);
  nor _14487_ (_06132_, _06131_, _06128_);
  and _14488_ (_06133_, _06132_, _06126_);
  not _14489_ (_06134_, _06133_);
  and _14490_ (_06135_, _06134_, _06111_);
  and _14491_ (_06136_, \oc8051_top_1.oc8051_decoder1.cy_sel [0], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor _14492_ (_06137_, _06136_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  nor _14493_ (_06138_, _06097_, ABINPUT[0]);
  nor _14494_ (_06139_, _06099_, \oc8051_top_1.oc8051_sfr1.bit_out );
  nor _14495_ (_06140_, _06139_, _06138_);
  nor _14496_ (_06141_, _06140_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  nor _14497_ (_06142_, _06141_, _06137_);
  not _14498_ (_06143_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [4]);
  or _14499_ (_06144_, _06077_, _06143_);
  not _14500_ (_06145_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [4]);
  or _14501_ (_06146_, _06082_, _06145_);
  and _14502_ (_06147_, _06146_, _06144_);
  not _14503_ (_06148_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  or _14504_ (_06149_, _06087_, _06148_);
  nand _14505_ (_06150_, _06090_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _14506_ (_06151_, _06150_, _06149_);
  and _14507_ (_06152_, _06151_, _06147_);
  or _14508_ (_06153_, _06097_, ABINPUT[5]);
  or _14509_ (_06154_, _06099_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  nand _14510_ (_06155_, _06154_, _06153_);
  or _14511_ (_06156_, _06155_, _06095_);
  not _14512_ (_06157_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or _14513_ (_06158_, _06105_, _06157_);
  nand _14514_ (_06159_, _06107_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [4]);
  and _14515_ (_06160_, _06159_, _06158_);
  and _14516_ (_06161_, _06160_, _06156_);
  nand _14517_ (_06162_, _06161_, _06152_);
  nor _14518_ (_06163_, _06162_, _06142_);
  not _14519_ (_06164_, _06162_);
  not _14520_ (_06165_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [3]);
  or _14521_ (_06166_, _06077_, _06165_);
  not _14522_ (_06167_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [3]);
  or _14523_ (_06168_, _06082_, _06167_);
  and _14524_ (_06169_, _06168_, _06166_);
  not _14525_ (_06170_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  or _14526_ (_06171_, _06087_, _06170_);
  nand _14527_ (_06172_, _06090_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and _14528_ (_06173_, _06172_, _06171_);
  and _14529_ (_06174_, _06173_, _06169_);
  or _14530_ (_06175_, _06097_, ABINPUT[4]);
  or _14531_ (_06176_, _06099_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  nand _14532_ (_06177_, _06176_, _06175_);
  or _14533_ (_06178_, _06177_, _06095_);
  not _14534_ (_06179_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or _14535_ (_06180_, _06105_, _06179_);
  nand _14536_ (_06181_, _06107_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [3]);
  and _14537_ (_06182_, _06181_, _06180_);
  and _14538_ (_06183_, _06182_, _06178_);
  nand _14539_ (_06184_, _06183_, _06174_);
  not _14540_ (_06185_, _06184_);
  not _14541_ (_06186_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [0]);
  nor _14542_ (_06187_, _06077_, _06186_);
  not _14543_ (_06188_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [0]);
  nor _14544_ (_06189_, _06082_, _06188_);
  nor _14545_ (_06190_, _06189_, _06187_);
  and _14546_ (_06191_, _06090_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  not _14547_ (_06192_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor _14548_ (_06193_, _06087_, _06192_);
  nor _14549_ (_06194_, _06193_, _06191_);
  and _14550_ (_06195_, _06194_, _06190_);
  or _14551_ (_06196_, _06097_, ABINPUT[1]);
  or _14552_ (_06197_, _06099_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  and _14553_ (_06198_, _06197_, _06196_);
  and _14554_ (_06199_, _06198_, _06094_);
  and _14555_ (_06200_, _06107_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [0]);
  not _14556_ (_06201_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor _14557_ (_06202_, _06105_, _06201_);
  nor _14558_ (_06203_, _06202_, _06200_);
  not _14559_ (_06204_, _06203_);
  nor _14560_ (_06205_, _06204_, _06199_);
  and _14561_ (_06206_, _06205_, _06195_);
  not _14562_ (_06207_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [2]);
  or _14563_ (_06208_, _06082_, _06207_);
  not _14564_ (_06209_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [2]);
  or _14565_ (_06210_, _06077_, _06209_);
  and _14566_ (_06211_, _06210_, _06208_);
  nand _14567_ (_06212_, _06107_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [2]);
  not _14568_ (_06213_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or _14569_ (_06214_, _06105_, _06213_);
  and _14570_ (_06215_, _06214_, _06212_);
  and _14571_ (_06216_, _06215_, _06211_);
  not _14572_ (_06217_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  or _14573_ (_06218_, _06089_, _06217_);
  not _14574_ (_06219_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  or _14575_ (_06220_, _06087_, _06219_);
  and _14576_ (_06221_, _06220_, _06218_);
  or _14577_ (_06222_, _06097_, ABINPUT[3]);
  or _14578_ (_06223_, _06099_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  nand _14579_ (_06224_, _06223_, _06222_);
  or _14580_ (_06225_, _06224_, _06095_);
  and _14581_ (_06226_, _06225_, _06221_);
  nand _14582_ (_06227_, _06226_, _06216_);
  not _14583_ (_06228_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [1]);
  or _14584_ (_06229_, _06077_, _06228_);
  not _14585_ (_06230_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [1]);
  or _14586_ (_06231_, _06082_, _06230_);
  and _14587_ (_06232_, _06231_, _06229_);
  not _14588_ (_06233_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  or _14589_ (_06234_, _06089_, _06233_);
  not _14590_ (_06235_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  or _14591_ (_06236_, _06087_, _06235_);
  and _14592_ (_06237_, _06236_, _06234_);
  and _14593_ (_06238_, _06237_, _06232_);
  or _14594_ (_06239_, _06097_, ABINPUT[2]);
  or _14595_ (_06240_, _06099_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  nand _14596_ (_06241_, _06240_, _06239_);
  or _14597_ (_06242_, _06241_, _06095_);
  not _14598_ (_06243_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or _14599_ (_06244_, _06105_, _06243_);
  nand _14600_ (_06245_, _06107_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [1]);
  and _14601_ (_06246_, _06245_, _06244_);
  and _14602_ (_06247_, _06246_, _06242_);
  nand _14603_ (_06248_, _06247_, _06238_);
  nor _14604_ (_06249_, _06248_, _06227_);
  and _14605_ (_06250_, _06249_, _06206_);
  and _14606_ (_06251_, _06250_, _06185_);
  and _14607_ (_06252_, _06251_, _06164_);
  not _14608_ (_06253_, _06142_);
  not _14609_ (_06254_, _06248_);
  nor _14610_ (_06255_, _06206_, _06254_);
  and _14611_ (_06256_, _06255_, _06227_);
  and _14612_ (_06257_, _06256_, _06184_);
  and _14613_ (_06258_, _06257_, _06253_);
  nor _14614_ (_06259_, _06258_, _06252_);
  nor _14615_ (_06260_, _06259_, _06163_);
  and _14616_ (_06261_, _06260_, _06111_);
  nor _14617_ (_06262_, _06260_, _06111_);
  not _14618_ (_06263_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and _14619_ (_06265_, _06116_, _06263_);
  and _14620_ (_06266_, _06127_, _06265_);
  not _14621_ (_06267_, _06266_);
  or _14622_ (_06268_, _06267_, _06262_);
  nor _14623_ (_06269_, _06268_, _06261_);
  nor _14624_ (_06270_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  not _14625_ (_06271_, _06270_);
  or _14626_ (_06272_, _06271_, _06101_);
  nand _14627_ (_06273_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  or _14628_ (_06274_, _06273_, _06074_);
  not _14629_ (_06275_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  nand _14630_ (_06276_, _06275_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  or _14631_ (_06277_, _06276_, _06103_);
  and _14632_ (_06278_, _06277_, _06274_);
  nand _14633_ (_06279_, _06278_, _06272_);
  nor _14634_ (_06280_, _06279_, _06111_);
  and _14635_ (_06281_, _06115_, _06121_);
  and _14636_ (_06282_, _06130_, _06281_);
  not _14637_ (_06283_, _06282_);
  nor _14638_ (_06284_, _06283_, _06280_);
  not _14639_ (_06285_, _06284_);
  and _14640_ (_06286_, _06279_, _06111_);
  and _14641_ (_06287_, _06116_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and _14642_ (_06288_, _06287_, _06123_);
  and _14643_ (_06289_, _06288_, _06286_);
  and _14644_ (_06290_, _06265_, _06123_);
  not _14645_ (_06291_, _06290_);
  nor _14646_ (_06292_, _06291_, _06111_);
  nor _14647_ (_06293_, _06292_, _06289_);
  nand _14648_ (_06294_, _06293_, _06285_);
  and _14649_ (_06295_, _06127_, _06287_);
  and _14650_ (_06296_, _06279_, _06142_);
  and _14651_ (_06297_, _06253_, _06111_);
  or _14652_ (_06298_, _06297_, _06296_);
  and _14653_ (_06299_, _06298_, _06295_);
  and _14654_ (_06300_, _06130_, _06117_);
  nor _14655_ (_06301_, _06286_, _06280_);
  and _14656_ (_06302_, _06301_, _06300_);
  or _14657_ (_06303_, _06302_, _06299_);
  or _14658_ (_06304_, _06303_, _06294_);
  or _14659_ (_06305_, _06304_, _06269_);
  nor _14660_ (_06306_, _06305_, _06135_);
  not _14661_ (_06307_, _06306_);
  and _14662_ (_06308_, _06056_, _06064_);
  and _14663_ (_06309_, _06308_, _06003_);
  and _14664_ (_06310_, _06309_, _06068_);
  and _14665_ (_06311_, _06310_, _06307_);
  or _14666_ (_06312_, _06311_, _06073_);
  and _14667_ (_10361_, _06312_, _05552_);
  not _14668_ (_06313_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and _14669_ (_06314_, _06123_, _06117_);
  and _14670_ (_06315_, _06314_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _14671_ (_06316_, _06315_, _06313_);
  and _14672_ (_06317_, _06315_, _06313_);
  or _14673_ (_06318_, _06317_, _06316_);
  and _14674_ (_10695_, _06318_, _05552_);
  not _14675_ (_06319_, _05586_);
  nor _14676_ (_06320_, _06319_, _05577_);
  nor _14677_ (_06321_, _06320_, _05556_);
  or _14678_ (_06322_, _06321_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  or _14679_ (_06323_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8], _05556_);
  or _14680_ (_06324_, _06323_, _05586_);
  and _14681_ (_06325_, _06324_, _05552_);
  and _14682_ (_11021_, _06325_, _06322_);
  nor _14683_ (_06326_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  nor _14684_ (_11823_, _06326_, rst);
  nor _14685_ (_06327_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  not _14686_ (_06328_, _06327_);
  and _14687_ (_06329_, _06328_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3]);
  not _14688_ (_06330_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  and _14689_ (_06331_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _06330_);
  not _14690_ (_06332_, _06331_);
  or _14691_ (_06333_, _06271_, _06177_);
  or _14692_ (_06334_, _06273_, _06165_);
  or _14693_ (_06335_, _06276_, _06179_);
  and _14694_ (_06336_, _06335_, _06334_);
  and _14695_ (_06337_, _06336_, _06333_);
  or _14696_ (_06339_, _06337_, _06332_);
  and _14697_ (_06340_, _06278_, _06272_);
  not _14698_ (_06341_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  and _14699_ (_06342_, _06341_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  not _14700_ (_06343_, _06342_);
  or _14701_ (_06344_, _06343_, _06340_);
  and _14702_ (_06345_, _06344_, _06339_);
  or _14703_ (_06346_, _06342_, _06331_);
  or _14704_ (_06347_, _06271_, _06241_);
  or _14705_ (_06348_, _06273_, _06228_);
  or _14706_ (_06349_, _06276_, _06243_);
  and _14707_ (_06350_, _06349_, _06348_);
  and _14708_ (_06351_, _06350_, _06347_);
  or _14709_ (_06352_, _06351_, _06346_);
  and _14710_ (_06353_, _06352_, _06328_);
  and _14711_ (_06354_, _06353_, _06345_);
  or _14712_ (_06355_, _06097_, ABINPUT[8]);
  or _14713_ (_06356_, _06099_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  nand _14714_ (_06357_, _06356_, _06355_);
  or _14715_ (_06358_, _06357_, _06271_);
  not _14716_ (_06359_, \oc8051_top_1.oc8051_memory_interface1.imm_r [7]);
  or _14717_ (_06360_, _06273_, _06359_);
  not _14718_ (_06361_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or _14719_ (_06362_, _06276_, _06361_);
  and _14720_ (_06363_, _06362_, _06360_);
  and _14721_ (_06364_, _06363_, _06358_);
  and _14722_ (_06365_, _06364_, _06327_);
  nor _14723_ (_06366_, _06365_, _06354_);
  and _14724_ (_06367_, _06366_, _06248_);
  not _14725_ (_06368_, _06206_);
  or _14726_ (_06369_, _06271_, _06224_);
  or _14727_ (_06370_, _06273_, _06209_);
  or _14728_ (_06371_, _06276_, _06213_);
  and _14729_ (_06372_, _06371_, _06370_);
  and _14730_ (_06373_, _06372_, _06369_);
  or _14731_ (_06374_, _06373_, _06332_);
  or _14732_ (_06375_, _06271_, _06155_);
  or _14733_ (_06376_, _06273_, _06143_);
  or _14734_ (_06377_, _06276_, _06157_);
  and _14735_ (_06378_, _06377_, _06376_);
  and _14736_ (_06379_, _06378_, _06375_);
  or _14737_ (_06380_, _06379_, _06343_);
  and _14738_ (_06381_, _06380_, _06374_);
  nand _14739_ (_06382_, _06270_, _06198_);
  or _14740_ (_06383_, _06273_, _06186_);
  or _14741_ (_06384_, _06276_, _06201_);
  and _14742_ (_06385_, _06384_, _06383_);
  and _14743_ (_06386_, _06385_, _06382_);
  or _14744_ (_06387_, _06386_, _06346_);
  and _14745_ (_06388_, _06387_, _06328_);
  nand _14746_ (_06389_, _06388_, _06381_);
  or _14747_ (_06390_, _06097_, ABINPUT[7]);
  or _14748_ (_06391_, _06099_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  nand _14749_ (_06392_, _06391_, _06390_);
  or _14750_ (_06393_, _06392_, _06271_);
  not _14751_ (_06394_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [6]);
  or _14752_ (_06395_, _06273_, _06394_);
  not _14753_ (_06396_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or _14754_ (_06397_, _06276_, _06396_);
  and _14755_ (_06398_, _06397_, _06395_);
  nand _14756_ (_06399_, _06398_, _06393_);
  or _14757_ (_06400_, _06399_, _06328_);
  and _14758_ (_06401_, _06400_, _06389_);
  and _14759_ (_06402_, _06401_, _06368_);
  and _14760_ (_06403_, _06402_, _06367_);
  and _14761_ (_06404_, _06401_, _06227_);
  nand _14762_ (_06405_, _06404_, _06367_);
  or _14763_ (_06406_, _06404_, _06367_);
  and _14764_ (_06407_, _06406_, _06405_);
  and _14765_ (_06408_, _06407_, _06403_);
  and _14766_ (_06409_, _06401_, _06184_);
  nand _14767_ (_06410_, _06400_, _06389_);
  or _14768_ (_06411_, _06410_, _06254_);
  and _14769_ (_06412_, _06366_, _06227_);
  and _14770_ (_06413_, _06412_, _06411_);
  nand _14771_ (_06414_, _06413_, _06409_);
  or _14772_ (_06415_, _06413_, _06409_);
  and _14773_ (_06416_, _06415_, _06414_);
  nand _14774_ (_06417_, _06416_, _06408_);
  not _14775_ (_06418_, _06417_);
  nand _14776_ (_06419_, _06414_, _06405_);
  or _14777_ (_06420_, _06365_, _06354_);
  or _14778_ (_06421_, _06420_, _06185_);
  or _14779_ (_06422_, _06410_, _06164_);
  or _14780_ (_06423_, _06422_, _06421_);
  nand _14781_ (_06424_, _06422_, _06421_);
  and _14782_ (_06425_, _06424_, _06423_);
  nand _14783_ (_06426_, _06425_, _06419_);
  or _14784_ (_06427_, _06425_, _06419_);
  and _14785_ (_06428_, _06427_, _06426_);
  and _14786_ (_06429_, _06428_, _06418_);
  and _14787_ (_06430_, _06425_, _06419_);
  and _14788_ (_06431_, _06366_, _06162_);
  and _14789_ (_06432_, _06431_, _06409_);
  not _14790_ (_06433_, _06111_);
  or _14791_ (_06434_, _06420_, _06433_);
  or _14792_ (_06435_, _06434_, _06422_);
  and _14793_ (_06436_, _06401_, _06111_);
  or _14794_ (_06437_, _06436_, _06431_);
  and _14795_ (_06438_, _06437_, _06435_);
  nand _14796_ (_06439_, _06438_, _06432_);
  or _14797_ (_06440_, _06438_, _06432_);
  and _14798_ (_06441_, _06440_, _06439_);
  nand _14799_ (_06442_, _06441_, _06430_);
  or _14800_ (_06443_, _06441_, _06430_);
  and _14801_ (_06444_, _06443_, _06442_);
  nand _14802_ (_06445_, _06444_, _06429_);
  or _14803_ (_06446_, _06444_, _06429_);
  and _14804_ (_06447_, _06446_, _06445_);
  and _14805_ (_06448_, _06447_, _06329_);
  nor _14806_ (_06449_, _06447_, _06329_);
  or _14807_ (_06450_, _06449_, _06448_);
  and _14808_ (_06451_, _06328_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1]);
  or _14809_ (_06452_, _06416_, _06408_);
  and _14810_ (_06453_, _06452_, _06417_);
  nand _14811_ (_06454_, _06453_, _06451_);
  and _14812_ (_06455_, _06328_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0]);
  not _14813_ (_06456_, _06455_);
  nor _14814_ (_06457_, _06407_, _06403_);
  or _14815_ (_06458_, _06457_, _06408_);
  or _14816_ (_06459_, _06458_, _06456_);
  or _14817_ (_06461_, _06453_, _06451_);
  nand _14818_ (_06462_, _06461_, _06454_);
  or _14819_ (_06463_, _06462_, _06459_);
  nand _14820_ (_06464_, _06463_, _06454_);
  and _14821_ (_06465_, _06328_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2]);
  nand _14822_ (_06466_, _06428_, _06418_);
  or _14823_ (_06467_, _06428_, _06418_);
  and _14824_ (_06469_, _06467_, _06466_);
  nand _14825_ (_06470_, _06469_, _06465_);
  or _14826_ (_06471_, _06469_, _06465_);
  and _14827_ (_06472_, _06471_, _06470_);
  nand _14828_ (_06473_, _06472_, _06464_);
  or _14829_ (_06474_, _06473_, _06450_);
  not _14830_ (_06475_, _06470_);
  nor _14831_ (_06476_, _06475_, _06448_);
  or _14832_ (_06477_, _06476_, _06449_);
  and _14833_ (_06478_, _06477_, _06474_);
  and _14834_ (_06479_, _06328_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4]);
  not _14835_ (_06480_, _06445_);
  not _14836_ (_06481_, _06434_);
  not _14837_ (_06482_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [6]);
  or _14838_ (_06483_, _06082_, _06482_);
  or _14839_ (_06485_, _06077_, _06394_);
  and _14840_ (_06486_, _06485_, _06483_);
  not _14841_ (_06487_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  or _14842_ (_06488_, _06087_, _06487_);
  not _14843_ (_06489_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  or _14844_ (_06490_, _06089_, _06489_);
  and _14845_ (_06491_, _06490_, _06488_);
  and _14846_ (_06492_, _06491_, _06486_);
  or _14847_ (_06493_, _06392_, _06095_);
  or _14848_ (_06494_, _06105_, _06396_);
  nand _14849_ (_06495_, _06107_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [6]);
  and _14850_ (_06496_, _06495_, _06494_);
  and _14851_ (_06497_, _06496_, _06493_);
  and _14852_ (_06498_, _06497_, _06492_);
  or _14853_ (_06499_, _06498_, _06435_);
  not _14854_ (_06500_, _06498_);
  and _14855_ (_06501_, _06500_, _06401_);
  not _14856_ (_06502_, _06501_);
  nand _14857_ (_06503_, _06502_, _06435_);
  and _14858_ (_06504_, _06503_, _06499_);
  nand _14859_ (_06505_, _06504_, _06481_);
  or _14860_ (_06506_, _06501_, _06481_);
  nand _14861_ (_06507_, _06506_, _06505_);
  and _14862_ (_06508_, _06442_, _06439_);
  nand _14863_ (_06509_, _06508_, _06507_);
  or _14864_ (_06510_, _06508_, _06507_);
  and _14865_ (_06511_, _06510_, _06509_);
  nand _14866_ (_06512_, _06511_, _06480_);
  or _14867_ (_06513_, _06511_, _06480_);
  and _14868_ (_06514_, _06513_, _06512_);
  nand _14869_ (_06515_, _06514_, _06479_);
  or _14870_ (_06516_, _06514_, _06479_);
  nand _14871_ (_06517_, _06516_, _06515_);
  or _14872_ (_06518_, _06517_, _06478_);
  not _14873_ (_06519_, _06518_);
  and _14874_ (_06520_, _06517_, _06478_);
  nor _14875_ (_06521_, _06520_, _06519_);
  and _14876_ (_12386_, _06521_, _05552_);
  and _14877_ (_06522_, _05934_, _05933_);
  not _14878_ (_06523_, _06522_);
  and _14879_ (_06524_, _06523_, _06068_);
  and _14880_ (_06525_, _06524_, _06020_);
  and _14881_ (_06526_, _06525_, _06060_);
  not _14882_ (_06527_, _05989_);
  and _14883_ (_06528_, _06001_, _06527_);
  nor _14884_ (_06529_, _05971_, _05958_);
  and _14885_ (_06530_, _06529_, _06528_);
  and _14886_ (_06531_, _06530_, _06526_);
  not _14887_ (_06532_, _06531_);
  and _14888_ (_06533_, _06532_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  nand _14889_ (_06534_, _06336_, _06333_);
  and _14890_ (_06535_, _06534_, _06295_);
  and _14891_ (_06536_, _06256_, _06253_);
  and _14892_ (_06537_, _06250_, _06142_);
  nor _14893_ (_06538_, _06537_, _06536_);
  nor _14894_ (_06539_, _06538_, _06185_);
  and _14895_ (_06540_, _06538_, _06185_);
  or _14896_ (_06541_, _06540_, _06267_);
  nor _14897_ (_06542_, _06541_, _06539_);
  nor _14898_ (_06543_, _06542_, _06535_);
  nor _14899_ (_06544_, _06534_, _06184_);
  nor _14900_ (_06545_, _06544_, _06283_);
  not _14901_ (_06546_, _06300_);
  and _14902_ (_06547_, _06534_, _06184_);
  or _14903_ (_06549_, _06547_, _06544_);
  nor _14904_ (_06550_, _06549_, _06546_);
  or _14905_ (_06551_, _06550_, _06545_);
  not _14906_ (_06552_, _06551_);
  and _14907_ (_06553_, _06547_, _06288_);
  nor _14908_ (_06554_, _06291_, _06184_);
  nor _14909_ (_06555_, _06554_, _06553_);
  and _14910_ (_06556_, _06184_, _06134_);
  not _14911_ (_06557_, _06556_);
  and _14912_ (_06558_, _06557_, _06555_);
  and _14913_ (_06559_, _06558_, _06552_);
  and _14914_ (_06560_, _06559_, _06543_);
  nor _14915_ (_06561_, _06560_, _06532_);
  nor _14916_ (_06562_, _06561_, _06533_);
  nor _14917_ (_13222_, _06562_, rst);
  or _14918_ (_06563_, _05550_, \oc8051_top_1.oc8051_rom1.data_o [26]);
  not _14919_ (_06564_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  nand _14920_ (_06565_, _05550_, _06564_);
  and _14921_ (_06566_, _06565_, _05552_);
  and _14922_ (_01193_, _06566_, _06563_);
  and _14923_ (_06567_, _05822_, _05669_);
  and _14924_ (_06568_, _06567_, _05839_);
  and _14925_ (_06569_, _05837_, _05812_);
  and _14926_ (_06570_, _06569_, _05738_);
  not _14927_ (_06571_, _06570_);
  nor _14928_ (_06572_, _05850_, _05822_);
  nor _14929_ (_06573_, _06572_, _06571_);
  nor _14930_ (_06574_, _06573_, _06568_);
  not _14931_ (_06575_, _06574_);
  and _14932_ (_06576_, _05547_, _05552_);
  nand _14933_ (_01436_, _06576_, _06575_);
  or _14934_ (_06577_, _06321_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  or _14935_ (_06578_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _05556_);
  or _14936_ (_06579_, _06578_, _05586_);
  and _14937_ (_06580_, _06579_, _05552_);
  and _14938_ (_01904_, _06580_, _06577_);
  and _14939_ (_06581_, _06265_, _06114_);
  not _14940_ (_06582_, _06581_);
  not _14941_ (_06583_, _06364_);
  not _14942_ (_06584_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [7]);
  or _14943_ (_06585_, _06082_, _06584_);
  or _14944_ (_06586_, _06077_, _06359_);
  and _14945_ (_06587_, _06586_, _06585_);
  not _14946_ (_06588_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  or _14947_ (_06589_, _06089_, _06588_);
  not _14948_ (_06590_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  or _14949_ (_06591_, _06087_, _06590_);
  and _14950_ (_06593_, _06591_, _06589_);
  and _14951_ (_06594_, _06593_, _06587_);
  or _14952_ (_06595_, _06357_, _06095_);
  or _14953_ (_06596_, _06105_, _06361_);
  nand _14954_ (_06597_, _06107_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [7]);
  and _14955_ (_06598_, _06597_, _06596_);
  and _14956_ (_06599_, _06598_, _06595_);
  and _14957_ (_06600_, _06599_, _06594_);
  and _14958_ (_06601_, _06600_, _06583_);
  and _14959_ (_06602_, _06600_, _06364_);
  nor _14960_ (_06603_, _06600_, _06364_);
  nor _14961_ (_06604_, _06603_, _06602_);
  nor _14962_ (_06605_, _06498_, _06399_);
  not _14963_ (_06606_, _06399_);
  nor _14964_ (_06608_, _06498_, _06606_);
  and _14965_ (_06609_, _06498_, _06606_);
  nor _14966_ (_06611_, _06609_, _06608_);
  and _14967_ (_06612_, _06340_, _06111_);
  nor _14968_ (_06613_, _06379_, _06162_);
  nor _14969_ (_06614_, _06613_, _06301_);
  nor _14970_ (_06615_, _06614_, _06612_);
  nor _14971_ (_06616_, _06615_, _06611_);
  nor _14972_ (_06617_, _06616_, _06605_);
  and _14973_ (_06618_, _06615_, _06611_);
  nor _14974_ (_06619_, _06618_, _06616_);
  not _14975_ (_06620_, _06619_);
  and _14976_ (_06621_, _06613_, _06301_);
  nor _14977_ (_06622_, _06621_, _06614_);
  not _14978_ (_06624_, _06622_);
  nand _14979_ (_06625_, _06378_, _06375_);
  and _14980_ (_06626_, _06625_, _06162_);
  nor _14981_ (_06627_, _06625_, _06162_);
  nor _14982_ (_06628_, _06627_, _06626_);
  not _14983_ (_06629_, _06628_);
  not _14984_ (_06630_, _06549_);
  nand _14985_ (_06631_, _06372_, _06369_);
  and _14986_ (_06632_, _06631_, _06227_);
  nor _14987_ (_06633_, _06631_, _06227_);
  nor _14988_ (_06634_, _06633_, _06632_);
  nand _14989_ (_06635_, _06350_, _06347_);
  and _14990_ (_06636_, _06635_, _06248_);
  nor _14991_ (_06637_, _06635_, _06248_);
  nor _14992_ (_06638_, _06637_, _06636_);
  nand _14993_ (_06639_, _06385_, _06382_);
  and _14994_ (_06640_, _06639_, _06206_);
  nor _14995_ (_06641_, _06640_, _06638_);
  and _14996_ (_06642_, _06351_, _06248_);
  nor _14997_ (_06643_, _06642_, _06641_);
  nor _14998_ (_06644_, _06643_, _06634_);
  and _14999_ (_06645_, _06373_, _06227_);
  nor _15000_ (_06646_, _06645_, _06644_);
  nor _15001_ (_06647_, _06646_, _06630_);
  and _15002_ (_06648_, _06646_, _06630_);
  nor _15003_ (_06649_, _06648_, _06647_);
  and _15004_ (_06650_, _06643_, _06634_);
  nor _15005_ (_06651_, _06650_, _06644_);
  not _15006_ (_06652_, _06651_);
  and _15007_ (_06653_, _06640_, _06638_);
  nor _15008_ (_06654_, _06653_, _06641_);
  not _15009_ (_06655_, _06654_);
  nor _15010_ (_06656_, _06386_, _06206_);
  and _15011_ (_06657_, _06386_, _06206_);
  nor _15012_ (_06658_, _06657_, _06656_);
  nor _15013_ (_06659_, _06658_, _06253_);
  and _15014_ (_06660_, _06659_, _06655_);
  and _15015_ (_06661_, _06660_, _06652_);
  not _15016_ (_06662_, _06661_);
  nor _15017_ (_06663_, _06662_, _06649_);
  nand _15018_ (_06664_, _06337_, _06184_);
  nor _15019_ (_06665_, _06337_, _06184_);
  or _15020_ (_06666_, _06646_, _06665_);
  and _15021_ (_06667_, _06666_, _06664_);
  or _15022_ (_06668_, _06667_, _06663_);
  and _15023_ (_06669_, _06668_, _06629_);
  and _15024_ (_06670_, _06669_, _06624_);
  and _15025_ (_06671_, _06670_, _06620_);
  nor _15026_ (_06672_, _06671_, _06617_);
  nor _15027_ (_06673_, _06672_, _06604_);
  nor _15028_ (_06674_, _06673_, _06601_);
  nor _15029_ (_06675_, _06674_, _06582_);
  not _15030_ (_06676_, _06675_);
  and _15031_ (_06677_, _06281_, _06114_);
  not _15032_ (_06678_, _06677_);
  not _15033_ (_06679_, _06603_);
  not _15034_ (_06680_, _06634_);
  and _15035_ (_06681_, _06656_, _06638_);
  nor _15036_ (_06682_, _06681_, _06636_);
  nor _15037_ (_06683_, _06682_, _06680_);
  nor _15038_ (_06684_, _06683_, _06632_);
  nor _15039_ (_06685_, _06684_, _06630_);
  and _15040_ (_06686_, _06684_, _06630_);
  nor _15041_ (_06687_, _06686_, _06685_);
  and _15042_ (_06688_, _06658_, _06142_);
  and _15043_ (_06689_, _06688_, _06638_);
  and _15044_ (_06690_, _06682_, _06680_);
  nor _15045_ (_06692_, _06690_, _06683_);
  and _15046_ (_06693_, _06692_, _06689_);
  not _15047_ (_06694_, _06693_);
  nor _15048_ (_06695_, _06694_, _06687_);
  nor _15049_ (_06696_, _06684_, _06544_);
  or _15050_ (_06697_, _06696_, _06547_);
  or _15051_ (_06698_, _06697_, _06695_);
  and _15052_ (_06699_, _06698_, _06628_);
  and _15053_ (_06700_, _06699_, _06301_);
  not _15054_ (_06701_, _06611_);
  and _15055_ (_06702_, _06626_, _06301_);
  nor _15056_ (_06703_, _06702_, _06286_);
  nor _15057_ (_06704_, _06703_, _06701_);
  and _15058_ (_06705_, _06703_, _06701_);
  nor _15059_ (_06706_, _06705_, _06704_);
  and _15060_ (_06707_, _06706_, _06700_);
  not _15061_ (_06708_, _06707_);
  nor _15062_ (_06709_, _06704_, _06608_);
  and _15063_ (_06710_, _06709_, _06708_);
  or _15064_ (_06711_, _06710_, _06602_);
  and _15065_ (_06712_, _06711_, _06679_);
  nor _15066_ (_06713_, _06712_, _06678_);
  nor _15067_ (_06714_, _06500_, _06111_);
  not _15068_ (_06715_, _06714_);
  and _15069_ (_06716_, _06281_, _06123_);
  nor _15070_ (_06717_, _06249_, _06185_);
  and _15071_ (_06718_, _06717_, _06716_);
  and _15072_ (_06719_, _06718_, _06162_);
  nor _15073_ (_06720_, _06719_, _06715_);
  nor _15074_ (_06721_, _06720_, _06600_);
  nor _15075_ (_06722_, _06721_, _06142_);
  not _15076_ (_06723_, _06722_);
  not _15077_ (_06724_, _06716_);
  nor _15078_ (_06725_, _06600_, _06253_);
  not _15079_ (_06726_, _06725_);
  nor _15080_ (_06727_, _06726_, _06720_);
  nor _15081_ (_06728_, _06727_, _06724_);
  and _15082_ (_06729_, _06728_, _06723_);
  not _15083_ (_06730_, _06718_);
  and _15084_ (_06731_, _06140_, _06137_);
  and _15085_ (_06732_, _06130_, _06265_);
  and _15086_ (_06733_, _06288_, _06140_);
  nor _15087_ (_06734_, _06733_, _06732_);
  nor _15088_ (_06735_, _06734_, _06731_);
  and _15089_ (_06736_, _06127_, _06281_);
  and _15090_ (_06737_, _06368_, _06736_);
  nor _15091_ (_06738_, _06737_, _06735_);
  nor _15092_ (_06739_, _06142_, _06140_);
  not _15093_ (_06740_, _06140_);
  nor _15094_ (_06741_, _06740_, _06137_);
  nor _15095_ (_06742_, _06741_, _06546_);
  nor _15096_ (_06743_, _06742_, _06282_);
  nor _15097_ (_06744_, _06743_, _06739_);
  not _15098_ (_06745_, _06744_);
  and _15099_ (_06746_, _06130_, _06287_);
  not _15100_ (_06747_, _06600_);
  and _15101_ (_06748_, _06747_, _06746_);
  or _15102_ (_06749_, _06290_, _06142_);
  and _15103_ (_06750_, _06127_, _06117_);
  and _15104_ (_06751_, _06740_, _06750_);
  nor _15105_ (_06752_, _06751_, _06118_);
  nand _15106_ (_06753_, _06752_, _06142_);
  and _15107_ (_06754_, _06753_, _06749_);
  nor _15108_ (_06755_, _06754_, _06748_);
  and _15109_ (_06756_, _06755_, _06745_);
  and _15110_ (_06757_, _06756_, _06738_);
  and _15111_ (_06758_, _06757_, _06730_);
  not _15112_ (_06759_, _06758_);
  nor _15113_ (_06760_, _06759_, _06729_);
  not _15114_ (_06761_, _06760_);
  nor _15115_ (_06762_, _06761_, _06713_);
  and _15116_ (_06763_, _06762_, _06676_);
  not _15117_ (_06764_, _06001_);
  and _15118_ (_06765_, _06764_, _05958_);
  nor _15119_ (_06766_, _06527_, _05971_);
  and _15120_ (_06767_, _06766_, _06020_);
  and _15121_ (_06768_, _06767_, _06765_);
  not _15122_ (_06769_, _06054_);
  nor _15123_ (_06770_, _06043_, _06030_);
  and _15124_ (_06771_, _06770_, _06769_);
  and _15125_ (_06772_, _06771_, _06768_);
  nand _15126_ (_06773_, _06772_, _06763_);
  and _15127_ (_06774_, _06523_, _06067_);
  and _15128_ (_06775_, _06774_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  or _15129_ (_06776_, _06772_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and _15130_ (_06777_, _06776_, _06775_);
  and _15131_ (_06778_, _06777_, _06773_);
  and _15132_ (_06779_, _06766_, _06765_);
  and _15133_ (_06781_, _06779_, _06061_);
  not _15134_ (_06782_, _06781_);
  and _15135_ (_06783_, _06600_, _06253_);
  not _15136_ (_06784_, _06783_);
  not _15137_ (_06785_, _06295_);
  and _15138_ (_06786_, _06364_, _06142_);
  nor _15139_ (_06787_, _06786_, _06785_);
  and _15140_ (_06788_, _06787_, _06784_);
  and _15141_ (_06789_, _06714_, _06252_);
  nor _15142_ (_06790_, _06789_, _06253_);
  and _15143_ (_06791_, _06162_, _06111_);
  and _15144_ (_06792_, _06791_, _06257_);
  and _15145_ (_06793_, _06792_, _06500_);
  nor _15146_ (_06794_, _06793_, _06142_);
  or _15147_ (_06795_, _06794_, _06790_);
  and _15148_ (_06796_, _06795_, _06600_);
  nor _15149_ (_06797_, _06795_, _06600_);
  nor _15150_ (_06798_, _06797_, _06796_);
  and _15151_ (_06799_, _06798_, _06266_);
  nor _15152_ (_06800_, _06799_, _06788_);
  nor _15153_ (_06801_, _06602_, _06283_);
  and _15154_ (_06802_, _06604_, _06300_);
  nor _15155_ (_06803_, _06802_, _06801_);
  and _15156_ (_06804_, _06603_, _06288_);
  and _15157_ (_06805_, _06600_, _06290_);
  nor _15158_ (_06806_, _06805_, _06804_);
  nor _15159_ (_06807_, _06600_, _06133_);
  not _15160_ (_06808_, _06807_);
  and _15161_ (_06809_, _06808_, _06806_);
  and _15162_ (_06810_, _06809_, _06803_);
  and _15163_ (_06811_, _06810_, _06800_);
  nor _15164_ (_06812_, _06811_, _06782_);
  and _15165_ (_06813_, _06782_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or _15166_ (_06814_, _06813_, _06812_);
  and _15167_ (_06815_, _06814_, _06524_);
  not _15168_ (_06816_, _06774_);
  and _15169_ (_06817_, _06816_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or _15170_ (_06818_, _06817_, rst);
  or _15171_ (_06819_, _06818_, _06815_);
  or _15172_ (_02004_, _06819_, _06778_);
  or _15173_ (_06820_, _06321_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  or _15174_ (_06821_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _05556_);
  or _15175_ (_06822_, _06821_, _05586_);
  and _15176_ (_06823_, _06822_, _05552_);
  and _15177_ (_02117_, _06823_, _06820_);
  or _15178_ (_06824_, _06321_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  or _15179_ (_06825_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _05556_);
  or _15180_ (_06826_, _06825_, _05586_);
  and _15181_ (_06827_, _06826_, _05552_);
  and _15182_ (_02328_, _06827_, _06824_);
  and _15183_ (_06828_, _06328_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7]);
  and _15184_ (_06829_, _06747_, _06366_);
  and _15185_ (_06830_, _06829_, _06502_);
  or _15186_ (_06831_, _06600_, _06410_);
  or _15187_ (_06832_, _06498_, _06420_);
  or _15188_ (_06833_, _06832_, _06831_);
  nand _15189_ (_06834_, _06832_, _06831_);
  and _15190_ (_06835_, _06834_, _06833_);
  not _15191_ (_06836_, _06835_);
  or _15192_ (_06837_, _06836_, _06505_);
  or _15193_ (_06838_, _06836_, _06499_);
  and _15194_ (_06839_, _06838_, _06837_);
  not _15195_ (_06840_, _06839_);
  nand _15196_ (_06841_, _06840_, _06830_);
  or _15197_ (_06842_, _06840_, _06830_);
  and _15198_ (_06843_, _06842_, _06841_);
  nor _15199_ (_06844_, _06507_, _06439_);
  nand _15200_ (_06845_, _06836_, _06505_);
  nand _15201_ (_06846_, _06845_, _06837_);
  nand _15202_ (_06847_, _06846_, _06499_);
  and _15203_ (_06848_, _06847_, _06838_);
  nand _15204_ (_06849_, _06848_, _06844_);
  or _15205_ (_06850_, _06848_, _06844_);
  and _15206_ (_06851_, _06850_, _06849_);
  or _15207_ (_06852_, _06507_, _06442_);
  nand _15208_ (_06853_, _06852_, _06512_);
  nand _15209_ (_06854_, _06853_, _06851_);
  nand _15210_ (_06855_, _06854_, _06849_);
  nand _15211_ (_06856_, _06855_, _06843_);
  and _15212_ (_06857_, _06841_, _06833_);
  nand _15213_ (_06858_, _06857_, _06856_);
  nand _15214_ (_06859_, _06858_, _06828_);
  or _15215_ (_06860_, _06858_, _06828_);
  nand _15216_ (_06861_, _06860_, _06859_);
  and _15217_ (_06862_, _06328_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6]);
  or _15218_ (_06863_, _06855_, _06843_);
  and _15219_ (_06864_, _06863_, _06856_);
  nand _15220_ (_06865_, _06864_, _06862_);
  or _15221_ (_06866_, _06865_, _06861_);
  nand _15222_ (_06867_, _06866_, _06859_);
  and _15223_ (_06868_, _06328_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8]);
  and _15224_ (_06869_, _06328_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  and _15225_ (_06870_, _06869_, _06868_);
  and _15226_ (_06871_, _06870_, _06867_);
  and _15227_ (_06872_, _06328_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5]);
  or _15228_ (_06873_, _06853_, _06851_);
  and _15229_ (_06874_, _06873_, _06854_);
  nand _15230_ (_06875_, _06874_, _06872_);
  or _15231_ (_06876_, _06874_, _06872_);
  nand _15232_ (_06877_, _06876_, _06875_);
  and _15233_ (_06878_, _06518_, _06515_);
  or _15234_ (_06879_, _06878_, _06877_);
  and _15235_ (_06880_, _06879_, _06875_);
  or _15236_ (_06881_, _06864_, _06862_);
  nand _15237_ (_06882_, _06881_, _06865_);
  nor _15238_ (_06883_, _06882_, _06861_);
  nand _15239_ (_06884_, _06870_, _06883_);
  nor _15240_ (_06885_, _06884_, _06880_);
  nor _15241_ (_06886_, _06885_, _06871_);
  or _15242_ (_06887_, _06882_, _06880_);
  and _15243_ (_06888_, _06887_, _06865_);
  or _15244_ (_06889_, _06888_, _06861_);
  nand _15245_ (_06890_, _06889_, _06859_);
  nand _15246_ (_06891_, _06890_, _06868_);
  not _15247_ (_06892_, _06869_);
  nand _15248_ (_06893_, _06892_, _06891_);
  and _15249_ (_06895_, _06893_, _06886_);
  and _15250_ (_03645_, _06895_, _05552_);
  or _15251_ (_06896_, _06885_, _06871_);
  and _15252_ (_06897_, _06328_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10]);
  and _15253_ (_06898_, _06328_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  and _15254_ (_06899_, _06898_, _06897_);
  nand _15255_ (_06901_, _06899_, _06896_);
  nand _15256_ (_06902_, _06897_, _06896_);
  not _15257_ (_06903_, _06898_);
  nand _15258_ (_06904_, _06903_, _06902_);
  and _15259_ (_06905_, _06904_, _06901_);
  and _15260_ (_03742_, _06905_, _05552_);
  or _15261_ (_06906_, _06897_, _06896_);
  and _15262_ (_06908_, _06906_, _06902_);
  and _15263_ (_04571_, _06908_, _05552_);
  and _15264_ (_06910_, _06001_, _05958_);
  not _15265_ (_06911_, _05971_);
  and _15266_ (_06913_, _06020_, _06527_);
  and _15267_ (_06915_, _06913_, _06911_);
  and _15268_ (_06916_, _06915_, _06910_);
  and _15269_ (_06918_, _06916_, _06771_);
  nand _15270_ (_06919_, _06918_, _06763_);
  or _15271_ (_06921_, _06918_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and _15272_ (_06922_, _06921_, _06775_);
  and _15273_ (_06924_, _06922_, _06919_);
  not _15274_ (_06925_, _05958_);
  nor _15275_ (_06926_, _05971_, _06925_);
  and _15276_ (_06927_, _06926_, _06528_);
  and _15277_ (_06928_, _06927_, _06061_);
  nand _15278_ (_06929_, _06928_, _06811_);
  or _15279_ (_06930_, _06928_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and _15280_ (_06931_, _06930_, _06524_);
  and _15281_ (_06932_, _06931_, _06929_);
  and _15282_ (_06933_, _06816_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  or _15283_ (_06934_, _06933_, rst);
  or _15284_ (_06935_, _06934_, _06932_);
  or _15285_ (_05142_, _06935_, _06924_);
  or _15286_ (_06936_, _06321_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2]);
  or _15287_ (_06937_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _05556_);
  or _15288_ (_06938_, _06937_, _05586_);
  and _15289_ (_06939_, _06938_, _05552_);
  and _15290_ (_05539_, _06939_, _06936_);
  or _15291_ (_06940_, _06321_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1]);
  or _15292_ (_06941_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2], _05556_);
  or _15293_ (_06942_, _06941_, _05586_);
  and _15294_ (_06943_, _06942_, _05552_);
  and _15295_ (_05540_, _06943_, _06940_);
  or _15296_ (_06944_, _06321_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  or _15297_ (_06945_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1], _05556_);
  or _15298_ (_06946_, _06945_, _05586_);
  and _15299_ (_06947_, _06946_, _05552_);
  and _15300_ (_05541_, _06947_, _06944_);
  and _15301_ (_06948_, _06065_, _06003_);
  and _15302_ (_06949_, _06948_, _06068_);
  nand _15303_ (_06950_, _06949_, _06306_);
  or _15304_ (_06951_, _06949_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  and _15305_ (_06952_, _06951_, _05552_);
  and _15306_ (_05578_, _06952_, _06950_);
  not _15307_ (_06953_, _06058_);
  nor _15308_ (_06954_, _06560_, _06953_);
  not _15309_ (_06955_, _06068_);
  and _15310_ (_06956_, _06953_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  or _15311_ (_06957_, _06956_, _06955_);
  or _15312_ (_06958_, _06957_, _06954_);
  or _15313_ (_06959_, _06068_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  and _15314_ (_06960_, _06959_, _05552_);
  and _15315_ (_05581_, _06960_, _06958_);
  not _15316_ (_06962_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1]);
  and _15317_ (_06963_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], _05545_);
  and _15318_ (_06965_, _06963_, _06962_);
  not _15319_ (_06966_, _06965_);
  not _15320_ (_06967_, _06524_);
  and _15321_ (_06968_, _06764_, _05989_);
  and _15322_ (_06969_, _06968_, _06529_);
  nand _15323_ (_06970_, _06969_, _06061_);
  or _15324_ (_06971_, _06970_, _06967_);
  and _15325_ (_06972_, _06971_, _06966_);
  not _15326_ (_06973_, _06972_);
  or _15327_ (_06974_, _06639_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  not _15328_ (_06975_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or _15329_ (_06976_, _06631_, _06975_);
  and _15330_ (_06977_, _06976_, _06974_);
  or _15331_ (_06978_, _06977_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or _15332_ (_06979_, _06625_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or _15333_ (_06980_, _06399_, _06975_);
  and _15334_ (_06981_, _06980_, _06979_);
  or _15335_ (_06982_, _06981_, _06313_);
  nand _15336_ (_06983_, _06982_, _06978_);
  and _15337_ (_06984_, _06982_, _06978_);
  nor _15338_ (_06985_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1], \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _15339_ (_06986_, _06985_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7]);
  not _15340_ (_06987_, _06986_);
  nand _15341_ (_06988_, _06985_, _06600_);
  and _15342_ (_06989_, _06988_, _06987_);
  not _15343_ (_06990_, _06989_);
  or _15344_ (_06991_, _06990_, _06984_);
  nor _15345_ (_06992_, _06985_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6]);
  not _15346_ (_06993_, _06992_);
  nand _15347_ (_06994_, _06985_, _06498_);
  and _15348_ (_06995_, _06994_, _06993_);
  not _15349_ (_06996_, _06995_);
  and _15350_ (_06997_, _06635_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or _15351_ (_06998_, _06997_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or _15352_ (_06999_, _06534_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or _15353_ (_07000_, _06279_, _06975_);
  and _15354_ (_07001_, _07000_, _06999_);
  or _15355_ (_07002_, _07001_, _06313_);
  and _15356_ (_07003_, _07002_, _06998_);
  or _15357_ (_07004_, _07003_, _06996_);
  or _15358_ (_07005_, _06989_, _06983_);
  and _15359_ (_07006_, _07005_, _06991_);
  not _15360_ (_07007_, _07006_);
  or _15361_ (_07008_, _07007_, _07004_);
  and _15362_ (_07009_, _07008_, _06991_);
  nand _15363_ (_07010_, _07002_, _06998_);
  or _15364_ (_07011_, _07010_, _06995_);
  and _15365_ (_07012_, _07011_, _07004_);
  and _15366_ (_07013_, _07012_, _07006_);
  not _15367_ (_07014_, _06985_);
  or _15368_ (_07015_, _07014_, _06111_);
  nor _15369_ (_07016_, _06985_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5]);
  not _15370_ (_07017_, _07016_);
  nand _15371_ (_07018_, _07017_, _07015_);
  and _15372_ (_07019_, _06639_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or _15373_ (_07020_, _07019_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or _15374_ (_07021_, _06631_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or _15375_ (_07022_, _06625_, _06975_);
  and _15376_ (_07023_, _07022_, _07021_);
  or _15377_ (_07024_, _07023_, _06313_);
  and _15378_ (_07025_, _07024_, _07020_);
  or _15379_ (_07026_, _07025_, _07018_);
  or _15380_ (_07027_, _06635_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or _15381_ (_07028_, _06534_, _06975_);
  and _15382_ (_07029_, _07028_, _07027_);
  and _15383_ (_07030_, _07029_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nor _15384_ (_07031_, _06985_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4]);
  not _15385_ (_07032_, _07031_);
  or _15386_ (_07033_, _07014_, _06162_);
  nand _15387_ (_07034_, _07033_, _07032_);
  or _15388_ (_07035_, _07034_, _07030_);
  and _15389_ (_07036_, _07017_, _07015_);
  nand _15390_ (_07037_, _07024_, _07020_);
  or _15391_ (_07038_, _07037_, _07036_);
  nand _15392_ (_07039_, _07038_, _07026_);
  or _15393_ (_07040_, _07039_, _07035_);
  nand _15394_ (_07041_, _07040_, _07026_);
  nand _15395_ (_07042_, _07041_, _07013_);
  and _15396_ (_07043_, _07042_, _07009_);
  and _15397_ (_07044_, _06977_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not _15398_ (_07045_, _07044_);
  nor _15399_ (_07046_, _06985_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3]);
  not _15400_ (_07047_, _07046_);
  or _15401_ (_07048_, _07014_, _06184_);
  and _15402_ (_07049_, _07048_, _07047_);
  nand _15403_ (_07050_, _07049_, _07045_);
  or _15404_ (_07051_, _07049_, _07045_);
  nand _15405_ (_07052_, _07051_, _07050_);
  nand _15406_ (_07053_, _06997_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or _15407_ (_07054_, _07014_, _06227_);
  nor _15408_ (_07055_, _06985_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2]);
  not _15409_ (_07056_, _07055_);
  and _15410_ (_07057_, _07056_, _07054_);
  nand _15411_ (_07058_, _07057_, _07053_);
  and _15412_ (_07059_, _07019_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or _15413_ (_07060_, _07014_, _06248_);
  nor _15414_ (_07061_, _06985_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1]);
  not _15415_ (_07062_, _07061_);
  nand _15416_ (_07063_, _07062_, _07060_);
  and _15417_ (_07064_, _07063_, _07059_);
  or _15418_ (_07065_, _07057_, _07053_);
  nand _15419_ (_07066_, _07065_, _07058_);
  or _15420_ (_07067_, _07066_, _07064_);
  and _15421_ (_07068_, _07067_, _07058_);
  or _15422_ (_07069_, _07068_, _07052_);
  nand _15423_ (_07070_, _07069_, _07050_);
  nand _15424_ (_07071_, _07034_, _07030_);
  and _15425_ (_07072_, _07071_, _07035_);
  and _15426_ (_07073_, _07038_, _07026_);
  and _15427_ (_07074_, _07073_, _07072_);
  and _15428_ (_07075_, _07074_, _07013_);
  nand _15429_ (_07076_, _07075_, _07070_);
  nand _15430_ (_07077_, _07076_, _07043_);
  nor _15431_ (_07078_, _07029_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or _15432_ (_07079_, _06279_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand _15433_ (_07081_, _06364_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand _15434_ (_07082_, _07081_, _07079_);
  and _15435_ (_07084_, _07082_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nor _15436_ (_07086_, _07084_, _07078_);
  not _15437_ (_07087_, _07086_);
  and _15438_ (_07088_, _06364_, _06606_);
  nor _15439_ (_07089_, _07088_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _15440_ (_07090_, _07001_, _06981_);
  not _15441_ (_07091_, _07023_);
  and _15442_ (_07092_, _07082_, _07091_);
  nand _15443_ (_07093_, _07092_, _07090_);
  and _15444_ (_07094_, _07093_, _06313_);
  nor _15445_ (_07095_, _07094_, _07089_);
  and _15446_ (_07096_, _07095_, _07087_);
  nand _15447_ (_07097_, _07096_, _07077_);
  not _15448_ (_07098_, _07012_);
  and _15449_ (_07099_, _07025_, _07018_);
  not _15450_ (_07100_, _07035_);
  and _15451_ (_07101_, _07072_, _07070_);
  nor _15452_ (_07102_, _07101_, _07100_);
  or _15453_ (_07103_, _07102_, _07099_);
  and _15454_ (_07104_, _07103_, _07026_);
  nor _15455_ (_07105_, _07104_, _07098_);
  and _15456_ (_07106_, _07104_, _07098_);
  nor _15457_ (_07108_, _07106_, _07105_);
  nor _15458_ (_07110_, _07108_, _07097_);
  and _15459_ (_07111_, _07097_, _06996_);
  nor _15460_ (_07112_, _07111_, _07110_);
  and _15461_ (_07114_, _07112_, _06983_);
  nor _15462_ (_07115_, _07112_, _06983_);
  nor _15463_ (_07116_, _07115_, _07114_);
  and _15464_ (_07117_, _07096_, _07077_);
  nand _15465_ (_07118_, _07039_, _07102_);
  or _15466_ (_07119_, _07039_, _07102_);
  nand _15467_ (_07120_, _07119_, _07118_);
  nand _15468_ (_07121_, _07120_, _07117_);
  and _15469_ (_07122_, _07097_, _07018_);
  not _15470_ (_07123_, _07122_);
  and _15471_ (_07124_, _07123_, _07121_);
  and _15472_ (_07125_, _07124_, _07010_);
  nor _15473_ (_07126_, _07072_, _07070_);
  or _15474_ (_07127_, _07126_, _07101_);
  and _15475_ (_07128_, _07127_, _07117_);
  and _15476_ (_07129_, _07097_, _07034_);
  nor _15477_ (_07130_, _07129_, _07128_);
  and _15478_ (_07131_, _07130_, _07037_);
  not _15479_ (_07132_, _07131_);
  nor _15480_ (_07133_, _07124_, _07010_);
  or _15481_ (_07134_, _07133_, _07125_);
  nor _15482_ (_07135_, _07134_, _07132_);
  nor _15483_ (_07136_, _07135_, _07125_);
  not _15484_ (_07137_, _07030_);
  and _15485_ (_07138_, _07068_, _07052_);
  not _15486_ (_07140_, _07138_);
  and _15487_ (_07141_, _07140_, _07069_);
  or _15488_ (_07142_, _07141_, _07097_);
  or _15489_ (_07143_, _07117_, _07049_);
  and _15490_ (_07144_, _07143_, _07142_);
  nor _15491_ (_07145_, _07144_, _07137_);
  not _15492_ (_07146_, _07145_);
  not _15493_ (_07147_, _07059_);
  or _15494_ (_07148_, _07097_, _07147_);
  nand _15495_ (_07149_, _07148_, _07063_);
  or _15496_ (_07150_, _07148_, _07063_);
  and _15497_ (_07151_, _07150_, _07149_);
  nand _15498_ (_07152_, _07151_, _07053_);
  or _15499_ (_07153_, _07151_, _07053_);
  and _15500_ (_07154_, _07153_, _07152_);
  and _15501_ (_07155_, _06985_, _06206_);
  nor _15502_ (_07156_, _06985_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0]);
  nor _15503_ (_07157_, _07156_, _07155_);
  nor _15504_ (_07158_, _07157_, _07147_);
  not _15505_ (_07159_, _07158_);
  nand _15506_ (_07160_, _07159_, _07154_);
  and _15507_ (_07161_, _07160_, _07152_);
  or _15508_ (_07162_, _07117_, _07057_);
  and _15509_ (_07163_, _07066_, _07064_);
  not _15510_ (_07164_, _07163_);
  and _15511_ (_07165_, _07164_, _07067_);
  or _15512_ (_07166_, _07165_, _07097_);
  and _15513_ (_07167_, _07166_, _07162_);
  nand _15514_ (_07168_, _07167_, _07045_);
  or _15515_ (_07169_, _07167_, _07045_);
  nand _15516_ (_07170_, _07169_, _07168_);
  or _15517_ (_07171_, _07170_, _07161_);
  and _15518_ (_07172_, _07144_, _07137_);
  not _15519_ (_07173_, _07172_);
  and _15520_ (_07174_, _07173_, _07168_);
  nand _15521_ (_07175_, _07174_, _07171_);
  and _15522_ (_07176_, _07175_, _07146_);
  nor _15523_ (_07177_, _07130_, _07037_);
  nor _15524_ (_07178_, _07177_, _07131_);
  not _15525_ (_07179_, _07178_);
  nor _15526_ (_07181_, _07134_, _07179_);
  nand _15527_ (_07182_, _07181_, _07176_);
  nand _15528_ (_07183_, _07182_, _07136_);
  nand _15529_ (_07184_, _07183_, _07116_);
  not _15530_ (_07185_, _07114_);
  and _15531_ (_07186_, _07097_, _06989_);
  not _15532_ (_07187_, _07105_);
  and _15533_ (_07188_, _07187_, _07004_);
  nand _15534_ (_07189_, _07188_, _07006_);
  or _15535_ (_07190_, _07188_, _07006_);
  nand _15536_ (_07191_, _07190_, _07189_);
  and _15537_ (_07192_, _07191_, _07117_);
  nor _15538_ (_07193_, _07192_, _07186_);
  or _15539_ (_07194_, _07193_, _07086_);
  and _15540_ (_07195_, _07194_, _07185_);
  nand _15541_ (_07196_, _07195_, _07184_);
  and _15542_ (_07197_, _07193_, _07086_);
  not _15543_ (_07198_, _07197_);
  and _15544_ (_07199_, _07198_, _07095_);
  and _15545_ (_07200_, _07199_, _07196_);
  and _15546_ (_07201_, _07198_, _07194_);
  nand _15547_ (_07202_, _07184_, _07185_);
  or _15548_ (_07203_, _07202_, _07201_);
  nand _15549_ (_07204_, _07202_, _07201_);
  and _15550_ (_07205_, _07204_, _07203_);
  nand _15551_ (_07206_, _07205_, _07200_);
  or _15552_ (_07208_, _07200_, _07193_);
  nand _15553_ (_07209_, _07208_, _07206_);
  nand _15554_ (_07210_, _07209_, _06314_);
  and _15555_ (_07211_, _06287_, _06114_);
  and _15556_ (_07212_, _06899_, _06896_);
  and _15557_ (_07213_, _06328_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12]);
  nand _15558_ (_07214_, _07213_, _07212_);
  and _15559_ (_07215_, _06328_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  nand _15560_ (_07216_, _07215_, _07214_);
  or _15561_ (_07217_, _07214_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  nand _15562_ (_07218_, _07217_, _07216_);
  nand _15563_ (_07219_, _07218_, _07211_);
  not _15564_ (_07220_, _06604_);
  and _15565_ (_07221_, _06672_, _07220_);
  nor _15566_ (_07222_, _06672_, _07220_);
  nor _15567_ (_07224_, _07222_, _07221_);
  and _15568_ (_07225_, _07224_, _06581_);
  not _15569_ (_07226_, _07225_);
  nor _15570_ (_07227_, _06710_, _06604_);
  and _15571_ (_07228_, _06710_, _06604_);
  or _15572_ (_07229_, _07228_, _07227_);
  and _15573_ (_07230_, _07229_, _06677_);
  nor _15574_ (_07231_, _06714_, _06600_);
  nor _15575_ (_07232_, _07231_, _06142_);
  and _15576_ (_07233_, _07232_, _06730_);
  nor _15577_ (_07234_, _07233_, _06720_);
  and _15578_ (_07235_, _07234_, _06600_);
  nor _15579_ (_07236_, _07234_, _06600_);
  nor _15580_ (_07237_, _07236_, _07235_);
  nor _15581_ (_07238_, _07237_, _06724_);
  and _15582_ (_07239_, _06368_, _06750_);
  and _15583_ (_07240_, _06142_, _06736_);
  nor _15584_ (_07241_, _07240_, _07239_);
  nor _15585_ (_07242_, _06600_, _06119_);
  and _15586_ (_07243_, _06500_, _06131_);
  nor _15587_ (_07244_, _07243_, _07242_);
  and _15588_ (_07245_, _07244_, _07241_);
  and _15589_ (_07246_, _07245_, _06806_);
  and _15590_ (_07247_, _07246_, _06803_);
  not _15591_ (_07248_, _07247_);
  nor _15592_ (_07249_, _07248_, _07238_);
  and _15593_ (_07250_, _07249_, _06800_);
  not _15594_ (_07251_, _07250_);
  nor _15595_ (_07252_, _07251_, _07230_);
  and _15596_ (_07253_, _07252_, _07226_);
  and _15597_ (_07254_, _07253_, _07219_);
  nand _15598_ (_07255_, _07254_, _07210_);
  nand _15599_ (_07257_, _07255_, _06973_);
  not _15600_ (_07258_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and _15601_ (_07259_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], _05545_);
  and _15602_ (_07260_, _07259_, _07258_);
  not _15603_ (_07261_, _07260_);
  nor _15604_ (_07262_, _06001_, _05958_);
  and _15605_ (_07263_, _07262_, _06775_);
  and _15606_ (_07264_, _07263_, _06767_);
  and _15607_ (_07265_, _07264_, _06771_);
  and _15608_ (_07266_, _07265_, _06763_);
  and _15609_ (_07267_, _07262_, _06767_);
  and _15610_ (_07269_, _07267_, _06775_);
  and _15611_ (_07270_, _07269_, _06771_);
  nor _15612_ (_07271_, _07270_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or _15613_ (_07272_, _07271_, _06973_);
  or _15614_ (_07273_, _07272_, _07266_);
  and _15615_ (_07274_, _07273_, _07261_);
  nand _15616_ (_07275_, _07274_, _07257_);
  nor _15617_ (_07276_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and _15618_ (_07277_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _06085_);
  nor _15619_ (_07278_, _07277_, _07276_);
  nor _15620_ (_07279_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and _15621_ (_07280_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _06170_);
  nor _15622_ (_07281_, _07280_, _07279_);
  nor _15623_ (_07282_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and _15624_ (_07283_, _06192_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _15625_ (_07284_, _07283_, _07282_);
  not _15626_ (_07285_, _07284_);
  nor _15627_ (_07286_, _07285_, _06712_);
  nor _15628_ (_07288_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  and _15629_ (_07289_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _06235_);
  nor _15630_ (_07290_, _07289_, _07288_);
  and _15631_ (_07291_, _07290_, _07286_);
  nor _15632_ (_07292_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  and _15633_ (_07293_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _06219_);
  nor _15634_ (_07294_, _07293_, _07292_);
  and _15635_ (_07295_, _07294_, _07291_);
  and _15636_ (_07296_, _07295_, _07281_);
  nor _15637_ (_07297_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and _15638_ (_07298_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _06148_);
  nor _15639_ (_07299_, _07298_, _07297_);
  and _15640_ (_07300_, _07299_, _07296_);
  and _15641_ (_07301_, _07300_, _07278_);
  nor _15642_ (_07302_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and _15643_ (_07303_, _06487_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _15644_ (_07304_, _07303_, _07302_);
  and _15645_ (_07305_, _07304_, _07301_);
  nor _15646_ (_07306_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  and _15647_ (_07308_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _06590_);
  nor _15648_ (_07309_, _07308_, _07306_);
  or _15649_ (_07310_, _07309_, _07305_);
  nand _15650_ (_07311_, _07309_, _07305_);
  and _15651_ (_07312_, _07311_, _07310_);
  nand _15652_ (_07313_, _07312_, _06677_);
  and _15653_ (_07314_, _06878_, _06877_);
  not _15654_ (_07315_, _07314_);
  and _15655_ (_07316_, _07315_, _06879_);
  and _15656_ (_07317_, _07316_, _07211_);
  nor _15657_ (_07318_, _06600_, _06386_);
  and _15658_ (_07319_, _07318_, _06793_);
  and _15659_ (_07320_, _07319_, _06635_);
  and _15660_ (_07321_, _07320_, _06631_);
  and _15661_ (_07322_, _07321_, _06534_);
  and _15662_ (_07323_, _07322_, _06625_);
  nor _15663_ (_07325_, _07323_, _06142_);
  and _15664_ (_07326_, _06789_, _06600_);
  and _15665_ (_07327_, _06351_, _06386_);
  and _15666_ (_07328_, _06337_, _06373_);
  and _15667_ (_07329_, _07328_, _07327_);
  and _15668_ (_07330_, _07329_, _07326_);
  and _15669_ (_07331_, _07330_, _06379_);
  nor _15670_ (_07332_, _07331_, _06253_);
  nor _15671_ (_07333_, _07332_, _07325_);
  nor _15672_ (_07334_, _06279_, _06142_);
  nor _15673_ (_07335_, _07334_, _06296_);
  and _15674_ (_07336_, _07335_, _07333_);
  nor _15675_ (_07337_, _06399_, _06142_);
  and _15676_ (_07339_, _06399_, _06142_);
  nor _15677_ (_07340_, _07339_, _07337_);
  and _15678_ (_07342_, _07340_, _07336_);
  and _15679_ (_07343_, _07342_, _06583_);
  nor _15680_ (_07344_, _07342_, _06583_);
  nor _15681_ (_07345_, _07344_, _07343_);
  and _15682_ (_07346_, _07345_, _06266_);
  and _15683_ (_07347_, _06314_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  nor _15684_ (_07348_, _06785_, _06142_);
  or _15685_ (_07349_, _07348_, _06118_);
  and _15686_ (_07350_, _07349_, _06583_);
  or _15687_ (_07351_, _07350_, _07347_);
  and _15688_ (_07352_, _06184_, _06746_);
  and _15689_ (_07353_, _06725_, _06295_);
  or _15690_ (_07354_, _07353_, _07352_);
  nor _15691_ (_07355_, _07354_, _07351_);
  not _15692_ (_07356_, _07355_);
  nor _15693_ (_07357_, _07356_, _07346_);
  not _15694_ (_07358_, _07357_);
  nor _15695_ (_07359_, _07358_, _07317_);
  nand _15696_ (_07360_, _07359_, _07313_);
  or _15697_ (_07362_, _07360_, _07261_);
  and _15698_ (_07363_, _07362_, _07275_);
  and _15699_ (_05610_, _07363_, _05552_);
  and _15700_ (_07364_, _06532_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and _15701_ (_07365_, _06251_, _06142_);
  nor _15702_ (_07366_, _07365_, _06258_);
  and _15703_ (_07367_, _07366_, _06164_);
  nor _15704_ (_07368_, _07366_, _06164_);
  nor _15705_ (_07369_, _07368_, _07367_);
  and _15706_ (_07370_, _07369_, _06266_);
  and _15707_ (_07371_, _06379_, _06142_);
  nor _15708_ (_07372_, _07371_, _06785_);
  not _15709_ (_07373_, _07372_);
  nor _15710_ (_07374_, _07373_, _06163_);
  nor _15711_ (_07375_, _07374_, _07370_);
  and _15712_ (_07376_, _06162_, _06134_);
  not _15713_ (_07377_, _07376_);
  and _15714_ (_07378_, _06628_, _06300_);
  not _15715_ (_07379_, _07378_);
  nor _15716_ (_07380_, _06627_, _06283_);
  not _15717_ (_07381_, _07380_);
  and _15718_ (_07382_, _06626_, _06288_);
  nor _15719_ (_07383_, _06291_, _06162_);
  nor _15720_ (_07384_, _07383_, _07382_);
  and _15721_ (_07385_, _07384_, _07381_);
  and _15722_ (_07386_, _07385_, _07379_);
  and _15723_ (_07387_, _07386_, _07377_);
  and _15724_ (_07388_, _07387_, _07375_);
  nor _15725_ (_07389_, _07388_, _06532_);
  nor _15726_ (_07390_, _07389_, _07364_);
  not _15727_ (_07391_, _07390_);
  and _15728_ (_07392_, _06562_, _05669_);
  and _15729_ (_07393_, _07392_, _07391_);
  and _15730_ (_07394_, _07393_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  and _15731_ (_07395_, _06562_, _05818_);
  and _15732_ (_07396_, _07395_, _07391_);
  and _15733_ (_07397_, _07396_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  nor _15734_ (_07398_, _07397_, _07394_);
  nor _15735_ (_07399_, _06562_, _05818_);
  and _15736_ (_07400_, _07399_, _07391_);
  and _15737_ (_07401_, _07400_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  nor _15738_ (_07402_, _06562_, _05669_);
  and _15739_ (_07403_, _07402_, _07391_);
  and _15740_ (_07404_, _07403_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  nor _15741_ (_07405_, _07404_, _07401_);
  and _15742_ (_07406_, _07405_, _07398_);
  and _15743_ (_07407_, _07395_, _07390_);
  and _15744_ (_07408_, _07407_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  and _15745_ (_07410_, _07392_, _07390_);
  and _15746_ (_07411_, _07410_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  nor _15747_ (_07412_, _07411_, _07408_);
  and _15748_ (_07413_, _07399_, _07390_);
  and _15749_ (_07414_, _07413_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  and _15750_ (_07416_, _07402_, _07390_);
  and _15751_ (_07417_, _07416_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  nor _15752_ (_07418_, _07417_, _07414_);
  and _15753_ (_07419_, _07418_, _07412_);
  and _15754_ (_07420_, _07419_, _07406_);
  nor _15755_ (_07421_, _07390_, _06527_);
  and _15756_ (_07422_, _07390_, _06527_);
  nor _15757_ (_07423_, _07422_, _07421_);
  and _15758_ (_07424_, _06562_, _06064_);
  nor _15759_ (_07425_, _06059_, _05669_);
  not _15760_ (_07426_, _07425_);
  and _15761_ (_07427_, _06068_, _06054_);
  and _15762_ (_07428_, _07427_, _06001_);
  and _15763_ (_07429_, _07428_, _05972_);
  nand _15764_ (_07430_, _07429_, _07426_);
  nor _15765_ (_07431_, _07430_, _07424_);
  nor _15766_ (_07432_, _06562_, _06064_);
  and _15767_ (_07433_, _06043_, _06031_);
  nor _15768_ (_07434_, _07433_, _05818_);
  nor _15769_ (_07435_, _07434_, _07432_);
  and _15770_ (_07436_, _07435_, _07431_);
  and _15771_ (_07437_, _07436_, _07423_);
  nor _15772_ (_07438_, _07437_, _07420_);
  not _15773_ (_07439_, _06811_);
  and _15774_ (_07440_, _07437_, _07439_);
  nor _15775_ (_07441_, _07440_, _07438_);
  nor _15776_ (_05672_, _07441_, rst);
  and _15777_ (_07442_, _06525_, _06054_);
  and _15778_ (_07443_, _06910_, _06766_);
  and _15779_ (_07444_, _07443_, _07442_);
  and _15780_ (_07445_, _07444_, _06770_);
  nand _15781_ (_07446_, _07199_, _07196_);
  or _15782_ (_07447_, _07172_, _07145_);
  and _15783_ (_07448_, _07171_, _07168_);
  nor _15784_ (_07449_, _07448_, _07447_);
  and _15785_ (_07450_, _07448_, _07447_);
  nor _15786_ (_07451_, _07450_, _07449_);
  or _15787_ (_07452_, _07451_, _07446_);
  or _15788_ (_07453_, _07200_, _07144_);
  and _15789_ (_07454_, _07453_, _07452_);
  nand _15790_ (_07455_, _07454_, _06314_);
  nand _15791_ (_07456_, _06895_, _07211_);
  and _15792_ (_07457_, _06694_, _06687_);
  or _15793_ (_07458_, _07457_, _06678_);
  nor _15794_ (_07459_, _07458_, _06695_);
  not _15795_ (_07460_, _07459_);
  and _15796_ (_07461_, _06662_, _06649_);
  nor _15797_ (_07462_, _07461_, _06663_);
  nor _15798_ (_07463_, _07462_, _06582_);
  and _15799_ (_07464_, _06184_, _06118_);
  and _15800_ (_07465_, _06227_, _06131_);
  nor _15801_ (_07466_, _07465_, _07464_);
  nor _15802_ (_07467_, _06717_, _06724_);
  not _15803_ (_07468_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor _15804_ (_07469_, _06249_, _07468_);
  or _15805_ (_07470_, _07469_, _06184_);
  nand _15806_ (_07471_, _07470_, _07467_);
  nand _15807_ (_07472_, _06162_, _06128_);
  and _15808_ (_07473_, _07472_, _06555_);
  and _15809_ (_07474_, _07473_, _07471_);
  and _15810_ (_07475_, _07474_, _07466_);
  and _15811_ (_07476_, _07475_, _06543_);
  and _15812_ (_07477_, _07476_, _06552_);
  not _15813_ (_07478_, _07477_);
  nor _15814_ (_07479_, _07478_, _07463_);
  and _15815_ (_07481_, _07479_, _07460_);
  and _15816_ (_07482_, _07481_, _07456_);
  nand _15817_ (_07483_, _07482_, _07455_);
  and _15818_ (_07484_, _07483_, _07445_);
  and _15819_ (_07485_, _07259_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  not _15820_ (_07486_, _07445_);
  and _15821_ (_07487_, _07486_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or _15822_ (_07488_, _07487_, _07485_);
  or _15823_ (_07489_, _07488_, _07484_);
  and _15824_ (_07490_, _06534_, _06118_);
  nor _15825_ (_07491_, _07321_, _06142_);
  and _15826_ (_07492_, _07327_, _07326_);
  and _15827_ (_07493_, _07492_, _06373_);
  nor _15828_ (_07494_, _07493_, _06253_);
  or _15829_ (_07495_, _07494_, _07491_);
  and _15830_ (_07496_, _07495_, _06337_);
  nor _15831_ (_07497_, _07495_, _06337_);
  nor _15832_ (_07498_, _07497_, _07496_);
  and _15833_ (_07499_, _07498_, _06266_);
  and _15834_ (_07500_, _06295_, _06184_);
  or _15835_ (_07501_, _07500_, _07499_);
  or _15836_ (_07503_, _07501_, _06748_);
  and _15837_ (_07504_, _06314_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  nor _15838_ (_07505_, _07295_, _07281_);
  nor _15839_ (_07506_, _07505_, _07296_);
  and _15840_ (_07507_, _07506_, _06677_);
  and _15841_ (_07508_, _06462_, _06459_);
  not _15842_ (_07509_, _07508_);
  and _15843_ (_07510_, _07509_, _06463_);
  and _15844_ (_07511_, _07510_, _07211_);
  or _15845_ (_07512_, _07511_, _07507_);
  or _15846_ (_07513_, _07512_, _07504_);
  or _15847_ (_07514_, _07513_, _07503_);
  nor _15848_ (_07515_, _07514_, _07490_);
  nand _15849_ (_07516_, _07515_, _07485_);
  and _15850_ (_07517_, _07516_, _05552_);
  and _15851_ (_05863_, _07517_, _07489_);
  or _15852_ (_07518_, _07183_, _07116_);
  nand _15853_ (_07519_, _07518_, _07184_);
  nand _15854_ (_07520_, _07519_, _07200_);
  or _15855_ (_07521_, _07200_, _07112_);
  and _15856_ (_07522_, _07521_, _07520_);
  nand _15857_ (_07523_, _07522_, _06314_);
  or _15858_ (_07524_, _07213_, _07212_);
  and _15859_ (_07525_, _07524_, _07214_);
  nand _15860_ (_07526_, _07525_, _07211_);
  nor _15861_ (_07527_, _06670_, _06620_);
  nor _15862_ (_07528_, _07527_, _06671_);
  nor _15863_ (_07529_, _07528_, _06582_);
  not _15864_ (_07530_, _07529_);
  nor _15865_ (_07531_, _06706_, _06700_);
  nor _15866_ (_07532_, _07531_, _06678_);
  and _15867_ (_07533_, _07532_, _06708_);
  nor _15868_ (_07534_, _06498_, _06142_);
  or _15869_ (_07535_, _07534_, _07339_);
  and _15870_ (_07536_, _07535_, _06295_);
  or _15871_ (_07537_, _06792_, _06500_);
  and _15872_ (_07538_, _07537_, _06794_);
  and _15873_ (_07539_, _06252_, _06433_);
  nor _15874_ (_07540_, _06498_, _07539_);
  or _15875_ (_07542_, _07540_, _06789_);
  and _15876_ (_07543_, _07542_, _06142_);
  or _15877_ (_07544_, _07543_, _07538_);
  and _15878_ (_07545_, _07544_, _06266_);
  nor _15879_ (_07546_, _07545_, _07536_);
  nor _15880_ (_07547_, _07233_, _06719_);
  and _15881_ (_07548_, _07547_, _06433_);
  and _15882_ (_07549_, _07548_, _06498_);
  nor _15883_ (_07550_, _07548_, _06498_);
  nor _15884_ (_07551_, _07550_, _07549_);
  nor _15885_ (_07552_, _07551_, _06724_);
  and _15886_ (_07553_, _06611_, _06300_);
  and _15887_ (_07554_, _06608_, _06288_);
  nor _15888_ (_07555_, _06609_, _06283_);
  and _15889_ (_07556_, _06498_, _06290_);
  or _15890_ (_07557_, _07556_, _07555_);
  or _15891_ (_07558_, _07557_, _07554_);
  nor _15892_ (_07559_, _07558_, _07553_);
  not _15893_ (_07560_, _06128_);
  or _15894_ (_07561_, _06600_, _07560_);
  and _15895_ (_07562_, _06131_, _06111_);
  nor _15896_ (_07563_, _06498_, _06119_);
  nor _15897_ (_07564_, _07563_, _07562_);
  and _15898_ (_07565_, _07564_, _07561_);
  and _15899_ (_07566_, _07565_, _07559_);
  not _15900_ (_07567_, _07566_);
  nor _15901_ (_07568_, _07567_, _07552_);
  and _15902_ (_07569_, _07568_, _07546_);
  not _15903_ (_07570_, _07569_);
  nor _15904_ (_07571_, _07570_, _07533_);
  and _15905_ (_07572_, _07571_, _07530_);
  and _15906_ (_07573_, _07572_, _07526_);
  nand _15907_ (_07574_, _07573_, _07523_);
  and _15908_ (_07575_, _07574_, _07445_);
  and _15909_ (_07576_, _07486_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or _15910_ (_07577_, _07576_, _07485_);
  or _15911_ (_07578_, _07577_, _07575_);
  not _15912_ (_07579_, _07485_);
  and _15913_ (_07580_, _06399_, _06118_);
  and _15914_ (_07581_, _06227_, _06746_);
  and _15915_ (_07582_, _07336_, _06606_);
  nor _15916_ (_07583_, _07336_, _06606_);
  or _15917_ (_07584_, _07583_, _07582_);
  and _15918_ (_07585_, _07584_, _06266_);
  and _15919_ (_07586_, _06498_, _06142_);
  not _15920_ (_07587_, _07586_);
  nor _15921_ (_07588_, _07337_, _06785_);
  and _15922_ (_07589_, _07588_, _07587_);
  or _15923_ (_07590_, _07589_, _07585_);
  or _15924_ (_07591_, _07590_, _07581_);
  and _15925_ (_07592_, _06314_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  nor _15926_ (_07593_, _07304_, _07301_);
  nor _15927_ (_07594_, _07593_, _07305_);
  and _15928_ (_07595_, _07594_, _06677_);
  and _15929_ (_07596_, _06521_, _07211_);
  or _15930_ (_07597_, _07596_, _07595_);
  or _15931_ (_07598_, _07597_, _07592_);
  or _15932_ (_07599_, _07598_, _07591_);
  or _15933_ (_07600_, _07599_, _07580_);
  or _15934_ (_07601_, _07600_, _07579_);
  and _15935_ (_07602_, _07601_, _05552_);
  and _15936_ (_05866_, _07602_, _07578_);
  nand _15937_ (_07603_, _07178_, _07176_);
  and _15938_ (_07604_, _07603_, _07132_);
  nand _15939_ (_07605_, _07134_, _07604_);
  or _15940_ (_07606_, _07134_, _07604_);
  and _15941_ (_07607_, _07606_, _07605_);
  or _15942_ (_07608_, _07607_, _07446_);
  or _15943_ (_07609_, _07200_, _07124_);
  and _15944_ (_07610_, _07609_, _07608_);
  and _15945_ (_07611_, _07610_, _06314_);
  and _15946_ (_07612_, _06905_, _07211_);
  nor _15947_ (_07613_, _06669_, _06624_);
  nor _15948_ (_07614_, _07613_, _06670_);
  nor _15949_ (_07616_, _07614_, _06582_);
  nor _15950_ (_07617_, _06626_, _06301_);
  nor _15951_ (_07618_, _07617_, _06702_);
  or _15952_ (_07619_, _07618_, _06699_);
  nor _15953_ (_07620_, _06700_, _06678_);
  and _15954_ (_07621_, _07620_, _07619_);
  nor _15955_ (_07622_, _07547_, _06433_);
  or _15956_ (_07623_, _07622_, _07548_);
  and _15957_ (_07624_, _07623_, _06716_);
  and _15958_ (_07625_, _06118_, _06111_);
  and _15959_ (_07626_, _06162_, _06131_);
  nor _15960_ (_07627_, _06498_, _07560_);
  or _15961_ (_07628_, _07627_, _07626_);
  or _15962_ (_07629_, _07628_, _07625_);
  or _15963_ (_07630_, _07629_, _07624_);
  or _15964_ (_07631_, _07630_, _06305_);
  or _15965_ (_07632_, _07631_, _07621_);
  or _15966_ (_07633_, _07632_, _07616_);
  or _15967_ (_07634_, _07633_, _07612_);
  or _15968_ (_07635_, _07634_, _07611_);
  and _15969_ (_07636_, _07635_, _07445_);
  and _15970_ (_07637_, _07486_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or _15971_ (_07638_, _07637_, _07485_);
  or _15972_ (_07639_, _07638_, _07636_);
  or _15973_ (_07640_, _07300_, _07278_);
  nor _15974_ (_07641_, _07301_, _06678_);
  and _15975_ (_07642_, _07641_, _07640_);
  and _15976_ (_07643_, _06473_, _06470_);
  nand _15977_ (_07644_, _07643_, _06450_);
  or _15978_ (_07645_, _07643_, _06450_);
  and _15979_ (_07646_, _07645_, _07644_);
  and _15980_ (_07647_, _07646_, _07211_);
  nand _15981_ (_07648_, _07333_, _06279_);
  or _15982_ (_07649_, _07333_, _06279_);
  and _15983_ (_07650_, _07649_, _06266_);
  and _15984_ (_07651_, _07650_, _07648_);
  and _15985_ (_07652_, _06248_, _06746_);
  or _15986_ (_07653_, _06253_, _06111_);
  nor _15987_ (_07654_, _07334_, _06785_);
  and _15988_ (_07655_, _07654_, _07653_);
  and _15989_ (_07656_, _06279_, _06118_);
  and _15990_ (_07657_, _06314_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  or _15991_ (_07658_, _07657_, _07656_);
  or _15992_ (_07659_, _07658_, _07655_);
  or _15993_ (_07660_, _07659_, _07652_);
  or _15994_ (_07661_, _07660_, _07651_);
  or _15995_ (_07662_, _07661_, _07647_);
  or _15996_ (_07663_, _07662_, _07642_);
  or _15997_ (_07664_, _07663_, _07579_);
  and _15998_ (_07665_, _07664_, _05552_);
  and _15999_ (_05871_, _07665_, _07639_);
  nor _16000_ (_07666_, _06043_, _06031_);
  and _16001_ (_07667_, _07444_, _07666_);
  nor _16002_ (_07668_, _07667_, _07485_);
  or _16003_ (_07669_, _07668_, _07483_);
  not _16004_ (_07670_, _07668_);
  or _16005_ (_07671_, _07670_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and _16006_ (_07672_, _07671_, _05552_);
  and _16007_ (_05899_, _07672_, _07669_);
  nand _16008_ (_07674_, _07200_, _07059_);
  and _16009_ (_07675_, _07674_, _07157_);
  nor _16010_ (_07676_, _07674_, _07157_);
  or _16011_ (_07677_, _07676_, _07675_);
  nand _16012_ (_07678_, _07677_, _06314_);
  nor _16013_ (_07679_, _06658_, _06142_);
  nor _16014_ (_07680_, _07679_, _06688_);
  nor _16015_ (_07681_, _06677_, _06581_);
  not _16016_ (_07682_, _07681_);
  and _16017_ (_07683_, _07682_, _07680_);
  not _16018_ (_07684_, _07683_);
  and _16019_ (_07685_, _06656_, _06288_);
  and _16020_ (_07686_, _06290_, _06206_);
  nor _16021_ (_07687_, _07686_, _07685_);
  and _16022_ (_07688_, _06639_, _06295_);
  and _16023_ (_07689_, _06266_, _06206_);
  nor _16024_ (_07690_, _07689_, _07688_);
  and _16025_ (_07691_, _06747_, _06732_);
  and _16026_ (_07692_, _06142_, _06746_);
  nor _16027_ (_07693_, _07692_, _07691_);
  and _16028_ (_07694_, _07693_, _07690_);
  and _16029_ (_07695_, _07694_, _07687_);
  not _16030_ (_07696_, _06887_);
  and _16031_ (_07697_, _06882_, _06880_);
  nor _16032_ (_07698_, _07697_, _07696_);
  and _16033_ (_07699_, _07698_, _07211_);
  nor _16034_ (_07700_, _06656_, _06546_);
  nor _16035_ (_07701_, _07700_, _06282_);
  or _16036_ (_07702_, _07701_, _06657_);
  and _16037_ (_07703_, _06248_, _06128_);
  nor _16038_ (_07704_, _06716_, _06118_);
  nor _16039_ (_07705_, _07704_, _06206_);
  nor _16040_ (_07706_, _07705_, _07703_);
  nand _16041_ (_07707_, _07706_, _07702_);
  nor _16042_ (_07708_, _07707_, _07699_);
  and _16043_ (_07709_, _07708_, _07695_);
  and _16044_ (_07710_, _07709_, _07684_);
  nand _16045_ (_07711_, _07710_, _07678_);
  or _16046_ (_07712_, _07711_, _07668_);
  or _16047_ (_07713_, _07670_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and _16048_ (_07714_, _07713_, _05552_);
  and _16049_ (_05929_, _07714_, _07712_);
  or _16050_ (_07715_, _07668_, _07574_);
  or _16051_ (_07716_, _07670_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and _16052_ (_07717_, _07716_, _05552_);
  and _16053_ (_05932_, _07717_, _07715_);
  and _16054_ (_06005_, _06402_, _05552_);
  or _16055_ (_07718_, _06472_, _06464_);
  and _16056_ (_07719_, _07718_, _06473_);
  and _16057_ (_06007_, _07719_, _05552_);
  and _16058_ (_06013_, _07510_, _05552_);
  and _16059_ (_07720_, _06458_, _06456_);
  not _16060_ (_07721_, _07720_);
  and _16061_ (_07722_, _07721_, _06459_);
  and _16062_ (_06017_, _07722_, _05552_);
  and _16063_ (_07723_, _06366_, _06368_);
  not _16064_ (_07724_, _07723_);
  and _16065_ (_07725_, _07724_, _06411_);
  nor _16066_ (_07726_, _07725_, _06403_);
  and _16067_ (_06036_, _07726_, _05552_);
  and _16068_ (_07727_, _05552_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  and _16069_ (_07728_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _05552_);
  and _16070_ (_07729_, _07728_, _05917_);
  or _16071_ (_06264_, _07729_, _07727_);
  nor _16072_ (_07730_, _05575_, _05562_);
  or _16073_ (_07731_, _07730_, _05556_);
  and _16074_ (_07732_, _07731_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  and _16075_ (_07733_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  nor _16076_ (_07734_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  nor _16077_ (_07735_, _07734_, _07733_);
  and _16078_ (_07736_, _05562_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and _16079_ (_07737_, _07736_, _07735_);
  or _16080_ (_07738_, _07737_, _07732_);
  and _16081_ (_06338_, _07738_, _05552_);
  and _16082_ (_07740_, _05585_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  or _16083_ (_06460_, _07740_, _05558_);
  nor _16084_ (_07741_, _05547_, _06584_);
  and _16085_ (_07742_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  not _16086_ (_07743_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nor _16087_ (_07744_, _05616_, _07743_);
  nor _16088_ (_07745_, _05624_, _05768_);
  or _16089_ (_07746_, _07745_, _07744_);
  and _16090_ (_07747_, _05725_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  nor _16091_ (_07748_, _05631_, _05762_);
  or _16092_ (_07749_, _07748_, _07747_);
  or _16093_ (_07750_, _07749_, _07746_);
  and _16094_ (_07751_, _05619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and _16095_ (_07752_, _05627_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  or _16096_ (_07753_, _07752_, _07751_);
  or _16097_ (_07754_, _07753_, _07750_);
  and _16098_ (_07755_, _07754_, _05671_);
  or _16099_ (_07756_, _07755_, _07742_);
  and _16100_ (_07757_, _07756_, _05547_);
  nor _16101_ (_07758_, _07757_, _07741_);
  nor _16102_ (_06468_, _07758_, rst);
  and _16103_ (_07759_, _05777_, _05729_);
  and _16104_ (_07760_, _05799_, _05752_);
  and _16105_ (_07761_, _07760_, _07759_);
  nor _16106_ (_07762_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , rst);
  and _16107_ (_07763_, _07762_, _05608_);
  and _16108_ (_07764_, _07763_, _05706_);
  and _16109_ (_07765_, _05660_, _05636_);
  and _16110_ (_07766_, _07765_, _07764_);
  and _16111_ (_07767_, _07766_, _05685_);
  and _16112_ (_06484_, _07767_, _07761_);
  and _16113_ (_06548_, _07316_, _05552_);
  not _16114_ (_07768_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  and _16115_ (_07769_, \oc8051_top_1.oc8051_memory_interface1.cdata [7], _07768_);
  and _16116_ (_07770_, \oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or _16117_ (_07771_, _07770_, _07769_);
  and _16118_ (_06592_, _07771_, _05552_);
  nor _16119_ (_07772_, _05710_, _05689_);
  not _16120_ (_07773_, _05665_);
  nor _16121_ (_07774_, _07773_, _05641_);
  and _16122_ (_07775_, _07774_, _07772_);
  not _16123_ (_07776_, _05781_);
  and _16124_ (_07777_, _05803_, _07776_);
  and _16125_ (_07778_, _05756_, _05733_);
  and _16126_ (_07779_, _07778_, _07777_);
  and _16127_ (_07780_, _07779_, _07775_);
  not _16128_ (_07781_, _05756_);
  and _16129_ (_07782_, _07781_, _05733_);
  nor _16130_ (_07783_, _05803_, _05781_);
  and _16131_ (_07784_, _07783_, _07782_);
  and _16132_ (_07785_, _07784_, _07775_);
  nor _16133_ (_07786_, _07785_, _07780_);
  not _16134_ (_07787_, _05803_);
  and _16135_ (_07788_, _07787_, _05781_);
  and _16136_ (_07789_, _05689_, _05641_);
  nor _16137_ (_07790_, _05733_, _05710_);
  and _16138_ (_07791_, _07790_, _07789_);
  and _16139_ (_07792_, _07791_, _07788_);
  not _16140_ (_07793_, _07792_);
  nor _16141_ (_07794_, _07781_, _05733_);
  and _16142_ (_07795_, _07794_, _07788_);
  and _16143_ (_07796_, _07795_, _05710_);
  nor _16144_ (_07797_, _05665_, _05641_);
  and _16145_ (_07798_, _07797_, _07772_);
  nor _16146_ (_07799_, _07798_, _07796_);
  and _16147_ (_07800_, _07799_, _07793_);
  and _16148_ (_07801_, _07800_, _07786_);
  nor _16149_ (_07802_, _05710_, _07773_);
  not _16150_ (_07803_, _05689_);
  nor _16151_ (_07804_, _07803_, _05641_);
  and _16152_ (_07805_, _07804_, _07802_);
  not _16153_ (_07806_, _07805_);
  and _16154_ (_07807_, _07782_, _07777_);
  not _16155_ (_07808_, _07807_);
  and _16156_ (_07809_, _07788_, _07778_);
  and _16157_ (_07810_, _07783_, _07781_);
  nor _16158_ (_07811_, _07810_, _07809_);
  and _16159_ (_07812_, _07811_, _07808_);
  nor _16160_ (_07813_, _07812_, _07806_);
  not _16161_ (_07814_, _05710_);
  and _16162_ (_07815_, _07804_, _07814_);
  and _16163_ (_07816_, _07815_, _07773_);
  not _16164_ (_07817_, _07816_);
  nor _16165_ (_07818_, _05756_, _05733_);
  and _16166_ (_07819_, _05803_, _05781_);
  and _16167_ (_07820_, _07819_, _07818_);
  and _16168_ (_07821_, _07783_, _05756_);
  nor _16169_ (_07823_, _07821_, _07820_);
  nor _16170_ (_07824_, _07823_, _07817_);
  nor _16171_ (_07825_, _07824_, _07813_);
  and _16172_ (_07826_, _07825_, _07801_);
  and _16173_ (_07827_, _07819_, _07782_);
  and _16174_ (_07828_, _07827_, _07816_);
  not _16175_ (_07830_, _07828_);
  and _16176_ (_07831_, _07803_, _05641_);
  nor _16177_ (_07832_, _07831_, _07804_);
  not _16178_ (_07833_, _07832_);
  and _16179_ (_07834_, _07777_, _07781_);
  and _16180_ (_07835_, _07834_, _07790_);
  and _16181_ (_07836_, _07835_, _07833_);
  and _16182_ (_07837_, _07816_, _07810_);
  nor _16183_ (_07838_, _07837_, _07836_);
  and _16184_ (_07839_, _07838_, _07830_);
  and _16185_ (_07840_, _07795_, _07775_);
  and _16186_ (_07841_, _05733_, _07814_);
  and _16187_ (_07842_, _07841_, _07789_);
  nor _16188_ (_07843_, _05803_, _05756_);
  and _16189_ (_07844_, _07843_, _05781_);
  or _16190_ (_07845_, _07834_, _07844_);
  and _16191_ (_07846_, _07845_, _07842_);
  nor _16192_ (_07847_, _07846_, _07840_);
  and _16193_ (_07848_, _07788_, _07782_);
  and _16194_ (_07849_, _07848_, _07775_);
  not _16195_ (_07850_, _07775_);
  and _16196_ (_07851_, _07794_, _07777_);
  nor _16197_ (_07852_, _07851_, _07834_);
  nor _16198_ (_07853_, _07852_, _07850_);
  nor _16199_ (_07854_, _07853_, _07849_);
  and _16200_ (_07855_, _07854_, _07847_);
  and _16201_ (_07856_, _07855_, _07839_);
  and _16202_ (_07857_, _07856_, _07826_);
  nor _16203_ (_07859_, _07794_, _07782_);
  and _16204_ (_07860_, _07859_, _07783_);
  and _16205_ (_07861_, _07860_, _07775_);
  and _16206_ (_07862_, _07819_, _07778_);
  and _16207_ (_07863_, _07862_, _07816_);
  nor _16208_ (_07864_, _07863_, _07861_);
  and _16209_ (_07865_, _07831_, _07802_);
  and _16210_ (_07866_, _07865_, _07821_);
  not _16211_ (_07867_, _07866_);
  or _16212_ (_07868_, _07807_, _07795_);
  and _16213_ (_07869_, _07868_, _07816_);
  and _16214_ (_07870_, _07848_, _07805_);
  nor _16215_ (_07871_, _07870_, _07869_);
  and _16216_ (_07872_, _07871_, _07867_);
  and _16217_ (_07873_, _07872_, _07864_);
  not _16218_ (_07874_, _07865_);
  and _16219_ (_07875_, _07819_, _07794_);
  nor _16220_ (_07876_, _07875_, _07848_);
  nor _16221_ (_07877_, _07876_, _07874_);
  and _16222_ (_07878_, _05803_, _05756_);
  and _16223_ (_07879_, _07878_, _05781_);
  and _16224_ (_07880_, _07818_, _07788_);
  nor _16225_ (_07881_, _07880_, _07879_);
  nor _16226_ (_07882_, _07881_, _07850_);
  nor _16227_ (_07883_, _07882_, _07877_);
  nor _16228_ (_07884_, _07875_, _07809_);
  nor _16229_ (_07885_, _07884_, _07817_);
  nor _16230_ (_07886_, _07862_, _07807_);
  nor _16231_ (_07887_, _07886_, _07874_);
  nor _16232_ (_07888_, _07887_, _07885_);
  and _16233_ (_07889_, _07888_, _07883_);
  and _16234_ (_07890_, _07889_, _07873_);
  and _16235_ (_07891_, _07890_, _07857_);
  and _16236_ (_07892_, _07833_, _07802_);
  nor _16237_ (_07893_, _07892_, _07816_);
  not _16238_ (_07894_, _07893_);
  and _16239_ (_07895_, _07894_, _07851_);
  not _16240_ (_07896_, _07895_);
  and _16241_ (_07897_, _07831_, _07814_);
  and _16242_ (_07898_, _07897_, _07773_);
  and _16243_ (_07899_, _07851_, _07898_);
  and _16244_ (_07900_, _07809_, _07775_);
  nor _16245_ (_07901_, _07900_, _07899_);
  not _16246_ (_07902_, _07901_);
  and _16247_ (_07903_, _07848_, _07816_);
  and _16248_ (_07904_, _07898_, _07779_);
  or _16249_ (_07905_, _07904_, _07903_);
  nor _16250_ (_07906_, _07905_, _07902_);
  and _16251_ (_07907_, _07906_, _07896_);
  and _16252_ (_07908_, _07865_, _07788_);
  and _16253_ (_07909_, _07908_, _07859_);
  and _16254_ (_07910_, _07908_, _07794_);
  nor _16255_ (_07911_, _07910_, _07909_);
  not _16256_ (_07912_, _07844_);
  and _16257_ (_07913_, _07886_, _07912_);
  nor _16258_ (_07914_, _07913_, _07814_);
  and _16259_ (_07915_, _07894_, _07779_);
  nor _16260_ (_07916_, _07915_, _07914_);
  and _16261_ (_07917_, _07916_, _07911_);
  and _16262_ (_07918_, _07917_, _07907_);
  and _16263_ (_07919_, _07918_, _07891_);
  and _16264_ (_07920_, _07818_, _07777_);
  and _16265_ (_07921_, _07920_, _07898_);
  or _16266_ (_07922_, _07789_, _05710_);
  and _16267_ (_07923_, _07922_, _07848_);
  or _16268_ (_07924_, _07923_, _07785_);
  nor _16269_ (_07925_, _07924_, _07921_);
  nand _16270_ (_07926_, _07925_, _07901_);
  nor _16271_ (_07928_, _07926_, _07905_);
  nand _16272_ (_07929_, _07928_, _07873_);
  nor _16273_ (_07930_, _07929_, _07919_);
  nor _16274_ (_07931_, _07930_, _05548_);
  nand _16275_ (_07932_, _07931_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor _16276_ (_07933_, rst, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _16277_ (_07934_, _07931_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _16278_ (_07935_, _07934_, _07933_);
  and _16279_ (_06607_, _07935_, _07932_);
  and _16280_ (_07936_, _06528_, _05972_);
  and _16281_ (_07937_, _07936_, _06057_);
  and _16282_ (_07938_, _07937_, _06068_);
  not _16283_ (_07939_, _07938_);
  and _16284_ (_07940_, _07939_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  nor _16285_ (_07941_, _06206_, _06133_);
  not _16286_ (_07942_, _07941_);
  and _16287_ (_07943_, _07942_, _07690_);
  and _16288_ (_07944_, _07943_, _07687_);
  and _16289_ (_07945_, _07944_, _07702_);
  nor _16290_ (_07946_, _07945_, _06955_);
  and _16291_ (_07947_, _07946_, _07937_);
  or _16292_ (_07948_, _07947_, _07940_);
  and _16293_ (_06610_, _07948_, _05552_);
  and _16294_ (_07949_, _07936_, _06061_);
  and _16295_ (_07950_, _07949_, _06068_);
  not _16296_ (_07951_, _07950_);
  and _16297_ (_07952_, _07951_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  and _16298_ (_07953_, _06635_, _06295_);
  and _16299_ (_07954_, _06206_, _06254_);
  nor _16300_ (_07955_, _06255_, _07954_);
  and _16301_ (_07956_, _07955_, _06253_);
  nor _16302_ (_07957_, _07955_, _06253_);
  or _16303_ (_07958_, _07957_, _07956_);
  and _16304_ (_07959_, _07958_, _06266_);
  nor _16305_ (_07960_, _07959_, _07953_);
  nor _16306_ (_07961_, _06254_, _06133_);
  not _16307_ (_07962_, _07961_);
  and _16308_ (_07963_, _06638_, _06300_);
  not _16309_ (_07964_, _07963_);
  nor _16310_ (_07965_, _06637_, _06283_);
  not _16311_ (_07966_, _07965_);
  and _16312_ (_07967_, _06636_, _06288_);
  nor _16313_ (_07969_, _06291_, _06248_);
  nor _16314_ (_07970_, _07969_, _07967_);
  and _16315_ (_07971_, _07970_, _07966_);
  and _16316_ (_07972_, _07971_, _07964_);
  and _16317_ (_07974_, _07972_, _07962_);
  and _16318_ (_07975_, _07974_, _07960_);
  nor _16319_ (_07976_, _07975_, _06955_);
  and _16320_ (_07977_, _07976_, _07949_);
  or _16321_ (_07978_, _07977_, _07952_);
  and _16322_ (_06623_, _07978_, _05552_);
  and _16323_ (_06691_, \oc8051_top_1.oc8051_memory_interface1.istb_t , _05552_);
  and _16324_ (_06780_, _05781_, _05552_);
  or _16325_ (_07979_, _06674_, _06672_);
  not _16326_ (_07980_, _06601_);
  nand _16327_ (_07981_, _06672_, _07980_);
  and _16328_ (_07982_, _07981_, _06581_);
  and _16329_ (_07983_, _07982_, _07979_);
  nand _16330_ (_07984_, _06710_, _06679_);
  and _16331_ (_07985_, _06711_, _06677_);
  and _16332_ (_07986_, _07985_, _07984_);
  and _16333_ (_07987_, _06379_, _06340_);
  and _16334_ (_07988_, _07987_, _07088_);
  and _16335_ (_07989_, _07988_, _07329_);
  nand _16336_ (_07990_, _07989_, _06314_);
  nand _16337_ (_07991_, _07990_, \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or _16338_ (_07992_, _07991_, _07986_);
  or _16339_ (_07993_, _07992_, _07983_);
  nand _16340_ (_07994_, _06888_, _06861_);
  and _16341_ (_07995_, _07994_, _06889_);
  or _16342_ (_07996_, _07995_, _07698_);
  or _16343_ (_07997_, _06890_, _06868_);
  and _16344_ (_07998_, _07997_, _06891_);
  or _16345_ (_07999_, _07998_, _07996_);
  or _16346_ (_08000_, _07999_, _06895_);
  or _16347_ (_08001_, _08000_, _06908_);
  or _16348_ (_08002_, _07525_, _06905_);
  or _16349_ (_08003_, _08002_, _07218_);
  or _16350_ (_08004_, _08003_, _08001_);
  and _16351_ (_08005_, _08004_, _07211_);
  or _16352_ (_08006_, _08005_, _07993_);
  nor _16353_ (_08007_, _06764_, _05958_);
  and _16354_ (_08008_, _08007_, _06775_);
  and _16355_ (_08009_, _08008_, _06915_);
  nor _16356_ (_08010_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  nor _16357_ (_08011_, _08010_, _08009_);
  and _16358_ (_08012_, _08011_, _08006_);
  and _16359_ (_08013_, _07666_, _06054_);
  not _16360_ (_08014_, _08013_);
  nor _16361_ (_08015_, _08014_, _06763_);
  and _16362_ (_08016_, _08014_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or _16363_ (_08017_, _08016_, _08015_);
  and _16364_ (_08018_, _08017_, _08009_);
  or _16365_ (_08019_, _08018_, _06531_);
  or _16366_ (_08020_, _08019_, _08012_);
  nor _16367_ (_08021_, _06255_, _06142_);
  nor _16368_ (_08022_, _07954_, _06253_);
  nor _16369_ (_08023_, _08022_, _08021_);
  nor _16370_ (_08024_, _08023_, _06227_);
  and _16371_ (_08025_, _08023_, _06227_);
  nor _16372_ (_08026_, _08025_, _08024_);
  and _16373_ (_08027_, _08026_, _06266_);
  and _16374_ (_08028_, _06631_, _06295_);
  nor _16375_ (_08029_, _08028_, _08027_);
  and _16376_ (_08030_, _06632_, _06288_);
  nor _16377_ (_08031_, _06291_, _06227_);
  nor _16378_ (_08033_, _08031_, _08030_);
  not _16379_ (_08034_, _06227_);
  nor _16380_ (_08035_, _08034_, _06133_);
  and _16381_ (_08036_, _06634_, _06300_);
  nor _16382_ (_08037_, _06633_, _06283_);
  or _16383_ (_08038_, _08037_, _08036_);
  nor _16384_ (_08039_, _08038_, _08035_);
  and _16385_ (_08040_, _08039_, _08033_);
  and _16386_ (_08041_, _08040_, _08029_);
  nand _16387_ (_08042_, _08041_, _06531_);
  and _16388_ (_08043_, _08042_, _05552_);
  and _16389_ (_06894_, _08043_, _08020_);
  not _16390_ (_08044_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and _16391_ (_08045_, _08009_, _06056_);
  nor _16392_ (_08046_, _08045_, _08044_);
  or _16393_ (_08047_, _08046_, _06531_);
  not _16394_ (_08048_, _06763_);
  and _16395_ (_08049_, _08045_, _08048_);
  or _16396_ (_08050_, _08049_, _08047_);
  nand _16397_ (_08051_, _07975_, _06531_);
  and _16398_ (_08052_, _08051_, _05552_);
  and _16399_ (_06900_, _08052_, _08050_);
  nor _16400_ (_06907_, _05665_, rst);
  and _16401_ (_06909_, _05641_, _05552_);
  and _16402_ (_06912_, _05689_, _05552_);
  and _16403_ (_06914_, _05710_, _05552_);
  and _16404_ (_06917_, _05733_, _05552_);
  nor _16405_ (_06920_, _05756_, rst);
  and _16406_ (_06923_, _05803_, _05552_);
  nand _16407_ (_08053_, _07975_, _06949_);
  or _16408_ (_08054_, _06949_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  and _16409_ (_08055_, _08054_, _08053_);
  and _16410_ (_06961_, _08055_, _05552_);
  not _16411_ (_08056_, _08009_);
  and _16412_ (_08057_, _06059_, _06769_);
  nor _16413_ (_08058_, _06059_, _06769_);
  nor _16414_ (_08059_, _08058_, _08057_);
  or _16415_ (_08060_, _08059_, _08056_);
  and _16416_ (_08061_, _08060_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and _16417_ (_08062_, _08057_, _08048_);
  and _16418_ (_08063_, _08058_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  or _16419_ (_08064_, _08063_, _08062_);
  and _16420_ (_08065_, _08064_, _08009_);
  or _16421_ (_08066_, _08065_, _08061_);
  and _16422_ (_08067_, _08066_, _06532_);
  or _16423_ (_08068_, _08067_, _07389_);
  and _16424_ (_06964_, _08068_, _05552_);
  or _16425_ (_08069_, _07159_, _07154_);
  and _16426_ (_08070_, _08069_, _07160_);
  or _16427_ (_08071_, _08070_, _07446_);
  or _16428_ (_08072_, _07200_, _07151_);
  and _16429_ (_08073_, _08072_, _08071_);
  nand _16430_ (_08074_, _08073_, _06314_);
  nand _16431_ (_08075_, _07995_, _07211_);
  nor _16432_ (_08076_, _06659_, _06655_);
  nor _16433_ (_08077_, _08076_, _06660_);
  nor _16434_ (_08078_, _08077_, _06582_);
  not _16435_ (_08079_, _08078_);
  nand _16436_ (_08080_, _06227_, _06128_);
  and _16437_ (_08081_, _06368_, _06131_);
  and _16438_ (_08082_, _06248_, _06118_);
  nor _16439_ (_08083_, _08082_, _08081_);
  and _16440_ (_08084_, _08083_, _08080_);
  and _16441_ (_08085_, _08084_, _07972_);
  and _16442_ (_08086_, _08085_, _07960_);
  nor _16443_ (_08087_, _06717_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and _16444_ (_08088_, _08087_, _06248_);
  nor _16445_ (_08089_, _08087_, _06248_);
  nor _16446_ (_08090_, _08089_, _08088_);
  nor _16447_ (_08091_, _08090_, _06724_);
  nor _16448_ (_08092_, _06656_, _06638_);
  or _16449_ (_08093_, _08092_, _06681_);
  and _16450_ (_08094_, _08093_, _06688_);
  nor _16451_ (_08095_, _08093_, _06688_);
  or _16452_ (_08096_, _08095_, _08094_);
  and _16453_ (_08097_, _08096_, _06677_);
  nor _16454_ (_08098_, _08097_, _08091_);
  and _16455_ (_08099_, _08098_, _08086_);
  and _16456_ (_08100_, _08099_, _08079_);
  and _16457_ (_08101_, _08100_, _08075_);
  nand _16458_ (_08102_, _08101_, _08074_);
  or _16459_ (_08103_, _08102_, _07668_);
  or _16460_ (_08104_, _07670_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and _16461_ (_08105_, _08104_, _05552_);
  and _16462_ (_07080_, _08105_, _08103_);
  and _16463_ (_08106_, _05917_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  or _16464_ (_08107_, _08106_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  and _16465_ (_07083_, _08107_, _05552_);
  and _16466_ (_08108_, _07170_, _07161_);
  not _16467_ (_08109_, _08108_);
  and _16468_ (_08110_, _08109_, _07171_);
  or _16469_ (_08111_, _08110_, _07446_);
  or _16470_ (_08112_, _07200_, _07167_);
  and _16471_ (_08113_, _08112_, _08111_);
  nand _16472_ (_08114_, _08113_, _06314_);
  nand _16473_ (_08115_, _07998_, _07211_);
  nor _16474_ (_08116_, _06660_, _06652_);
  nor _16475_ (_08117_, _08116_, _06661_);
  nor _16476_ (_08118_, _08117_, _06582_);
  not _16477_ (_08120_, _08118_);
  nor _16478_ (_08121_, _06692_, _06689_);
  not _16479_ (_08122_, _08121_);
  nor _16480_ (_08123_, _06693_, _06678_);
  and _16481_ (_08124_, _08123_, _08122_);
  not _16482_ (_08125_, _08124_);
  and _16483_ (_08126_, _06249_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor _16484_ (_08127_, _08089_, _08034_);
  nor _16485_ (_08128_, _08127_, _08126_);
  nor _16486_ (_08129_, _08128_, _06724_);
  nor _16487_ (_08130_, _08129_, _08038_);
  nand _16488_ (_08131_, _06184_, _06128_);
  and _16489_ (_08132_, _06248_, _06131_);
  not _16490_ (_08133_, _08132_);
  and _16491_ (_08134_, _08133_, _08131_);
  and _16492_ (_08135_, _06227_, _06118_);
  not _16493_ (_08136_, _08135_);
  and _16494_ (_08137_, _08136_, _08033_);
  and _16495_ (_08138_, _08137_, _08134_);
  and _16496_ (_08139_, _08138_, _08029_);
  and _16497_ (_08140_, _08139_, _08130_);
  and _16498_ (_08141_, _08140_, _08125_);
  and _16499_ (_08142_, _08141_, _08120_);
  and _16500_ (_08143_, _08142_, _08115_);
  nand _16501_ (_08144_, _08143_, _08114_);
  or _16502_ (_08145_, _08144_, _07668_);
  or _16503_ (_08146_, _07670_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and _16504_ (_08147_, _08146_, _05552_);
  and _16505_ (_07085_, _08147_, _08145_);
  and _16506_ (_08148_, _08102_, _07445_);
  and _16507_ (_08149_, _07486_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or _16508_ (_08150_, _08149_, _07485_);
  or _16509_ (_08151_, _08150_, _08148_);
  and _16510_ (_08152_, _06635_, _06118_);
  and _16511_ (_08153_, _06746_, _06111_);
  and _16512_ (_08154_, _07326_, _06386_);
  nor _16513_ (_08155_, _08154_, _06253_);
  nor _16514_ (_08156_, _07319_, _06142_);
  nor _16515_ (_08157_, _08156_, _08155_);
  nor _16516_ (_08158_, _08157_, _06635_);
  and _16517_ (_08159_, _08157_, _06635_);
  or _16518_ (_08160_, _08159_, _06267_);
  nor _16519_ (_08161_, _08160_, _08158_);
  and _16520_ (_08162_, _06295_, _06248_);
  or _16521_ (_08163_, _08162_, _08161_);
  or _16522_ (_08164_, _08163_, _08153_);
  and _16523_ (_08165_, _07117_, _06314_);
  nor _16524_ (_08166_, _07290_, _07286_);
  nor _16525_ (_08167_, _08166_, _07291_);
  and _16526_ (_08168_, _08167_, _06677_);
  and _16527_ (_08169_, _07726_, _07211_);
  or _16528_ (_08170_, _08169_, _08168_);
  or _16529_ (_08171_, _08170_, _08165_);
  or _16530_ (_08172_, _08171_, _08164_);
  nor _16531_ (_08173_, _08172_, _08152_);
  nand _16532_ (_08174_, _08173_, _07485_);
  and _16533_ (_08175_, _08174_, _05552_);
  and _16534_ (_07107_, _08175_, _08151_);
  and _16535_ (_08176_, _08144_, _07445_);
  and _16536_ (_08177_, _07486_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or _16537_ (_08178_, _08177_, _07485_);
  or _16538_ (_08179_, _08178_, _08176_);
  and _16539_ (_08180_, _06631_, _06118_);
  and _16540_ (_08181_, _06500_, _06746_);
  nor _16541_ (_08182_, _07492_, _06253_);
  nor _16542_ (_08183_, _07320_, _06142_);
  nor _16543_ (_08184_, _08183_, _08182_);
  and _16544_ (_08185_, _08184_, _06373_);
  nor _16545_ (_08186_, _08184_, _06373_);
  nor _16546_ (_08187_, _08186_, _08185_);
  nor _16547_ (_08188_, _08187_, _06267_);
  and _16548_ (_08189_, _06295_, _06227_);
  or _16549_ (_08190_, _08189_, _08188_);
  or _16550_ (_08191_, _08190_, _08181_);
  and _16551_ (_08192_, _06314_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  nor _16552_ (_08193_, _07294_, _07291_);
  nor _16553_ (_08194_, _08193_, _07295_);
  and _16554_ (_08195_, _08194_, _06677_);
  and _16555_ (_08196_, _07722_, _07211_);
  or _16556_ (_08197_, _08196_, _08195_);
  or _16557_ (_08198_, _08197_, _08192_);
  or _16558_ (_08199_, _08198_, _08191_);
  nor _16559_ (_08200_, _08199_, _08180_);
  nand _16560_ (_08201_, _08200_, _07485_);
  and _16561_ (_08202_, _08201_, _05552_);
  and _16562_ (_07109_, _08202_, _08179_);
  and _16563_ (_08203_, _07711_, _07445_);
  and _16564_ (_08204_, _07486_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or _16565_ (_08205_, _08204_, _07485_);
  or _16566_ (_08206_, _08205_, _08203_);
  and _16567_ (_08207_, _07285_, _06712_);
  nor _16568_ (_08208_, _08207_, _07286_);
  and _16569_ (_08209_, _08208_, _06677_);
  nand _16570_ (_08210_, _07200_, _06314_);
  nor _16571_ (_08211_, _06783_, _06725_);
  not _16572_ (_08212_, _08211_);
  nor _16573_ (_08213_, _08212_, _06795_);
  nor _16574_ (_08214_, _08213_, _06639_);
  and _16575_ (_08215_, _08213_, _06639_);
  nor _16576_ (_08216_, _08215_, _08214_);
  and _16577_ (_08217_, _08216_, _06266_);
  and _16578_ (_08218_, _06639_, _06118_);
  and _16579_ (_08219_, _06402_, _07211_);
  and _16580_ (_08220_, _06162_, _06746_);
  nor _16581_ (_08221_, _06785_, _06206_);
  or _16582_ (_08222_, _08221_, _08220_);
  or _16583_ (_08223_, _08222_, _08219_);
  nor _16584_ (_08224_, _08223_, _08218_);
  not _16585_ (_08225_, _08224_);
  nor _16586_ (_08226_, _08225_, _08217_);
  nand _16587_ (_08227_, _08226_, _08210_);
  or _16588_ (_08228_, _08227_, _08209_);
  or _16589_ (_08229_, _08228_, _07579_);
  and _16590_ (_08230_, _08229_, _05552_);
  and _16591_ (_07113_, _08230_, _08206_);
  nor _16592_ (_08232_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor _16593_ (_08233_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _07768_);
  nor _16594_ (_08234_, _08233_, _08232_);
  not _16595_ (_08235_, \oc8051_symbolic_cxrom1.regvalid [5]);
  not _16596_ (_08236_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor _16597_ (_08237_, _05550_, _08236_);
  and _16598_ (_08238_, _08237_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor _16599_ (_08239_, _08237_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor _16600_ (_08240_, _08239_, _08238_);
  nor _16601_ (_08241_, _08240_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor _16602_ (_08242_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _07768_);
  nor _16603_ (_08243_, _08242_, _08241_);
  nor _16604_ (_08244_, _08243_, _08235_);
  and _16605_ (_08245_, _08243_, \oc8051_symbolic_cxrom1.regvalid [13]);
  nor _16606_ (_08246_, _08245_, _08244_);
  not _16607_ (_08247_, _08246_);
  nor _16608_ (_08248_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor _16609_ (_08249_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _07768_);
  nor _16610_ (_08250_, _08249_, _08248_);
  not _16611_ (_08251_, _08250_);
  and _16612_ (_08252_, _05550_, _08236_);
  nor _16613_ (_08253_, _08252_, _08237_);
  nor _16614_ (_08254_, _08253_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor _16615_ (_08255_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _07768_);
  nor _16616_ (_08256_, _08255_, _08254_);
  and _16617_ (_08257_, _08256_, _08251_);
  nand _16618_ (_08258_, _08257_, _08247_);
  and _16619_ (_08259_, _08258_, _08234_);
  nor _16620_ (_08260_, _08256_, _08251_);
  not _16621_ (_08261_, _08260_);
  not _16622_ (_08262_, \oc8051_symbolic_cxrom1.regvalid [3]);
  nor _16623_ (_08263_, _08243_, _08262_);
  and _16624_ (_08264_, _08243_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor _16625_ (_08265_, _08264_, _08263_);
  nor _16626_ (_08266_, _08265_, _08261_);
  and _16627_ (_08267_, _08256_, _08250_);
  not _16628_ (_08268_, _08267_);
  nor _16629_ (_08269_, _08243_, \oc8051_symbolic_cxrom1.regvalid [7]);
  not _16630_ (_08270_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and _16631_ (_08271_, _08243_, _08270_);
  or _16632_ (_08272_, _08271_, _08269_);
  nor _16633_ (_08273_, _08272_, _08268_);
  nor _16634_ (_08274_, _08273_, _08266_);
  and _16635_ (_08275_, _08243_, \oc8051_symbolic_cxrom1.regvalid [9]);
  not _16636_ (_08276_, \oc8051_symbolic_cxrom1.regvalid [1]);
  nor _16637_ (_08277_, _08243_, _08276_);
  nor _16638_ (_08278_, _08277_, _08275_);
  nor _16639_ (_08279_, _08256_, _08250_);
  not _16640_ (_08280_, _08279_);
  or _16641_ (_08281_, _08280_, _08278_);
  and _16642_ (_08282_, _08281_, _08274_);
  and _16643_ (_08283_, _08282_, _08259_);
  and _16644_ (_08284_, _08243_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and _16645_ (_08285_, _08284_, _08260_);
  not _16646_ (_08286_, _08243_);
  and _16647_ (_08288_, _08260_, _08286_);
  and _16648_ (_08289_, _08288_, \oc8051_symbolic_cxrom1.regvalid [2]);
  or _16649_ (_08290_, _08289_, _08234_);
  or _16650_ (_08291_, _08290_, _08285_);
  and _16651_ (_08292_, _08243_, \oc8051_symbolic_cxrom1.regvalid [8]);
  not _16652_ (_08293_, \oc8051_symbolic_cxrom1.regvalid [0]);
  nor _16653_ (_08294_, _08243_, _08293_);
  nor _16654_ (_08295_, _08294_, _08292_);
  nor _16655_ (_08296_, _08295_, _08280_);
  nor _16656_ (_08297_, _08243_, \oc8051_symbolic_cxrom1.regvalid [6]);
  not _16657_ (_08298_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and _16658_ (_08299_, _08243_, _08298_);
  or _16659_ (_08300_, _08299_, _08297_);
  nor _16660_ (_08301_, _08300_, _08268_);
  not _16661_ (_08302_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and _16662_ (_08303_, _08243_, _08302_);
  nor _16663_ (_08304_, _08243_, \oc8051_symbolic_cxrom1.regvalid [4]);
  or _16664_ (_08305_, _08304_, _08303_);
  not _16665_ (_08306_, _08305_);
  and _16666_ (_08307_, _08306_, _08257_);
  or _16667_ (_08308_, _08307_, _08301_);
  or _16668_ (_08309_, _08308_, _08296_);
  nor _16669_ (_08310_, _08309_, _08291_);
  nor _16670_ (_08311_, _08310_, _08283_);
  not _16671_ (_08312_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  nand _16672_ (_08313_, _08234_, _08312_);
  or _16673_ (_08314_, _08234_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  and _16674_ (_08315_, _08314_, _08313_);
  and _16675_ (_08316_, _08315_, _08267_);
  not _16676_ (_08317_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  nand _16677_ (_08318_, _08234_, _08317_);
  or _16678_ (_08319_, _08234_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  and _16679_ (_08320_, _08319_, _08318_);
  and _16680_ (_08321_, _08320_, _08260_);
  or _16681_ (_08322_, _08321_, _08316_);
  not _16682_ (_08323_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  nand _16683_ (_08324_, _08234_, _08323_);
  or _16684_ (_08325_, _08234_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  and _16685_ (_08326_, _08325_, _08324_);
  and _16686_ (_08327_, _08326_, _08257_);
  not _16687_ (_08328_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  nand _16688_ (_08329_, _08234_, _08328_);
  or _16689_ (_08330_, _08234_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  and _16690_ (_08331_, _08330_, _08329_);
  and _16691_ (_08332_, _08331_, _08279_);
  or _16692_ (_08333_, _08332_, _08327_);
  or _16693_ (_08334_, _08333_, _08322_);
  and _16694_ (_08335_, _08334_, _08243_);
  not _16695_ (_08336_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  nand _16696_ (_08337_, _08234_, _08336_);
  or _16697_ (_08338_, _08234_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  and _16698_ (_08339_, _08338_, _08337_);
  and _16699_ (_08340_, _08339_, _08260_);
  not _16700_ (_08341_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  nand _16701_ (_08342_, _08234_, _08341_);
  or _16702_ (_08343_, _08234_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  and _16703_ (_08344_, _08343_, _08342_);
  and _16704_ (_08345_, _08344_, _08267_);
  or _16705_ (_08346_, _08345_, _08340_);
  not _16706_ (_08347_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  nand _16707_ (_08348_, _08234_, _08347_);
  or _16708_ (_08349_, _08234_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  and _16709_ (_08350_, _08349_, _08348_);
  and _16710_ (_08351_, _08350_, _08257_);
  not _16711_ (_08352_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  nand _16712_ (_08353_, _08234_, _08352_);
  or _16713_ (_08354_, _08234_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  and _16714_ (_08355_, _08354_, _08353_);
  and _16715_ (_08356_, _08355_, _08279_);
  or _16716_ (_08357_, _08356_, _08351_);
  or _16717_ (_08358_, _08357_, _08346_);
  and _16718_ (_08359_, _08358_, _08286_);
  or _16719_ (_08360_, _08359_, _08335_);
  and _16720_ (_08361_, _08360_, _08311_);
  not _16721_ (_08362_, _08311_);
  and _16722_ (_08363_, _08362_, word_in[7]);
  or _16723_ (\oc8051_symbolic_cxrom1.cxrom_data_out [7], _08363_, _08361_);
  nor _16724_ (_08364_, _06054_, _06043_);
  and _16725_ (_08365_, _08364_, _06030_);
  not _16726_ (_08366_, _08365_);
  nor _16727_ (_08367_, _08366_, _06763_);
  or _16728_ (_08368_, _08365_, _07468_);
  nand _16729_ (_08369_, _08368_, _08009_);
  or _16730_ (_08370_, _08369_, _08367_);
  and _16731_ (_08371_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  or _16732_ (_08372_, _08371_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and _16733_ (_08373_, _06668_, _06581_);
  and _16734_ (_08374_, _06698_, _06677_);
  nand _16735_ (_08375_, _06118_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nand _16736_ (_08376_, _08375_, _08371_);
  or _16737_ (_08377_, _08376_, _08374_);
  or _16738_ (_08378_, _08377_, _08373_);
  and _16739_ (_08379_, _08378_, _08372_);
  or _16740_ (_08380_, _08379_, _08009_);
  and _16741_ (_08381_, _08380_, _08370_);
  or _16742_ (_08382_, _08381_, _06531_);
  nor _16743_ (_08383_, _06498_, _06133_);
  not _16744_ (_08384_, _08383_);
  and _16745_ (_08385_, _08384_, _07559_);
  and _16746_ (_08386_, _08385_, _07546_);
  nand _16747_ (_08387_, _08386_, _06531_);
  and _16748_ (_08388_, _08387_, _05552_);
  and _16749_ (_07139_, _08388_, _08382_);
  not _16750_ (_08389_, _08234_);
  and _16751_ (_08390_, _08250_, _08389_);
  not _16752_ (_08391_, _08390_);
  and _16753_ (_08392_, _08250_, _08234_);
  nor _16754_ (_08393_, _08392_, _08256_);
  and _16755_ (_08394_, _08392_, _08256_);
  nor _16756_ (_08395_, _08394_, _08393_);
  not _16757_ (_08396_, _08395_);
  nor _16758_ (_08397_, _08396_, _08272_);
  and _16759_ (_08398_, _08394_, _08286_);
  or _16760_ (_08399_, _08394_, _08286_);
  not _16761_ (_08400_, _08399_);
  nor _16762_ (_08401_, _08400_, _08398_);
  nor _16763_ (_08402_, _08401_, _08395_);
  and _16764_ (_08403_, _08402_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and _16765_ (_08404_, _08393_, _08286_);
  and _16766_ (_08405_, _08394_, _08243_);
  nor _16767_ (_08406_, _08405_, _08404_);
  nor _16768_ (_08407_, _08406_, _08262_);
  or _16769_ (_08408_, _08407_, _08403_);
  nor _16770_ (_08409_, _08408_, _08397_);
  nor _16771_ (_08410_, _08409_, _08391_);
  not _16772_ (_08411_, _08392_);
  nor _16773_ (_08412_, _08396_, _08305_);
  nor _16774_ (_08413_, _08406_, _08293_);
  nor _16775_ (_08414_, _08413_, _08412_);
  or _16776_ (_08415_, _08414_, _08411_);
  nand _16777_ (_08416_, _08398_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and _16778_ (_08417_, _08416_, _08415_);
  not _16779_ (_08418_, _08417_);
  nor _16780_ (_08419_, _08418_, _08410_);
  and _16781_ (_08420_, _08251_, _08234_);
  not _16782_ (_08421_, _08420_);
  nor _16783_ (_08422_, _08396_, _08300_);
  and _16784_ (_08423_, _08402_, \oc8051_symbolic_cxrom1.regvalid [10]);
  not _16785_ (_08424_, \oc8051_symbolic_cxrom1.regvalid [2]);
  nor _16786_ (_08425_, _08406_, _08424_);
  or _16787_ (_08426_, _08425_, _08423_);
  nor _16788_ (_08427_, _08426_, _08422_);
  nor _16789_ (_08428_, _08427_, _08421_);
  nor _16790_ (_08429_, _08250_, _08234_);
  not _16791_ (_08430_, _08429_);
  nor _16792_ (_08431_, _08396_, _08246_);
  and _16793_ (_08432_, _08402_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor _16794_ (_08433_, _08406_, _08276_);
  or _16795_ (_08434_, _08433_, _08432_);
  nor _16796_ (_08436_, _08434_, _08431_);
  nor _16797_ (_08437_, _08436_, _08430_);
  nor _16798_ (_08438_, _08437_, _08428_);
  and _16799_ (_08439_, _08438_, _08419_);
  or _16800_ (_08440_, _08429_, _08392_);
  not _16801_ (_08441_, _08440_);
  not _16802_ (_08442_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  nand _16803_ (_08443_, _08234_, _08442_);
  or _16804_ (_08445_, _08234_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  and _16805_ (_08446_, _08445_, _08443_);
  and _16806_ (_08447_, _08446_, _08441_);
  not _16807_ (_08448_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  nand _16808_ (_08449_, _08234_, _08448_);
  or _16809_ (_08450_, _08234_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  and _16810_ (_08451_, _08450_, _08449_);
  and _16811_ (_08452_, _08451_, _08440_);
  or _16812_ (_08453_, _08452_, _08447_);
  and _16813_ (_08454_, _08453_, _08402_);
  not _16814_ (_08455_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  nand _16815_ (_08456_, _08234_, _08455_);
  or _16816_ (_08457_, _08234_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  and _16817_ (_08458_, _08457_, _08456_);
  and _16818_ (_08459_, _08458_, _08441_);
  not _16819_ (_08460_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  nand _16820_ (_08461_, _08234_, _08460_);
  or _16821_ (_08462_, _08234_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  and _16822_ (_08463_, _08462_, _08461_);
  and _16823_ (_08464_, _08463_, _08440_);
  nor _16824_ (_08465_, _08464_, _08459_);
  nor _16825_ (_08466_, _08465_, _08406_);
  and _16826_ (_08467_, _08395_, _08286_);
  not _16827_ (_08468_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  nand _16828_ (_08469_, _08234_, _08468_);
  or _16829_ (_08470_, _08234_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  and _16830_ (_08471_, _08470_, _08469_);
  and _16831_ (_08472_, _08471_, _08441_);
  not _16832_ (_08473_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  nand _16833_ (_08474_, _08234_, _08473_);
  or _16834_ (_08475_, _08234_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  and _16835_ (_08476_, _08475_, _08474_);
  and _16836_ (_08477_, _08476_, _08440_);
  or _16837_ (_08478_, _08477_, _08472_);
  and _16838_ (_08479_, _08478_, _08467_);
  and _16839_ (_08480_, _08395_, _08243_);
  not _16840_ (_08481_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  nand _16841_ (_08482_, _08234_, _08481_);
  or _16842_ (_08483_, _08234_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  and _16843_ (_08484_, _08483_, _08482_);
  and _16844_ (_08485_, _08484_, _08441_);
  not _16845_ (_08486_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  nand _16846_ (_08487_, _08234_, _08486_);
  or _16847_ (_08488_, _08234_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  and _16848_ (_08489_, _08488_, _08487_);
  and _16849_ (_08490_, _08489_, _08440_);
  or _16850_ (_08491_, _08490_, _08485_);
  and _16851_ (_08492_, _08491_, _08480_);
  or _16852_ (_08493_, _08492_, _08479_);
  or _16853_ (_08494_, _08493_, _08466_);
  nor _16854_ (_08495_, _08494_, _08454_);
  nor _16855_ (_08496_, _08495_, _08439_);
  and _16856_ (_08497_, _08439_, word_in[15]);
  or _16857_ (\oc8051_symbolic_cxrom1.cxrom_data_out [15], _08497_, _08496_);
  nor _16858_ (_08498_, _08279_, _08267_);
  not _16859_ (_08499_, _08498_);
  and _16860_ (_08500_, _08268_, _08243_);
  and _16861_ (_08501_, _08267_, _08286_);
  nor _16862_ (_08502_, _08501_, _08500_);
  and _16863_ (_08503_, _08502_, _08499_);
  and _16864_ (_08504_, _08503_, \oc8051_symbolic_cxrom1.regvalid [1]);
  not _16865_ (_08505_, _08504_);
  nor _16866_ (_08506_, _08499_, _08246_);
  nor _16867_ (_08507_, _08502_, _08498_);
  and _16868_ (_08508_, _08507_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor _16869_ (_08509_, _08508_, _08506_);
  and _16870_ (_08510_, _08509_, _08505_);
  nor _16871_ (_08511_, _08510_, _08411_);
  and _16872_ (_08512_, _08503_, \oc8051_symbolic_cxrom1.regvalid [3]);
  not _16873_ (_08513_, _08512_);
  nor _16874_ (_08514_, _08499_, _08272_);
  and _16875_ (_08515_, _08507_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor _16876_ (_08516_, _08515_, _08514_);
  and _16877_ (_08517_, _08516_, _08513_);
  nor _16878_ (_08518_, _08517_, _08421_);
  nor _16879_ (_08519_, _08518_, _08511_);
  nor _16880_ (_08520_, _08499_, _08300_);
  and _16881_ (_08521_, _08507_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and _16882_ (_08522_, _08503_, \oc8051_symbolic_cxrom1.regvalid [2]);
  or _16883_ (_08523_, _08522_, _08521_);
  nor _16884_ (_08524_, _08523_, _08520_);
  nor _16885_ (_08525_, _08524_, _08430_);
  nor _16886_ (_08526_, _08499_, _08305_);
  and _16887_ (_08527_, _08507_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and _16888_ (_08528_, _08503_, \oc8051_symbolic_cxrom1.regvalid [0]);
  or _16889_ (_08529_, _08528_, _08527_);
  nor _16890_ (_08530_, _08529_, _08526_);
  nor _16891_ (_08531_, _08530_, _08391_);
  nor _16892_ (_08532_, _08531_, _08525_);
  and _16893_ (_08533_, _08532_, _08519_);
  and _16894_ (_08534_, _08344_, _08257_);
  and _16895_ (_08535_, _08355_, _08267_);
  or _16896_ (_08536_, _08535_, _08534_);
  and _16897_ (_08537_, _08350_, _08260_);
  and _16898_ (_08538_, _08339_, _08279_);
  or _16899_ (_08539_, _08538_, _08537_);
  or _16900_ (_08540_, _08539_, _08536_);
  and _16901_ (_08541_, _08540_, _08502_);
  and _16902_ (_08542_, _08320_, _08279_);
  and _16903_ (_08543_, _08331_, _08267_);
  or _16904_ (_08544_, _08543_, _08542_);
  and _16905_ (_08545_, _08315_, _08257_);
  and _16906_ (_08546_, _08326_, _08260_);
  or _16907_ (_08547_, _08546_, _08545_);
  nor _16908_ (_08548_, _08547_, _08544_);
  nor _16909_ (_08549_, _08548_, _08502_);
  nor _16910_ (_08550_, _08549_, _08541_);
  nor _16911_ (_08552_, _08550_, _08533_);
  and _16912_ (_08553_, _08533_, word_in[23]);
  or _16913_ (\oc8051_symbolic_cxrom1.cxrom_data_out [23], _08553_, _08552_);
  and _16914_ (_08554_, _08256_, _08243_);
  and _16915_ (_08555_, _08554_, _08420_);
  and _16916_ (_08556_, _08555_, \oc8051_symbolic_cxrom1.regvalid [0]);
  nor _16917_ (_08557_, _08430_, _08256_);
  not _16918_ (_08558_, _08557_);
  nand _16919_ (_08559_, _08430_, _08256_);
  and _16920_ (_08561_, _08559_, _08558_);
  not _16921_ (_08562_, _08561_);
  nor _16922_ (_08563_, _08305_, _08562_);
  and _16923_ (_08564_, _08559_, _08243_);
  nor _16924_ (_08565_, _08559_, _08243_);
  nor _16925_ (_08566_, _08565_, _08564_);
  nor _16926_ (_08567_, _08566_, _08561_);
  and _16927_ (_08568_, _08567_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor _16928_ (_08569_, _08568_, _08563_);
  nor _16929_ (_08570_, _08569_, _08421_);
  nor _16930_ (_08571_, _08300_, _08562_);
  and _16931_ (_08572_, _08566_, _08562_);
  and _16932_ (_08573_, _08572_, \oc8051_symbolic_cxrom1.regvalid [2]);
  and _16933_ (_08574_, _08567_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or _16934_ (_08575_, _08574_, _08573_);
  nor _16935_ (_08576_, _08575_, _08571_);
  nor _16936_ (_08577_, _08576_, _08411_);
  or _16937_ (_08578_, _08577_, _08570_);
  nor _16938_ (_08579_, _08578_, _08556_);
  nor _16939_ (_08580_, _08562_, _08246_);
  and _16940_ (_08581_, _08567_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and _16941_ (_08582_, _08572_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or _16942_ (_08583_, _08582_, _08581_);
  nor _16943_ (_08584_, _08583_, _08580_);
  nor _16944_ (_08585_, _08584_, _08391_);
  nor _16945_ (_08587_, _08562_, _08272_);
  and _16946_ (_08588_, _08567_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor _16947_ (_08589_, _08588_, _08587_);
  nor _16948_ (_08590_, _08589_, _08430_);
  and _16949_ (_08592_, _08557_, _08263_);
  or _16950_ (_08593_, _08592_, _08590_);
  nor _16951_ (_08594_, _08593_, _08585_);
  and _16952_ (_08595_, _08594_, _08579_);
  and _16953_ (_08596_, _08451_, _08441_);
  and _16954_ (_08598_, _08446_, _08440_);
  or _16955_ (_08599_, _08598_, _08596_);
  and _16956_ (_08601_, _08599_, _08567_);
  and _16957_ (_08602_, _08463_, _08441_);
  and _16958_ (_08603_, _08458_, _08440_);
  or _16959_ (_08604_, _08603_, _08602_);
  and _16960_ (_08605_, _08604_, _08572_);
  and _16961_ (_08607_, _08561_, _08286_);
  and _16962_ (_08608_, _08476_, _08441_);
  and _16963_ (_08609_, _08471_, _08440_);
  or _16964_ (_08610_, _08609_, _08608_);
  and _16965_ (_08611_, _08610_, _08607_);
  and _16966_ (_08613_, _08561_, _08243_);
  and _16967_ (_08615_, _08489_, _08441_);
  and _16968_ (_08616_, _08484_, _08440_);
  or _16969_ (_08618_, _08616_, _08615_);
  and _16970_ (_08620_, _08618_, _08613_);
  or _16971_ (_08621_, _08620_, _08611_);
  or _16972_ (_08622_, _08621_, _08605_);
  nor _16973_ (_08623_, _08622_, _08601_);
  nor _16974_ (_08624_, _08623_, _08595_);
  and _16975_ (_08625_, _08595_, word_in[31]);
  or _16976_ (\oc8051_symbolic_cxrom1.cxrom_data_out [31], _08625_, _08624_);
  and _16977_ (_08626_, _07731_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and _16978_ (_08627_, _07733_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  nor _16979_ (_08628_, _08627_, _05593_);
  or _16980_ (_08629_, _08628_, _08626_);
  and _16981_ (_08630_, _07733_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _16982_ (_08631_, _08630_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and _16983_ (_08632_, _08631_, _05552_);
  and _16984_ (_07180_, _08632_, _08629_);
  or _16985_ (_08633_, _08554_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and _16986_ (_07207_, _08633_, _05552_);
  not _16987_ (_08634_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and _16988_ (_08635_, _07433_, _06769_);
  and _16989_ (_08636_, _08009_, _08635_);
  nor _16990_ (_08637_, _08636_, _08634_);
  or _16991_ (_08638_, _08637_, _06531_);
  and _16992_ (_08639_, _08636_, _08048_);
  or _16993_ (_08640_, _08639_, _08638_);
  nand _16994_ (_08641_, _06531_, _06306_);
  and _16995_ (_08642_, _08641_, _05552_);
  and _16996_ (_07223_, _08642_, _08640_);
  and _16997_ (_08643_, _08498_, _08243_);
  and _16998_ (_08644_, _08533_, _05552_);
  and _16999_ (_08645_, _08644_, _08420_);
  and _17000_ (_08646_, _08645_, _08643_);
  not _17001_ (_08647_, _08646_);
  and _17002_ (_08648_, _08439_, _05552_);
  and _17003_ (_08649_, _08648_, _08390_);
  and _17004_ (_08650_, _08649_, _08480_);
  and _17005_ (_08651_, _08283_, _05552_);
  and _17006_ (_08652_, _08651_, _08250_);
  nor _17007_ (_08653_, _08311_, rst);
  and _17008_ (_08654_, _08653_, _08554_);
  and _17009_ (_08655_, _08654_, _08652_);
  and _17010_ (_08656_, _08653_, word_in[7]);
  and _17011_ (_08657_, _08656_, _08655_);
  nor _17012_ (_08658_, _08655_, _08312_);
  nor _17013_ (_08659_, _08658_, _08657_);
  nor _17014_ (_08660_, _08659_, _08650_);
  and _17015_ (_08661_, _08650_, word_in[15]);
  or _17016_ (_08662_, _08661_, _08660_);
  and _17017_ (_08663_, _08662_, _08647_);
  and _17018_ (_08664_, _08595_, _05552_);
  and _17019_ (_08665_, _08664_, _08429_);
  and _17020_ (_08666_, _08665_, _08554_);
  and _17021_ (_08667_, _08644_, word_in[23]);
  and _17022_ (_08668_, _08667_, _08646_);
  or _17023_ (_08669_, _08668_, _08666_);
  or _17024_ (_08670_, _08669_, _08663_);
  not _17025_ (_08671_, _08666_);
  and _17026_ (_08672_, _08664_, word_in[31]);
  or _17027_ (_08673_, _08672_, _08671_);
  and _17028_ (_13877_, _08673_, _08670_);
  or _17029_ (_08674_, _08572_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and _17030_ (_07256_, _08674_, _05552_);
  not _17031_ (_08675_, _05546_);
  or _17032_ (_08676_, _05641_, _08675_);
  or _17033_ (_08677_, _05546_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and _17034_ (_08678_, _08677_, _05552_);
  and _17035_ (_07268_, _08678_, _08676_);
  or _17036_ (_08679_, _08280_, _08243_);
  not _17037_ (_08680_, _08679_);
  nor _17038_ (_08681_, _08405_, _08680_);
  and _17039_ (_08682_, _08554_, _08390_);
  nor _17040_ (_08683_, _08682_, \oc8051_symbolic_cxrom1.regvalid [1]);
  nand _17041_ (_08684_, _08683_, _08681_);
  and _17042_ (_07287_, _08684_, _05552_);
  and _17043_ (_08685_, _08404_, _08250_);
  nor _17044_ (_08686_, _08685_, \oc8051_symbolic_cxrom1.regvalid [2]);
  nand _17045_ (_08687_, _08686_, _08681_);
  and _17046_ (_07324_, _08687_, _05552_);
  or _17047_ (_08688_, _05550_, \oc8051_top_1.oc8051_rom1.data_o [18]);
  not _17048_ (_08689_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  nand _17049_ (_08690_, _05550_, _08689_);
  and _17050_ (_08691_, _08690_, _05552_);
  and _17051_ (_07338_, _08691_, _08688_);
  or _17052_ (_08692_, _05733_, _08675_);
  or _17053_ (_08693_, _05546_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and _17054_ (_08694_, _08693_, _05552_);
  and _17055_ (_07341_, _08694_, _08692_);
  or _17056_ (_08695_, _08411_, _08243_);
  nor _17057_ (_08696_, _08695_, _08256_);
  or _17058_ (_08697_, _08256_, _08243_);
  or _17059_ (_08698_, _08697_, _08390_);
  and _17060_ (_08699_, _08698_, \oc8051_symbolic_cxrom1.regvalid [3]);
  or _17061_ (_08700_, _08699_, _08696_);
  and _17062_ (_08701_, _08700_, _08406_);
  and _17063_ (_08702_, _08279_, _08263_);
  or _17064_ (_08703_, _08702_, _08685_);
  or _17065_ (_08704_, _08703_, _08701_);
  and _17066_ (_08706_, _08704_, _08681_);
  or _17067_ (_08707_, _08702_, _08700_);
  and _17068_ (_08708_, _08707_, _08405_);
  or _17069_ (_08710_, _08708_, _08680_);
  or _17070_ (_08711_, _08710_, _08706_);
  and _17071_ (_07361_, _08711_, _05552_);
  nand _17072_ (_08713_, _05665_, _05546_);
  or _17073_ (_08714_, _05546_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and _17074_ (_08716_, _08714_, _05552_);
  and _17075_ (_07409_, _08716_, _08713_);
  not _17076_ (_08718_, _08256_);
  nor _17077_ (_08720_, _08718_, _08243_);
  and _17078_ (_08722_, _08720_, _08429_);
  or _17079_ (_08723_, _08696_, \oc8051_symbolic_cxrom1.regvalid [4]);
  or _17080_ (_08725_, _08723_, _08722_);
  and _17081_ (_08726_, _08725_, _08406_);
  or _17082_ (_08727_, _08722_, \oc8051_symbolic_cxrom1.regvalid [4]);
  and _17083_ (_08728_, _08727_, _08405_);
  and _17084_ (_08729_, _08420_, _08607_);
  and _17085_ (_08730_, _08557_, _08286_);
  and _17086_ (_08731_, _08730_, \oc8051_symbolic_cxrom1.regvalid [4]);
  or _17087_ (_08732_, _08731_, _08729_);
  or _17088_ (_08733_, _08732_, _08728_);
  or _17089_ (_08734_, _08733_, _08685_);
  or _17090_ (_08735_, _08734_, _08726_);
  and _17091_ (_07415_, _08735_, _05552_);
  nor _17092_ (_08736_, _08267_, _08243_);
  not _17093_ (_08737_, _08736_);
  or _17094_ (_08738_, _08722_, _08696_);
  or _17095_ (_08739_, _08738_, _08737_);
  and _17096_ (_08740_, _08739_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and _17097_ (_08741_, _08420_, _08720_);
  and _17098_ (_08742_, _08393_, _08244_);
  or _17099_ (_08743_, _08742_, _08741_);
  or _17100_ (_08744_, _08743_, _08740_);
  or _17101_ (_08745_, _08400_, _08565_);
  and _17102_ (_08746_, _08745_, _08744_);
  and _17103_ (_08747_, _08561_, _08244_);
  or _17104_ (_08748_, _08747_, _08722_);
  or _17105_ (_08749_, _08748_, _08746_);
  and _17106_ (_08750_, _08749_, _08682_);
  or _17107_ (_08751_, _08720_, _08500_);
  and _17108_ (_08752_, _08749_, _08751_);
  and _17109_ (_08753_, _08744_, _08405_);
  nor _17110_ (_08754_, _08679_, _08235_);
  or _17111_ (_08755_, _08754_, _08685_);
  or _17112_ (_08756_, _08755_, _08696_);
  or _17113_ (_08757_, _08756_, _08753_);
  or _17114_ (_08758_, _08757_, _08752_);
  or _17115_ (_08759_, _08758_, _08750_);
  and _17116_ (_07480_, _08759_, _05552_);
  and _17117_ (_08760_, _06569_, _05822_);
  and _17118_ (_08761_, _06569_, _05737_);
  nand _17119_ (_08762_, _06576_, _08761_);
  or _17120_ (_08763_, _08762_, _06572_);
  and _17121_ (_08764_, _08763_, _01436_);
  or _17122_ (_07502_, _08764_, _08760_);
  and _17123_ (_08765_, _08720_, _08390_);
  or _17124_ (_08766_, _08765_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or _17125_ (_08767_, _08765_, _08243_);
  and _17126_ (_08768_, _08256_, _08234_);
  and _17127_ (_08769_, _08404_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or _17128_ (_08770_, _08769_, _08768_);
  or _17129_ (_08771_, _08770_, _08767_);
  and _17130_ (_08772_, _08771_, _08766_);
  and _17131_ (_08773_, _08772_, _08737_);
  and _17132_ (_08774_, _08738_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or _17133_ (_08775_, _08774_, _08741_);
  or _17134_ (_08776_, _08775_, _08773_);
  and _17135_ (_08777_, _08776_, _08745_);
  and _17136_ (_08778_, _08766_, _08405_);
  or _17137_ (_08779_, _08769_, _08696_);
  or _17138_ (_08780_, _08779_, _08722_);
  or _17139_ (_08781_, _08780_, _08778_);
  or _17140_ (_08782_, _08781_, _08777_);
  and _17141_ (_07541_, _08782_, _05552_);
  and _17142_ (_08783_, _08243_, \oc8051_symbolic_cxrom1.regvalid [7]);
  and _17143_ (_08784_, _08730_, \oc8051_symbolic_cxrom1.regvalid [7]);
  and _17144_ (_08785_, _08607_, \oc8051_symbolic_cxrom1.regvalid [7]);
  or _17145_ (_08786_, _08785_, _08722_);
  or _17146_ (_08787_, _08786_, _08784_);
  or _17147_ (_08788_, _08741_, _08765_);
  or _17148_ (_08789_, _08788_, _08787_);
  or _17149_ (_08790_, _08789_, _08398_);
  or _17150_ (_08791_, _08790_, _08783_);
  and _17151_ (_07615_, _08791_, _05552_);
  nor _17152_ (_08792_, _08607_, _08567_);
  or _17153_ (_08793_, _08792_, _08398_);
  and _17154_ (_08794_, _08793_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and _17155_ (_08795_, _08557_, _08243_);
  not _17156_ (_08796_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor _17157_ (_08797_, _08440_, _08796_);
  and _17158_ (_08798_, _08797_, _08607_);
  and _17159_ (_08799_, _08738_, \oc8051_symbolic_cxrom1.regvalid [8]);
  or _17160_ (_08800_, _08799_, _08798_);
  or _17161_ (_08802_, _08800_, _08795_);
  or _17162_ (_08803_, _08802_, _08794_);
  and _17163_ (_08804_, _08803_, _08243_);
  not _17164_ (_08806_, _08768_);
  and _17165_ (_08807_, _08736_, _08806_);
  and _17166_ (_08808_, _08807_, \oc8051_symbolic_cxrom1.regvalid [8]);
  or _17167_ (_08809_, _08741_, _08398_);
  or _17168_ (_08811_, _08809_, _08808_);
  or _17169_ (_08812_, _08811_, _08765_);
  or _17170_ (_08813_, _08812_, _08804_);
  and _17171_ (_07673_, _08813_, _05552_);
  nor _17172_ (_08815_, _08399_, _08557_);
  and _17173_ (_08816_, _08501_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and _17174_ (_08818_, _08420_, _08613_);
  or _17175_ (_08819_, _08818_, _08275_);
  or _17176_ (_08820_, _08819_, _08816_);
  and _17177_ (_08821_, _08820_, _08815_);
  or _17178_ (_08823_, _08741_, _08607_);
  and _17179_ (_08824_, _08823_, \oc8051_symbolic_cxrom1.regvalid [9]);
  or _17180_ (_08826_, _08816_, _08795_);
  or _17181_ (_08827_, _08826_, _08824_);
  or _17182_ (_08828_, _08827_, _08821_);
  and _17183_ (_08829_, _08828_, _08400_);
  and _17184_ (_08830_, _08736_, \oc8051_symbolic_cxrom1.regvalid [9]);
  or _17185_ (_08831_, _08830_, _08765_);
  and _17186_ (_08832_, _08820_, _08405_);
  or _17187_ (_08833_, _08832_, _08398_);
  or _17188_ (_08834_, _08833_, _08831_);
  or _17189_ (_08835_, _08834_, _08829_);
  and _17190_ (_07739_, _08835_, _05552_);
  not _17191_ (_08836_, rxd_i);
  and _17192_ (_08837_, _07734_, _05564_);
  and _17193_ (_08838_, _07736_, _08837_);
  nand _17194_ (_08839_, _08838_, _08836_);
  or _17195_ (_08840_, _08838_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  and _17196_ (_08841_, _08840_, _05552_);
  and _17197_ (_07822_, _08841_, _08839_);
  and _17198_ (_08842_, _08280_, _08243_);
  and _17199_ (_08843_, _08765_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or _17200_ (_08844_, _08738_, _08741_);
  and _17201_ (_08846_, _08844_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or _17202_ (_08847_, _08846_, _08843_);
  and _17203_ (_08848_, _08730_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and _17204_ (_08849_, _08643_, _08390_);
  or _17205_ (_08850_, _08256_, _08234_);
  and _17206_ (_08851_, _08850_, _08284_);
  or _17207_ (_08852_, _08851_, _08849_);
  or _17208_ (_08853_, _08852_, _08848_);
  and _17209_ (_08854_, _08441_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and _17210_ (_08855_, _08854_, _08607_);
  or _17211_ (_08856_, _08795_, _08398_);
  and _17212_ (_08857_, _08856_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or _17213_ (_08858_, _08857_, _08855_);
  or _17214_ (_08859_, _08858_, _08853_);
  or _17215_ (_08860_, _08859_, _08847_);
  and _17216_ (_08861_, _08860_, _08842_);
  and _17217_ (_08862_, _08498_, _08286_);
  and _17218_ (_08863_, _08862_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and _17219_ (_08864_, _08680_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or _17220_ (_08865_, _08864_, _08398_);
  or _17221_ (_08866_, _08865_, _08843_);
  or _17222_ (_08867_, _08866_, _08863_);
  or _17223_ (_08868_, _08867_, _08818_);
  or _17224_ (_08869_, _08868_, _08861_);
  or _17225_ (_08870_, _08869_, _08795_);
  and _17226_ (_07829_, _08870_, _05552_);
  or _17227_ (_08871_, _08628_, _07731_);
  and _17228_ (_08872_, _08871_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  and _17229_ (_08873_, _08627_, _05563_);
  and _17230_ (_08874_, _07736_, _08873_);
  or _17231_ (_08875_, _08874_, _08872_);
  and _17232_ (_07858_, _08875_, _05552_);
  and _17233_ (_08876_, _08730_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and _17234_ (_08877_, _08467_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and _17235_ (_08878_, _08398_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor _17236_ (_08879_, _08440_, _08697_);
  and _17237_ (_08880_, _08879_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or _17238_ (_08881_, _08880_, _08878_);
  or _17239_ (_08882_, _08881_, _08877_);
  or _17240_ (_08883_, _08882_, _08795_);
  or _17241_ (_08884_, _08883_, _08876_);
  or _17242_ (_08885_, _08405_, _08480_);
  and _17243_ (_08886_, _08680_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and _17244_ (_08887_, _08720_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or _17245_ (_08888_, _08887_, _08886_);
  and _17246_ (_08889_, _08288_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and _17247_ (_08890_, _08260_, _08243_);
  or _17248_ (_08891_, _08234_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and _17249_ (_08892_, _08891_, _08890_);
  and _17250_ (_08893_, _08264_, _08261_);
  or _17251_ (_08894_, _08893_, _08892_);
  or _17252_ (_08895_, _08894_, _08889_);
  or _17253_ (_08896_, _08895_, _08888_);
  and _17254_ (_08897_, _08896_, _08885_);
  or _17255_ (_08898_, _08897_, _08884_);
  or _17256_ (_08900_, _08898_, _08818_);
  or _17257_ (_08901_, _08900_, _08849_);
  and _17258_ (_07927_, _08901_, _05552_);
  nand _17259_ (_08903_, _07600_, _07260_);
  or _17260_ (_08904_, _07574_, _06972_);
  nor _17261_ (_08905_, _07264_, _06396_);
  nor _17262_ (_08906_, _08905_, _06973_);
  nor _17263_ (_08908_, _08365_, _06396_);
  nor _17264_ (_08909_, _08908_, _08367_);
  and _17265_ (_08910_, _07261_, _06972_);
  and _17266_ (_08911_, _08910_, _07269_);
  not _17267_ (_08913_, _08911_);
  or _17268_ (_08914_, _08913_, _08909_);
  and _17269_ (_08915_, _08914_, _08906_);
  nor _17270_ (_08917_, _08915_, _07260_);
  nand _17271_ (_08918_, _08917_, _08904_);
  nand _17272_ (_08920_, _08918_, _08903_);
  and _17273_ (_07968_, _08920_, _05552_);
  nand _17274_ (_08921_, _08102_, _06973_);
  and _17275_ (_08923_, _08910_, _07264_);
  not _17276_ (_08924_, _08923_);
  not _17277_ (_08925_, _06056_);
  nor _17278_ (_08926_, _06763_, _08925_);
  nor _17279_ (_08927_, _06056_, _06243_);
  nor _17280_ (_08928_, _08927_, _08926_);
  or _17281_ (_08929_, _08928_, _08924_);
  and _17282_ (_08930_, _06020_, _05989_);
  and _17283_ (_08931_, _07262_, _08930_);
  and _17284_ (_08932_, _08931_, _06911_);
  and _17285_ (_08933_, _08932_, _06775_);
  not _17286_ (_08934_, _08933_);
  and _17287_ (_08935_, _08934_, _08910_);
  and _17288_ (_08936_, _08935_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor _17289_ (_08937_, _08936_, _07260_);
  and _17290_ (_08938_, _08937_, _08929_);
  nand _17291_ (_08939_, _08938_, _08921_);
  and _17292_ (_08940_, _08173_, _07260_);
  not _17293_ (_08941_, _08940_);
  and _17294_ (_08942_, _08941_, _08939_);
  and _17295_ (_07973_, _08942_, _05552_);
  and _17296_ (_08943_, _08554_, _08430_);
  and _17297_ (_08944_, _08943_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and _17298_ (_08945_, _08795_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and _17299_ (_08946_, _08643_, _08806_);
  or _17300_ (_08947_, _08946_, _08945_);
  and _17301_ (_08948_, _08250_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and _17302_ (_08949_, _08948_, _08607_);
  nor _17303_ (_08950_, _08679_, _08302_);
  and _17304_ (_08951_, _08720_, \oc8051_symbolic_cxrom1.regvalid [12]);
  or _17305_ (_08952_, _08951_, _08818_);
  or _17306_ (_08953_, _08952_, _08950_);
  or _17307_ (_08954_, _08953_, _08949_);
  or _17308_ (_08955_, _08954_, _08947_);
  or _17309_ (_08956_, _08955_, _08944_);
  and _17310_ (_08032_, _08956_, _05552_);
  nand _17311_ (_08957_, _08411_, _08243_);
  and _17312_ (_08958_, _08957_, _08695_);
  nor _17313_ (_08959_, _08958_, _08806_);
  nor _17314_ (_08960_, _08959_, _08393_);
  and _17315_ (_08961_, _08718_, _08243_);
  or _17316_ (_08962_, _08961_, _08398_);
  or _17317_ (_08963_, _08962_, _08960_);
  and _17318_ (_08964_, _08963_, \oc8051_symbolic_cxrom1.regvalid [13]);
  or _17319_ (_08965_, _08964_, _08251_);
  and _17320_ (_08966_, _08965_, _08554_);
  not _17321_ (_08967_, \oc8051_symbolic_cxrom1.regvalid [13]);
  nor _17322_ (_08968_, _08842_, _08967_);
  or _17323_ (_08969_, _08968_, _08890_);
  or _17324_ (_08970_, _08969_, _08966_);
  and _17325_ (_08119_, _08970_, _05552_);
  or _17326_ (_08971_, _08480_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and _17327_ (_08231_, _08971_, _05552_);
  not _17328_ (_08972_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and _17329_ (_08973_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  nor _17330_ (_08974_, _08973_, _08972_);
  and _17331_ (_08975_, _08973_, _08972_);
  nor _17332_ (_08976_, _08975_, _08974_);
  not _17333_ (_08977_, _08976_);
  and _17334_ (_08978_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and _17335_ (_08979_, _08978_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor _17336_ (_08980_, _08978_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor _17337_ (_08981_, _08980_, _08979_);
  or _17338_ (_08982_, _08981_, _08973_);
  and _17339_ (_08983_, _08982_, _08977_);
  nor _17340_ (_08984_, _08974_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and _17341_ (_08985_, _08974_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  or _17342_ (_08986_, _08985_, _08984_);
  or _17343_ (_08987_, _08979_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  and _17344_ (_10089_, _08987_, _05552_);
  and _17345_ (_08988_, _10089_, _08986_);
  and _17346_ (_08435_, _08988_, _08983_);
  nor _17347_ (_08989_, _06967_, _06020_);
  and _17348_ (_08990_, _08989_, _06060_);
  and _17349_ (_08991_, _08990_, _07443_);
  not _17350_ (_08992_, _08991_);
  not _17351_ (_08993_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff );
  and _17352_ (_08994_, _08993_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  not _17353_ (_08995_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  not _17354_ (_08996_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  and _17355_ (_08997_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  not _17356_ (_08998_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and _17357_ (_08999_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _08998_);
  nor _17358_ (_09000_, _08999_, _08997_);
  nor _17359_ (_09001_, _09000_, _08996_);
  or _17360_ (_09002_, _09001_, _08995_);
  and _17361_ (_09003_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], _08998_);
  and _17362_ (_09004_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _17363_ (_09005_, _09004_, _09003_);
  nor _17364_ (_09006_, _09005_, _08996_);
  not _17365_ (_09007_, _09006_);
  and _17366_ (_09008_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and _17367_ (_09009_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _08998_);
  nor _17368_ (_09010_, _09009_, _09008_);
  nor _17369_ (_09012_, _09010_, _08996_);
  nand _17370_ (_09013_, _09012_, _09007_);
  or _17371_ (_09014_, _09013_, _09002_);
  and _17372_ (_09015_, _09014_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or _17373_ (_09017_, _09015_, _08994_);
  nor _17374_ (_09018_, _06054_, _06020_);
  and _17375_ (_09019_, _09018_, _07433_);
  and _17376_ (_09020_, _09019_, _07443_);
  and _17377_ (_09021_, _09020_, _06775_);
  or _17378_ (_09022_, _09021_, _09017_);
  and _17379_ (_09023_, _09022_, _08992_);
  nand _17380_ (_09024_, _09021_, _06763_);
  and _17381_ (_09025_, _09024_, _09023_);
  nor _17382_ (_09026_, _08992_, _06306_);
  or _17383_ (_09027_, _09026_, _09025_);
  and _17384_ (_08444_, _09027_, _05552_);
  and _17385_ (_09028_, _07936_, _06308_);
  and _17386_ (_09029_, _09028_, _06068_);
  not _17387_ (_09030_, _09029_);
  and _17388_ (_09031_, _09030_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  and _17389_ (_09032_, _09028_, _07946_);
  or _17390_ (_09033_, _09032_, _09031_);
  and _17391_ (_08551_, _09033_, _05552_);
  and _17392_ (_09035_, _05552_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  and _17393_ (_09036_, _09035_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and _17394_ (_09038_, _05547_, _05671_);
  not _17395_ (_09039_, _09038_);
  not _17396_ (_09040_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor _17397_ (_09041_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13], \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  not _17398_ (_09042_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  not _17399_ (_09043_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  not _17400_ (_09044_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  not _17401_ (_09045_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  not _17402_ (_09046_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  not _17403_ (_09047_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  not _17404_ (_09048_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor _17405_ (_09049_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4], \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and _17406_ (_09050_, _09049_, _09048_);
  and _17407_ (_09051_, _09050_, _09047_);
  and _17408_ (_09052_, _09051_, _09046_);
  and _17409_ (_09053_, _09052_, _09045_);
  and _17410_ (_09054_, _09053_, _09044_);
  and _17411_ (_09055_, _09054_, _09043_);
  and _17412_ (_09056_, _09055_, _09042_);
  and _17413_ (_09057_, _09056_, _09041_);
  and _17414_ (_09058_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and _17415_ (_09059_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and _17416_ (_09060_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor _17417_ (_09061_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  nor _17418_ (_09062_, _09061_, _09059_);
  and _17419_ (_09063_, _09062_, _09060_);
  nor _17420_ (_09064_, _09063_, _09059_);
  nor _17421_ (_09065_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor _17422_ (_09066_, _09065_, _09058_);
  not _17423_ (_09067_, _09066_);
  nor _17424_ (_09068_, _09067_, _09064_);
  nor _17425_ (_09069_, _09068_, _09058_);
  and _17426_ (_09070_, _09069_, _09057_);
  and _17427_ (_09071_, _09070_, _09040_);
  nor _17428_ (_09072_, _09071_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and _17429_ (_09073_, _09071_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nor _17430_ (_09074_, _09073_, _09072_);
  not _17431_ (_09075_, _09074_);
  nor _17432_ (_09076_, _09070_, _09040_);
  nor _17433_ (_09077_, _09076_, _09071_);
  not _17434_ (_09078_, _09077_);
  not _17435_ (_09079_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and _17436_ (_09080_, _09069_, _09054_);
  and _17437_ (_09081_, _09080_, _09043_);
  and _17438_ (_09082_, _09081_, _09042_);
  and _17439_ (_09083_, _09082_, _09079_);
  nor _17440_ (_09084_, _09083_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and _17441_ (_09085_, _09083_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor _17442_ (_09086_, _09085_, _09084_);
  nor _17443_ (_09087_, _09082_, _09079_);
  nor _17444_ (_09088_, _09087_, _09083_);
  not _17445_ (_09089_, _09088_);
  nor _17446_ (_09090_, _09081_, _09042_);
  or _17447_ (_09091_, _09090_, _09082_);
  nor _17448_ (_09092_, _09080_, _09043_);
  nor _17449_ (_09093_, _09092_, _09081_);
  not _17450_ (_09094_, _09093_);
  and _17451_ (_09095_, _09069_, _09053_);
  nor _17452_ (_09096_, _09095_, _09044_);
  nor _17453_ (_09097_, _09096_, _09080_);
  not _17454_ (_09098_, _09097_);
  and _17455_ (_09099_, _09069_, _09051_);
  nor _17456_ (_09100_, _09099_, _09046_);
  and _17457_ (_09101_, _09069_, _09052_);
  or _17458_ (_09102_, _09101_, _09100_);
  and _17459_ (_09103_, _09069_, _09050_);
  nor _17460_ (_09104_, _09103_, _09047_);
  or _17461_ (_09105_, _09104_, _09099_);
  not _17462_ (_09106_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  not _17463_ (_09107_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and _17464_ (_09108_, _09069_, _09048_);
  and _17465_ (_09109_, _09108_, _09107_);
  nor _17466_ (_09111_, _09109_, _09106_);
  or _17467_ (_09112_, _09111_, _09103_);
  nor _17468_ (_09113_, _09069_, _09048_);
  nor _17469_ (_09114_, _09113_, _09108_);
  not _17470_ (_09116_, _09114_);
  nor _17471_ (_09117_, _09062_, _09060_);
  nor _17472_ (_09118_, _09117_, _09063_);
  not _17473_ (_09119_, _09118_);
  nor _17474_ (_09121_, _09119_, _07919_);
  not _17475_ (_09122_, _09121_);
  not _17476_ (_09123_, _07930_);
  nor _17477_ (_09124_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor _17478_ (_09126_, _09124_, _09060_);
  and _17479_ (_09127_, _09126_, _09123_);
  and _17480_ (_09128_, _09119_, _07919_);
  nor _17481_ (_09130_, _09128_, _09121_);
  nand _17482_ (_09131_, _09130_, _09127_);
  and _17483_ (_09132_, _09131_, _09122_);
  not _17484_ (_09133_, _09132_);
  and _17485_ (_09135_, _09067_, _09064_);
  nor _17486_ (_09136_, _09135_, _09068_);
  and _17487_ (_09137_, _09136_, _09133_);
  and _17488_ (_09139_, _09137_, _09116_);
  nor _17489_ (_09140_, _09108_, _09107_);
  or _17490_ (_09142_, _09140_, _09109_);
  and _17491_ (_09143_, _09142_, _09139_);
  and _17492_ (_09144_, _09143_, _09112_);
  and _17493_ (_09145_, _09144_, _09105_);
  and _17494_ (_09146_, _09145_, _09102_);
  nor _17495_ (_09147_, _09101_, _09045_);
  or _17496_ (_09148_, _09147_, _09095_);
  and _17497_ (_09149_, _09148_, _09146_);
  and _17498_ (_09150_, _09149_, _09098_);
  and _17499_ (_09151_, _09150_, _09094_);
  and _17500_ (_09152_, _09151_, _09091_);
  and _17501_ (_09153_, _09152_, _09089_);
  and _17502_ (_09154_, _09153_, _09086_);
  and _17503_ (_09155_, _09154_, _09078_);
  nor _17504_ (_09156_, _09155_, _09075_);
  and _17505_ (_09157_, _09155_, _09075_);
  or _17506_ (_09158_, _09157_, _09156_);
  or _17507_ (_09159_, _09158_, _09039_);
  or _17508_ (_09160_, _09038_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and _17509_ (_09161_, _09160_, _07933_);
  and _17510_ (_09162_, _09161_, _09159_);
  or _17511_ (_08560_, _09162_, _09036_);
  and _17512_ (_09163_, _08653_, _08250_);
  nor _17513_ (_09165_, _09163_, _08651_);
  and _17514_ (_09166_, _08653_, _08697_);
  not _17515_ (_09167_, _09166_);
  and _17516_ (_09168_, _09167_, _09165_);
  and _17517_ (_09169_, _09168_, _08653_);
  not _17518_ (_09170_, _09169_);
  and _17519_ (_09171_, _09170_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  and _17520_ (_09172_, _08653_, word_in[0]);
  and _17521_ (_09173_, _09172_, _09168_);
  or _17522_ (_09174_, _09173_, _09171_);
  and _17523_ (_09175_, _08648_, _08405_);
  not _17524_ (_09176_, _09175_);
  and _17525_ (_09177_, _09176_, _09174_);
  and _17526_ (_09178_, _08644_, _08682_);
  and _17527_ (_09179_, _08405_, word_in[8]);
  and _17528_ (_09180_, _09179_, _08648_);
  or _17529_ (_09181_, _09180_, _09178_);
  or _17530_ (_09182_, _09181_, _09177_);
  and _17531_ (_09183_, _08664_, _08555_);
  not _17532_ (_09184_, _09183_);
  not _17533_ (_09185_, _09178_);
  or _17534_ (_09186_, _09185_, word_in[16]);
  and _17535_ (_09187_, _09186_, _09184_);
  and _17536_ (_09188_, _09187_, _09182_);
  and _17537_ (_09189_, _08664_, word_in[24]);
  and _17538_ (_09190_, _09189_, _08555_);
  or _17539_ (_08586_, _09190_, _09188_);
  and _17540_ (_09191_, _08664_, word_in[25]);
  and _17541_ (_09192_, _09191_, _08555_);
  and _17542_ (_09193_, _09178_, word_in[17]);
  and _17543_ (_09194_, _09170_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  and _17544_ (_09195_, _08653_, word_in[1]);
  and _17545_ (_09196_, _09195_, _09168_);
  or _17546_ (_09197_, _09196_, _09194_);
  or _17547_ (_09198_, _09197_, _09175_);
  or _17548_ (_09199_, _09176_, word_in[9]);
  and _17549_ (_09200_, _09199_, _09185_);
  and _17550_ (_09201_, _09200_, _09198_);
  or _17551_ (_09202_, _09201_, _09193_);
  and _17552_ (_09203_, _09202_, _09184_);
  or _17553_ (_08591_, _09203_, _09192_);
  and _17554_ (_09204_, _08664_, word_in[26]);
  and _17555_ (_09205_, _09204_, _08555_);
  and _17556_ (_09206_, _09178_, word_in[18]);
  and _17557_ (_09207_, _08653_, word_in[2]);
  and _17558_ (_09208_, _09207_, _09168_);
  and _17559_ (_09209_, _09170_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  or _17560_ (_09210_, _09209_, _09208_);
  or _17561_ (_09211_, _09210_, _09175_);
  or _17562_ (_09212_, _09176_, word_in[10]);
  and _17563_ (_09213_, _09212_, _09185_);
  and _17564_ (_09214_, _09213_, _09211_);
  or _17565_ (_09215_, _09214_, _09206_);
  and _17566_ (_09216_, _09215_, _09184_);
  or _17567_ (_08597_, _09216_, _09205_);
  and _17568_ (_09218_, _08664_, word_in[27]);
  and _17569_ (_09219_, _09218_, _08555_);
  and _17570_ (_09221_, _09178_, word_in[19]);
  and _17571_ (_09222_, _09170_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  and _17572_ (_09223_, _08653_, word_in[3]);
  and _17573_ (_09225_, _09223_, _09168_);
  or _17574_ (_09226_, _09225_, _09222_);
  or _17575_ (_09227_, _09226_, _09175_);
  or _17576_ (_09228_, _09176_, word_in[11]);
  and _17577_ (_09230_, _09228_, _09185_);
  and _17578_ (_09231_, _09230_, _09227_);
  or _17579_ (_09232_, _09231_, _09221_);
  and _17580_ (_09234_, _09232_, _09184_);
  or _17581_ (_08600_, _09234_, _09219_);
  and _17582_ (_09236_, _08664_, word_in[28]);
  and _17583_ (_09237_, _09236_, _08555_);
  and _17584_ (_09239_, _09178_, word_in[20]);
  and _17585_ (_09240_, _09170_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  and _17586_ (_09241_, _08653_, word_in[4]);
  and _17587_ (_09243_, _09241_, _09169_);
  or _17588_ (_09244_, _09243_, _09240_);
  or _17589_ (_09245_, _09244_, _09175_);
  or _17590_ (_09246_, _09176_, word_in[12]);
  and _17591_ (_09247_, _09246_, _09185_);
  and _17592_ (_09248_, _09247_, _09245_);
  or _17593_ (_09249_, _09248_, _09239_);
  and _17594_ (_09250_, _09249_, _09184_);
  or _17595_ (_08606_, _09250_, _09237_);
  and _17596_ (_09251_, _08664_, word_in[29]);
  and _17597_ (_09252_, _09251_, _08555_);
  and _17598_ (_09253_, _08653_, word_in[5]);
  and _17599_ (_09254_, _09253_, _09168_);
  and _17600_ (_09255_, _09170_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  or _17601_ (_09256_, _09255_, _09254_);
  or _17602_ (_09257_, _09256_, _09175_);
  or _17603_ (_09258_, _09176_, word_in[13]);
  and _17604_ (_09259_, _09258_, _09185_);
  and _17605_ (_09260_, _09259_, _09257_);
  and _17606_ (_09261_, _09178_, word_in[21]);
  or _17607_ (_09262_, _09261_, _09260_);
  and _17608_ (_09263_, _09262_, _09184_);
  or _17609_ (_08612_, _09263_, _09252_);
  and _17610_ (_09264_, _09030_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  and _17611_ (_09265_, _09028_, _07976_);
  or _17612_ (_09266_, _09265_, _09264_);
  and _17613_ (_08614_, _09266_, _05552_);
  and _17614_ (_09267_, _08664_, word_in[30]);
  and _17615_ (_09268_, _09267_, _08555_);
  and _17616_ (_09269_, _08653_, word_in[6]);
  and _17617_ (_09270_, _09269_, _09168_);
  and _17618_ (_09271_, _09170_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  or _17619_ (_09272_, _09271_, _09270_);
  or _17620_ (_09273_, _09272_, _09175_);
  or _17621_ (_09274_, _09176_, word_in[14]);
  and _17622_ (_09275_, _09274_, _09185_);
  and _17623_ (_09276_, _09275_, _09273_);
  and _17624_ (_09277_, _09178_, word_in[22]);
  or _17625_ (_09278_, _09277_, _09276_);
  and _17626_ (_09279_, _09278_, _09184_);
  or _17627_ (_08617_, _09279_, _09268_);
  and _17628_ (_09280_, _09178_, word_in[23]);
  not _17629_ (_09281_, word_in[15]);
  nand _17630_ (_09282_, _09175_, _09281_);
  and _17631_ (_09283_, _09282_, _09185_);
  and _17632_ (_09284_, _09169_, word_in[7]);
  nor _17633_ (_09285_, _09169_, _08460_);
  or _17634_ (_09286_, _09285_, _09284_);
  or _17635_ (_09287_, _09286_, _09175_);
  and _17636_ (_09288_, _09287_, _09283_);
  or _17637_ (_09289_, _09288_, _09280_);
  and _17638_ (_09290_, _09289_, _09184_);
  and _17639_ (_09291_, _09183_, word_in[31]);
  or _17640_ (_08619_, _09291_, _09290_);
  and _17641_ (_09292_, _08664_, _08682_);
  not _17642_ (_09293_, _09292_);
  and _17643_ (_09294_, _08644_, _08392_);
  and _17644_ (_09295_, _09294_, _08503_);
  not _17645_ (_09296_, _09295_);
  not _17646_ (_09297_, _08406_);
  and _17647_ (_09298_, _08648_, _08429_);
  and _17648_ (_09299_, _09298_, _09297_);
  and _17649_ (_09300_, _08651_, _08251_);
  not _17650_ (_09301_, _09300_);
  nor _17651_ (_09302_, _09301_, _09166_);
  and _17652_ (_09303_, _09302_, _09172_);
  not _17653_ (_09304_, _09302_);
  and _17654_ (_09305_, _09304_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  nor _17655_ (_09306_, _09305_, _09303_);
  nor _17656_ (_09307_, _09306_, _09299_);
  and _17657_ (_09308_, _09299_, word_in[8]);
  or _17658_ (_09309_, _09308_, _09307_);
  and _17659_ (_09310_, _09309_, _09296_);
  and _17660_ (_09311_, _08644_, word_in[16]);
  and _17661_ (_09312_, _09295_, _09311_);
  or _17662_ (_09313_, _09312_, _09310_);
  and _17663_ (_09314_, _09313_, _09293_);
  and _17664_ (_09315_, _09292_, word_in[24]);
  or _17665_ (_08705_, _09315_, _09314_);
  and _17666_ (_09316_, _08644_, word_in[17]);
  and _17667_ (_09317_, _09295_, _09316_);
  and _17668_ (_09318_, _09302_, _09195_);
  and _17669_ (_09319_, _09304_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  nor _17670_ (_09320_, _09319_, _09318_);
  nor _17671_ (_09321_, _09320_, _09299_);
  and _17672_ (_09322_, _09299_, word_in[9]);
  or _17673_ (_09323_, _09322_, _09321_);
  and _17674_ (_09324_, _09323_, _09296_);
  or _17675_ (_09325_, _09324_, _09317_);
  and _17676_ (_09326_, _09325_, _09293_);
  and _17677_ (_09327_, _09292_, word_in[25]);
  or _17678_ (_08709_, _09327_, _09326_);
  and _17679_ (_09328_, _09302_, _09207_);
  and _17680_ (_09329_, _09304_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  nor _17681_ (_09330_, _09329_, _09328_);
  nor _17682_ (_09331_, _09330_, _09299_);
  and _17683_ (_09332_, _09299_, word_in[10]);
  or _17684_ (_09333_, _09332_, _09331_);
  and _17685_ (_09334_, _09333_, _09296_);
  and _17686_ (_09335_, _08644_, word_in[18]);
  and _17687_ (_09336_, _09295_, _09335_);
  or _17688_ (_09337_, _09336_, _09334_);
  and _17689_ (_09338_, _09337_, _09293_);
  and _17690_ (_09339_, _09292_, word_in[26]);
  or _17691_ (_08712_, _09339_, _09338_);
  and _17692_ (_09340_, _08644_, word_in[19]);
  and _17693_ (_09341_, _09295_, _09340_);
  and _17694_ (_09342_, _09302_, _09223_);
  and _17695_ (_09343_, _09304_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  nor _17696_ (_09344_, _09343_, _09342_);
  nor _17697_ (_09345_, _09344_, _09299_);
  and _17698_ (_09346_, _09299_, word_in[11]);
  or _17699_ (_09347_, _09346_, _09345_);
  and _17700_ (_09348_, _09347_, _09296_);
  or _17701_ (_09349_, _09348_, _09341_);
  and _17702_ (_09350_, _09349_, _09293_);
  and _17703_ (_09351_, _09292_, word_in[27]);
  or _17704_ (_08715_, _09351_, _09350_);
  and _17705_ (_09352_, _09302_, _09241_);
  and _17706_ (_09353_, _09304_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  nor _17707_ (_09354_, _09353_, _09352_);
  nor _17708_ (_09355_, _09354_, _09299_);
  and _17709_ (_09356_, _09299_, word_in[12]);
  or _17710_ (_09357_, _09356_, _09355_);
  and _17711_ (_09358_, _09357_, _09296_);
  and _17712_ (_09359_, _08644_, word_in[20]);
  and _17713_ (_09360_, _09295_, _09359_);
  or _17714_ (_09361_, _09360_, _09358_);
  and _17715_ (_09362_, _09361_, _09293_);
  and _17716_ (_09363_, _09292_, word_in[28]);
  or _17717_ (_08717_, _09363_, _09362_);
  and _17718_ (_09364_, _08644_, word_in[21]);
  and _17719_ (_09365_, _09295_, _09364_);
  and _17720_ (_09366_, _09302_, _09253_);
  and _17721_ (_09367_, _09304_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  nor _17722_ (_09368_, _09367_, _09366_);
  nor _17723_ (_09369_, _09368_, _09299_);
  and _17724_ (_09370_, _09299_, word_in[13]);
  or _17725_ (_09371_, _09370_, _09369_);
  and _17726_ (_09372_, _09371_, _09296_);
  or _17727_ (_09373_, _09372_, _09365_);
  and _17728_ (_09374_, _09373_, _09293_);
  and _17729_ (_09375_, _09292_, word_in[29]);
  or _17730_ (_08719_, _09375_, _09374_);
  and _17731_ (_09376_, _09302_, _09269_);
  and _17732_ (_09377_, _09304_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  nor _17733_ (_09378_, _09377_, _09376_);
  nor _17734_ (_09379_, _09378_, _09299_);
  and _17735_ (_09380_, _09299_, word_in[14]);
  or _17736_ (_09381_, _09380_, _09379_);
  and _17737_ (_09382_, _09381_, _09296_);
  and _17738_ (_09383_, _08644_, word_in[22]);
  and _17739_ (_09384_, _09295_, _09383_);
  or _17740_ (_09385_, _09384_, _09382_);
  and _17741_ (_09386_, _09385_, _09293_);
  and _17742_ (_09387_, _09292_, word_in[30]);
  or _17743_ (_08721_, _09387_, _09386_);
  nor _17744_ (_09388_, _09302_, _08352_);
  and _17745_ (_09389_, _09302_, _08656_);
  or _17746_ (_09390_, _09389_, _09388_);
  or _17747_ (_09391_, _09390_, _09299_);
  nand _17748_ (_09392_, _09299_, _09281_);
  and _17749_ (_09393_, _09392_, _09391_);
  or _17750_ (_09394_, _09393_, _09295_);
  or _17751_ (_09395_, _09296_, _08667_);
  and _17752_ (_09396_, _09395_, _09293_);
  and _17753_ (_09397_, _09396_, _09394_);
  and _17754_ (_09398_, _09292_, word_in[31]);
  or _17755_ (_08724_, _09398_, _09397_);
  and _17756_ (_09399_, _08664_, _08392_);
  and _17757_ (_09400_, _09399_, _08572_);
  and _17758_ (_09401_, _08644_, _08429_);
  and _17759_ (_09402_, _09401_, _08503_);
  not _17760_ (_09404_, _09402_);
  and _17761_ (_09405_, _08648_, _08420_);
  and _17762_ (_09406_, _09405_, _09297_);
  not _17763_ (_09407_, _08697_);
  not _17764_ (_09409_, _08651_);
  and _17765_ (_09410_, _09163_, _09409_);
  and _17766_ (_09411_, _09410_, _09407_);
  or _17767_ (_09412_, _09411_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  not _17768_ (_09413_, _09411_);
  or _17769_ (_09414_, _09413_, _09172_);
  and _17770_ (_09415_, _09414_, _09412_);
  or _17771_ (_09416_, _09415_, _09406_);
  not _17772_ (_09417_, _09406_);
  or _17773_ (_09418_, _09417_, word_in[8]);
  and _17774_ (_09419_, _09418_, _09416_);
  and _17775_ (_09420_, _09419_, _09404_);
  and _17776_ (_09421_, _09402_, _09311_);
  or _17777_ (_09422_, _09421_, _09420_);
  or _17778_ (_09423_, _09422_, _09400_);
  not _17779_ (_09424_, _09400_);
  or _17780_ (_09425_, _09424_, word_in[24]);
  and _17781_ (_08801_, _09425_, _09423_);
  and _17782_ (_09426_, _09411_, _09195_);
  and _17783_ (_09427_, _09413_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  or _17784_ (_09428_, _09427_, _09426_);
  and _17785_ (_09429_, _09428_, _09417_);
  and _17786_ (_09430_, _09406_, word_in[9]);
  or _17787_ (_09431_, _09430_, _09429_);
  and _17788_ (_09432_, _09431_, _09404_);
  and _17789_ (_09433_, _09402_, _09316_);
  or _17790_ (_09434_, _09433_, _09400_);
  or _17791_ (_09435_, _09434_, _09432_);
  or _17792_ (_09436_, _09424_, word_in[25]);
  and _17793_ (_08805_, _09436_, _09435_);
  and _17794_ (_09437_, _09402_, _09335_);
  and _17795_ (_09438_, _09411_, _09207_);
  and _17796_ (_09439_, _09413_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  or _17797_ (_09440_, _09439_, _09438_);
  or _17798_ (_09441_, _09440_, _09406_);
  or _17799_ (_09442_, _09417_, word_in[10]);
  and _17800_ (_09443_, _09442_, _09404_);
  and _17801_ (_09444_, _09443_, _09441_);
  or _17802_ (_09445_, _09444_, _09437_);
  and _17803_ (_09446_, _09445_, _09424_);
  and _17804_ (_09447_, _09400_, word_in[26]);
  or _17805_ (_08810_, _09447_, _09446_);
  and _17806_ (_09448_, _09411_, _09223_);
  and _17807_ (_09449_, _09413_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  or _17808_ (_09450_, _09449_, _09448_);
  or _17809_ (_09451_, _09450_, _09406_);
  or _17810_ (_09452_, _09417_, word_in[11]);
  and _17811_ (_09453_, _09452_, _09404_);
  and _17812_ (_09454_, _09453_, _09451_);
  and _17813_ (_09455_, _09402_, _09340_);
  or _17814_ (_09456_, _09455_, _09454_);
  and _17815_ (_09457_, _09456_, _09424_);
  and _17816_ (_09458_, _09400_, word_in[27]);
  or _17817_ (_08814_, _09458_, _09457_);
  and _17818_ (_09459_, _09411_, _09241_);
  and _17819_ (_09460_, _09413_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  or _17820_ (_09461_, _09460_, _09459_);
  or _17821_ (_09462_, _09461_, _09406_);
  or _17822_ (_09463_, _09417_, word_in[12]);
  and _17823_ (_09464_, _09463_, _09404_);
  and _17824_ (_09465_, _09464_, _09462_);
  and _17825_ (_09466_, _09402_, _09359_);
  or _17826_ (_09467_, _09466_, _09400_);
  or _17827_ (_09468_, _09467_, _09465_);
  or _17828_ (_09469_, _09424_, word_in[28]);
  and _17829_ (_08817_, _09469_, _09468_);
  and _17830_ (_09470_, _09411_, _09253_);
  and _17831_ (_09471_, _09413_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  or _17832_ (_09472_, _09471_, _09470_);
  or _17833_ (_09473_, _09472_, _09406_);
  or _17834_ (_09474_, _09417_, word_in[13]);
  and _17835_ (_09475_, _09474_, _09404_);
  and _17836_ (_09476_, _09475_, _09473_);
  and _17837_ (_09477_, _09402_, _09364_);
  or _17838_ (_09478_, _09477_, _09400_);
  or _17839_ (_09479_, _09478_, _09476_);
  or _17840_ (_09480_, _09424_, word_in[29]);
  and _17841_ (_13878_, _09480_, _09479_);
  and _17842_ (_09481_, _09411_, _09269_);
  and _17843_ (_09482_, _09413_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  or _17844_ (_09483_, _09482_, _09481_);
  or _17845_ (_09484_, _09483_, _09406_);
  or _17846_ (_09485_, _09417_, word_in[14]);
  and _17847_ (_09486_, _09485_, _09404_);
  and _17848_ (_09487_, _09486_, _09484_);
  and _17849_ (_09488_, _09402_, _09383_);
  or _17850_ (_09489_, _09488_, _09400_);
  or _17851_ (_09490_, _09489_, _09487_);
  or _17852_ (_09491_, _09424_, word_in[30]);
  and _17853_ (_08822_, _09491_, _09490_);
  and _17854_ (_09492_, _09402_, _08667_);
  and _17855_ (_09493_, _09411_, _08656_);
  nor _17856_ (_09494_, _09411_, _08455_);
  or _17857_ (_09495_, _09494_, _09493_);
  or _17858_ (_09496_, _09495_, _09406_);
  nand _17859_ (_09497_, _09406_, _09281_);
  and _17860_ (_09498_, _09497_, _09404_);
  and _17861_ (_09499_, _09498_, _09496_);
  or _17862_ (_09500_, _09499_, _09492_);
  and _17863_ (_09501_, _09500_, _09424_);
  and _17864_ (_09502_, _09400_, word_in[31]);
  or _17865_ (_08825_, _09502_, _09501_);
  nor _17866_ (_09503_, _07949_, _07937_);
  and _17867_ (_09504_, _07936_, _06065_);
  not _17868_ (_09505_, _09504_);
  nand _17869_ (_09506_, _09505_, _09503_);
  nor _17870_ (_09507_, _09506_, _06069_);
  or _17871_ (_09508_, _09507_, _06955_);
  and _17872_ (_09509_, _09508_, _09030_);
  or _17873_ (_09510_, _09509_, _06069_);
  and _17874_ (_09511_, _09510_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  nor _17875_ (_09512_, _09030_, _06306_);
  and _17876_ (_09513_, _06068_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  and _17877_ (_09514_, _09513_, _09506_);
  or _17878_ (_09515_, _09514_, _09512_);
  or _17879_ (_09516_, _09515_, _09511_);
  and _17880_ (_08845_, _09516_, _05552_);
  and _17881_ (_09517_, _08645_, _08503_);
  not _17882_ (_09518_, _09517_);
  and _17883_ (_09519_, _08649_, _09297_);
  not _17884_ (_09520_, _08652_);
  nor _17885_ (_09521_, _09166_, _09520_);
  and _17886_ (_09522_, _09521_, _09172_);
  not _17887_ (_09523_, _09521_);
  and _17888_ (_09524_, _09523_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  nor _17889_ (_09525_, _09524_, _09522_);
  nor _17890_ (_09526_, _09525_, _09519_);
  and _17891_ (_09527_, _09519_, word_in[8]);
  or _17892_ (_09528_, _09527_, _09526_);
  and _17893_ (_09529_, _09528_, _09518_);
  and _17894_ (_09530_, _08665_, _08572_);
  and _17895_ (_09531_, _09517_, _09311_);
  or _17896_ (_09532_, _09531_, _09530_);
  or _17897_ (_09533_, _09532_, _09529_);
  not _17898_ (_09534_, _09530_);
  or _17899_ (_09535_, _09534_, word_in[24]);
  and _17900_ (_13879_, _09535_, _09533_);
  and _17901_ (_09536_, _09521_, _09195_);
  and _17902_ (_09537_, _09523_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  nor _17903_ (_09538_, _09537_, _09536_);
  nor _17904_ (_09539_, _09538_, _09519_);
  and _17905_ (_09540_, _09519_, word_in[9]);
  or _17906_ (_09541_, _09540_, _09539_);
  and _17907_ (_09542_, _09541_, _09518_);
  and _17908_ (_09543_, _09517_, _09316_);
  or _17909_ (_09544_, _09543_, _09530_);
  or _17910_ (_09545_, _09544_, _09542_);
  or _17911_ (_09546_, _09534_, word_in[25]);
  and _17912_ (_08899_, _09546_, _09545_);
  and _17913_ (_09547_, _09521_, _09207_);
  and _17914_ (_09548_, _09523_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  nor _17915_ (_09549_, _09548_, _09547_);
  nor _17916_ (_09550_, _09549_, _09519_);
  and _17917_ (_09551_, _09519_, word_in[10]);
  or _17918_ (_09552_, _09551_, _09550_);
  and _17919_ (_09553_, _09552_, _09518_);
  and _17920_ (_09554_, _09517_, _09335_);
  or _17921_ (_09555_, _09554_, _09530_);
  or _17922_ (_09556_, _09555_, _09553_);
  or _17923_ (_09557_, _09534_, word_in[26]);
  and _17924_ (_08902_, _09557_, _09556_);
  and _17925_ (_09558_, _09521_, _09223_);
  and _17926_ (_09559_, _09523_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  nor _17927_ (_09560_, _09559_, _09558_);
  nor _17928_ (_09561_, _09560_, _09519_);
  and _17929_ (_09562_, _09519_, word_in[11]);
  or _17930_ (_09563_, _09562_, _09561_);
  and _17931_ (_09564_, _09563_, _09518_);
  and _17932_ (_09565_, _09517_, _09340_);
  or _17933_ (_09566_, _09565_, _09564_);
  and _17934_ (_09567_, _09566_, _09534_);
  and _17935_ (_09568_, _09530_, word_in[27]);
  or _17936_ (_08907_, _09568_, _09567_);
  and _17937_ (_09569_, _09521_, _09241_);
  and _17938_ (_09570_, _09523_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  nor _17939_ (_09571_, _09570_, _09569_);
  nor _17940_ (_09572_, _09571_, _09519_);
  and _17941_ (_09573_, _09519_, word_in[12]);
  or _17942_ (_09574_, _09573_, _09572_);
  and _17943_ (_09575_, _09574_, _09518_);
  and _17944_ (_09576_, _09517_, _09359_);
  or _17945_ (_09577_, _09576_, _09530_);
  or _17946_ (_09578_, _09577_, _09575_);
  or _17947_ (_09579_, _09534_, word_in[28]);
  and _17948_ (_08912_, _09579_, _09578_);
  or _17949_ (_09580_, _09521_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  or _17950_ (_09581_, _09523_, _09253_);
  and _17951_ (_09582_, _09581_, _09580_);
  or _17952_ (_09583_, _09582_, _09519_);
  not _17953_ (_09584_, word_in[13]);
  nand _17954_ (_09585_, _09519_, _09584_);
  and _17955_ (_09586_, _09585_, _09583_);
  and _17956_ (_09587_, _09586_, _09518_);
  and _17957_ (_09588_, _09517_, _09364_);
  or _17958_ (_09589_, _09588_, _09530_);
  or _17959_ (_09590_, _09589_, _09587_);
  or _17960_ (_09591_, _09534_, word_in[29]);
  and _17961_ (_08916_, _09591_, _09590_);
  and _17962_ (_09592_, _09521_, _09269_);
  and _17963_ (_09593_, _09523_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  nor _17964_ (_09594_, _09593_, _09592_);
  nor _17965_ (_09595_, _09594_, _09519_);
  and _17966_ (_09596_, _09519_, word_in[14]);
  or _17967_ (_09597_, _09596_, _09595_);
  and _17968_ (_09598_, _09597_, _09518_);
  and _17969_ (_09599_, _09517_, _09383_);
  or _17970_ (_09600_, _09599_, _09530_);
  or _17971_ (_09601_, _09600_, _09598_);
  or _17972_ (_09602_, _09534_, word_in[30]);
  and _17973_ (_08919_, _09602_, _09601_);
  nor _17974_ (_09603_, _09521_, _08336_);
  and _17975_ (_09604_, _09521_, _08656_);
  or _17976_ (_09605_, _09604_, _09603_);
  or _17977_ (_09606_, _09605_, _09519_);
  nand _17978_ (_09607_, _09519_, _09281_);
  and _17979_ (_09608_, _09607_, _09606_);
  or _17980_ (_09609_, _09608_, _09517_);
  or _17981_ (_09610_, _09518_, _08667_);
  and _17982_ (_09611_, _09610_, _09534_);
  and _17983_ (_09612_, _09611_, _09609_);
  and _17984_ (_09613_, _09530_, word_in[31]);
  or _17985_ (_08922_, _09613_, _09612_);
  and _17986_ (_09614_, _08644_, _08685_);
  not _17987_ (_09615_, _09614_);
  and _17988_ (_09616_, _08648_, _08696_);
  not _17989_ (_09617_, _09616_);
  and _17990_ (_09618_, _08653_, _08720_);
  and _17991_ (_09619_, _09618_, _09165_);
  not _17992_ (_09620_, _09619_);
  and _17993_ (_09621_, _09620_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  and _17994_ (_09622_, _09619_, word_in[0]);
  or _17995_ (_09623_, _09622_, _09621_);
  and _17996_ (_09624_, _09623_, _09617_);
  and _17997_ (_09625_, _09616_, word_in[8]);
  or _17998_ (_09626_, _09625_, _09624_);
  and _17999_ (_09627_, _09626_, _09615_);
  and _18000_ (_09628_, _08664_, _08561_);
  and _18001_ (_09629_, _09628_, _08566_);
  and _18002_ (_09630_, _09629_, _08420_);
  and _18003_ (_09631_, _09614_, _09311_);
  or _18004_ (_09632_, _09631_, _09630_);
  or _18005_ (_09633_, _09632_, _09627_);
  not _18006_ (_09634_, _09630_);
  or _18007_ (_09635_, _09634_, _09189_);
  and _18008_ (_09011_, _09635_, _09633_);
  and _18009_ (_09636_, _09620_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  and _18010_ (_09637_, _09619_, word_in[1]);
  or _18011_ (_09638_, _09637_, _09636_);
  and _18012_ (_09639_, _09638_, _09617_);
  and _18013_ (_09640_, _09616_, word_in[9]);
  or _18014_ (_09641_, _09640_, _09639_);
  or _18015_ (_09642_, _09641_, _09614_);
  nor _18016_ (_09643_, _09615_, _09316_);
  nor _18017_ (_09644_, _09643_, _09630_);
  and _18018_ (_09645_, _09644_, _09642_);
  and _18019_ (_09646_, _09630_, _09191_);
  or _18020_ (_09016_, _09646_, _09645_);
  and _18021_ (_09647_, _09620_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  and _18022_ (_09648_, _09619_, word_in[2]);
  or _18023_ (_09649_, _09648_, _09647_);
  and _18024_ (_09650_, _09649_, _09617_);
  and _18025_ (_09651_, _09616_, word_in[10]);
  or _18026_ (_09652_, _09651_, _09650_);
  and _18027_ (_09653_, _09652_, _09615_);
  and _18028_ (_09654_, _09614_, _09335_);
  or _18029_ (_09655_, _09654_, _09630_);
  or _18030_ (_09656_, _09655_, _09653_);
  or _18031_ (_09657_, _09634_, _09204_);
  and _18032_ (_13880_, _09657_, _09656_);
  and _18033_ (_09658_, _09620_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  and _18034_ (_09659_, _09619_, word_in[3]);
  or _18035_ (_09660_, _09659_, _09658_);
  and _18036_ (_09661_, _09660_, _09617_);
  and _18037_ (_09662_, _09616_, word_in[11]);
  or _18038_ (_09663_, _09662_, _09661_);
  and _18039_ (_09664_, _09663_, _09615_);
  and _18040_ (_09665_, _09614_, _09340_);
  or _18041_ (_09666_, _09665_, _09630_);
  or _18042_ (_09667_, _09666_, _09664_);
  or _18043_ (_09668_, _09634_, _09218_);
  and _18044_ (_13881_, _09668_, _09667_);
  and _18045_ (_09669_, _09620_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  and _18046_ (_09670_, _09619_, word_in[4]);
  or _18047_ (_09671_, _09670_, _09669_);
  and _18048_ (_09672_, _09671_, _09617_);
  and _18049_ (_09673_, _09616_, word_in[12]);
  or _18050_ (_09674_, _09673_, _09672_);
  and _18051_ (_09675_, _09674_, _09615_);
  and _18052_ (_09676_, _09614_, _09359_);
  or _18053_ (_09677_, _09676_, _09630_);
  or _18054_ (_09678_, _09677_, _09675_);
  or _18055_ (_09679_, _09634_, _09236_);
  and _18056_ (_13882_, _09679_, _09678_);
  and _18057_ (_09680_, _09620_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  and _18058_ (_09681_, _09619_, word_in[5]);
  or _18059_ (_09682_, _09681_, _09680_);
  and _18060_ (_09683_, _09682_, _09617_);
  and _18061_ (_09684_, _09616_, word_in[13]);
  or _18062_ (_09685_, _09684_, _09683_);
  and _18063_ (_09686_, _09685_, _09615_);
  and _18064_ (_09687_, _09614_, _09364_);
  or _18065_ (_09688_, _09687_, _09630_);
  or _18066_ (_09689_, _09688_, _09686_);
  or _18067_ (_09690_, _09634_, _09251_);
  and _18068_ (_13883_, _09690_, _09689_);
  and _18069_ (_09691_, _09620_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  and _18070_ (_09692_, _09619_, word_in[6]);
  or _18071_ (_09693_, _09692_, _09691_);
  and _18072_ (_09694_, _09693_, _09617_);
  and _18073_ (_09695_, _09616_, word_in[14]);
  or _18074_ (_09696_, _09695_, _09694_);
  and _18075_ (_09697_, _09696_, _09615_);
  and _18076_ (_09698_, _09614_, _09383_);
  or _18077_ (_09699_, _09698_, _09630_);
  or _18078_ (_09700_, _09699_, _09697_);
  or _18079_ (_09701_, _09634_, _09267_);
  and _18080_ (_09034_, _09701_, _09700_);
  nor _18081_ (_09702_, _09619_, _08473_);
  and _18082_ (_09703_, _09619_, word_in[7]);
  or _18083_ (_09704_, _09703_, _09702_);
  or _18084_ (_09705_, _09704_, _09616_);
  nand _18085_ (_09706_, _09616_, _09281_);
  and _18086_ (_09707_, _09706_, _09705_);
  or _18087_ (_09708_, _09707_, _09614_);
  or _18088_ (_09709_, _09615_, _08667_);
  and _18089_ (_09710_, _09709_, _09708_);
  or _18090_ (_09711_, _09710_, _09630_);
  or _18091_ (_09712_, _09634_, _08672_);
  and _18092_ (_09037_, _09712_, _09711_);
  and _18093_ (_09713_, _09629_, _08390_);
  not _18094_ (_09714_, _09713_);
  and _18095_ (_09715_, _09294_, _08862_);
  and _18096_ (_09716_, _09715_, _09311_);
  not _18097_ (_09717_, _09715_);
  and _18098_ (_09718_, _09298_, _08467_);
  and _18099_ (_09719_, _09618_, _09300_);
  and _18100_ (_09720_, _09719_, _09172_);
  not _18101_ (_09721_, _09719_);
  and _18102_ (_09722_, _09721_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  nor _18103_ (_09723_, _09722_, _09720_);
  nor _18104_ (_09724_, _09723_, _09718_);
  and _18105_ (_09725_, _09718_, word_in[8]);
  or _18106_ (_09726_, _09725_, _09724_);
  and _18107_ (_09727_, _09726_, _09717_);
  or _18108_ (_09728_, _09727_, _09716_);
  and _18109_ (_09729_, _09728_, _09714_);
  and _18110_ (_09730_, _09713_, word_in[24]);
  or _18111_ (_09110_, _09730_, _09729_);
  and _18112_ (_09731_, _09715_, _09316_);
  and _18113_ (_09732_, _09719_, _09195_);
  and _18114_ (_09733_, _09721_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  nor _18115_ (_09734_, _09733_, _09732_);
  nor _18116_ (_09735_, _09734_, _09718_);
  and _18117_ (_09736_, _09718_, word_in[9]);
  or _18118_ (_09737_, _09736_, _09735_);
  and _18119_ (_09738_, _09737_, _09717_);
  or _18120_ (_09739_, _09738_, _09731_);
  and _18121_ (_09740_, _09739_, _09714_);
  and _18122_ (_09741_, _09713_, word_in[25]);
  or _18123_ (_09115_, _09741_, _09740_);
  or _18124_ (_09742_, _09719_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  or _18125_ (_09743_, _09721_, _09207_);
  and _18126_ (_09744_, _09743_, _09742_);
  or _18127_ (_09745_, _09744_, _09718_);
  not _18128_ (_09746_, _09718_);
  or _18129_ (_09747_, _09746_, word_in[10]);
  and _18130_ (_09748_, _09747_, _09745_);
  or _18131_ (_09749_, _09748_, _09715_);
  or _18132_ (_09750_, _09717_, _09335_);
  and _18133_ (_09752_, _09750_, _09749_);
  or _18134_ (_09753_, _09752_, _09713_);
  or _18135_ (_09754_, _09714_, word_in[26]);
  and _18136_ (_09120_, _09754_, _09753_);
  or _18137_ (_09756_, _09717_, _09340_);
  or _18138_ (_09757_, _09719_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  or _18139_ (_09759_, _09721_, _09223_);
  and _18140_ (_09761_, _09759_, _09757_);
  or _18141_ (_09763_, _09761_, _09718_);
  or _18142_ (_09764_, _09746_, word_in[11]);
  and _18143_ (_09766_, _09764_, _09763_);
  or _18144_ (_09767_, _09766_, _09715_);
  and _18145_ (_09768_, _09767_, _09756_);
  or _18146_ (_09770_, _09768_, _09713_);
  or _18147_ (_09771_, _09714_, word_in[27]);
  and _18148_ (_09125_, _09771_, _09770_);
  and _18149_ (_09773_, _09719_, _09241_);
  and _18150_ (_09774_, _09721_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  nor _18151_ (_09775_, _09774_, _09773_);
  nor _18152_ (_09776_, _09775_, _09718_);
  and _18153_ (_09777_, _09718_, word_in[12]);
  or _18154_ (_09778_, _09777_, _09776_);
  and _18155_ (_09779_, _09778_, _09717_);
  and _18156_ (_09780_, _09715_, _09359_);
  or _18157_ (_09781_, _09780_, _09713_);
  or _18158_ (_09782_, _09781_, _09779_);
  or _18159_ (_09783_, _09714_, word_in[28]);
  and _18160_ (_09129_, _09783_, _09782_);
  or _18161_ (_09784_, _09719_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  or _18162_ (_09785_, _09721_, _09253_);
  and _18163_ (_09786_, _09785_, _09784_);
  or _18164_ (_09787_, _09786_, _09718_);
  nand _18165_ (_09788_, _09718_, _09584_);
  and _18166_ (_09789_, _09788_, _09787_);
  or _18167_ (_09790_, _09789_, _09715_);
  or _18168_ (_09791_, _09717_, _09364_);
  and _18169_ (_09792_, _09791_, _09790_);
  or _18170_ (_09793_, _09792_, _09713_);
  or _18171_ (_09794_, _09714_, word_in[29]);
  and _18172_ (_09134_, _09794_, _09793_);
  or _18173_ (_09795_, _09717_, _09383_);
  or _18174_ (_09796_, _09719_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  or _18175_ (_09797_, _09721_, _09269_);
  and _18176_ (_09798_, _09797_, _09796_);
  or _18177_ (_09799_, _09798_, _09718_);
  or _18178_ (_09800_, _09746_, word_in[14]);
  and _18179_ (_09801_, _09800_, _09799_);
  or _18180_ (_09802_, _09801_, _09715_);
  and _18181_ (_09803_, _09802_, _09795_);
  or _18182_ (_09804_, _09803_, _09713_);
  or _18183_ (_09805_, _09714_, word_in[30]);
  and _18184_ (_09138_, _09805_, _09804_);
  or _18185_ (_09806_, _09717_, _08667_);
  nor _18186_ (_09807_, _09719_, _08347_);
  and _18187_ (_09808_, _09719_, _08656_);
  or _18188_ (_09809_, _09808_, _09807_);
  or _18189_ (_09810_, _09809_, _09718_);
  nand _18190_ (_09811_, _09718_, _09281_);
  and _18191_ (_09812_, _09811_, _09810_);
  or _18192_ (_09813_, _09812_, _09715_);
  and _18193_ (_09814_, _09813_, _09806_);
  or _18194_ (_09815_, _09814_, _09713_);
  or _18195_ (_09816_, _09714_, word_in[31]);
  and _18196_ (_09141_, _09816_, _09815_);
  and _18197_ (_09817_, _05552_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  nand _18198_ (_09818_, _09817_, _05556_);
  nand _18199_ (_09819_, _05585_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  nand _18200_ (_09164_, _09819_, _09818_);
  and _18201_ (_09820_, _09401_, _08862_);
  not _18202_ (_09821_, _09820_);
  and _18203_ (_09822_, _09405_, _08467_);
  not _18204_ (_09823_, _09822_);
  and _18205_ (_09824_, _09618_, _09410_);
  not _18206_ (_09825_, _09824_);
  and _18207_ (_09826_, _09825_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  and _18208_ (_09827_, _09824_, word_in[0]);
  or _18209_ (_09828_, _09827_, _09826_);
  and _18210_ (_09829_, _09828_, _09823_);
  and _18211_ (_09830_, _09822_, word_in[8]);
  or _18212_ (_09831_, _09830_, _09829_);
  and _18213_ (_09833_, _09831_, _09821_);
  and _18214_ (_09834_, _09629_, _08392_);
  and _18215_ (_09835_, _09820_, _09311_);
  or _18216_ (_09837_, _09835_, _09834_);
  or _18217_ (_09838_, _09837_, _09833_);
  not _18218_ (_09839_, _09834_);
  or _18219_ (_09841_, _09839_, word_in[24]);
  and _18220_ (_09217_, _09841_, _09838_);
  and _18221_ (_09843_, _09824_, word_in[1]);
  and _18222_ (_09844_, _09825_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  or _18223_ (_09846_, _09844_, _09843_);
  and _18224_ (_09848_, _09846_, _09823_);
  and _18225_ (_09849_, _09822_, word_in[9]);
  or _18226_ (_09851_, _09849_, _09848_);
  and _18227_ (_09852_, _09851_, _09821_);
  and _18228_ (_09853_, _09820_, _09316_);
  or _18229_ (_09854_, _09853_, _09834_);
  or _18230_ (_09855_, _09854_, _09852_);
  or _18231_ (_09856_, _09839_, word_in[25]);
  and _18232_ (_09220_, _09856_, _09855_);
  or _18233_ (_09857_, _09821_, _09335_);
  or _18234_ (_09858_, _09824_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  or _18235_ (_09859_, _09825_, word_in[2]);
  and _18236_ (_09860_, _09859_, _09858_);
  or _18237_ (_09861_, _09860_, _09822_);
  or _18238_ (_09862_, _09823_, word_in[10]);
  and _18239_ (_09863_, _09862_, _09861_);
  or _18240_ (_09864_, _09863_, _09820_);
  and _18241_ (_09865_, _09864_, _09857_);
  or _18242_ (_09866_, _09865_, _09834_);
  or _18243_ (_09867_, _09839_, word_in[26]);
  and _18244_ (_09224_, _09867_, _09866_);
  and _18245_ (_09868_, _09825_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  and _18246_ (_09869_, _09824_, word_in[3]);
  or _18247_ (_09870_, _09869_, _09868_);
  and _18248_ (_09871_, _09870_, _09823_);
  and _18249_ (_09872_, _09822_, word_in[11]);
  or _18250_ (_09873_, _09872_, _09871_);
  and _18251_ (_09874_, _09873_, _09821_);
  and _18252_ (_09875_, _09820_, _09340_);
  or _18253_ (_09876_, _09875_, _09834_);
  or _18254_ (_09877_, _09876_, _09874_);
  or _18255_ (_09878_, _09839_, word_in[27]);
  and _18256_ (_09229_, _09878_, _09877_);
  and _18257_ (_09879_, _09825_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  and _18258_ (_09880_, _09824_, word_in[4]);
  or _18259_ (_09881_, _09880_, _09879_);
  and _18260_ (_09882_, _09881_, _09823_);
  and _18261_ (_09883_, _09822_, word_in[12]);
  or _18262_ (_09884_, _09883_, _09882_);
  and _18263_ (_09885_, _09884_, _09821_);
  and _18264_ (_09886_, _09820_, _09359_);
  or _18265_ (_09887_, _09886_, _09834_);
  or _18266_ (_09888_, _09887_, _09885_);
  or _18267_ (_09889_, _09839_, word_in[28]);
  and _18268_ (_09233_, _09889_, _09888_);
  or _18269_ (_09890_, _09821_, _09364_);
  and _18270_ (_09891_, _09825_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  and _18271_ (_09892_, _09824_, word_in[5]);
  or _18272_ (_09893_, _09892_, _09891_);
  or _18273_ (_09894_, _09893_, _09822_);
  nand _18274_ (_09895_, _09822_, _09584_);
  and _18275_ (_09896_, _09895_, _09894_);
  or _18276_ (_09897_, _09896_, _09820_);
  and _18277_ (_09898_, _09897_, _09890_);
  or _18278_ (_09899_, _09898_, _09834_);
  or _18279_ (_09900_, _09839_, word_in[29]);
  and _18280_ (_09235_, _09900_, _09899_);
  and _18281_ (_09901_, _09824_, word_in[6]);
  and _18282_ (_09902_, _09825_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  or _18283_ (_09903_, _09902_, _09901_);
  and _18284_ (_09904_, _09903_, _09823_);
  and _18285_ (_09905_, _09822_, word_in[14]);
  or _18286_ (_09906_, _09905_, _09904_);
  and _18287_ (_09907_, _09906_, _09821_);
  and _18288_ (_09908_, _09820_, _09383_);
  or _18289_ (_09909_, _09908_, _09834_);
  or _18290_ (_09911_, _09909_, _09907_);
  or _18291_ (_09912_, _09839_, word_in[30]);
  and _18292_ (_09238_, _09912_, _09911_);
  nor _18293_ (_09913_, _09824_, _08468_);
  and _18294_ (_09914_, _09824_, word_in[7]);
  or _18295_ (_09915_, _09914_, _09913_);
  or _18296_ (_09916_, _09915_, _09822_);
  nand _18297_ (_09917_, _09822_, _09281_);
  and _18298_ (_09918_, _09917_, _09916_);
  and _18299_ (_09919_, _09918_, _09821_);
  and _18300_ (_09920_, _09820_, _08667_);
  or _18301_ (_09921_, _09920_, _09834_);
  or _18302_ (_09922_, _09921_, _09919_);
  or _18303_ (_09924_, _09839_, word_in[31]);
  and _18304_ (_09242_, _09924_, _09922_);
  and _18305_ (_09927_, _08664_, _08722_);
  and _18306_ (_09928_, _08649_, _08467_);
  and _18307_ (_09930_, _09618_, _08652_);
  or _18308_ (_09931_, _09930_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  not _18309_ (_09933_, _09930_);
  or _18310_ (_09934_, _09933_, _09172_);
  and _18311_ (_09936_, _09934_, _09931_);
  or _18312_ (_09937_, _09936_, _09928_);
  not _18313_ (_09938_, _09928_);
  or _18314_ (_09940_, _09938_, word_in[8]);
  and _18315_ (_09942_, _09940_, _09937_);
  and _18316_ (_09943_, _08644_, _08498_);
  and _18317_ (_09944_, _09943_, _08502_);
  and _18318_ (_09945_, _09944_, _08420_);
  or _18319_ (_09946_, _09945_, _09942_);
  nand _18320_ (_09947_, _08862_, _08645_);
  or _18321_ (_09948_, _09947_, _09311_);
  and _18322_ (_09949_, _09948_, _09946_);
  or _18323_ (_09950_, _09949_, _09927_);
  not _18324_ (_09951_, _09927_);
  or _18325_ (_09952_, _09951_, word_in[24]);
  and _18326_ (_13884_, _09952_, _09950_);
  or _18327_ (_09953_, _09930_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  or _18328_ (_09954_, _09933_, _09195_);
  and _18329_ (_09955_, _09954_, _09953_);
  or _18330_ (_09956_, _09955_, _09928_);
  or _18331_ (_09957_, _09938_, word_in[9]);
  and _18332_ (_09958_, _09957_, _09956_);
  or _18333_ (_09959_, _09958_, _09945_);
  or _18334_ (_09960_, _09947_, _09316_);
  and _18335_ (_09961_, _09960_, _09959_);
  or _18336_ (_09962_, _09961_, _09927_);
  or _18337_ (_09963_, _09951_, word_in[25]);
  and _18338_ (_13885_, _09963_, _09962_);
  or _18339_ (_09964_, _09930_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  or _18340_ (_09965_, _09933_, _09207_);
  and _18341_ (_09966_, _09965_, _09964_);
  or _18342_ (_09967_, _09966_, _09928_);
  or _18343_ (_09968_, _09938_, word_in[10]);
  and _18344_ (_09969_, _09968_, _09967_);
  or _18345_ (_09970_, _09969_, _09945_);
  or _18346_ (_09971_, _09947_, _09335_);
  and _18347_ (_09972_, _09971_, _09970_);
  or _18348_ (_09973_, _09972_, _09927_);
  or _18349_ (_09974_, _09951_, word_in[26]);
  and _18350_ (_13886_, _09974_, _09973_);
  or _18351_ (_09975_, _09930_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  or _18352_ (_09976_, _09933_, _09223_);
  and _18353_ (_09977_, _09976_, _09975_);
  or _18354_ (_09978_, _09977_, _09928_);
  or _18355_ (_09979_, _09938_, word_in[11]);
  and _18356_ (_09980_, _09979_, _09978_);
  or _18357_ (_09981_, _09980_, _09945_);
  or _18358_ (_09982_, _09947_, _09340_);
  and _18359_ (_09983_, _09982_, _09981_);
  or _18360_ (_09984_, _09983_, _09927_);
  or _18361_ (_09985_, _09951_, word_in[27]);
  and _18362_ (_13887_, _09985_, _09984_);
  and _18363_ (_09986_, _09933_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  and _18364_ (_09987_, _09930_, _09241_);
  nor _18365_ (_09988_, _09987_, _09986_);
  nor _18366_ (_09989_, _09988_, _09928_);
  and _18367_ (_09990_, _09928_, word_in[12]);
  or _18368_ (_09991_, _09990_, _09989_);
  and _18369_ (_09992_, _09991_, _09947_);
  and _18370_ (_09993_, _09945_, _09359_);
  or _18371_ (_09994_, _09993_, _09992_);
  and _18372_ (_09995_, _09994_, _09951_);
  and _18373_ (_09996_, _09927_, word_in[28]);
  or _18374_ (_13888_, _09996_, _09995_);
  or _18375_ (_09997_, _09947_, _09364_);
  or _18376_ (_09998_, _09930_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  or _18377_ (_09999_, _09933_, _09253_);
  and _18378_ (_10000_, _09999_, _09998_);
  or _18379_ (_10001_, _10000_, _09928_);
  nand _18380_ (_10002_, _09928_, _09584_);
  and _18381_ (_10003_, _10002_, _10001_);
  or _18382_ (_10004_, _10003_, _09945_);
  and _18383_ (_10005_, _10004_, _09997_);
  or _18384_ (_10006_, _10005_, _09927_);
  or _18385_ (_10007_, _09951_, word_in[29]);
  and _18386_ (_13889_, _10007_, _10006_);
  or _18387_ (_10008_, _09930_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  or _18388_ (_10009_, _09933_, _09269_);
  and _18389_ (_10010_, _10009_, _10008_);
  or _18390_ (_10011_, _10010_, _09928_);
  or _18391_ (_10012_, _09938_, word_in[14]);
  and _18392_ (_10013_, _10012_, _10011_);
  or _18393_ (_10014_, _10013_, _09945_);
  or _18394_ (_10015_, _09947_, _09383_);
  and _18395_ (_10016_, _10015_, _10014_);
  or _18396_ (_10017_, _10016_, _09927_);
  or _18397_ (_10018_, _09951_, word_in[30]);
  and _18398_ (_13890_, _10018_, _10017_);
  nand _18399_ (_10019_, _09928_, _09281_);
  nor _18400_ (_10020_, _09930_, _08341_);
  and _18401_ (_10021_, _09930_, _08656_);
  or _18402_ (_10022_, _10021_, _10020_);
  nor _18403_ (_10023_, _10022_, _09928_);
  nor _18404_ (_10024_, _10023_, _09945_);
  and _18405_ (_10025_, _10024_, _10019_);
  and _18406_ (_10026_, _09945_, _08667_);
  or _18407_ (_10027_, _10026_, _10025_);
  and _18408_ (_10028_, _10027_, _09951_);
  and _18409_ (_10029_, _09927_, word_in[31]);
  or _18410_ (_13891_, _10029_, _10028_);
  and _18411_ (_10030_, _08664_, _08741_);
  not _18412_ (_10031_, _10030_);
  and _18413_ (_10032_, _08644_, _08765_);
  and _18414_ (_10034_, _10032_, word_in[16]);
  not _18415_ (_10035_, _10032_);
  and _18416_ (_10036_, _08648_, _08398_);
  not _18417_ (_10037_, _10036_);
  and _18418_ (_10038_, _08653_, _08961_);
  and _18419_ (_10039_, _10038_, _09165_);
  and _18420_ (_10040_, _10039_, word_in[0]);
  not _18421_ (_10041_, _10039_);
  and _18422_ (_10042_, _10041_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  or _18423_ (_10043_, _10042_, _10040_);
  and _18424_ (_10044_, _10043_, _10037_);
  and _18425_ (_10045_, _10036_, word_in[8]);
  or _18426_ (_10046_, _10045_, _10044_);
  and _18427_ (_10047_, _10046_, _10035_);
  or _18428_ (_10048_, _10047_, _10034_);
  and _18429_ (_10049_, _10048_, _10031_);
  and _18430_ (_10050_, _10030_, word_in[24]);
  or _18431_ (_09403_, _10050_, _10049_);
  and _18432_ (_10051_, _10032_, word_in[17]);
  and _18433_ (_10052_, _10041_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  and _18434_ (_10053_, _10039_, word_in[1]);
  or _18435_ (_10054_, _10053_, _10052_);
  and _18436_ (_10055_, _10054_, _10037_);
  and _18437_ (_10056_, _10036_, word_in[9]);
  or _18438_ (_10057_, _10056_, _10055_);
  and _18439_ (_10058_, _10057_, _10035_);
  or _18440_ (_10059_, _10058_, _10051_);
  and _18441_ (_10060_, _10059_, _10031_);
  and _18442_ (_10061_, _10030_, word_in[25]);
  or _18443_ (_09408_, _10061_, _10060_);
  and _18444_ (_10062_, _10032_, word_in[18]);
  and _18445_ (_10063_, _10041_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  and _18446_ (_10064_, _10039_, word_in[2]);
  or _18447_ (_10065_, _10064_, _10063_);
  and _18448_ (_10066_, _10065_, _10037_);
  and _18449_ (_10067_, _10036_, word_in[10]);
  or _18450_ (_10068_, _10067_, _10066_);
  and _18451_ (_10069_, _10068_, _10035_);
  or _18452_ (_10070_, _10069_, _10062_);
  and _18453_ (_10071_, _10070_, _10031_);
  and _18454_ (_10072_, _10030_, word_in[26]);
  or _18455_ (_13892_, _10072_, _10071_);
  and _18456_ (_10073_, _10032_, word_in[19]);
  and _18457_ (_10074_, _10041_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  and _18458_ (_10075_, _10039_, word_in[3]);
  or _18459_ (_10076_, _10075_, _10074_);
  and _18460_ (_10077_, _10076_, _10037_);
  and _18461_ (_10078_, _10036_, word_in[11]);
  or _18462_ (_10079_, _10078_, _10077_);
  and _18463_ (_10080_, _10079_, _10035_);
  or _18464_ (_10081_, _10080_, _10073_);
  and _18465_ (_10082_, _10081_, _10031_);
  and _18466_ (_10083_, _10030_, word_in[27]);
  or _18467_ (_13893_, _10083_, _10082_);
  and _18468_ (_10084_, _10032_, word_in[20]);
  and _18469_ (_10085_, _10041_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  and _18470_ (_10086_, _10039_, word_in[4]);
  or _18471_ (_10087_, _10086_, _10085_);
  and _18472_ (_10088_, _10087_, _10037_);
  and _18473_ (_10090_, _10036_, word_in[12]);
  or _18474_ (_10091_, _10090_, _10088_);
  and _18475_ (_10092_, _10091_, _10035_);
  or _18476_ (_10093_, _10092_, _10084_);
  and _18477_ (_10094_, _10093_, _10031_);
  and _18478_ (_10095_, _10030_, word_in[28]);
  or _18479_ (_13894_, _10095_, _10094_);
  and _18480_ (_10096_, _10032_, word_in[21]);
  and _18481_ (_10097_, _10041_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  and _18482_ (_10098_, _10039_, word_in[5]);
  or _18483_ (_10099_, _10098_, _10097_);
  and _18484_ (_10100_, _10099_, _10037_);
  and _18485_ (_10101_, _10036_, word_in[13]);
  or _18486_ (_10102_, _10101_, _10100_);
  and _18487_ (_10103_, _10102_, _10035_);
  or _18488_ (_10104_, _10103_, _10096_);
  and _18489_ (_10105_, _10104_, _10031_);
  and _18490_ (_10106_, _10030_, word_in[29]);
  or _18491_ (_13895_, _10106_, _10105_);
  and _18492_ (_10107_, _10032_, word_in[22]);
  and _18493_ (_10108_, _10041_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  and _18494_ (_10109_, _10039_, word_in[6]);
  or _18495_ (_10110_, _10109_, _10108_);
  and _18496_ (_10111_, _10110_, _10037_);
  and _18497_ (_10112_, _10036_, word_in[14]);
  or _18498_ (_10113_, _10112_, _10111_);
  and _18499_ (_10114_, _10113_, _10035_);
  or _18500_ (_10115_, _10114_, _10107_);
  and _18501_ (_10116_, _10115_, _10031_);
  and _18502_ (_10117_, _10030_, word_in[30]);
  or _18503_ (_13896_, _10117_, _10116_);
  nor _18504_ (_10118_, _10039_, _08448_);
  and _18505_ (_10120_, _10039_, word_in[7]);
  or _18506_ (_10121_, _10120_, _10118_);
  and _18507_ (_10122_, _10121_, _10037_);
  and _18508_ (_10123_, _10036_, word_in[15]);
  or _18509_ (_10124_, _10123_, _10122_);
  and _18510_ (_10125_, _10124_, _10035_);
  and _18511_ (_10126_, _10032_, word_in[23]);
  or _18512_ (_10127_, _10126_, _10125_);
  and _18513_ (_10128_, _10127_, _10031_);
  and _18514_ (_10129_, _10030_, word_in[31]);
  or _18515_ (_13897_, _10129_, _10128_);
  and _18516_ (_10130_, _09294_, _08507_);
  and _18517_ (_10131_, _09298_, _08402_);
  and _18518_ (_10132_, _10038_, _09300_);
  or _18519_ (_10133_, _10132_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  not _18520_ (_10134_, _10132_);
  or _18521_ (_10135_, _10134_, word_in[0]);
  and _18522_ (_10136_, _10135_, _10133_);
  or _18523_ (_10137_, _10136_, _10131_);
  not _18524_ (_10138_, _10131_);
  or _18525_ (_10139_, _10138_, word_in[8]);
  and _18526_ (_10140_, _10139_, _10137_);
  or _18527_ (_10141_, _10140_, _10130_);
  and _18528_ (_10142_, _08664_, _08567_);
  and _18529_ (_10143_, _10142_, _08390_);
  not _18530_ (_10144_, _10143_);
  not _18531_ (_10145_, _10130_);
  or _18532_ (_10146_, _10145_, _09311_);
  and _18533_ (_10147_, _10146_, _10144_);
  and _18534_ (_10148_, _10147_, _10141_);
  and _18535_ (_10149_, _10143_, word_in[24]);
  or _18536_ (_13898_, _10149_, _10148_);
  and _18537_ (_10150_, _10130_, _09316_);
  and _18538_ (_10151_, _10134_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  and _18539_ (_10152_, _10132_, word_in[1]);
  nor _18540_ (_10153_, _10152_, _10151_);
  nor _18541_ (_10154_, _10153_, _10131_);
  and _18542_ (_10155_, _10131_, word_in[9]);
  or _18543_ (_10156_, _10155_, _10154_);
  and _18544_ (_10157_, _10156_, _10145_);
  or _18545_ (_10158_, _10157_, _10150_);
  and _18546_ (_10159_, _10158_, _10144_);
  and _18547_ (_10160_, _10143_, word_in[25]);
  or _18548_ (_13899_, _10160_, _10159_);
  and _18549_ (_10161_, _10134_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  and _18550_ (_10162_, _10132_, word_in[2]);
  nor _18551_ (_10163_, _10162_, _10161_);
  nor _18552_ (_10164_, _10163_, _10131_);
  and _18553_ (_10165_, _10131_, word_in[10]);
  or _18554_ (_10166_, _10165_, _10164_);
  and _18555_ (_10167_, _10166_, _10145_);
  and _18556_ (_10168_, _10130_, _09335_);
  or _18557_ (_10169_, _10168_, _10167_);
  and _18558_ (_10170_, _10169_, _10144_);
  and _18559_ (_10171_, _10143_, word_in[26]);
  or _18560_ (_13900_, _10171_, _10170_);
  and _18561_ (_10172_, _10132_, word_in[3]);
  and _18562_ (_10173_, _10134_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  nor _18563_ (_10174_, _10173_, _10172_);
  nor _18564_ (_10175_, _10174_, _10131_);
  and _18565_ (_10176_, _10131_, word_in[11]);
  or _18566_ (_10177_, _10176_, _10175_);
  and _18567_ (_10178_, _10177_, _10145_);
  and _18568_ (_10179_, _10130_, _09340_);
  or _18569_ (_10180_, _10179_, _10143_);
  or _18570_ (_10181_, _10180_, _10178_);
  or _18571_ (_10182_, _10144_, word_in[27]);
  and _18572_ (_13901_, _10182_, _10181_);
  and _18573_ (_10183_, _10132_, word_in[4]);
  and _18574_ (_10184_, _10134_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  nor _18575_ (_10185_, _10184_, _10183_);
  nor _18576_ (_10186_, _10185_, _10131_);
  and _18577_ (_10187_, _10131_, word_in[12]);
  or _18578_ (_10188_, _10187_, _10186_);
  and _18579_ (_10189_, _10188_, _10145_);
  and _18580_ (_10190_, _10130_, _09359_);
  or _18581_ (_10191_, _10190_, _10189_);
  and _18582_ (_10192_, _10191_, _10144_);
  and _18583_ (_10193_, _10143_, word_in[28]);
  or _18584_ (_13902_, _10193_, _10192_);
  and _18585_ (_10194_, _10132_, word_in[5]);
  and _18586_ (_10195_, _10134_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  nor _18587_ (_10196_, _10195_, _10194_);
  nor _18588_ (_10197_, _10196_, _10131_);
  and _18589_ (_10198_, _10131_, word_in[13]);
  or _18590_ (_10199_, _10198_, _10197_);
  and _18591_ (_10200_, _10199_, _10145_);
  and _18592_ (_10201_, _10130_, _09364_);
  or _18593_ (_10202_, _10201_, _10200_);
  and _18594_ (_10203_, _10202_, _10144_);
  and _18595_ (_10204_, _10143_, word_in[29]);
  or _18596_ (_13903_, _10204_, _10203_);
  or _18597_ (_10205_, _10132_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  or _18598_ (_10206_, _10134_, word_in[6]);
  and _18599_ (_10207_, _10206_, _10205_);
  or _18600_ (_10208_, _10207_, _10131_);
  or _18601_ (_10209_, _10138_, word_in[14]);
  and _18602_ (_10210_, _10209_, _10208_);
  or _18603_ (_10211_, _10210_, _10130_);
  or _18604_ (_10212_, _10145_, _09383_);
  and _18605_ (_10213_, _10212_, _10144_);
  and _18606_ (_10214_, _10213_, _10211_);
  and _18607_ (_10215_, _10143_, word_in[30]);
  or _18608_ (_13904_, _10215_, _10214_);
  and _18609_ (_10216_, _10132_, word_in[7]);
  nor _18610_ (_10217_, _10132_, _08328_);
  nor _18611_ (_10218_, _10217_, _10216_);
  nor _18612_ (_10219_, _10218_, _10131_);
  and _18613_ (_10220_, _10131_, word_in[15]);
  or _18614_ (_10221_, _10220_, _10219_);
  and _18615_ (_10222_, _10221_, _10145_);
  and _18616_ (_10223_, _10130_, _08667_);
  or _18617_ (_10224_, _10223_, _10222_);
  and _18618_ (_10225_, _10224_, _10144_);
  and _18619_ (_10226_, _10143_, word_in[31]);
  or _18620_ (_13905_, _10226_, _10225_);
  and _18621_ (_10227_, _09401_, _08507_);
  and _18622_ (_10228_, _09405_, _08402_);
  and _18623_ (_10229_, _09410_, _08961_);
  not _18624_ (_10230_, _10229_);
  and _18625_ (_10231_, _10230_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and _18626_ (_10232_, _10229_, word_in[0]);
  or _18627_ (_10233_, _10232_, _10231_);
  or _18628_ (_10234_, _10233_, _10228_);
  not _18629_ (_10235_, _10228_);
  or _18630_ (_10236_, _10235_, word_in[8]);
  and _18631_ (_10237_, _10236_, _10234_);
  or _18632_ (_10238_, _10237_, _10227_);
  and _18633_ (_10239_, _10142_, _08392_);
  not _18634_ (_10240_, _10239_);
  not _18635_ (_10241_, _10227_);
  or _18636_ (_10242_, _10241_, _09311_);
  and _18637_ (_10243_, _10242_, _10240_);
  and _18638_ (_10244_, _10243_, _10238_);
  and _18639_ (_10245_, _10239_, word_in[24]);
  or _18640_ (_13853_, _10245_, _10244_);
  or _18641_ (_10246_, _10229_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  or _18642_ (_10248_, _10230_, word_in[1]);
  and _18643_ (_10249_, _10248_, _10246_);
  or _18644_ (_10250_, _10249_, _10228_);
  or _18645_ (_10251_, _10235_, word_in[9]);
  and _18646_ (_10252_, _10251_, _10250_);
  or _18647_ (_10253_, _10252_, _10227_);
  or _18648_ (_10255_, _10241_, _09316_);
  and _18649_ (_10256_, _10255_, _10253_);
  and _18650_ (_10258_, _10256_, _10240_);
  and _18651_ (_10259_, _10239_, word_in[25]);
  or _18652_ (_13854_, _10259_, _10258_);
  or _18653_ (_10260_, _10229_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  or _18654_ (_10261_, _10230_, word_in[2]);
  and _18655_ (_10262_, _10261_, _10260_);
  or _18656_ (_10264_, _10262_, _10228_);
  or _18657_ (_10265_, _10235_, word_in[10]);
  and _18658_ (_10266_, _10265_, _10264_);
  or _18659_ (_10267_, _10266_, _10227_);
  or _18660_ (_10268_, _10241_, _09335_);
  and _18661_ (_10270_, _10268_, _10240_);
  and _18662_ (_10271_, _10270_, _10267_);
  and _18663_ (_10272_, _10239_, word_in[26]);
  or _18664_ (_13855_, _10272_, _10271_);
  and _18665_ (_10273_, _10230_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  and _18666_ (_10274_, _10229_, word_in[3]);
  or _18667_ (_10275_, _10274_, _10273_);
  or _18668_ (_10276_, _10275_, _10228_);
  or _18669_ (_10277_, _10235_, word_in[11]);
  and _18670_ (_10278_, _10277_, _10276_);
  or _18671_ (_10279_, _10278_, _10227_);
  or _18672_ (_10280_, _10241_, _09340_);
  and _18673_ (_10281_, _10280_, _10240_);
  and _18674_ (_10283_, _10281_, _10279_);
  and _18675_ (_10284_, _10239_, word_in[27]);
  or _18676_ (_13856_, _10284_, _10283_);
  and _18677_ (_10285_, _10227_, _09359_);
  and _18678_ (_10286_, _10229_, word_in[4]);
  and _18679_ (_10287_, _10230_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  or _18680_ (_10288_, _10287_, _10286_);
  or _18681_ (_10289_, _10288_, _10228_);
  or _18682_ (_10290_, _10235_, word_in[12]);
  and _18683_ (_10291_, _10290_, _10241_);
  and _18684_ (_10292_, _10291_, _10289_);
  or _18685_ (_10293_, _10292_, _10285_);
  and _18686_ (_10294_, _10293_, _10240_);
  and _18687_ (_10295_, _10239_, word_in[28]);
  or _18688_ (_13857_, _10295_, _10294_);
  and _18689_ (_10296_, _10230_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  and _18690_ (_10297_, _10229_, word_in[5]);
  or _18691_ (_10299_, _10297_, _10296_);
  or _18692_ (_10300_, _10299_, _10228_);
  nand _18693_ (_10301_, _10228_, _09584_);
  and _18694_ (_10303_, _10301_, _10300_);
  or _18695_ (_10304_, _10303_, _10227_);
  or _18696_ (_10305_, _10241_, _09364_);
  and _18697_ (_10306_, _10305_, _10240_);
  and _18698_ (_10307_, _10306_, _10304_);
  and _18699_ (_10308_, _10239_, word_in[29]);
  or _18700_ (_13858_, _10308_, _10307_);
  or _18701_ (_10309_, _10229_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  or _18702_ (_10310_, _10230_, word_in[6]);
  and _18703_ (_10311_, _10310_, _10309_);
  or _18704_ (_10312_, _10311_, _10228_);
  or _18705_ (_10313_, _10235_, word_in[14]);
  and _18706_ (_10314_, _10313_, _10312_);
  or _18707_ (_10315_, _10314_, _10227_);
  or _18708_ (_10316_, _10241_, _09383_);
  and _18709_ (_10317_, _10316_, _10240_);
  and _18710_ (_10318_, _10317_, _10315_);
  and _18711_ (_10319_, _10239_, word_in[30]);
  or _18712_ (_13859_, _10319_, _10318_);
  nor _18713_ (_10320_, _10229_, _08442_);
  and _18714_ (_10321_, _10229_, word_in[7]);
  or _18715_ (_10322_, _10321_, _10320_);
  or _18716_ (_10323_, _10322_, _10228_);
  nand _18717_ (_10324_, _10228_, _09281_);
  and _18718_ (_10325_, _10324_, _10323_);
  or _18719_ (_10326_, _10325_, _10227_);
  or _18720_ (_10327_, _10241_, _08667_);
  and _18721_ (_10328_, _10327_, _10240_);
  and _18722_ (_10329_, _10328_, _10326_);
  and _18723_ (_10330_, _10239_, word_in[31]);
  or _18724_ (_13860_, _10330_, _10329_);
  and _18725_ (_10331_, _08645_, _08507_);
  not _18726_ (_10332_, _10331_);
  and _18727_ (_10333_, _08649_, _08402_);
  and _18728_ (_10334_, _10038_, _08652_);
  and _18729_ (_10335_, _10334_, word_in[0]);
  not _18730_ (_10336_, _10334_);
  and _18731_ (_10337_, _10336_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  nor _18732_ (_10338_, _10337_, _10335_);
  nor _18733_ (_10339_, _10338_, _10333_);
  and _18734_ (_10340_, _10333_, word_in[8]);
  or _18735_ (_10341_, _10340_, _10339_);
  and _18736_ (_10342_, _10341_, _10332_);
  and _18737_ (_10343_, _10142_, _08429_);
  and _18738_ (_10344_, _10331_, _09311_);
  or _18739_ (_10345_, _10344_, _10343_);
  or _18740_ (_10346_, _10345_, _10342_);
  not _18741_ (_10347_, _10343_);
  or _18742_ (_10348_, _10347_, _09189_);
  and _18743_ (_13861_, _10348_, _10346_);
  and _18744_ (_10349_, _10334_, word_in[1]);
  and _18745_ (_10350_, _10336_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  nor _18746_ (_10351_, _10350_, _10349_);
  nor _18747_ (_10352_, _10351_, _10333_);
  and _18748_ (_10353_, _10333_, word_in[9]);
  or _18749_ (_10354_, _10353_, _10352_);
  and _18750_ (_10355_, _10354_, _10332_);
  and _18751_ (_10356_, _10331_, _09316_);
  or _18752_ (_10357_, _10356_, _10343_);
  or _18753_ (_10358_, _10357_, _10355_);
  or _18754_ (_10359_, _10347_, _09191_);
  and _18755_ (_13862_, _10359_, _10358_);
  and _18756_ (_10360_, _10331_, _09335_);
  and _18757_ (_10362_, _10334_, word_in[2]);
  and _18758_ (_10363_, _10336_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  nor _18759_ (_10364_, _10363_, _10362_);
  nor _18760_ (_10365_, _10364_, _10333_);
  and _18761_ (_10366_, _10333_, word_in[10]);
  or _18762_ (_10367_, _10366_, _10365_);
  and _18763_ (_10368_, _10367_, _10332_);
  or _18764_ (_10369_, _10368_, _10360_);
  and _18765_ (_10370_, _10369_, _10347_);
  and _18766_ (_10371_, _10343_, word_in[26]);
  or _18767_ (_13863_, _10371_, _10370_);
  or _18768_ (_10372_, _10334_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  or _18769_ (_10373_, _10336_, word_in[3]);
  and _18770_ (_10374_, _10373_, _10372_);
  or _18771_ (_10375_, _10374_, _10333_);
  not _18772_ (_10376_, word_in[11]);
  nand _18773_ (_10377_, _10333_, _10376_);
  and _18774_ (_10378_, _10377_, _10375_);
  or _18775_ (_10379_, _10378_, _10331_);
  or _18776_ (_10380_, _10332_, _09340_);
  and _18777_ (_10381_, _10380_, _10347_);
  and _18778_ (_10382_, _10381_, _10379_);
  and _18779_ (_10383_, _10343_, _09218_);
  or _18780_ (_13864_, _10383_, _10382_);
  and _18781_ (_10384_, _10334_, word_in[4]);
  and _18782_ (_10385_, _10336_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  nor _18783_ (_10386_, _10385_, _10384_);
  nor _18784_ (_10387_, _10386_, _10333_);
  and _18785_ (_10388_, _10333_, word_in[12]);
  or _18786_ (_10389_, _10388_, _10387_);
  and _18787_ (_10390_, _10389_, _10332_);
  and _18788_ (_10391_, _10331_, _09359_);
  or _18789_ (_10392_, _10391_, _10390_);
  and _18790_ (_10393_, _10392_, _10347_);
  and _18791_ (_10394_, _10343_, word_in[28]);
  or _18792_ (_13865_, _10394_, _10393_);
  and _18793_ (_10395_, _10334_, word_in[5]);
  and _18794_ (_10396_, _10336_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  nor _18795_ (_10397_, _10396_, _10395_);
  nor _18796_ (_10398_, _10397_, _10333_);
  and _18797_ (_10399_, _10333_, word_in[13]);
  or _18798_ (_10400_, _10399_, _10398_);
  and _18799_ (_10401_, _10400_, _10332_);
  and _18800_ (_10402_, _10331_, _09364_);
  or _18801_ (_10403_, _10402_, _10343_);
  or _18802_ (_10404_, _10403_, _10401_);
  or _18803_ (_10405_, _10347_, _09251_);
  and _18804_ (_13866_, _10405_, _10404_);
  and _18805_ (_10406_, _10334_, word_in[6]);
  and _18806_ (_10407_, _10336_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  nor _18807_ (_10408_, _10407_, _10406_);
  nor _18808_ (_10409_, _10408_, _10333_);
  and _18809_ (_10410_, _10333_, word_in[14]);
  or _18810_ (_10411_, _10410_, _10409_);
  and _18811_ (_10412_, _10411_, _10332_);
  and _18812_ (_10413_, _10331_, _09383_);
  or _18813_ (_10414_, _10413_, _10412_);
  and _18814_ (_10415_, _10414_, _10347_);
  and _18815_ (_10416_, _10343_, word_in[30]);
  or _18816_ (_13867_, _10416_, _10415_);
  and _18817_ (_10417_, _10334_, word_in[7]);
  nor _18818_ (_10418_, _10334_, _08317_);
  nor _18819_ (_10419_, _10418_, _10417_);
  nor _18820_ (_10420_, _10419_, _10333_);
  and _18821_ (_10421_, _10333_, word_in[15]);
  or _18822_ (_10422_, _10421_, _10420_);
  and _18823_ (_10423_, _10422_, _10332_);
  and _18824_ (_10424_, _10331_, _08667_);
  or _18825_ (_10425_, _10424_, _10343_);
  or _18826_ (_10426_, _10425_, _10423_);
  or _18827_ (_10427_, _10347_, _08672_);
  and _18828_ (_13868_, _10427_, _10426_);
  and _18829_ (_10428_, _08644_, _08849_);
  not _18830_ (_10429_, _10428_);
  and _18831_ (_10430_, _08613_, _08392_);
  and _18832_ (_10431_, _08648_, _10430_);
  not _18833_ (_10432_, _10431_);
  and _18834_ (_10433_, _09165_, _08654_);
  and _18835_ (_10434_, _10433_, word_in[0]);
  not _18836_ (_10435_, _10433_);
  and _18837_ (_10436_, _10435_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  or _18838_ (_10437_, _10436_, _10434_);
  and _18839_ (_10438_, _10437_, _10432_);
  and _18840_ (_10439_, _10431_, word_in[8]);
  or _18841_ (_10440_, _10439_, _10438_);
  and _18842_ (_10441_, _10440_, _10429_);
  not _18843_ (_10442_, _08566_);
  and _18844_ (_10443_, _09628_, _10442_);
  and _18845_ (_10444_, _10443_, _08420_);
  and _18846_ (_10445_, _10428_, word_in[16]);
  or _18847_ (_10446_, _10445_, _10444_);
  or _18848_ (_10447_, _10446_, _10441_);
  not _18849_ (_10448_, _10444_);
  or _18850_ (_10449_, _10448_, _09189_);
  and _18851_ (_09751_, _10449_, _10447_);
  and _18852_ (_10450_, _10435_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  and _18853_ (_10451_, _10433_, word_in[1]);
  or _18854_ (_10452_, _10451_, _10450_);
  and _18855_ (_10453_, _10452_, _10432_);
  and _18856_ (_10454_, _10431_, word_in[9]);
  or _18857_ (_10455_, _10454_, _10453_);
  and _18858_ (_10456_, _10455_, _10429_);
  and _18859_ (_10457_, _10428_, word_in[17]);
  or _18860_ (_10458_, _10457_, _10444_);
  or _18861_ (_10459_, _10458_, _10456_);
  or _18862_ (_10460_, _10448_, _09191_);
  and _18863_ (_09755_, _10460_, _10459_);
  and _18864_ (_10461_, _10433_, word_in[2]);
  and _18865_ (_10462_, _10435_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  or _18866_ (_10463_, _10462_, _10461_);
  and _18867_ (_10464_, _10463_, _10432_);
  and _18868_ (_10465_, _10431_, word_in[10]);
  or _18869_ (_10466_, _10465_, _10464_);
  and _18870_ (_10467_, _10466_, _10429_);
  and _18871_ (_10468_, _10428_, word_in[18]);
  or _18872_ (_10469_, _10468_, _10444_);
  or _18873_ (_10470_, _10469_, _10467_);
  or _18874_ (_10471_, _10448_, _09204_);
  and _18875_ (_09758_, _10471_, _10470_);
  and _18876_ (_10472_, _10433_, word_in[3]);
  and _18877_ (_10473_, _10435_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  or _18878_ (_10474_, _10473_, _10472_);
  and _18879_ (_10475_, _10474_, _10432_);
  and _18880_ (_10476_, _10431_, word_in[11]);
  or _18881_ (_10477_, _10476_, _10475_);
  and _18882_ (_10478_, _10477_, _10429_);
  and _18883_ (_10479_, _10428_, word_in[19]);
  or _18884_ (_10480_, _10479_, _10444_);
  or _18885_ (_10481_, _10480_, _10478_);
  or _18886_ (_10482_, _10448_, _09218_);
  and _18887_ (_09760_, _10482_, _10481_);
  and _18888_ (_10483_, _10433_, word_in[4]);
  and _18889_ (_10484_, _10435_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  or _18890_ (_10485_, _10484_, _10483_);
  and _18891_ (_10486_, _10485_, _10432_);
  and _18892_ (_10487_, _10431_, word_in[12]);
  or _18893_ (_10488_, _10487_, _10486_);
  and _18894_ (_10489_, _10488_, _10429_);
  and _18895_ (_10490_, _10428_, word_in[20]);
  or _18896_ (_10491_, _10490_, _10444_);
  or _18897_ (_10492_, _10491_, _10489_);
  or _18898_ (_10493_, _10448_, _09236_);
  and _18899_ (_09762_, _10493_, _10492_);
  and _18900_ (_10494_, _10433_, word_in[5]);
  and _18901_ (_10495_, _10435_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  or _18902_ (_10496_, _10495_, _10494_);
  and _18903_ (_10497_, _10496_, _10432_);
  and _18904_ (_10498_, _10431_, word_in[13]);
  or _18905_ (_10499_, _10498_, _10497_);
  and _18906_ (_10500_, _10499_, _10429_);
  and _18907_ (_10501_, _10428_, word_in[21]);
  or _18908_ (_10502_, _10501_, _10444_);
  or _18909_ (_10503_, _10502_, _10500_);
  or _18910_ (_10504_, _10448_, _09251_);
  and _18911_ (_09765_, _10504_, _10503_);
  and _18912_ (_10505_, _10435_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  and _18913_ (_10506_, _10433_, word_in[6]);
  or _18914_ (_10507_, _10506_, _10505_);
  and _18915_ (_10508_, _10507_, _10432_);
  and _18916_ (_10509_, _10431_, word_in[14]);
  or _18917_ (_10510_, _10509_, _10508_);
  and _18918_ (_10511_, _10510_, _10429_);
  and _18919_ (_10512_, _10428_, word_in[22]);
  or _18920_ (_10513_, _10512_, _10444_);
  or _18921_ (_10514_, _10513_, _10511_);
  or _18922_ (_10515_, _10448_, _09267_);
  and _18923_ (_09769_, _10515_, _10514_);
  nor _18924_ (_10516_, _10433_, _08486_);
  and _18925_ (_10517_, _10433_, word_in[7]);
  or _18926_ (_10518_, _10517_, _10516_);
  and _18927_ (_10519_, _10518_, _10432_);
  and _18928_ (_10520_, _10431_, word_in[15]);
  or _18929_ (_10521_, _10520_, _10519_);
  and _18930_ (_10522_, _10521_, _10429_);
  and _18931_ (_10523_, _10428_, word_in[23]);
  or _18932_ (_10524_, _10523_, _10444_);
  or _18933_ (_10525_, _10524_, _10522_);
  or _18934_ (_10526_, _10448_, _08672_);
  and _18935_ (_09772_, _10526_, _10525_);
  and _18936_ (_10527_, _10443_, _08390_);
  and _18937_ (_10528_, _09294_, _08643_);
  not _18938_ (_10529_, _10528_);
  or _18939_ (_10530_, _10529_, _09311_);
  and _18940_ (_10531_, _09298_, _08480_);
  and _18941_ (_10532_, _09300_, _08654_);
  not _18942_ (_10533_, _10532_);
  and _18943_ (_10534_, _10533_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  and _18944_ (_10535_, _10532_, word_in[0]);
  or _18945_ (_10536_, _10535_, _10534_);
  or _18946_ (_10537_, _10536_, _10531_);
  not _18947_ (_10538_, _10531_);
  or _18948_ (_10539_, _10538_, word_in[8]);
  and _18949_ (_10540_, _10539_, _10537_);
  or _18950_ (_10541_, _10540_, _10528_);
  and _18951_ (_10542_, _10541_, _10530_);
  or _18952_ (_10543_, _10542_, _10527_);
  not _18953_ (_10544_, _10527_);
  or _18954_ (_10545_, _10544_, word_in[24]);
  and _18955_ (_13869_, _10545_, _10543_);
  or _18956_ (_10546_, _10529_, _09316_);
  or _18957_ (_10547_, _10532_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  or _18958_ (_10548_, _10533_, word_in[1]);
  and _18959_ (_10549_, _10548_, _10547_);
  or _18960_ (_10550_, _10549_, _10531_);
  or _18961_ (_10551_, _10538_, word_in[9]);
  and _18962_ (_10552_, _10551_, _10550_);
  or _18963_ (_10553_, _10552_, _10528_);
  and _18964_ (_10554_, _10553_, _10546_);
  or _18965_ (_10555_, _10554_, _10527_);
  or _18966_ (_10556_, _10544_, word_in[25]);
  and _18967_ (_09832_, _10556_, _10555_);
  or _18968_ (_10557_, _10529_, _09335_);
  or _18969_ (_10558_, _10532_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  or _18970_ (_10559_, _10533_, word_in[2]);
  and _18971_ (_10560_, _10559_, _10558_);
  or _18972_ (_10561_, _10560_, _10531_);
  or _18973_ (_10562_, _10538_, word_in[10]);
  and _18974_ (_10563_, _10562_, _10561_);
  or _18975_ (_10564_, _10563_, _10528_);
  and _18976_ (_10565_, _10564_, _10557_);
  or _18977_ (_10566_, _10565_, _10527_);
  or _18978_ (_10567_, _10544_, word_in[26]);
  and _18979_ (_09836_, _10567_, _10566_);
  and _18980_ (_10568_, _10533_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  and _18981_ (_10569_, _10532_, word_in[3]);
  nor _18982_ (_10570_, _10569_, _10568_);
  nor _18983_ (_10571_, _10570_, _10531_);
  and _18984_ (_10572_, _10531_, word_in[11]);
  or _18985_ (_10573_, _10572_, _10571_);
  and _18986_ (_10574_, _10573_, _10529_);
  and _18987_ (_10575_, _10528_, _09340_);
  or _18988_ (_10576_, _10575_, _10527_);
  or _18989_ (_10577_, _10576_, _10574_);
  or _18990_ (_10578_, _10544_, word_in[27]);
  and _18991_ (_09840_, _10578_, _10577_);
  and _18992_ (_10579_, _10533_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  and _18993_ (_10580_, _10532_, word_in[4]);
  nor _18994_ (_10581_, _10580_, _10579_);
  nor _18995_ (_10582_, _10581_, _10531_);
  and _18996_ (_10583_, _10531_, word_in[12]);
  or _18997_ (_10584_, _10583_, _10582_);
  and _18998_ (_10585_, _10584_, _10529_);
  and _18999_ (_10586_, _10528_, _09359_);
  or _19000_ (_10587_, _10586_, _10527_);
  or _19001_ (_10588_, _10587_, _10585_);
  or _19002_ (_10589_, _10544_, word_in[28]);
  and _19003_ (_09842_, _10589_, _10588_);
  and _19004_ (_10590_, _10533_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  and _19005_ (_10591_, _10532_, word_in[5]);
  nor _19006_ (_10592_, _10591_, _10590_);
  nor _19007_ (_10593_, _10592_, _10531_);
  and _19008_ (_10594_, _10531_, word_in[13]);
  or _19009_ (_10595_, _10594_, _10593_);
  and _19010_ (_10596_, _10595_, _10529_);
  and _19011_ (_10597_, _10528_, _09364_);
  or _19012_ (_10598_, _10597_, _10527_);
  or _19013_ (_10599_, _10598_, _10596_);
  or _19014_ (_10600_, _10544_, word_in[29]);
  and _19015_ (_09845_, _10600_, _10599_);
  and _19016_ (_10601_, _10533_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  and _19017_ (_10602_, _10532_, word_in[6]);
  nor _19018_ (_10603_, _10602_, _10601_);
  nor _19019_ (_10605_, _10603_, _10531_);
  and _19020_ (_10606_, _10531_, word_in[14]);
  or _19021_ (_10607_, _10606_, _10605_);
  and _19022_ (_10608_, _10607_, _10529_);
  and _19023_ (_10609_, _10528_, _09383_);
  or _19024_ (_10610_, _10609_, _10527_);
  or _19025_ (_10611_, _10610_, _10608_);
  or _19026_ (_10612_, _10544_, word_in[30]);
  and _19027_ (_09847_, _10612_, _10611_);
  nor _19028_ (_10613_, _10532_, _08323_);
  and _19029_ (_10614_, _10532_, word_in[7]);
  nor _19030_ (_10615_, _10614_, _10613_);
  nor _19031_ (_10616_, _10615_, _10531_);
  and _19032_ (_10617_, _10531_, word_in[15]);
  or _19033_ (_10618_, _10617_, _10616_);
  and _19034_ (_10619_, _10618_, _10529_);
  and _19035_ (_10620_, _10528_, _08667_);
  or _19036_ (_10621_, _10620_, _10527_);
  or _19037_ (_10622_, _10621_, _10619_);
  or _19038_ (_10624_, _10544_, word_in[31]);
  and _19039_ (_09850_, _10624_, _10622_);
  and _19040_ (_10626_, _08007_, _06766_);
  and _19041_ (_10627_, _08989_, _08013_);
  and _19042_ (_10629_, _10627_, _10626_);
  nand _19043_ (_10630_, _10629_, _06811_);
  and _19044_ (_10632_, _06770_, _06054_);
  and _19045_ (_10633_, _08989_, _10632_);
  and _19046_ (_10635_, _10633_, _10626_);
  not _19047_ (_10636_, _10635_);
  and _19048_ (_10638_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  nor _19049_ (_10639_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and _19050_ (_10641_, _10639_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and _19051_ (_10642_, _10641_, _10638_);
  not _19052_ (_10643_, _10642_);
  and _19053_ (_10644_, _10643_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and _19054_ (_10645_, _10642_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or _19055_ (_10646_, _10645_, _10644_);
  or _19056_ (_10647_, _10629_, _10646_);
  and _19057_ (_10648_, _10647_, _10636_);
  and _19058_ (_10649_, _10648_, _10630_);
  and _19059_ (_10650_, _10635_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  or _19060_ (_10651_, _10650_, _10649_);
  and _19061_ (_09910_, _10651_, _05552_);
  and _19062_ (_10652_, _09401_, _08643_);
  not _19063_ (_10653_, _10652_);
  and _19064_ (_10654_, _09405_, _08480_);
  not _19065_ (_10655_, _10654_);
  and _19066_ (_10656_, _09410_, _08654_);
  not _19067_ (_10657_, _10656_);
  and _19068_ (_10658_, _10657_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and _19069_ (_10659_, _10656_, word_in[0]);
  or _19070_ (_10660_, _10659_, _10658_);
  and _19071_ (_10661_, _10660_, _10655_);
  and _19072_ (_10662_, _10654_, word_in[8]);
  or _19073_ (_10663_, _10662_, _10661_);
  and _19074_ (_10664_, _10663_, _10653_);
  and _19075_ (_10665_, _10443_, _08392_);
  and _19076_ (_10666_, _10652_, _09311_);
  or _19077_ (_10667_, _10666_, _10665_);
  or _19078_ (_10668_, _10667_, _10664_);
  not _19079_ (_10669_, _10665_);
  or _19080_ (_10670_, _10669_, word_in[24]);
  and _19081_ (_09923_, _10670_, _10668_);
  and _19082_ (_10671_, _10656_, word_in[1]);
  and _19083_ (_10672_, _10657_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  or _19084_ (_10673_, _10672_, _10671_);
  and _19085_ (_10674_, _10673_, _10655_);
  and _19086_ (_10675_, _10654_, word_in[9]);
  or _19087_ (_10676_, _10675_, _10674_);
  and _19088_ (_10677_, _10676_, _10653_);
  and _19089_ (_10678_, _10652_, _09316_);
  or _19090_ (_10679_, _10678_, _10665_);
  or _19091_ (_10680_, _10679_, _10677_);
  or _19092_ (_10681_, _10669_, word_in[25]);
  and _19093_ (_09925_, _10681_, _10680_);
  and _19094_ (_10682_, _10656_, word_in[2]);
  and _19095_ (_10683_, _10657_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  or _19096_ (_10684_, _10683_, _10682_);
  and _19097_ (_10685_, _10684_, _10655_);
  and _19098_ (_10686_, _10654_, word_in[10]);
  or _19099_ (_10687_, _10686_, _10685_);
  and _19100_ (_10688_, _10687_, _10653_);
  and _19101_ (_10689_, _10652_, _09335_);
  or _19102_ (_10690_, _10689_, _10688_);
  and _19103_ (_10691_, _10690_, _10669_);
  and _19104_ (_10692_, _10665_, word_in[26]);
  or _19105_ (_09926_, _10692_, _10691_);
  and _19106_ (_10694_, _10657_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  and _19107_ (_10696_, _10656_, word_in[3]);
  or _19108_ (_10697_, _10696_, _10694_);
  and _19109_ (_10698_, _10697_, _10655_);
  and _19110_ (_10699_, _10654_, word_in[11]);
  or _19111_ (_10700_, _10699_, _10698_);
  and _19112_ (_10701_, _10700_, _10653_);
  and _19113_ (_10702_, _10652_, _09340_);
  or _19114_ (_10703_, _10702_, _10665_);
  or _19115_ (_10704_, _10703_, _10701_);
  or _19116_ (_10705_, _10669_, word_in[27]);
  and _19117_ (_09929_, _10705_, _10704_);
  and _19118_ (_10706_, _10657_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  and _19119_ (_10707_, _10656_, word_in[4]);
  or _19120_ (_10708_, _10707_, _10706_);
  and _19121_ (_10709_, _10708_, _10655_);
  and _19122_ (_10710_, _10654_, word_in[12]);
  or _19123_ (_10711_, _10710_, _10709_);
  and _19124_ (_10712_, _10711_, _10653_);
  and _19125_ (_10713_, _10652_, _09359_);
  or _19126_ (_10714_, _10713_, _10665_);
  or _19127_ (_10715_, _10714_, _10712_);
  or _19128_ (_10716_, _10669_, word_in[28]);
  and _19129_ (_09932_, _10716_, _10715_);
  or _19130_ (_10717_, _10653_, _09364_);
  or _19131_ (_10718_, _10656_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  or _19132_ (_10719_, _10657_, word_in[5]);
  and _19133_ (_10720_, _10719_, _10718_);
  or _19134_ (_10721_, _10720_, _10654_);
  nand _19135_ (_10722_, _10654_, _09584_);
  and _19136_ (_10723_, _10722_, _10721_);
  or _19137_ (_10724_, _10723_, _10652_);
  and _19138_ (_10725_, _10724_, _10717_);
  or _19139_ (_10726_, _10725_, _10665_);
  or _19140_ (_10727_, _10669_, word_in[29]);
  and _19141_ (_09935_, _10727_, _10726_);
  and _19142_ (_10728_, _10656_, word_in[6]);
  and _19143_ (_10729_, _10657_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  or _19144_ (_10730_, _10729_, _10728_);
  and _19145_ (_10732_, _10730_, _10655_);
  and _19146_ (_10733_, _10654_, word_in[14]);
  or _19147_ (_10734_, _10733_, _10732_);
  and _19148_ (_10735_, _10734_, _10653_);
  and _19149_ (_10736_, _10652_, _09383_);
  or _19150_ (_10737_, _10736_, _10665_);
  or _19151_ (_10738_, _10737_, _10735_);
  or _19152_ (_10739_, _10669_, word_in[30]);
  and _19153_ (_09939_, _10739_, _10738_);
  nor _19154_ (_10740_, _10656_, _08481_);
  and _19155_ (_10741_, _10656_, word_in[7]);
  or _19156_ (_10742_, _10741_, _10740_);
  or _19157_ (_10743_, _10742_, _10654_);
  nand _19158_ (_10744_, _10654_, _09281_);
  and _19159_ (_10745_, _10744_, _10743_);
  or _19160_ (_10746_, _10745_, _10652_);
  or _19161_ (_10747_, _10653_, _08667_);
  and _19162_ (_10748_, _10747_, _10746_);
  or _19163_ (_10749_, _10748_, _10665_);
  or _19164_ (_10750_, _10669_, word_in[31]);
  and _19165_ (_09941_, _10750_, _10749_);
  not _19166_ (_10751_, _08655_);
  and _19167_ (_10752_, _10751_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  and _19168_ (_10753_, _08655_, word_in[0]);
  nor _19169_ (_10754_, _10753_, _10752_);
  nor _19170_ (_10755_, _10754_, _08650_);
  and _19171_ (_10756_, _08650_, word_in[8]);
  or _19172_ (_10757_, _10756_, _10755_);
  and _19173_ (_10758_, _10757_, _08647_);
  and _19174_ (_10759_, _09311_, _08646_);
  or _19175_ (_10760_, _10759_, _08666_);
  or _19176_ (_10761_, _10760_, _10758_);
  or _19177_ (_10762_, _08671_, word_in[24]);
  and _19178_ (_13870_, _10762_, _10761_);
  and _19179_ (_10763_, _10751_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  and _19180_ (_10764_, _08655_, word_in[1]);
  nor _19181_ (_10765_, _10764_, _10763_);
  nor _19182_ (_10766_, _10765_, _08650_);
  and _19183_ (_10767_, _08650_, word_in[9]);
  or _19184_ (_10768_, _10767_, _10766_);
  and _19185_ (_10769_, _10768_, _08647_);
  and _19186_ (_10770_, _09316_, _08646_);
  or _19187_ (_10771_, _10770_, _08666_);
  or _19188_ (_10772_, _10771_, _10769_);
  or _19189_ (_10773_, _08671_, word_in[25]);
  and _19190_ (_13871_, _10773_, _10772_);
  and _19191_ (_10774_, _10751_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  and _19192_ (_10775_, _08655_, word_in[2]);
  nor _19193_ (_10776_, _10775_, _10774_);
  nor _19194_ (_10777_, _10776_, _08650_);
  and _19195_ (_10778_, _08650_, word_in[10]);
  or _19196_ (_10779_, _10778_, _10777_);
  and _19197_ (_10780_, _10779_, _08647_);
  and _19198_ (_10781_, _09335_, _08646_);
  or _19199_ (_10782_, _10781_, _08666_);
  or _19200_ (_10783_, _10782_, _10780_);
  or _19201_ (_10784_, _08671_, word_in[26]);
  and _19202_ (_13872_, _10784_, _10783_);
  and _19203_ (_10785_, _10751_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  and _19204_ (_10786_, _08655_, word_in[3]);
  nor _19205_ (_10787_, _10786_, _10785_);
  nor _19206_ (_10788_, _10787_, _08650_);
  and _19207_ (_10789_, _08650_, word_in[11]);
  or _19208_ (_10790_, _10789_, _10788_);
  and _19209_ (_10791_, _10790_, _08647_);
  and _19210_ (_10792_, _09340_, _08646_);
  or _19211_ (_10793_, _10792_, _08666_);
  or _19212_ (_10794_, _10793_, _10791_);
  or _19213_ (_10795_, _08671_, word_in[27]);
  and _19214_ (_13873_, _10795_, _10794_);
  and _19215_ (_10796_, _10751_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  and _19216_ (_10797_, _08655_, word_in[4]);
  nor _19217_ (_10798_, _10797_, _10796_);
  nor _19218_ (_10799_, _10798_, _08650_);
  and _19219_ (_10800_, _08650_, word_in[12]);
  or _19220_ (_10801_, _10800_, _10799_);
  and _19221_ (_10802_, _10801_, _08647_);
  and _19222_ (_10803_, _09359_, _08646_);
  or _19223_ (_10804_, _10803_, _08666_);
  or _19224_ (_10805_, _10804_, _10802_);
  or _19225_ (_10806_, _08671_, word_in[28]);
  and _19226_ (_13874_, _10806_, _10805_);
  or _19227_ (_10808_, _09364_, _08647_);
  or _19228_ (_10809_, _08655_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  or _19229_ (_10811_, _10751_, word_in[5]);
  and _19230_ (_10812_, _10811_, _10809_);
  or _19231_ (_10814_, _10812_, _08650_);
  nand _19232_ (_10815_, _08650_, _09584_);
  and _19233_ (_10817_, _10815_, _10814_);
  or _19234_ (_10818_, _10817_, _08646_);
  and _19235_ (_10819_, _10818_, _10808_);
  or _19236_ (_10820_, _10819_, _08666_);
  or _19237_ (_10821_, _08671_, word_in[29]);
  and _19238_ (_13875_, _10821_, _10820_);
  and _19239_ (_10822_, _10751_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  and _19240_ (_10823_, _08655_, word_in[6]);
  nor _19241_ (_10824_, _10823_, _10822_);
  nor _19242_ (_10825_, _10824_, _08650_);
  and _19243_ (_10826_, _08650_, word_in[14]);
  or _19244_ (_10827_, _10826_, _10825_);
  and _19245_ (_10828_, _10827_, _08647_);
  and _19246_ (_10829_, _09383_, _08646_);
  or _19247_ (_10830_, _10829_, _08666_);
  or _19248_ (_10831_, _10830_, _10828_);
  or _19249_ (_10832_, _08671_, word_in[30]);
  and _19250_ (_13876_, _10832_, _10831_);
  and _19251_ (_10833_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  nor _19252_ (_10834_, _05550_, _05677_);
  or _19253_ (_10835_, _10834_, _10833_);
  and _19254_ (_10033_, _10835_, _05552_);
  and _19255_ (_10836_, _08009_, _10632_);
  nand _19256_ (_10837_, _10836_, _06763_);
  or _19257_ (_10838_, _10836_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and _19258_ (_10839_, _10838_, _06532_);
  and _19259_ (_10841_, _10839_, _10837_);
  or _19260_ (_10842_, _10841_, _06561_);
  and _19261_ (_10119_, _10842_, _05552_);
  and _19262_ (_10843_, _05715_, _05819_);
  and _19263_ (_10844_, _10843_, _05737_);
  and _19264_ (_10845_, _10844_, _05837_);
  and _19265_ (_10846_, _05875_, _05827_);
  and _19266_ (_10847_, _10843_, _05809_);
  or _19267_ (_10848_, _10847_, _10846_);
  or _19268_ (_10849_, _10848_, _10845_);
  and _19269_ (_10850_, _05851_, _05738_);
  and _19270_ (_10851_, _10843_, _05814_);
  or _19271_ (_10852_, _10851_, _10850_);
  or _19272_ (_10853_, _10852_, _10849_);
  or _19273_ (_10854_, _10853_, _05889_);
  and _19274_ (_10855_, _10854_, _05547_);
  and _19275_ (_10856_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _19276_ (_10857_, _10856_, _10855_);
  or _19277_ (_10858_, _10857_, _05902_);
  and _19278_ (_10247_, _10858_, _05552_);
  not _19279_ (_10859_, _06775_);
  nor _19280_ (_10860_, _10859_, _06020_);
  and _19281_ (_10861_, _10860_, _07443_);
  nand _19282_ (_10862_, _10861_, _06030_);
  and _19283_ (_10863_, _10862_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or _19284_ (_10864_, _10863_, _08991_);
  nand _19285_ (_10865_, _06030_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  nor _19286_ (_10866_, _10865_, _08364_);
  or _19287_ (_10867_, _10866_, _08367_);
  and _19288_ (_10868_, _10867_, _10861_);
  or _19289_ (_10869_, _10868_, _10864_);
  nand _19290_ (_10870_, _08991_, _08386_);
  and _19291_ (_10871_, _10870_, _05552_);
  and _19292_ (_10254_, _10871_, _10869_);
  and _19293_ (_10872_, _10861_, _06771_);
  nand _19294_ (_10873_, _10872_, _06763_);
  nor _19295_ (_10874_, _06326_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf );
  nand _19296_ (_10875_, _09010_, _09006_);
  or _19297_ (_10876_, _10875_, _09002_);
  and _19298_ (_10877_, _10876_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or _19299_ (_10878_, _10877_, _10874_);
  or _19300_ (_10879_, _10878_, _10872_);
  and _19301_ (_10880_, _10879_, _10873_);
  or _19302_ (_10881_, _10880_, _08991_);
  nand _19303_ (_10882_, _08991_, _06811_);
  and _19304_ (_10883_, _10882_, _05552_);
  and _19305_ (_10257_, _10883_, _10881_);
  nor _19306_ (_10884_, _09153_, _09086_);
  nor _19307_ (_10885_, _10884_, _09154_);
  or _19308_ (_10886_, _10885_, _09039_);
  or _19309_ (_10887_, _09038_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and _19310_ (_10888_, _10887_, _05605_);
  and _19311_ (_10890_, _10888_, _10886_);
  and _19312_ (_10891_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or _19313_ (_10892_, _10891_, _10890_);
  and _19314_ (_10263_, _10892_, _05552_);
  and _19315_ (_10893_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  nor _19316_ (_10894_, _05550_, _05611_);
  or _19317_ (_10895_, _10894_, _10893_);
  and _19318_ (_10269_, _10895_, _05552_);
  and _19319_ (_10896_, _05894_, _05830_);
  and _19320_ (_10897_, _06567_, _05808_);
  and _19321_ (_10898_, _05715_, _05646_);
  and _19322_ (_10899_, _10898_, _05840_);
  or _19323_ (_10901_, _10899_, _10897_);
  or _19324_ (_10902_, _10901_, _10896_);
  not _19325_ (_10904_, _05716_);
  and _19326_ (_10905_, _05808_, _05760_);
  nor _19327_ (_10906_, _10905_, _05877_);
  nor _19328_ (_10907_, _10906_, _10904_);
  nor _19329_ (_10908_, _10906_, _05714_);
  and _19330_ (_10909_, _05852_, _05738_);
  and _19331_ (_10910_, _10909_, _06567_);
  or _19332_ (_10911_, _10910_, _10908_);
  or _19333_ (_10912_, _10911_, _10907_);
  and _19334_ (_10913_, _05850_, _05840_);
  or _19335_ (_10914_, _05896_, _05878_);
  or _19336_ (_10915_, _10914_, _10913_);
  and _19337_ (_10917_, _05853_, _05737_);
  and _19338_ (_10918_, _06567_, _10917_);
  or _19339_ (_10919_, _10918_, _05838_);
  or _19340_ (_10920_, _10919_, _10915_);
  or _19341_ (_10921_, _10920_, _10912_);
  or _19342_ (_10922_, _10921_, _10902_);
  nand _19343_ (_10923_, _05894_, _05828_);
  not _19344_ (_10924_, _10923_);
  and _19345_ (_10925_, _05827_, _05815_);
  nor _19346_ (_10926_, _10925_, _10924_);
  not _19347_ (_10927_, _10926_);
  and _19348_ (_10929_, _05894_, _06569_);
  or _19349_ (_10930_, _10929_, _10927_);
  and _19350_ (_10931_, _05894_, _05810_);
  or _19351_ (_10932_, _05846_, _05824_);
  and _19352_ (_10933_, _10932_, _05894_);
  or _19353_ (_10934_, _10933_, _10931_);
  or _19354_ (_10935_, _10934_, _05897_);
  or _19355_ (_10936_, _10935_, _10930_);
  and _19356_ (_10937_, _10843_, _05877_);
  and _19357_ (_10938_, _05737_, _05820_);
  and _19358_ (_10939_, _10938_, _05839_);
  and _19359_ (_10940_, _10905_, _10843_);
  or _19360_ (_10941_, _10940_, _10939_);
  or _19361_ (_10942_, _10941_, _10937_);
  and _19362_ (_10943_, _10843_, _05840_);
  or _19363_ (_10944_, _10943_, _06569_);
  or _19364_ (_10945_, _10938_, _10844_);
  and _19365_ (_10946_, _10945_, _10944_);
  and _19366_ (_10947_, _06568_, _05737_);
  or _19367_ (_10948_, _10947_, _10946_);
  or _19368_ (_10949_, _10948_, _10942_);
  or _19369_ (_10950_, _10949_, _10936_);
  or _19370_ (_10952_, _10950_, _10922_);
  and _19371_ (_10953_, _10952_, _05547_);
  and _19372_ (_10955_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and _19373_ (_10956_, _06575_, _05893_);
  and _19374_ (_10957_, _05896_, _05545_);
  and _19375_ (_10958_, _05897_, _05545_);
  nor _19376_ (_10959_, _10958_, _10957_);
  nor _19377_ (_10960_, _10959_, _05546_);
  or _19378_ (_10961_, _10960_, _10956_);
  or _19379_ (_10962_, _10961_, _10955_);
  or _19380_ (_10963_, _10962_, _10953_);
  and _19381_ (_10282_, _10963_, _05552_);
  nor _19382_ (_10964_, _09154_, _09078_);
  nor _19383_ (_10965_, _10964_, _09155_);
  or _19384_ (_10966_, _10965_, _09039_);
  or _19385_ (_10967_, _09038_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and _19386_ (_10968_, _10967_, _05605_);
  and _19387_ (_10969_, _10968_, _10966_);
  and _19388_ (_10970_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or _19389_ (_10971_, _10970_, _10969_);
  and _19390_ (_10298_, _10971_, _05552_);
  nor _19391_ (_10972_, _09152_, _09089_);
  nor _19392_ (_10973_, _10972_, _09153_);
  or _19393_ (_10974_, _10973_, _09039_);
  or _19394_ (_10975_, _09038_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _19395_ (_10976_, _10975_, _05605_);
  and _19396_ (_10977_, _10976_, _10974_);
  and _19397_ (_10978_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  or _19398_ (_10979_, _10978_, _10977_);
  and _19399_ (_10302_, _10979_, _05552_);
  nor _19400_ (_10980_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  and _19401_ (_10981_, _10980_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  not _19402_ (_10982_, _10981_);
  or _19403_ (_10983_, _10982_, _08144_);
  or _19404_ (_10984_, _10981_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2]);
  and _19405_ (_10986_, _10984_, _05552_);
  and _19406_ (_10604_, _10986_, _10983_);
  and _19407_ (_10987_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor _19408_ (_10988_, _05550_, _05921_);
  or _19409_ (_10989_, _10988_, _10987_);
  and _19410_ (_10623_, _10989_, _05552_);
  and _19411_ (_10990_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  not _19412_ (_10991_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  nor _19413_ (_10992_, _05550_, _10991_);
  or _19414_ (_10993_, _10992_, _10990_);
  and _19415_ (_10625_, _10993_, _05552_);
  and _19416_ (_10994_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  not _19417_ (_10995_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  nor _19418_ (_10996_, _05550_, _10995_);
  or _19419_ (_10997_, _10996_, _10994_);
  and _19420_ (_10628_, _10997_, _05552_);
  and _19421_ (_10998_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor _19422_ (_10999_, _05550_, _05553_);
  or _19423_ (_11000_, _10999_, _10998_);
  and _19424_ (_10631_, _11000_, _05552_);
  and _19425_ (_11001_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  not _19426_ (_11002_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nor _19427_ (_11003_, _05550_, _11002_);
  or _19428_ (_11004_, _11003_, _11001_);
  and _19429_ (_10634_, _11004_, _05552_);
  and _19430_ (_11005_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  not _19431_ (_11006_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nor _19432_ (_11007_, _05550_, _11006_);
  or _19433_ (_11008_, _11007_, _11005_);
  and _19434_ (_10637_, _11008_, _05552_);
  and _19435_ (_11009_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  nor _19436_ (_11010_, _05550_, _05748_);
  or _19437_ (_11011_, _11010_, _11009_);
  and _19438_ (_10640_, _11011_, _05552_);
  or _19439_ (_11012_, _10918_, _10908_);
  and _19440_ (_11014_, _05878_, _05818_);
  and _19441_ (_11015_, _10898_, _10905_);
  and _19442_ (_11016_, _11015_, _05738_);
  or _19443_ (_11017_, _11016_, _11014_);
  or _19444_ (_11018_, _11017_, _11012_);
  or _19445_ (_11019_, _11018_, _05889_);
  and _19446_ (_11020_, _11015_, _05737_);
  and _19447_ (_11022_, _10898_, _05877_);
  or _19448_ (_11023_, _11022_, _05896_);
  or _19449_ (_11024_, _11023_, _06568_);
  or _19450_ (_11025_, _11024_, _11020_);
  or _19451_ (_11026_, _11025_, _10902_);
  or _19452_ (_11027_, _11026_, _11019_);
  and _19453_ (_11028_, _05894_, _05860_);
  and _19454_ (_11029_, _05894_, _05853_);
  or _19455_ (_11030_, _11029_, _11028_);
  and _19456_ (_11031_, _08761_, _05716_);
  or _19457_ (_11032_, _11031_, _11030_);
  and _19458_ (_11033_, _10938_, _05837_);
  or _19459_ (_11035_, _11033_, _10943_);
  or _19460_ (_11036_, _11035_, _10845_);
  or _19461_ (_11037_, _11036_, _11032_);
  or _19462_ (_11038_, _11037_, _10942_);
  or _19463_ (_11039_, _11038_, _10936_);
  or _19464_ (_11040_, _11039_, _11027_);
  and _19465_ (_11041_, _11040_, _05547_);
  and _19466_ (_11042_, \oc8051_top_1.oc8051_sfr1.wait_data , \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  or _19467_ (_11043_, _11042_, _10961_);
  or _19468_ (_11045_, _11043_, _11041_);
  and _19469_ (_10693_, _11045_, _05552_);
  or _19470_ (_11046_, _10982_, _07483_);
  or _19471_ (_11048_, _10981_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3]);
  and _19472_ (_11050_, _11048_, _05552_);
  and _19473_ (_10731_, _11050_, _11046_);
  and _19474_ (_11051_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  not _19475_ (_11052_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  nor _19476_ (_11053_, _05550_, _11052_);
  or _19477_ (_11054_, _11053_, _11051_);
  and _19478_ (_10807_, _11054_, _05552_);
  and _19479_ (_11056_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  not _19480_ (_11057_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  nor _19481_ (_11058_, _05550_, _11057_);
  or _19482_ (_11059_, _11058_, _11056_);
  and _19483_ (_10810_, _11059_, _05552_);
  and _19484_ (_11060_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  not _19485_ (_11061_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nor _19486_ (_11062_, _05550_, _11061_);
  or _19487_ (_11063_, _11062_, _11060_);
  and _19488_ (_10813_, _11063_, _05552_);
  nand _19489_ (_11064_, _07388_, _06949_);
  or _19490_ (_11065_, _06949_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  and _19491_ (_11066_, _11065_, _05552_);
  and _19492_ (_10816_, _11066_, _11064_);
  nor _19493_ (_11067_, _07211_, _06341_);
  and _19494_ (_11068_, _06346_, _07211_);
  or _19495_ (_11069_, _11068_, _11067_);
  and _19496_ (_10840_, _11069_, _05552_);
  and _19497_ (_11070_, _05852_, _05850_);
  and _19498_ (_11071_, _11070_, _05886_);
  not _19499_ (_11072_, _11071_);
  and _19500_ (_11073_, _05850_, _05738_);
  and _19501_ (_11074_, _11073_, _10905_);
  and _19502_ (_11075_, _05850_, _05737_);
  and _19503_ (_11076_, _11075_, _05808_);
  nor _19504_ (_11077_, _11076_, _11074_);
  not _19505_ (_11078_, _11077_);
  and _19506_ (_11079_, _11071_, _05761_);
  nor _19507_ (_11080_, _11079_, _11078_);
  nor _19508_ (_11081_, _11080_, _05892_);
  and _19509_ (_11082_, _11081_, _11072_);
  and _19510_ (_11083_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _19511_ (_11084_, _05546_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not _19512_ (_11085_, _11084_);
  and _19513_ (_11086_, _06567_, _05840_);
  not _19514_ (_11087_, _11086_);
  and _19515_ (_11088_, _05895_, _06567_);
  nor _19516_ (_11089_, _11088_, _10918_);
  and _19517_ (_11090_, _11089_, _11087_);
  and _19518_ (_11091_, _11090_, _05898_);
  nor _19519_ (_11092_, _11091_, _11085_);
  nor _19520_ (_11093_, _11071_, _10960_);
  not _19521_ (_11094_, _11093_);
  nor _19522_ (_11095_, _11094_, _11092_);
  nor _19523_ (_11097_, _11095_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _19524_ (_11098_, _11097_, _11083_);
  and _19525_ (_11099_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  and _19526_ (_11100_, _10905_, _05823_);
  nand _19527_ (_11101_, _11100_, _05885_);
  or _19528_ (_11102_, _11101_, _05884_);
  or _19529_ (_11103_, _10940_, _10937_);
  and _19530_ (_11105_, _05850_, _05846_);
  or _19531_ (_11106_, _11105_, _05876_);
  nor _19532_ (_11107_, _11106_, _11103_);
  not _19533_ (_11108_, _10847_);
  nand _19534_ (_11109_, _10843_, _05828_);
  and _19535_ (_11111_, _11109_, _11108_);
  nor _19536_ (_11112_, _10943_, _10851_);
  and _19537_ (_11113_, _11112_, _11111_);
  or _19538_ (_11114_, _10909_, _06570_);
  and _19539_ (_11115_, _11114_, _10843_);
  nor _19540_ (_11116_, _11115_, _11100_);
  and _19541_ (_11117_, _11116_, _11113_);
  and _19542_ (_11118_, _11117_, _11107_);
  and _19543_ (_11119_, _11090_, _11118_);
  nor _19544_ (_11120_, _11119_, _11085_);
  and _19545_ (_11121_, _10905_, _05738_);
  nand _19546_ (_11122_, _11121_, _05850_);
  and _19547_ (_11123_, _10905_, _05737_);
  and _19548_ (_11124_, _11123_, _05850_);
  nor _19549_ (_11125_, _11124_, _05887_);
  and _19550_ (_11126_, _11125_, _11122_);
  and _19551_ (_11127_, _05859_, _05850_);
  and _19552_ (_11128_, _11127_, _05886_);
  not _19553_ (_11129_, _11128_);
  and _19554_ (_11130_, _11129_, _11126_);
  nor _19555_ (_11131_, _11130_, _05892_);
  not _19556_ (_11132_, _05886_);
  and _19557_ (_11133_, _05853_, _05850_);
  nor _19558_ (_11134_, _11133_, _11127_);
  nor _19559_ (_11135_, _11134_, _11132_);
  not _19560_ (_11136_, _11135_);
  nor _19561_ (_11137_, _11136_, _11131_);
  nor _19562_ (_11138_, _11137_, _11120_);
  and _19563_ (_11139_, _11138_, _11102_);
  nor _19564_ (_11140_, _11139_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _19565_ (_11141_, _11140_, _11099_);
  not _19566_ (_11142_, _11141_);
  and _19567_ (_11144_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  not _19568_ (_11145_, _05816_);
  nor _19569_ (_11147_, _05861_, _05842_);
  and _19570_ (_11148_, _11147_, _11145_);
  and _19571_ (_11149_, _10898_, _05860_);
  and _19572_ (_11150_, _11149_, _05669_);
  and _19573_ (_11151_, _11075_, _05827_);
  or _19574_ (_11152_, _11151_, _11150_);
  and _19575_ (_11153_, _10917_, _05823_);
  and _19576_ (_11154_, _11073_, _05827_);
  or _19577_ (_11155_, _11154_, _11153_);
  or _19578_ (_11157_, _11155_, _05833_);
  nor _19579_ (_11158_, _11157_, _11152_);
  and _19580_ (_11159_, _11158_, _11148_);
  and _19581_ (_11160_, _05857_, _05823_);
  nor _19582_ (_11161_, _11160_, _05878_);
  and _19583_ (_11163_, _11161_, _11077_);
  and _19584_ (_11164_, _05854_, _05716_);
  nor _19585_ (_11166_, _11164_, _05845_);
  and _19586_ (_11167_, _05846_, _05822_);
  and _19587_ (_11169_, _11167_, _05818_);
  nor _19588_ (_11170_, _11169_, _05841_);
  and _19589_ (_11171_, _11170_, _11166_);
  and _19590_ (_11172_, _11171_, _11163_);
  nor _19591_ (_11173_, _11100_, _10907_);
  and _19592_ (_11174_, _05895_, _05823_);
  and _19593_ (_11175_, _05826_, _05815_);
  nor _19594_ (_11176_, _11175_, _11174_);
  and _19595_ (_11177_, _11176_, _11173_);
  and _19596_ (_11178_, _06570_, _05716_);
  not _19597_ (_11179_, _11178_);
  and _19598_ (_11180_, _05895_, _05820_);
  nor _19599_ (_11181_, _11180_, _10846_);
  and _19600_ (_11182_, _11181_, _11179_);
  nor _19601_ (_11183_, _05858_, _05811_);
  and _19602_ (_11185_, _11183_, _05856_);
  and _19603_ (_11186_, _11185_, _11182_);
  and _19604_ (_11187_, _11186_, _11177_);
  and _19605_ (_11188_, _11187_, _11172_);
  and _19606_ (_11189_, _11188_, _11159_);
  nor _19607_ (_11190_, _11189_, _11085_);
  nor _19608_ (_11192_, _11190_, _11135_);
  and _19609_ (_11193_, _11192_, _11102_);
  nor _19610_ (_11194_, _11193_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _19611_ (_11195_, _11194_, _11144_);
  and _19612_ (_11196_, _11195_, _11142_);
  and _19613_ (_11197_, _11196_, _11098_);
  and _19614_ (_11198_, _07393_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  and _19615_ (_11199_, _07396_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  nor _19616_ (_11200_, _11199_, _11198_);
  and _19617_ (_11201_, _07400_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  and _19618_ (_11202_, _07403_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  nor _19619_ (_11203_, _11202_, _11201_);
  and _19620_ (_11204_, _11203_, _11200_);
  and _19621_ (_11205_, _07407_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  and _19622_ (_11206_, _07410_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  nor _19623_ (_11207_, _11206_, _11205_);
  and _19624_ (_11208_, _07413_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  and _19625_ (_11209_, _07416_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  nor _19626_ (_11210_, _11209_, _11208_);
  and _19627_ (_11211_, _11210_, _11207_);
  and _19628_ (_11212_, _11211_, _11204_);
  nor _19629_ (_11213_, _11212_, _07437_);
  not _19630_ (_11214_, _06560_);
  and _19631_ (_11216_, _07437_, _11214_);
  nor _19632_ (_11217_, _11216_, _11213_);
  not _19633_ (_11218_, _11217_);
  and _19634_ (_11219_, _11218_, _11197_);
  not _19635_ (_11220_, _11219_);
  nor _19636_ (_11221_, _11195_, _11141_);
  and _19637_ (_11222_, _11098_, _11221_);
  and _19638_ (_11223_, _07443_, _06057_);
  and _19639_ (_11224_, _11223_, _06524_);
  not _19640_ (_11225_, _11224_);
  nor _19641_ (_11226_, _11225_, _06560_);
  and _19642_ (_11227_, _11225_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor _19643_ (_11228_, _11226_, _11227_);
  and _19644_ (_11230_, _11225_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor _19645_ (_11231_, _11225_, _08041_);
  nor _19646_ (_11232_, _11231_, _11230_);
  and _19647_ (_11233_, _11225_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  not _19648_ (_11234_, _07975_);
  and _19649_ (_11235_, _11224_, _11234_);
  nor _19650_ (_11236_, _11235_, _11233_);
  nor _19651_ (_11237_, _11224_, _06025_);
  not _19652_ (_11238_, _07945_);
  and _19653_ (_11239_, _11224_, _11238_);
  nor _19654_ (_11240_, _11239_, _11237_);
  and _19655_ (_11241_, _11240_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and _19656_ (_11242_, _11241_, _11236_);
  and _19657_ (_11243_, _11242_, _11232_);
  and _19658_ (_11244_, _11243_, _11228_);
  nor _19659_ (_11245_, _11243_, _11228_);
  nor _19660_ (_11246_, _11245_, _11244_);
  nor _19661_ (_11247_, _11246_, _05936_);
  nor _19662_ (_11248_, _11247_, _06012_);
  nor _19663_ (_11249_, _11248_, _11224_);
  nor _19664_ (_11250_, _11249_, _11226_);
  not _19665_ (_11251_, _11250_);
  and _19666_ (_11252_, _11251_, _11222_);
  not _19667_ (_11253_, _11252_);
  not _19668_ (_11254_, _06562_);
  and _19669_ (_11255_, _11098_, _11141_);
  and _19670_ (_11256_, _11255_, _11195_);
  and _19671_ (_11257_, _11256_, _11254_);
  not _19672_ (_11258_, _11195_);
  and _19673_ (_11260_, _11255_, _11258_);
  nor _19674_ (_11261_, _05547_, _06165_);
  nor _19675_ (_11262_, _05616_, _05699_);
  and _19676_ (_11263_, _05632_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor _19677_ (_11264_, _11263_, _11262_);
  and _19678_ (_11265_, _05619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and _19679_ (_11266_, _05627_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor _19680_ (_11267_, _11266_, _11265_);
  nor _19681_ (_11268_, _05613_, _11002_);
  nor _19682_ (_11269_, _05624_, _05695_);
  nor _19683_ (_11270_, _11269_, _11268_);
  and _19684_ (_11271_, _11270_, _11267_);
  and _19685_ (_11272_, _11271_, _11264_);
  nor _19686_ (_11273_, _11272_, _09039_);
  nor _19687_ (_11274_, _11273_, _11261_);
  not _19688_ (_11275_, _11274_);
  and _19689_ (_11276_, _11275_, _11260_);
  nor _19690_ (_11277_, _11276_, _11257_);
  and _19691_ (_11278_, _11277_, _11253_);
  and _19692_ (_11279_, _11278_, _11220_);
  nor _19693_ (_11280_, _11279_, _06064_);
  and _19694_ (_11281_, _11279_, _06064_);
  nor _19695_ (_11282_, _11281_, _11280_);
  and _19696_ (_11283_, _11224_, _06811_);
  and _19697_ (_11284_, _11225_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  nor _19698_ (_11285_, _11225_, _07388_);
  nor _19699_ (_11286_, _11285_, _11284_);
  and _19700_ (_11287_, _11286_, _11244_);
  and _19701_ (_11288_, _11225_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor _19702_ (_11289_, _11225_, _06306_);
  nor _19703_ (_11290_, _11289_, _11288_);
  and _19704_ (_11291_, _11290_, _11287_);
  and _19705_ (_11292_, _11225_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor _19706_ (_11294_, _11225_, _08386_);
  nor _19707_ (_11296_, _11294_, _11292_);
  and _19708_ (_11297_, _11296_, _11291_);
  nor _19709_ (_11299_, _11224_, _05959_);
  nor _19710_ (_11300_, _11299_, _11297_);
  and _19711_ (_11301_, _11299_, _11297_);
  or _19712_ (_11303_, _11301_, _11300_);
  nor _19713_ (_11304_, _11303_, _05936_);
  nor _19714_ (_11305_, _11224_, _05963_);
  not _19715_ (_11306_, _11305_);
  nor _19716_ (_11307_, _11306_, _11304_);
  nor _19717_ (_11308_, _11307_, _11283_);
  and _19718_ (_11309_, _11308_, _11221_);
  not _19719_ (_11310_, _11309_);
  nor _19720_ (_11311_, _11195_, _11142_);
  nor _19721_ (_11312_, _05547_, _06359_);
  nor _19722_ (_11313_, _05616_, _05762_);
  nor _19723_ (_11315_, _05631_, _05768_);
  nor _19724_ (_11316_, _11315_, _11313_);
  and _19725_ (_11317_, _05619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and _19726_ (_11318_, _05627_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  nor _19727_ (_11320_, _11318_, _11317_);
  nor _19728_ (_11321_, _05613_, _07743_);
  nor _19729_ (_11322_, _05624_, _05770_);
  nor _19730_ (_11323_, _11322_, _11321_);
  and _19731_ (_11324_, _11323_, _11320_);
  and _19732_ (_11325_, _11324_, _11316_);
  nor _19733_ (_11326_, _11325_, _09039_);
  nor _19734_ (_11327_, _11326_, _11312_);
  not _19735_ (_11328_, _11327_);
  and _19736_ (_11329_, _11328_, _11311_);
  not _19737_ (_11330_, _11098_);
  not _19738_ (_11331_, _07441_);
  and _19739_ (_11332_, _11196_, _11331_);
  or _19740_ (_11333_, _11332_, _11330_);
  nor _19741_ (_11334_, _11333_, _11329_);
  and _19742_ (_11335_, _11334_, _11310_);
  nor _19743_ (_11336_, _11335_, _06911_);
  and _19744_ (_11337_, _11335_, _06911_);
  nor _19745_ (_11338_, _11337_, _11336_);
  nor _19746_ (_11339_, _11296_, _11291_);
  nor _19747_ (_11340_, _11339_, _11297_);
  nor _19748_ (_11341_, _11340_, _05936_);
  nor _19749_ (_11342_, _11341_, _05940_);
  nor _19750_ (_11343_, _11342_, _11224_);
  nor _19751_ (_11344_, _11343_, _11294_);
  not _19752_ (_11345_, _11344_);
  and _19753_ (_11346_, _11345_, _11222_);
  not _19754_ (_11347_, _11346_);
  and _19755_ (_11348_, _07416_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  and _19756_ (_11349_, _07410_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  nor _19757_ (_11351_, _11349_, _11348_);
  and _19758_ (_11352_, _07393_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  and _19759_ (_11353_, _07407_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  nor _19760_ (_11354_, _11353_, _11352_);
  and _19761_ (_11356_, _11354_, _11351_);
  and _19762_ (_11358_, _07400_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  and _19763_ (_11359_, _07396_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  nor _19764_ (_11360_, _11359_, _11358_);
  and _19765_ (_11361_, _07403_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  and _19766_ (_11362_, _07413_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  nor _19767_ (_11363_, _11362_, _11361_);
  and _19768_ (_11364_, _11363_, _11360_);
  and _19769_ (_11365_, _11364_, _11356_);
  nor _19770_ (_11366_, _11365_, _07437_);
  not _19771_ (_11367_, _08386_);
  and _19772_ (_11368_, _11367_, _07437_);
  nor _19773_ (_11370_, _11368_, _11366_);
  not _19774_ (_11371_, _11370_);
  and _19775_ (_11372_, _11371_, _11197_);
  not _19776_ (_11373_, _11372_);
  nor _19777_ (_11374_, _11196_, _11098_);
  nor _19778_ (_11376_, _05547_, _06394_);
  nor _19779_ (_11377_, _05616_, _05786_);
  nor _19780_ (_11378_, _05631_, _05791_);
  nor _19781_ (_11379_, _11378_, _11377_);
  and _19782_ (_11380_, _05619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and _19783_ (_11381_, _05627_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor _19784_ (_11382_, _11381_, _11380_);
  not _19785_ (_11383_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nor _19786_ (_11384_, _05613_, _11383_);
  and _19787_ (_11385_, _05625_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor _19788_ (_11386_, _11385_, _11384_);
  and _19789_ (_11387_, _11386_, _11382_);
  and _19790_ (_11388_, _11387_, _11379_);
  nor _19791_ (_11389_, _11388_, _09039_);
  nor _19792_ (_11390_, _11389_, _11376_);
  not _19793_ (_11391_, _11390_);
  and _19794_ (_11392_, _11391_, _11260_);
  nor _19795_ (_11393_, _11392_, _11374_);
  and _19796_ (_11394_, _11393_, _11373_);
  and _19797_ (_11395_, _11394_, _11347_);
  nor _19798_ (_11396_, _11395_, _06925_);
  and _19799_ (_11397_, _11395_, _06925_);
  nor _19800_ (_11398_, _11397_, _11396_);
  and _19801_ (_11399_, _11398_, _11338_);
  and _19802_ (_11400_, _07400_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  and _19803_ (_11401_, _07413_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  nor _19804_ (_11402_, _11401_, _11400_);
  and _19805_ (_11403_, _07403_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  and _19806_ (_11404_, _07416_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  nor _19807_ (_11405_, _11404_, _11403_);
  and _19808_ (_11406_, _11405_, _11402_);
  and _19809_ (_11407_, _07393_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  and _19810_ (_11408_, _07396_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  nor _19811_ (_11409_, _11408_, _11407_);
  and _19812_ (_11410_, _07407_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  and _19813_ (_11411_, _07410_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  nor _19814_ (_11412_, _11411_, _11410_);
  and _19815_ (_11413_, _11412_, _11409_);
  and _19816_ (_11414_, _11413_, _11406_);
  nor _19817_ (_11415_, _11414_, _07437_);
  and _19818_ (_11416_, _07437_, _06307_);
  nor _19819_ (_11418_, _11416_, _11415_);
  not _19820_ (_11419_, _11418_);
  and _19821_ (_11420_, _11419_, _11197_);
  not _19822_ (_11421_, _11311_);
  and _19823_ (_11422_, _11374_, _11421_);
  nor _19824_ (_11423_, _11422_, _11420_);
  nor _19825_ (_11424_, _11290_, _11287_);
  nor _19826_ (_11425_, _11424_, _11291_);
  nor _19827_ (_11426_, _11425_, _05936_);
  nor _19828_ (_11427_, _11426_, _05993_);
  nor _19829_ (_11428_, _11427_, _11224_);
  nor _19830_ (_11429_, _11428_, _11289_);
  not _19831_ (_11430_, _11429_);
  and _19832_ (_11431_, _11430_, _11222_);
  nor _19833_ (_11432_, _05547_, _06074_);
  nor _19834_ (_11433_, _05616_, _05748_);
  nor _19835_ (_11434_, _05631_, _05743_);
  nor _19836_ (_11436_, _11434_, _11433_);
  and _19837_ (_11437_, _05619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and _19838_ (_11439_, _05627_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor _19839_ (_11440_, _11439_, _11437_);
  not _19840_ (_11441_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  nor _19841_ (_11442_, _05613_, _11441_);
  and _19842_ (_11443_, _05625_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor _19843_ (_11444_, _11443_, _11442_);
  and _19844_ (_11445_, _11444_, _11440_);
  and _19845_ (_11446_, _11445_, _11436_);
  nor _19846_ (_11447_, _11446_, _09039_);
  nor _19847_ (_11448_, _11447_, _11432_);
  not _19848_ (_11449_, _11448_);
  and _19849_ (_11450_, _11449_, _11260_);
  nor _19850_ (_11451_, _11450_, _11431_);
  and _19851_ (_11452_, _11451_, _11423_);
  nor _19852_ (_11453_, _11452_, _06764_);
  and _19853_ (_11454_, _11452_, _06764_);
  nor _19854_ (_11455_, _11454_, _11453_);
  nor _19855_ (_11456_, _05547_, _06143_);
  and _19856_ (_11457_, _05650_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and _19857_ (_11458_, _05632_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor _19858_ (_11459_, _11458_, _11457_);
  and _19859_ (_11460_, _05619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and _19860_ (_11461_, _05627_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  nor _19861_ (_11462_, _11461_, _11460_);
  nor _19862_ (_11463_, _05613_, _11061_);
  and _19863_ (_11464_, _05625_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor _19864_ (_11465_, _11464_, _11463_);
  and _19865_ (_11466_, _11465_, _11462_);
  and _19866_ (_11467_, _11466_, _11459_);
  nor _19867_ (_11468_, _11467_, _09039_);
  nor _19868_ (_11469_, _11468_, _11456_);
  not _19869_ (_11470_, _11469_);
  and _19870_ (_11471_, _11470_, _11260_);
  and _19871_ (_11472_, _11256_, _07391_);
  nor _19872_ (_11473_, _11472_, _11471_);
  and _19873_ (_11474_, _07393_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  and _19874_ (_11475_, _07396_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  nor _19875_ (_11476_, _11475_, _11474_);
  and _19876_ (_11477_, _07400_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  and _19877_ (_11478_, _07413_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  nor _19878_ (_11479_, _11478_, _11477_);
  and _19879_ (_11480_, _11479_, _11476_);
  and _19880_ (_11481_, _07407_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  and _19881_ (_11482_, _07410_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  nor _19882_ (_11483_, _11482_, _11481_);
  and _19883_ (_11484_, _07403_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  and _19884_ (_11485_, _07416_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  nor _19885_ (_11486_, _11485_, _11484_);
  and _19886_ (_11487_, _11486_, _11483_);
  and _19887_ (_11488_, _11487_, _11480_);
  nor _19888_ (_11489_, _11488_, _07437_);
  not _19889_ (_11490_, _07388_);
  and _19890_ (_11491_, _07437_, _11490_);
  nor _19891_ (_11492_, _11491_, _11489_);
  not _19892_ (_11493_, _11492_);
  and _19893_ (_11494_, _11493_, _11197_);
  not _19894_ (_11495_, _11494_);
  nor _19895_ (_11496_, _11286_, _11244_);
  nor _19896_ (_11497_, _11496_, _11287_);
  nor _19897_ (_11499_, _11497_, _05936_);
  nor _19898_ (_11500_, _11499_, _05976_);
  nor _19899_ (_11501_, _11500_, _11224_);
  nor _19900_ (_11502_, _11501_, _11285_);
  not _19901_ (_11503_, _11502_);
  and _19902_ (_11505_, _11503_, _11222_);
  and _19903_ (_11506_, _11330_, _11141_);
  nor _19904_ (_11507_, _11506_, _11505_);
  and _19905_ (_11508_, _11507_, _11495_);
  and _19906_ (_11509_, _11508_, _11473_);
  nor _19907_ (_11510_, _11509_, _06527_);
  and _19908_ (_11511_, _11509_, _06527_);
  nor _19909_ (_11512_, _11511_, _11510_);
  and _19910_ (_11513_, _11512_, _11455_);
  and _19911_ (_11514_, _11513_, _11399_);
  and _19912_ (_11515_, _11514_, _11282_);
  nor _19913_ (_11516_, _06771_, _06967_);
  and _19914_ (_11518_, _11516_, _11515_);
  and _19915_ (_11519_, _11518_, _11082_);
  not _19916_ (_11520_, _11519_);
  not _19917_ (_11521_, _07224_);
  not _19918_ (_11522_, _11131_);
  nor _19919_ (_11523_, _06668_, _06628_);
  and _19920_ (_11524_, _06668_, _06628_);
  nor _19921_ (_11525_, _11524_, _11523_);
  nor _19922_ (_11526_, _07680_, _06654_);
  nand _19923_ (_11527_, _11526_, _08117_);
  nor _19924_ (_11528_, _11527_, _11071_);
  and _19925_ (_11529_, _11528_, _07462_);
  not _19926_ (_11530_, _11529_);
  nor _19927_ (_11531_, _11530_, _11525_);
  and _19928_ (_11532_, _11531_, _07614_);
  and _19929_ (_11533_, _11532_, _11522_);
  and _19930_ (_11534_, _11533_, _07528_);
  and _19931_ (_11535_, _11534_, _11521_);
  and _19932_ (_11536_, _11082_, _06140_);
  and _19933_ (_11537_, _11079_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor _19934_ (_11538_, _11081_, _11072_);
  nor _19935_ (_11539_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor _19936_ (_11540_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and _19937_ (_11541_, _11540_, _11539_);
  nor _19938_ (_11542_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor _19939_ (_11543_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and _19940_ (_11544_, _11543_, _11542_);
  and _19941_ (_11545_, _11544_, _11541_);
  and _19942_ (_11546_, _11545_, _11538_);
  or _19943_ (_11547_, _11546_, _11537_);
  or _19944_ (_11548_, _11547_, _11536_);
  nor _19945_ (_11549_, _11548_, _11535_);
  and _19946_ (_11550_, _10938_, _05814_);
  not _19947_ (_11552_, _11550_);
  nand _19948_ (_11553_, _05846_, _05716_);
  nand _19949_ (_11555_, _05828_, _05716_);
  and _19950_ (_11556_, _11555_, _10923_);
  and _19951_ (_11557_, _11556_, _11553_);
  and _19952_ (_11558_, _11557_, _11552_);
  and _19953_ (_11559_, _10938_, _05827_);
  not _19954_ (_11560_, _11559_);
  and _19955_ (_11561_, _11560_, _11109_);
  or _19956_ (_11562_, _05877_, _10917_);
  nand _19957_ (_11563_, _11562_, _05850_);
  and _19958_ (_11564_, _11563_, _11561_);
  nand _19959_ (_11565_, _11564_, _11558_);
  nor _19960_ (_11566_, _11565_, _11124_);
  not _19961_ (_11567_, _11566_);
  and _19962_ (_11568_, _11567_, _11549_);
  not _19963_ (_11569_, _11568_);
  and _19964_ (_11570_, _05857_, _05850_);
  nor _19965_ (_11571_, _11570_, _10918_);
  not _19966_ (_11572_, _11122_);
  or _19967_ (_11573_, _11572_, _05887_);
  nor _19968_ (_11574_, _11134_, _05737_);
  nor _19969_ (_11575_, _11574_, _11573_);
  or _19970_ (_11576_, _11575_, _11549_);
  and _19971_ (_11577_, _11576_, _11571_);
  and _19972_ (_11578_, _11577_, _11569_);
  nor _19973_ (_11579_, _11578_, _11132_);
  not _19974_ (_11580_, _11101_);
  and _19975_ (_11581_, _05823_, _05809_);
  nor _19976_ (_11582_, _05869_, _11581_);
  nor _19977_ (_11583_, _11085_, _11582_);
  nor _19978_ (_11584_, _11583_, _11580_);
  not _19979_ (_11585_, _11584_);
  nor _19980_ (_11586_, _11585_, _11579_);
  not _19981_ (_11587_, _08935_);
  and _19982_ (_11589_, _11538_, _11587_);
  nor _19983_ (_11590_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  not _19984_ (_11591_, _11590_);
  nor _19985_ (_11592_, _11591_, _08009_);
  and _19986_ (_11593_, _11592_, _06532_);
  not _19987_ (_11594_, _11593_);
  and _19988_ (_11595_, _11594_, _11079_);
  nor _19989_ (_11596_, _11595_, _11589_);
  not _19990_ (_11597_, _11596_);
  nor _19991_ (_11598_, _11597_, _11586_);
  and _19992_ (_11599_, _11196_, _11330_);
  not _19993_ (_11600_, _11599_);
  and _19994_ (_11601_, _11256_, _05819_);
  nor _19995_ (_11602_, _05547_, _06228_);
  nor _19996_ (_11603_, _05616_, _05611_);
  nor _19997_ (_11604_, _05631_, _05615_);
  nor _19998_ (_11605_, _11604_, _11603_);
  and _19999_ (_11606_, _05619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and _20000_ (_11607_, _05627_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor _20001_ (_11608_, _11607_, _11606_);
  not _20002_ (_11609_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor _20003_ (_11610_, _05613_, _11609_);
  and _20004_ (_11611_, _05625_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor _20005_ (_11612_, _11611_, _11610_);
  and _20006_ (_11613_, _11612_, _11608_);
  and _20007_ (_11614_, _11613_, _11605_);
  nor _20008_ (_11615_, _11614_, _09039_);
  nor _20009_ (_11616_, _11615_, _11602_);
  not _20010_ (_11617_, _11616_);
  and _20011_ (_11618_, _11617_, _11260_);
  nor _20012_ (_11619_, _11618_, _11601_);
  and _20013_ (_11620_, _11619_, _11600_);
  nor _20014_ (_11621_, _11241_, _11236_);
  nor _20015_ (_11622_, _11621_, _11242_);
  nor _20016_ (_11623_, _11622_, _05936_);
  nor _20017_ (_11624_, _11623_, _06034_);
  nor _20018_ (_11625_, _11624_, _11224_);
  nor _20019_ (_11626_, _11625_, _11235_);
  not _20020_ (_11627_, _11626_);
  and _20021_ (_11628_, _11627_, _11222_);
  and _20022_ (_11629_, _07400_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  and _20023_ (_11630_, _07407_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  nor _20024_ (_11631_, _11630_, _11629_);
  and _20025_ (_11632_, _07393_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  and _20026_ (_11633_, _07416_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  nor _20027_ (_11634_, _11633_, _11632_);
  and _20028_ (_11635_, _11634_, _11631_);
  and _20029_ (_11636_, _07396_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  and _20030_ (_11637_, _07410_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  nor _20031_ (_11638_, _11637_, _11636_);
  and _20032_ (_11639_, _07403_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  and _20033_ (_11640_, _07413_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  nor _20034_ (_11641_, _11640_, _11639_);
  and _20035_ (_11642_, _11641_, _11638_);
  and _20036_ (_11643_, _11642_, _11635_);
  nor _20037_ (_11644_, _11643_, _07437_);
  and _20038_ (_11645_, _11234_, _07437_);
  nor _20039_ (_11646_, _11645_, _11644_);
  not _20040_ (_11647_, _11646_);
  and _20041_ (_11648_, _11647_, _11197_);
  nor _20042_ (_11649_, _11648_, _11628_);
  and _20043_ (_11650_, _11649_, _11620_);
  nor _20044_ (_11651_, _11650_, _06043_);
  and _20045_ (_11652_, _11650_, _06043_);
  nor _20046_ (_11653_, _11652_, _11651_);
  and _20047_ (_11654_, _07400_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  and _20048_ (_11655_, _07416_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  nor _20049_ (_11656_, _11655_, _11654_);
  and _20050_ (_11657_, _07403_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  and _20051_ (_11658_, _07410_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  nor _20052_ (_11660_, _11658_, _11657_);
  and _20053_ (_11661_, _11660_, _11656_);
  and _20054_ (_11662_, _07413_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  and _20055_ (_11663_, _07407_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  nor _20056_ (_11664_, _11663_, _11662_);
  and _20057_ (_11665_, _07393_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  and _20058_ (_11666_, _07396_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  nor _20059_ (_11667_, _11666_, _11665_);
  and _20060_ (_11668_, _11667_, _11664_);
  and _20061_ (_11669_, _11668_, _11661_);
  nor _20062_ (_11670_, _11669_, _07437_);
  and _20063_ (_11671_, _11238_, _07437_);
  nor _20064_ (_11672_, _11671_, _11670_);
  not _20065_ (_11673_, _11672_);
  and _20066_ (_11674_, _11673_, _11197_);
  nor _20067_ (_11675_, _05547_, _06186_);
  nor _20068_ (_11676_, _05616_, _05656_);
  and _20069_ (_11677_, _05632_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor _20070_ (_11678_, _11677_, _11676_);
  and _20071_ (_11679_, _05619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  nor _20072_ (_11680_, _05624_, _05652_);
  nor _20073_ (_11682_, _11680_, _11679_);
  and _20074_ (_11683_, _05627_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor _20075_ (_11684_, _05613_, _11006_);
  nor _20076_ (_11686_, _11684_, _11683_);
  and _20077_ (_11687_, _11686_, _11682_);
  and _20078_ (_11688_, _11687_, _11678_);
  nor _20079_ (_11689_, _11688_, _09039_);
  nor _20080_ (_11690_, _11689_, _11675_);
  not _20081_ (_11691_, _11690_);
  and _20082_ (_11692_, _11691_, _11260_);
  nor _20083_ (_11693_, _11692_, _11674_);
  nor _20084_ (_11694_, _11240_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  nor _20085_ (_11695_, _11694_, _11241_);
  nor _20086_ (_11696_, _11695_, _05936_);
  nor _20087_ (_11697_, _11696_, _06026_);
  nor _20088_ (_11698_, _11697_, _11224_);
  nor _20089_ (_11699_, _11698_, _11239_);
  not _20090_ (_11700_, _11699_);
  and _20091_ (_11701_, _11700_, _11222_);
  and _20092_ (_11702_, _11256_, _05669_);
  nor _20093_ (_11703_, _11702_, _11701_);
  and _20094_ (_11704_, _11703_, _11693_);
  and _20095_ (_11705_, _11704_, _06031_);
  nor _20096_ (_11706_, _11704_, _06031_);
  or _20097_ (_11707_, _11706_, _11705_);
  nor _20098_ (_11708_, _11707_, _11653_);
  and _20099_ (_11709_, _07407_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  and _20100_ (_11710_, _07410_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  nor _20101_ (_11711_, _11710_, _11709_);
  and _20102_ (_11712_, _07413_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  and _20103_ (_11713_, _07416_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  nor _20104_ (_11714_, _11713_, _11712_);
  and _20105_ (_11715_, _11714_, _11711_);
  and _20106_ (_11716_, _07403_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  and _20107_ (_11717_, _07396_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  nor _20108_ (_11718_, _11717_, _11716_);
  and _20109_ (_11719_, _07400_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  and _20110_ (_11721_, _07393_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  nor _20111_ (_11722_, _11721_, _11719_);
  and _20112_ (_11723_, _11722_, _11718_);
  and _20113_ (_11724_, _11723_, _11715_);
  nor _20114_ (_11725_, _11724_, _07437_);
  not _20115_ (_11726_, _08041_);
  and _20116_ (_11727_, _11726_, _07437_);
  nor _20117_ (_11728_, _11727_, _11725_);
  not _20118_ (_11729_, _11728_);
  and _20119_ (_11730_, _11729_, _11197_);
  nor _20120_ (_11731_, _05547_, _06209_);
  nor _20121_ (_11732_, _05616_, _05677_);
  and _20122_ (_11733_, _05632_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor _20123_ (_11734_, _11733_, _11732_);
  and _20124_ (_11735_, _05619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and _20125_ (_11736_, _05625_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor _20126_ (_11737_, _11736_, _11735_);
  and _20127_ (_11738_, _05627_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  not _20128_ (_11739_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nor _20129_ (_11740_, _05613_, _11739_);
  nor _20130_ (_11742_, _11740_, _11738_);
  and _20131_ (_11743_, _11742_, _11737_);
  and _20132_ (_11744_, _11743_, _11734_);
  nor _20133_ (_11745_, _11744_, _09039_);
  nor _20134_ (_11746_, _11745_, _11731_);
  not _20135_ (_11747_, _11746_);
  and _20136_ (_11749_, _11747_, _11260_);
  nor _20137_ (_11750_, _11749_, _11730_);
  nor _20138_ (_11751_, _11242_, _11232_);
  nor _20139_ (_11752_, _11751_, _11243_);
  nor _20140_ (_11753_, _11752_, _05936_);
  nor _20141_ (_11754_, _11753_, _06046_);
  nor _20142_ (_11756_, _11754_, _11224_);
  nor _20143_ (_11757_, _11756_, _11231_);
  not _20144_ (_11759_, _11757_);
  and _20145_ (_11760_, _11759_, _11222_);
  and _20146_ (_11761_, _11256_, _05693_);
  nor _20147_ (_11762_, _11761_, _11760_);
  and _20148_ (_11763_, _11762_, _11750_);
  nor _20149_ (_11764_, _11763_, _06054_);
  and _20150_ (_11765_, _11763_, _06054_);
  nor _20151_ (_11766_, _11765_, _11764_);
  nor _20152_ (_11767_, _11766_, _06816_);
  and _20153_ (_11768_, _11767_, _11708_);
  and _20154_ (_11769_, _11768_, _11515_);
  nor _20155_ (_11770_, _05971_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and _20156_ (_11771_, _11770_, _11769_);
  not _20157_ (_11772_, _11771_);
  and _20158_ (_11773_, _11772_, _11598_);
  and _20159_ (_11774_, _11773_, _11520_);
  and _20160_ (_11775_, _11557_, _11126_);
  nand _20161_ (_11776_, _11775_, _11561_);
  nand _20162_ (_11777_, _11776_, _05886_);
  and _20163_ (_11778_, _10905_, _11084_);
  and _20164_ (_11779_, _11778_, _05850_);
  and _20165_ (_11780_, _11084_, _11581_);
  nor _20166_ (_11781_, _11780_, _11779_);
  and _20167_ (_11782_, _11781_, _11102_);
  nand _20168_ (_11783_, _11782_, _11777_);
  and _20169_ (_11784_, _10918_, _05886_);
  nor _20170_ (_11785_, _11784_, _11583_);
  nor _20171_ (_11786_, _11785_, _11783_);
  not _20172_ (_11787_, _11786_);
  nor _20173_ (_11788_, _11550_, _11070_);
  nand _20174_ (_11789_, _11788_, _11571_);
  nand _20175_ (_11790_, _11789_, _05886_);
  nand _20176_ (_11791_, _11790_, _11777_);
  nor _20177_ (_11792_, _11791_, _11787_);
  and _20178_ (_11793_, \oc8051_top_1.oc8051_memory_interface1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and _20179_ (_11794_, \oc8051_top_1.oc8051_memory_interface1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and _20180_ (_11795_, _11794_, _11793_);
  and _20181_ (_11796_, \oc8051_top_1.oc8051_memory_interface1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and _20182_ (_11797_, _11796_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and _20183_ (_11799_, \oc8051_top_1.oc8051_memory_interface1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and _20184_ (_11800_, _11799_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and _20185_ (_11801_, _11800_, _11797_);
  and _20186_ (_11802_, _11801_, _11795_);
  and _20187_ (_11803_, _11802_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _20188_ (_11804_, _11803_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _20189_ (_11805_, _11804_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and _20190_ (_11806_, _11805_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  or _20191_ (_11807_, _11806_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nand _20192_ (_11808_, _11806_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and _20193_ (_11809_, _11808_, _11807_);
  and _20194_ (_11810_, _11809_, _11792_);
  not _20195_ (_11811_, _11102_);
  and _20196_ (_11812_, _11811_, _07255_);
  and _20197_ (_11813_, _11784_, _07360_);
  and _20198_ (_11814_, _11780_, _11328_);
  and _20199_ (_11815_, _11782_, _11777_);
  nand _20200_ (_11816_, _11785_, _11815_);
  nor _20201_ (_11817_, _11816_, _11791_);
  and _20202_ (_11818_, _11817_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  or _20203_ (_11819_, _11818_, _11814_);
  or _20204_ (_11820_, _11819_, _11813_);
  or _20205_ (_11821_, _11820_, _11812_);
  nor _20206_ (_11822_, _11821_, _11810_);
  nand _20207_ (_11824_, _11822_, _11774_);
  and _20208_ (_11825_, _11783_, _07758_);
  and _20209_ (_11827_, _11815_, _11327_);
  nor _20210_ (_11828_, _11827_, _11825_);
  nor _20211_ (_11829_, _11828_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and _20212_ (_11830_, _11828_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor _20213_ (_11831_, _05547_, _06482_);
  and _20214_ (_11832_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _20215_ (_11833_, _05616_, _11383_);
  nor _20216_ (_11834_, _05624_, _05791_);
  or _20217_ (_11835_, _11834_, _11833_);
  nor _20218_ (_11836_, _05613_, _05907_);
  nor _20219_ (_11837_, _05631_, _05786_);
  or _20220_ (_11838_, _11837_, _11836_);
  or _20221_ (_11839_, _11838_, _11835_);
  and _20222_ (_11840_, _05619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and _20223_ (_11842_, _05627_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  or _20224_ (_11843_, _11842_, _11840_);
  or _20225_ (_11844_, _11843_, _11839_);
  and _20226_ (_11845_, _11844_, _05671_);
  or _20227_ (_11846_, _11845_, _11832_);
  and _20228_ (_11847_, _11846_, _05547_);
  nor _20229_ (_11848_, _11847_, _11831_);
  and _20230_ (_11849_, _11848_, _11783_);
  and _20231_ (_11850_, _11815_, _11390_);
  nor _20232_ (_11851_, _11850_, _11849_);
  and _20233_ (_11852_, _11851_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor _20234_ (_11853_, _11851_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor _20235_ (_11854_, _11853_, _11852_);
  nor _20236_ (_11855_, _05547_, _06079_);
  and _20237_ (_11856_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _20238_ (_11857_, _05613_, _11057_);
  nor _20239_ (_11858_, _05624_, _05743_);
  nor _20240_ (_11859_, _11858_, _11857_);
  and _20241_ (_11860_, _05619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  nor _20242_ (_11861_, _05631_, _05748_);
  nor _20243_ (_11862_, _11861_, _11860_);
  and _20244_ (_11863_, _05627_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor _20245_ (_11864_, _05616_, _11441_);
  nor _20246_ (_11865_, _11864_, _11863_);
  and _20247_ (_11866_, _11865_, _11862_);
  and _20248_ (_11867_, _11866_, _11859_);
  nor _20249_ (_11868_, _11867_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _20250_ (_11870_, _11868_, _11856_);
  nor _20251_ (_11871_, _11870_, _05548_);
  nor _20252_ (_11872_, _11871_, _11855_);
  and _20253_ (_11873_, _11872_, _11783_);
  and _20254_ (_11874_, _11815_, _11448_);
  nor _20255_ (_11875_, _11874_, _11873_);
  nor _20256_ (_11876_, _11875_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and _20257_ (_11877_, _11875_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nor _20258_ (_11878_, _05547_, _06145_);
  and _20259_ (_11879_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _20260_ (_11881_, _05616_, _11061_);
  and _20261_ (_11883_, _05625_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  or _20262_ (_11884_, _11883_, _11881_);
  nor _20263_ (_11886_, _05613_, _10995_);
  and _20264_ (_11887_, _05632_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  or _20265_ (_11889_, _11887_, _11886_);
  or _20266_ (_11890_, _11889_, _11884_);
  and _20267_ (_11891_, _05619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and _20268_ (_11892_, _05627_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  or _20269_ (_11893_, _11892_, _11891_);
  or _20270_ (_11895_, _11893_, _11890_);
  and _20271_ (_11896_, _11895_, _05671_);
  or _20272_ (_11898_, _11896_, _11879_);
  and _20273_ (_11899_, _11898_, _05547_);
  nor _20274_ (_11900_, _11899_, _11878_);
  and _20275_ (_11901_, _11900_, _11783_);
  and _20276_ (_11902_, _11815_, _11469_);
  nor _20277_ (_11903_, _11902_, _11901_);
  nand _20278_ (_11904_, _11903_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nor _20279_ (_11905_, _05547_, _06167_);
  and _20280_ (_11906_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _20281_ (_11907_, _05616_, _11002_);
  and _20282_ (_11908_, _05625_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  or _20283_ (_11909_, _11908_, _11907_);
  and _20284_ (_11910_, _05725_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  nor _20285_ (_11911_, _05631_, _05699_);
  or _20286_ (_11912_, _11911_, _11910_);
  or _20287_ (_11913_, _11912_, _11909_);
  and _20288_ (_11914_, _05619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and _20289_ (_11915_, _05627_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  or _20290_ (_11916_, _11915_, _11914_);
  or _20291_ (_11917_, _11916_, _11913_);
  and _20292_ (_11918_, _11917_, _05671_);
  or _20293_ (_11919_, _11918_, _11906_);
  and _20294_ (_11920_, _11919_, _05547_);
  nor _20295_ (_11921_, _11920_, _11905_);
  and _20296_ (_11922_, _11921_, _11783_);
  and _20297_ (_11923_, _11815_, _11274_);
  nor _20298_ (_11924_, _11923_, _11922_);
  nor _20299_ (_11925_, _11924_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and _20300_ (_11926_, _11924_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nor _20301_ (_11927_, _05547_, _06207_);
  and _20302_ (_11928_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and _20303_ (_11929_, _05619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and _20304_ (_11930_, _05625_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor _20305_ (_11931_, _11930_, _11929_);
  nor _20306_ (_11932_, _05616_, _11739_);
  and _20307_ (_11933_, _05627_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor _20308_ (_11934_, _11933_, _11932_);
  nor _20309_ (_11935_, _05613_, _08689_);
  nor _20310_ (_11936_, _05631_, _05677_);
  nor _20311_ (_11937_, _11936_, _11935_);
  and _20312_ (_11938_, _11937_, _11934_);
  and _20313_ (_11939_, _11938_, _11931_);
  nor _20314_ (_11940_, _11939_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _20315_ (_11941_, _11940_, _11928_);
  nor _20316_ (_11942_, _11941_, _05548_);
  nor _20317_ (_11943_, _11942_, _11927_);
  not _20318_ (_11944_, _11943_);
  or _20319_ (_11945_, _11944_, _11815_);
  or _20320_ (_11946_, _11783_, _11747_);
  nand _20321_ (_11947_, _11946_, _11945_);
  or _20322_ (_11948_, _11947_, _06217_);
  not _20323_ (_11949_, _11948_);
  nor _20324_ (_11950_, _05547_, _06230_);
  and _20325_ (_11951_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _20326_ (_11952_, _05613_, _05553_);
  nor _20327_ (_11953_, _05624_, _05615_);
  nor _20328_ (_11954_, _11953_, _11952_);
  and _20329_ (_11955_, _05619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  nor _20330_ (_11956_, _05631_, _05611_);
  nor _20331_ (_11957_, _11956_, _11955_);
  and _20332_ (_11958_, _05627_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor _20333_ (_11959_, _05616_, _11609_);
  nor _20334_ (_11960_, _11959_, _11958_);
  and _20335_ (_11961_, _11960_, _11957_);
  and _20336_ (_11962_, _11961_, _11954_);
  nor _20337_ (_11964_, _11962_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _20338_ (_11965_, _11964_, _11951_);
  nor _20339_ (_11966_, _11965_, _05548_);
  nor _20340_ (_11967_, _11966_, _11950_);
  not _20341_ (_11968_, _11967_);
  or _20342_ (_11969_, _11968_, _11815_);
  or _20343_ (_11970_, _11783_, _11617_);
  and _20344_ (_11971_, _11970_, _11969_);
  nand _20345_ (_11972_, _11971_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nor _20346_ (_11973_, _05547_, _06188_);
  and _20347_ (_11975_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _20348_ (_11976_, _05616_, _11006_);
  and _20349_ (_11977_, _05625_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  or _20350_ (_11978_, _11977_, _11976_);
  and _20351_ (_11979_, _05725_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  nor _20352_ (_11980_, _05631_, _05656_);
  or _20353_ (_11982_, _11980_, _11979_);
  or _20354_ (_11983_, _11982_, _11978_);
  and _20355_ (_11985_, _05619_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and _20356_ (_11986_, _05627_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  or _20357_ (_11987_, _11986_, _11985_);
  or _20358_ (_11988_, _11987_, _11983_);
  and _20359_ (_11989_, _11988_, _05671_);
  or _20360_ (_11990_, _11989_, _11975_);
  and _20361_ (_11991_, _11990_, _05547_);
  nor _20362_ (_11993_, _11991_, _11973_);
  not _20363_ (_11994_, _11993_);
  or _20364_ (_11995_, _11994_, _11815_);
  or _20365_ (_11996_, _11783_, _11691_);
  and _20366_ (_11997_, _11996_, _11995_);
  and _20367_ (_11998_, _11997_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  or _20368_ (_11999_, _11971_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and _20369_ (_12000_, _11999_, _11972_);
  and _20370_ (_12001_, _12000_, _11998_);
  not _20371_ (_12002_, _12001_);
  nand _20372_ (_12004_, _12002_, _11972_);
  nand _20373_ (_12005_, _11947_, _06217_);
  and _20374_ (_12006_, _12005_, _11948_);
  and _20375_ (_12007_, _12006_, _12004_);
  or _20376_ (_12008_, _12007_, _11949_);
  nor _20377_ (_12009_, _12008_, _11926_);
  nor _20378_ (_12010_, _12009_, _11925_);
  or _20379_ (_12012_, _11903_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _20380_ (_12013_, _12012_, _11904_);
  nand _20381_ (_12014_, _12013_, _12010_);
  nand _20382_ (_12015_, _12014_, _11904_);
  nor _20383_ (_12016_, _12015_, _11877_);
  nor _20384_ (_12017_, _12016_, _11876_);
  and _20385_ (_12018_, _12017_, _11854_);
  or _20386_ (_12019_, _12018_, _11852_);
  nor _20387_ (_12020_, _12019_, _11830_);
  nor _20388_ (_12021_, _12020_, _11829_);
  or _20389_ (_12022_, _12021_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  or _20390_ (_12024_, _12022_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  or _20391_ (_12025_, _12024_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  or _20392_ (_12027_, _12025_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor _20393_ (_12028_, _12027_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _20394_ (_12029_, _12028_, _06085_);
  nand _20395_ (_12030_, _12029_, _06487_);
  nand _20396_ (_12031_, _12030_, _11828_);
  not _20397_ (_12032_, _11828_);
  and _20398_ (_12034_, _12021_, _11797_);
  nand _20399_ (_12035_, _12034_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  or _20400_ (_12036_, _12035_, _06148_);
  nor _20401_ (_12037_, _12036_, _06085_);
  nand _20402_ (_12038_, _12037_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand _20403_ (_12039_, _12038_, _12032_);
  nand _20404_ (_12040_, _12039_, _12031_);
  nand _20405_ (_12041_, _12040_, _06590_);
  or _20406_ (_12043_, _12040_, _06590_);
  and _20407_ (_12044_, _12043_, _12041_);
  and _20408_ (_12045_, _11084_, _05850_);
  and _20409_ (_12046_, _12045_, _10905_);
  and _20410_ (_12047_, _11561_, _11134_);
  and _20411_ (_12048_, _12047_, _11126_);
  and _20412_ (_12050_, _11571_, _11558_);
  and _20413_ (_12051_, _12050_, _12048_);
  nor _20414_ (_12052_, _12051_, _11132_);
  nor _20415_ (_12053_, _12052_, _12046_);
  nor _20416_ (_12054_, _12053_, _11786_);
  and _20417_ (_12056_, _12054_, _12044_);
  or _20418_ (_12057_, _12056_, _11824_);
  and _20419_ (_12059_, _08238_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and _20420_ (_12060_, _12059_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and _20421_ (_12061_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7], \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and _20422_ (_12062_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10], \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and _20423_ (_12063_, _12062_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and _20424_ (_12064_, _12063_, _12061_);
  and _20425_ (_12066_, _12064_, _12060_);
  and _20426_ (_12068_, _12066_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and _20427_ (_12069_, _12068_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and _20428_ (_12071_, _12069_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and _20429_ (_12072_, _12071_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or _20430_ (_12073_, _12072_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nand _20431_ (_12074_, _12072_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and _20432_ (_12075_, _12074_, _12073_);
  or _20433_ (_12076_, _12075_, _11774_);
  and _20434_ (_12077_, _12076_, _05552_);
  and _20435_ (_10889_, _12077_, _12057_);
  and _20436_ (_12080_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _05556_);
  and _20437_ (_12081_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _20438_ (_12082_, _12081_, _12080_);
  and _20439_ (_10900_, _12082_, _05552_);
  or _20440_ (_12083_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  nand _20441_ (_12085_, _05550_, _05743_);
  and _20442_ (_12086_, _12085_, _05552_);
  and _20443_ (_10903_, _12086_, _12083_);
  and _20444_ (_12088_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor _20445_ (_12089_, _05550_, _11441_);
  or _20446_ (_12090_, _12089_, _12088_);
  and _20447_ (_10916_, _12090_, _05552_);
  and _20448_ (_12091_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  nor _20449_ (_12092_, _05550_, _05656_);
  or _20450_ (_12093_, _12092_, _12091_);
  and _20451_ (_10928_, _12093_, _05552_);
  and _20452_ (_10951_, _05552_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  not _20453_ (_12094_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  and _20454_ (_12095_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  not _20455_ (_12096_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and _20456_ (_12097_, _10874_, _12096_);
  not _20457_ (_12098_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  nor _20458_ (_12099_, _12098_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  or _20459_ (_12100_, _12099_, _12097_);
  nor _20460_ (_12101_, _12100_, _12095_);
  nand _20461_ (_12103_, _12101_, _12094_);
  nor _20462_ (_12104_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  nor _20463_ (_12106_, _12104_, _12101_);
  nand _20464_ (_12107_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  nand _20465_ (_12108_, _12107_, _12106_);
  and _20466_ (_12109_, _12108_, _05552_);
  and _20467_ (_10954_, _12109_, _12103_);
  and _20468_ (_12111_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor _20469_ (_12112_, _05550_, _11383_);
  or _20470_ (_12114_, _12112_, _12111_);
  and _20471_ (_10985_, _12114_, _05552_);
  nor _20472_ (_12116_, _09136_, _09133_);
  nor _20473_ (_12117_, _12116_, _09137_);
  or _20474_ (_12118_, _12117_, _09039_);
  or _20475_ (_12119_, _09038_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and _20476_ (_12120_, _12119_, _05605_);
  and _20477_ (_12121_, _12120_, _12118_);
  and _20478_ (_12122_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  or _20479_ (_12123_, _12122_, _12121_);
  and _20480_ (_11013_, _12123_, _05552_);
  and _20481_ (_12124_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], _07768_);
  and _20482_ (_12125_, \oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or _20483_ (_12126_, _12125_, _12124_);
  and _20484_ (_11034_, _12126_, _05552_);
  nor _20485_ (_11044_, _11921_, rst);
  nor _20486_ (_11047_, _11746_, rst);
  nand _20487_ (_12127_, _07483_, _06973_);
  and _20488_ (_12128_, _08935_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and _20489_ (_12129_, _10632_, _08048_);
  nor _20490_ (_12130_, _10632_, _06179_);
  nor _20491_ (_12131_, _12130_, _12129_);
  nor _20492_ (_12132_, _12131_, _08924_);
  nor _20493_ (_12133_, _12132_, _12128_);
  and _20494_ (_12134_, _12133_, _07261_);
  and _20495_ (_12136_, _12134_, _12127_);
  and _20496_ (_12137_, _07515_, _07260_);
  nor _20497_ (_12138_, _12137_, _12136_);
  and _20498_ (_11049_, _12138_, _05552_);
  and _20499_ (_12139_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  not _20500_ (_12140_, _05550_);
  and _20501_ (_12141_, _12140_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  or _20502_ (_12142_, _12141_, _12139_);
  and _20503_ (_11055_, _12142_, _05552_);
  nor _20504_ (_12143_, _09151_, _09091_);
  nor _20505_ (_12144_, _12143_, _09152_);
  or _20506_ (_12145_, _12144_, _09039_);
  or _20507_ (_12146_, _09038_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _20508_ (_12147_, _12146_, _07933_);
  and _20509_ (_12148_, _12147_, _12145_);
  and _20510_ (_12149_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and _20511_ (_12150_, _12149_, _05552_);
  or _20512_ (_11096_, _12150_, _12148_);
  and _20513_ (_12152_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  nor _20514_ (_12153_, _05550_, _05699_);
  or _20515_ (_12154_, _12153_, _12152_);
  and _20516_ (_11104_, _12154_, _05552_);
  nand _20517_ (_12155_, _12027_, _11828_);
  nand _20518_ (_12156_, _12035_, _12032_);
  and _20519_ (_12157_, _12156_, _12155_);
  nand _20520_ (_12159_, _12157_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor _20521_ (_12160_, _11791_, _11779_);
  nor _20522_ (_12161_, _12160_, _11786_);
  or _20523_ (_12162_, _12157_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _20524_ (_12163_, _12162_, _12161_);
  and _20525_ (_12164_, _12163_, _12159_);
  or _20526_ (_12165_, _07178_, _07176_);
  and _20527_ (_12166_, _12165_, _07603_);
  or _20528_ (_12167_, _12166_, _07446_);
  or _20529_ (_12168_, _07200_, _07130_);
  and _20530_ (_12169_, _12168_, _12167_);
  and _20531_ (_12170_, _12169_, _06314_);
  and _20532_ (_12171_, _06908_, _07211_);
  and _20533_ (_12172_, _11525_, _06581_);
  or _20534_ (_12173_, _06698_, _06628_);
  nor _20535_ (_12174_, _06699_, _06678_);
  and _20536_ (_12175_, _12174_, _12173_);
  nor _20537_ (_12176_, _07467_, _06118_);
  nor _20538_ (_12177_, _12176_, _06164_);
  and _20539_ (_12178_, _06718_, _06164_);
  and _20540_ (_12179_, _06128_, _06111_);
  and _20541_ (_12180_, _06184_, _06131_);
  or _20542_ (_12181_, _12180_, _12179_);
  nor _20543_ (_12182_, _12181_, _12178_);
  nand _20544_ (_12183_, _12182_, _07386_);
  nor _20545_ (_12184_, _12183_, _12177_);
  nand _20546_ (_12185_, _12184_, _07375_);
  or _20547_ (_12186_, _12185_, _12175_);
  or _20548_ (_12187_, _12186_, _12172_);
  or _20549_ (_12188_, _12187_, _12171_);
  or _20550_ (_12189_, _12188_, _12170_);
  and _20551_ (_12190_, _12189_, _11811_);
  or _20552_ (_12192_, _07299_, _07296_);
  nor _20553_ (_12193_, _07300_, _06678_);
  and _20554_ (_12194_, _12193_, _12192_);
  and _20555_ (_12195_, _07719_, _07211_);
  nor _20556_ (_12196_, _07322_, _06142_);
  nor _20557_ (_12197_, _07330_, _06253_);
  or _20558_ (_12198_, _12197_, _12196_);
  nand _20559_ (_12199_, _12198_, _06379_);
  or _20560_ (_12200_, _12198_, _06379_);
  and _20561_ (_12201_, _12200_, _06266_);
  and _20562_ (_12202_, _12201_, _12199_);
  or _20563_ (_12203_, _06162_, _06253_);
  or _20564_ (_12204_, _06625_, _06142_);
  and _20565_ (_12205_, _12204_, _06295_);
  and _20566_ (_12206_, _12205_, _12203_);
  and _20567_ (_12207_, _06368_, _06746_);
  and _20568_ (_12208_, _06625_, _06118_);
  and _20569_ (_12209_, _06314_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  or _20570_ (_12210_, _12209_, _12208_);
  or _20571_ (_12211_, _12210_, _12207_);
  or _20572_ (_12212_, _12211_, _12206_);
  or _20573_ (_12213_, _12212_, _12202_);
  or _20574_ (_12214_, _12213_, _12195_);
  or _20575_ (_12215_, _12214_, _12194_);
  and _20576_ (_12216_, _12215_, _11784_);
  nor _20577_ (_12217_, _11803_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor _20578_ (_12218_, _12217_, _11804_);
  and _20579_ (_12219_, _12218_, _11792_);
  and _20580_ (_12220_, _11780_, _11470_);
  or _20581_ (_12221_, _12220_, _12219_);
  and _20582_ (_12222_, _11817_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  or _20583_ (_12223_, _12222_, _12221_);
  nor _20584_ (_12224_, _12223_, _12216_);
  nand _20585_ (_12225_, _12224_, _11774_);
  or _20586_ (_12226_, _12225_, _12190_);
  or _20587_ (_12227_, _12226_, _12164_);
  nor _20588_ (_12228_, _12068_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor _20589_ (_12229_, _12228_, _12069_);
  or _20590_ (_12230_, _12229_, _11774_);
  and _20591_ (_12231_, _12230_, _05552_);
  and _20592_ (_11110_, _12231_, _12227_);
  nor _20593_ (_11143_, _11690_, rst);
  or _20594_ (_12232_, _09130_, _09127_);
  and _20595_ (_12233_, _12232_, _09131_);
  or _20596_ (_12234_, _12233_, _09039_);
  or _20597_ (_12235_, _09038_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and _20598_ (_12236_, _12235_, _05605_);
  and _20599_ (_12237_, _12236_, _12234_);
  and _20600_ (_12238_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _20601_ (_12239_, _12238_, _12237_);
  and _20602_ (_11146_, _12239_, _05552_);
  nor _20603_ (_11156_, _11728_, rst);
  or _20604_ (_12240_, _05550_, \oc8051_top_1.oc8051_rom1.data_o [24]);
  nand _20605_ (_12241_, _05550_, _10991_);
  and _20606_ (_12242_, _12241_, _05552_);
  and _20607_ (_11162_, _12242_, _12240_);
  or _20608_ (_12243_, _05550_, \oc8051_top_1.oc8051_rom1.data_o [7]);
  nand _20609_ (_12244_, _05550_, _05762_);
  and _20610_ (_12245_, _12244_, _05552_);
  and _20611_ (_11165_, _12245_, _12243_);
  or _20612_ (_12246_, _09126_, _09123_);
  nor _20613_ (_12247_, _09039_, _09127_);
  and _20614_ (_12248_, _12247_, _12246_);
  and _20615_ (_12249_, _09039_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  or _20616_ (_12250_, _12249_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _20617_ (_12251_, _12250_, _12248_);
  or _20618_ (_12252_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], _05605_);
  and _20619_ (_12253_, _12252_, _05552_);
  and _20620_ (_11168_, _12253_, _12251_);
  and _20621_ (_11184_, _05693_, _05552_);
  nor _20622_ (_12254_, _06306_, _06953_);
  and _20623_ (_12255_, _06953_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  or _20624_ (_12256_, _12255_, _06955_);
  or _20625_ (_12257_, _12256_, _12254_);
  or _20626_ (_12258_, _06068_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  and _20627_ (_12259_, _12258_, _05552_);
  and _20628_ (_11191_, _12259_, _12257_);
  and _20629_ (_12260_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  nor _20630_ (_12261_, _05550_, _05762_);
  or _20631_ (_12262_, _12261_, _12260_);
  and _20632_ (_11215_, _12262_, _05552_);
  not _20633_ (_12263_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  and _20634_ (_12264_, _09504_, _06068_);
  nor _20635_ (_12265_, _12264_, _12263_);
  and _20636_ (_12266_, _09504_, _07976_);
  or _20637_ (_12267_, _12266_, _12265_);
  and _20638_ (_11229_, _12267_, _05552_);
  nor _20639_ (_11259_, _11335_, rst);
  nand _20640_ (_12268_, _11161_, _11089_);
  or _20641_ (_12269_, _11028_, _05861_);
  or _20642_ (_12270_, _12269_, _11153_);
  and _20643_ (_12271_, _06567_, _05809_);
  and _20644_ (_12272_, _12271_, _05737_);
  or _20645_ (_12273_, _12272_, _12270_);
  or _20646_ (_12274_, _12273_, _12268_);
  or _20647_ (_12276_, _05860_, _05814_);
  and _20648_ (_12277_, _12276_, _10843_);
  or _20649_ (_12278_, _11150_, _11016_);
  or _20650_ (_12279_, _12278_, _12277_);
  and _20651_ (_12280_, _10898_, _05830_);
  and _20652_ (_12282_, _05894_, _05846_);
  nor _20653_ (_12283_, _05737_, _05714_);
  and _20654_ (_12284_, _12283_, _05813_);
  or _20655_ (_12285_, _12284_, _12282_);
  or _20656_ (_12287_, _12285_, _12280_);
  or _20657_ (_12288_, _11103_, _10908_);
  or _20658_ (_12289_, _12288_, _12287_);
  or _20659_ (_12290_, _12289_, _12279_);
  and _20660_ (_12291_, _11123_, _06567_);
  or _20661_ (_12292_, _11025_, _12291_);
  or _20662_ (_12293_, _12292_, _12290_);
  or _20663_ (_12295_, _12293_, _12274_);
  and _20664_ (_12296_, _12295_, _06576_);
  nor _20665_ (_12297_, _11084_, rst);
  and _20666_ (_12298_, _12297_, _05896_);
  and _20667_ (_12299_, _05552_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and _20668_ (_12300_, _12299_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  or _20669_ (_12301_, _12300_, _12298_);
  or _20670_ (_11293_, _12301_, _12296_);
  and _20671_ (_12302_, \oc8051_top_1.oc8051_decoder1.alu_op [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _20672_ (_12303_, _12302_, _10957_);
  and _20673_ (_12304_, _12303_, _05552_);
  not _20674_ (_12305_, _11112_);
  or _20675_ (_12306_, _12305_, _10899_);
  not _20676_ (_12307_, _11561_);
  and _20677_ (_12308_, _12283_, _05814_);
  or _20678_ (_12309_, _12308_, _10939_);
  or _20679_ (_12310_, _12309_, _12307_);
  or _20680_ (_12311_, _12310_, _12306_);
  nand _20681_ (_12312_, _10905_, _06567_);
  and _20682_ (_12313_, _10938_, _05859_);
  nor _20683_ (_12314_, _12313_, _10937_);
  and _20684_ (_12315_, _12314_, _11108_);
  nand _20685_ (_12316_, _12315_, _12312_);
  or _20686_ (_12317_, _12316_, _12311_);
  not _20687_ (_12318_, _11022_);
  and _20688_ (_12319_, _11161_, _12318_);
  not _20689_ (_12320_, _12319_);
  or _20690_ (_12321_, _12320_, _10930_);
  or _20691_ (_12322_, _12321_, _12317_);
  and _20692_ (_12324_, _10898_, _05824_);
  or _20693_ (_12325_, _10931_, _05817_);
  or _20694_ (_12327_, _12325_, _12324_);
  and _20695_ (_12328_, _06567_, _05828_);
  or _20696_ (_12329_, _12328_, _05829_);
  and _20697_ (_12330_, _05810_, _05820_);
  and _20698_ (_12331_, _10932_, _05820_);
  or _20699_ (_12332_, _12331_, _12330_);
  or _20700_ (_12333_, _12280_, _11154_);
  or _20701_ (_12334_, _12333_, _12332_);
  or _20702_ (_12335_, _12334_, _12329_);
  or _20703_ (_12336_, _12335_, _12327_);
  or _20704_ (_12337_, _12336_, _12322_);
  and _20705_ (_12338_, _12337_, _06576_);
  or _20706_ (_11295_, _12338_, _12304_);
  nor _20707_ (_12339_, _07939_, _06560_);
  and _20708_ (_12340_, _07939_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  or _20709_ (_12341_, _12340_, _12339_);
  and _20710_ (_11298_, _12341_, _05552_);
  nor _20711_ (_12342_, _07939_, _06306_);
  and _20712_ (_12344_, _07939_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  or _20713_ (_12345_, _12344_, _12342_);
  and _20714_ (_11302_, _12345_, _05552_);
  and _20715_ (_12347_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], _07768_);
  and _20716_ (_12348_, \oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or _20717_ (_12349_, _12348_, _12347_);
  and _20718_ (_11314_, _12349_, _05552_);
  nor _20719_ (_11319_, _11274_, rst);
  nor _20720_ (_11350_, _11616_, rst);
  or _20721_ (_12350_, _05550_, \oc8051_top_1.oc8051_rom1.data_o [8]);
  nand _20722_ (_12351_, _05550_, _11006_);
  and _20723_ (_12352_, _12351_, _05552_);
  and _20724_ (_11355_, _12352_, _12350_);
  or _20725_ (_12353_, _07731_, _05565_);
  or _20726_ (_12354_, _07736_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and _20727_ (_12355_, _12354_, _05552_);
  and _20728_ (_11357_, _12355_, _12353_);
  nor _20729_ (_12357_, _09143_, _09112_);
  nor _20730_ (_12359_, _12357_, _09144_);
  or _20731_ (_12360_, _12359_, _09039_);
  or _20732_ (_12362_, _09038_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and _20733_ (_12363_, _12362_, _07933_);
  and _20734_ (_12364_, _12363_, _12360_);
  and _20735_ (_12365_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and _20736_ (_12366_, _12365_, _05552_);
  or _20737_ (_11369_, _12366_, _12364_);
  nor _20738_ (_11375_, _07390_, rst);
  or _20739_ (_12367_, _09149_, _09098_);
  nor _20740_ (_12368_, _09039_, _09150_);
  and _20741_ (_12369_, _12368_, _12367_);
  nor _20742_ (_12371_, _09038_, _06235_);
  or _20743_ (_12372_, _12371_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _20744_ (_12373_, _12372_, _12369_);
  or _20745_ (_12374_, _05605_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and _20746_ (_12375_, _12374_, _05552_);
  and _20747_ (_11417_, _12375_, _12373_);
  and _20748_ (_12376_, _08362_, word_in[0]);
  or _20749_ (_12377_, _08389_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  or _20750_ (_12378_, _08234_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  and _20751_ (_12379_, _12378_, _12377_);
  and _20752_ (_12380_, _12379_, _08279_);
  or _20753_ (_12381_, _08389_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  or _20754_ (_12382_, _08234_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and _20755_ (_12384_, _12382_, _12381_);
  and _20756_ (_12385_, _12384_, _08260_);
  or _20757_ (_12387_, _08389_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  or _20758_ (_12388_, _08234_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  and _20759_ (_12389_, _12388_, _12387_);
  and _20760_ (_12390_, _12389_, _08257_);
  or _20761_ (_12391_, _12390_, _12385_);
  or _20762_ (_12392_, _12391_, _12380_);
  or _20763_ (_12393_, _08389_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  or _20764_ (_12394_, _08234_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and _20765_ (_12395_, _12394_, _12393_);
  and _20766_ (_12396_, _12395_, _08267_);
  or _20767_ (_12397_, _12396_, _08286_);
  or _20768_ (_12398_, _12397_, _12392_);
  or _20769_ (_12399_, _08389_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  or _20770_ (_12400_, _08234_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  and _20771_ (_12401_, _12400_, _12399_);
  and _20772_ (_12402_, _12401_, _08279_);
  or _20773_ (_12403_, _08389_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  or _20774_ (_12404_, _08234_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  and _20775_ (_12405_, _12404_, _12403_);
  and _20776_ (_12406_, _12405_, _08260_);
  or _20777_ (_12407_, _08389_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  or _20778_ (_12408_, _08234_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  and _20779_ (_12409_, _12408_, _12407_);
  and _20780_ (_12410_, _12409_, _08257_);
  or _20781_ (_12411_, _12410_, _12406_);
  or _20782_ (_12412_, _12411_, _12402_);
  or _20783_ (_12413_, _08389_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  or _20784_ (_12414_, _08234_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  and _20785_ (_12415_, _12414_, _12413_);
  and _20786_ (_12416_, _12415_, _08267_);
  or _20787_ (_12417_, _12416_, _08243_);
  or _20788_ (_12418_, _12417_, _12412_);
  and _20789_ (_12419_, _12418_, _12398_);
  and _20790_ (_12420_, _12419_, _08311_);
  or _20791_ (\oc8051_symbolic_cxrom1.cxrom_data_out [0], _12420_, _12376_);
  and _20792_ (_12421_, _08362_, word_in[1]);
  or _20793_ (_12422_, _08389_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  or _20794_ (_12423_, _08234_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  and _20795_ (_12424_, _12423_, _12422_);
  and _20796_ (_12425_, _12424_, _08279_);
  or _20797_ (_12426_, _08389_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  or _20798_ (_12427_, _08234_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  and _20799_ (_12428_, _12427_, _12426_);
  and _20800_ (_12429_, _12428_, _08260_);
  or _20801_ (_12430_, _08389_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  or _20802_ (_12431_, _08234_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  and _20803_ (_12432_, _12431_, _12430_);
  and _20804_ (_12433_, _12432_, _08257_);
  or _20805_ (_12434_, _12433_, _12429_);
  or _20806_ (_12435_, _12434_, _12425_);
  or _20807_ (_12436_, _08389_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  or _20808_ (_12437_, _08234_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  and _20809_ (_12438_, _12437_, _12436_);
  and _20810_ (_12439_, _12438_, _08267_);
  or _20811_ (_12441_, _12439_, _08286_);
  or _20812_ (_12442_, _12441_, _12435_);
  or _20813_ (_12443_, _08389_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  or _20814_ (_12444_, _08234_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  and _20815_ (_12445_, _12444_, _12443_);
  and _20816_ (_12446_, _12445_, _08279_);
  or _20817_ (_12447_, _08389_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  or _20818_ (_12448_, _08234_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  and _20819_ (_12449_, _12448_, _12447_);
  and _20820_ (_12450_, _12449_, _08260_);
  or _20821_ (_12451_, _08389_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  or _20822_ (_12452_, _08234_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  and _20823_ (_12453_, _12452_, _12451_);
  and _20824_ (_12454_, _12453_, _08257_);
  or _20825_ (_12456_, _12454_, _12450_);
  or _20826_ (_12457_, _12456_, _12446_);
  or _20827_ (_12458_, _08389_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  or _20828_ (_12459_, _08234_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  and _20829_ (_12460_, _12459_, _12458_);
  and _20830_ (_12461_, _12460_, _08267_);
  or _20831_ (_12462_, _12461_, _08243_);
  or _20832_ (_12463_, _12462_, _12457_);
  and _20833_ (_12464_, _12463_, _12442_);
  and _20834_ (_12465_, _12464_, _08311_);
  or _20835_ (\oc8051_symbolic_cxrom1.cxrom_data_out [1], _12465_, _12421_);
  and _20836_ (_12466_, _08362_, word_in[2]);
  or _20837_ (_12468_, _08389_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  or _20838_ (_12469_, _08234_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  and _20839_ (_12470_, _12469_, _12468_);
  and _20840_ (_12471_, _12470_, _08279_);
  or _20841_ (_12472_, _08389_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  or _20842_ (_12473_, _08234_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  and _20843_ (_12474_, _12473_, _12472_);
  and _20844_ (_12475_, _12474_, _08260_);
  or _20845_ (_12476_, _08389_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  or _20846_ (_12477_, _08234_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  and _20847_ (_12478_, _12477_, _12476_);
  and _20848_ (_12479_, _12478_, _08257_);
  or _20849_ (_12480_, _12479_, _12475_);
  or _20850_ (_12481_, _12480_, _12471_);
  or _20851_ (_12482_, _08389_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  or _20852_ (_12483_, _08234_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  and _20853_ (_12484_, _12483_, _12482_);
  and _20854_ (_12485_, _12484_, _08267_);
  or _20855_ (_12486_, _12485_, _08286_);
  or _20856_ (_12487_, _12486_, _12481_);
  or _20857_ (_12488_, _08389_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  or _20858_ (_12489_, _08234_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  and _20859_ (_12490_, _12489_, _12488_);
  and _20860_ (_12491_, _12490_, _08279_);
  or _20861_ (_12492_, _08389_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  or _20862_ (_12493_, _08234_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  and _20863_ (_12494_, _12493_, _12492_);
  and _20864_ (_12495_, _12494_, _08260_);
  or _20865_ (_12496_, _08389_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  or _20866_ (_12497_, _08234_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  and _20867_ (_12498_, _12497_, _12496_);
  and _20868_ (_12499_, _12498_, _08257_);
  or _20869_ (_12500_, _12499_, _12495_);
  or _20870_ (_12501_, _12500_, _12491_);
  or _20871_ (_12502_, _08389_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  or _20872_ (_12503_, _08234_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  and _20873_ (_12504_, _12503_, _12502_);
  and _20874_ (_12505_, _12504_, _08267_);
  or _20875_ (_12506_, _12505_, _08243_);
  or _20876_ (_12507_, _12506_, _12501_);
  and _20877_ (_12508_, _12507_, _12487_);
  and _20878_ (_12509_, _12508_, _08311_);
  or _20879_ (\oc8051_symbolic_cxrom1.cxrom_data_out [2], _12509_, _12466_);
  and _20880_ (_12510_, _08362_, word_in[3]);
  or _20881_ (_12511_, _08389_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  or _20882_ (_12512_, _08234_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  and _20883_ (_12513_, _12512_, _12511_);
  and _20884_ (_12514_, _12513_, _08279_);
  or _20885_ (_12515_, _08389_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  or _20886_ (_12516_, _08234_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  and _20887_ (_12517_, _12516_, _12515_);
  and _20888_ (_12518_, _12517_, _08260_);
  or _20889_ (_12519_, _12518_, _12514_);
  or _20890_ (_12521_, _08389_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  or _20891_ (_12522_, _08234_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  and _20892_ (_12524_, _12522_, _12521_);
  and _20893_ (_12525_, _12524_, _08267_);
  or _20894_ (_12526_, _08389_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  or _20895_ (_12527_, _08234_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  and _20896_ (_12528_, _12527_, _12526_);
  and _20897_ (_12529_, _12528_, _08257_);
  or _20898_ (_12530_, _12529_, _12525_);
  or _20899_ (_12531_, _12530_, _12519_);
  and _20900_ (_12532_, _12531_, _08243_);
  or _20901_ (_12533_, _08389_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  or _20902_ (_12534_, _08234_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  and _20903_ (_12535_, _12534_, _12533_);
  and _20904_ (_12536_, _12535_, _08260_);
  or _20905_ (_12537_, _08389_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  or _20906_ (_12538_, _08234_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  and _20907_ (_12539_, _12538_, _12537_);
  and _20908_ (_12540_, _12539_, _08279_);
  or _20909_ (_12541_, _12540_, _12536_);
  or _20910_ (_12542_, _08389_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  or _20911_ (_12543_, _08234_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  and _20912_ (_12544_, _12543_, _12542_);
  and _20913_ (_12545_, _12544_, _08267_);
  or _20914_ (_12546_, _08389_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  or _20915_ (_12547_, _08234_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  and _20916_ (_12548_, _12547_, _12546_);
  and _20917_ (_12549_, _12548_, _08257_);
  or _20918_ (_12550_, _12549_, _12545_);
  or _20919_ (_12551_, _12550_, _12541_);
  and _20920_ (_12552_, _12551_, _08286_);
  or _20921_ (_12553_, _12552_, _12532_);
  and _20922_ (_12554_, _12553_, _08311_);
  or _20923_ (\oc8051_symbolic_cxrom1.cxrom_data_out [3], _12554_, _12510_);
  and _20924_ (_12555_, _08362_, word_in[4]);
  or _20925_ (_12556_, _08389_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  or _20926_ (_12557_, _08234_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  and _20927_ (_12558_, _12557_, _12556_);
  and _20928_ (_12559_, _12558_, _08279_);
  or _20929_ (_12560_, _08389_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  or _20930_ (_12561_, _08234_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  and _20931_ (_12562_, _12561_, _12560_);
  and _20932_ (_12563_, _12562_, _08257_);
  or _20933_ (_12564_, _08389_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  or _20934_ (_12565_, _08234_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  and _20935_ (_12566_, _12565_, _12564_);
  and _20936_ (_12567_, _12566_, _08260_);
  or _20937_ (_12568_, _12567_, _12563_);
  or _20938_ (_12569_, _12568_, _12559_);
  or _20939_ (_12570_, _08389_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  or _20940_ (_12571_, _08234_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  and _20941_ (_12572_, _12571_, _12570_);
  and _20942_ (_12573_, _12572_, _08267_);
  or _20943_ (_12574_, _12573_, _08286_);
  or _20944_ (_12575_, _12574_, _12569_);
  or _20945_ (_12576_, _08389_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  or _20946_ (_12577_, _08234_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  and _20947_ (_12578_, _12577_, _12576_);
  and _20948_ (_12579_, _12578_, _08279_);
  or _20949_ (_12580_, _08389_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  or _20950_ (_12581_, _08234_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  and _20951_ (_12582_, _12581_, _12580_);
  and _20952_ (_12583_, _12582_, _08260_);
  or _20953_ (_12584_, _08389_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  or _20954_ (_12585_, _08234_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  and _20955_ (_12586_, _12585_, _12584_);
  and _20956_ (_12587_, _12586_, _08257_);
  or _20957_ (_12588_, _12587_, _12583_);
  or _20958_ (_12589_, _12588_, _12579_);
  or _20959_ (_12590_, _08389_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  or _20960_ (_12591_, _08234_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  and _20961_ (_12592_, _12591_, _12590_);
  and _20962_ (_12593_, _12592_, _08267_);
  or _20963_ (_12594_, _12593_, _08243_);
  or _20964_ (_12595_, _12594_, _12589_);
  and _20965_ (_12596_, _12595_, _12575_);
  and _20966_ (_12597_, _12596_, _08311_);
  or _20967_ (\oc8051_symbolic_cxrom1.cxrom_data_out [4], _12597_, _12555_);
  and _20968_ (_12599_, _08362_, word_in[5]);
  or _20969_ (_12600_, _08389_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  or _20970_ (_12601_, _08234_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  and _20971_ (_12602_, _12601_, _12600_);
  and _20972_ (_12603_, _12602_, _08279_);
  or _20973_ (_12604_, _08389_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  or _20974_ (_12605_, _08234_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  and _20975_ (_12606_, _12605_, _12604_);
  and _20976_ (_12607_, _12606_, _08260_);
  or _20977_ (_12608_, _08389_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  or _20978_ (_12609_, _08234_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  and _20979_ (_12610_, _12609_, _12608_);
  and _20980_ (_12611_, _12610_, _08257_);
  or _20981_ (_12612_, _12611_, _12607_);
  or _20982_ (_12613_, _12612_, _12603_);
  or _20983_ (_12614_, _08389_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  or _20984_ (_12615_, _08234_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  and _20985_ (_12616_, _12615_, _12614_);
  and _20986_ (_12617_, _12616_, _08267_);
  or _20987_ (_12618_, _12617_, _08286_);
  or _20988_ (_12619_, _12618_, _12613_);
  or _20989_ (_12620_, _08389_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  or _20990_ (_12621_, _08234_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  and _20991_ (_12622_, _12621_, _12620_);
  and _20992_ (_12623_, _12622_, _08279_);
  or _20993_ (_12624_, _08389_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  or _20994_ (_12625_, _08234_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  and _20995_ (_12626_, _12625_, _12624_);
  and _20996_ (_12627_, _12626_, _08260_);
  or _20997_ (_12628_, _08389_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  or _20998_ (_12629_, _08234_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  and _20999_ (_12630_, _12629_, _12628_);
  and _21000_ (_12631_, _12630_, _08257_);
  or _21001_ (_12632_, _12631_, _12627_);
  or _21002_ (_12633_, _12632_, _12623_);
  or _21003_ (_12634_, _08389_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  or _21004_ (_12635_, _08234_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  and _21005_ (_12636_, _12635_, _12634_);
  and _21006_ (_12637_, _12636_, _08267_);
  or _21007_ (_12638_, _12637_, _08243_);
  or _21008_ (_12639_, _12638_, _12633_);
  and _21009_ (_12640_, _12639_, _12619_);
  and _21010_ (_12641_, _12640_, _08311_);
  or _21011_ (\oc8051_symbolic_cxrom1.cxrom_data_out [5], _12641_, _12599_);
  and _21012_ (_12642_, _08362_, word_in[6]);
  or _21013_ (_12643_, _08389_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  or _21014_ (_12644_, _08234_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  and _21015_ (_12645_, _12644_, _12643_);
  and _21016_ (_12646_, _12645_, _08260_);
  or _21017_ (_12647_, _08389_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  or _21018_ (_12648_, _08234_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  and _21019_ (_12649_, _12648_, _12647_);
  and _21020_ (_12650_, _12649_, _08257_);
  or _21021_ (_12651_, _08389_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  or _21022_ (_12652_, _08234_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  and _21023_ (_12653_, _12652_, _12651_);
  and _21024_ (_12654_, _12653_, _08279_);
  or _21025_ (_12655_, _12654_, _12650_);
  or _21026_ (_12656_, _12655_, _12646_);
  or _21027_ (_12657_, _08389_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  or _21028_ (_12658_, _08234_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  and _21029_ (_12659_, _12658_, _12657_);
  and _21030_ (_12660_, _12659_, _08267_);
  or _21031_ (_12661_, _12660_, _08286_);
  or _21032_ (_12662_, _12661_, _12656_);
  or _21033_ (_12663_, _08389_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  or _21034_ (_12664_, _08234_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  and _21035_ (_12665_, _12664_, _12663_);
  and _21036_ (_12666_, _12665_, _08260_);
  or _21037_ (_12667_, _08389_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  or _21038_ (_12668_, _08234_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  and _21039_ (_12669_, _12668_, _12667_);
  and _21040_ (_12670_, _12669_, _08279_);
  or _21041_ (_12671_, _08389_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  or _21042_ (_12672_, _08234_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  and _21043_ (_12673_, _12672_, _12671_);
  and _21044_ (_12674_, _12673_, _08257_);
  or _21045_ (_12675_, _12674_, _12670_);
  or _21046_ (_12676_, _12675_, _12666_);
  or _21047_ (_12677_, _08389_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  or _21048_ (_12678_, _08234_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  and _21049_ (_12679_, _12678_, _12677_);
  and _21050_ (_12680_, _12679_, _08267_);
  or _21051_ (_12681_, _12680_, _08243_);
  or _21052_ (_12682_, _12681_, _12676_);
  and _21053_ (_12683_, _12682_, _12662_);
  and _21054_ (_12684_, _12683_, _08311_);
  or _21055_ (\oc8051_symbolic_cxrom1.cxrom_data_out [6], _12684_, _12642_);
  nor _21056_ (_12685_, _09148_, _09146_);
  nor _21057_ (_12686_, _12685_, _09149_);
  or _21058_ (_12687_, _12686_, _09039_);
  or _21059_ (_12688_, _09038_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and _21060_ (_12689_, _12688_, _05605_);
  and _21061_ (_12690_, _12689_, _12687_);
  and _21062_ (_12691_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  or _21063_ (_12692_, _12691_, _12690_);
  and _21064_ (_11435_, _12692_, _05552_);
  or _21065_ (_12693_, _09145_, _09102_);
  nor _21066_ (_12694_, _09039_, _09146_);
  and _21067_ (_12695_, _12694_, _12693_);
  nor _21068_ (_12696_, _09038_, _06588_);
  or _21069_ (_12697_, _12696_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _21070_ (_12698_, _12697_, _12695_);
  or _21071_ (_12699_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7], _05605_);
  and _21072_ (_12700_, _12699_, _05552_);
  and _21073_ (_11438_, _12700_, _12698_);
  and _21074_ (_12701_, _08439_, word_in[8]);
  or _21075_ (_12702_, _08389_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  or _21076_ (_12703_, _08234_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and _21077_ (_12704_, _12703_, _12702_);
  and _21078_ (_12705_, _12704_, _08441_);
  or _21079_ (_12706_, _08389_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  or _21080_ (_12707_, _08234_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  and _21081_ (_12708_, _12707_, _12706_);
  and _21082_ (_12709_, _12708_, _08440_);
  or _21083_ (_12710_, _12709_, _12705_);
  and _21084_ (_12711_, _12710_, _08402_);
  or _21085_ (_12712_, _08389_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  or _21086_ (_12713_, _08234_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  and _21087_ (_12714_, _12713_, _12712_);
  and _21088_ (_12715_, _12714_, _08441_);
  or _21089_ (_12716_, _08389_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  or _21090_ (_12717_, _08234_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  and _21091_ (_12718_, _12717_, _12716_);
  and _21092_ (_12719_, _12718_, _08440_);
  nor _21093_ (_12720_, _12719_, _12715_);
  nor _21094_ (_12721_, _12720_, _08406_);
  or _21095_ (_12722_, _08389_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  or _21096_ (_12723_, _08234_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  and _21097_ (_12724_, _12723_, _12722_);
  and _21098_ (_12725_, _12724_, _08441_);
  or _21099_ (_12726_, _08389_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  or _21100_ (_12727_, _08234_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  and _21101_ (_12728_, _12727_, _12726_);
  and _21102_ (_12729_, _12728_, _08440_);
  or _21103_ (_12730_, _12729_, _12725_);
  and _21104_ (_12731_, _12730_, _08467_);
  or _21105_ (_12732_, _08389_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  or _21106_ (_12733_, _08234_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  and _21107_ (_12734_, _12733_, _12732_);
  and _21108_ (_12735_, _12734_, _08441_);
  or _21109_ (_12736_, _08389_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  or _21110_ (_12737_, _08234_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  and _21111_ (_12738_, _12737_, _12736_);
  and _21112_ (_12739_, _12738_, _08440_);
  or _21113_ (_12740_, _12739_, _12735_);
  and _21114_ (_12741_, _12740_, _08480_);
  or _21115_ (_12742_, _12741_, _12731_);
  or _21116_ (_12743_, _12742_, _12721_);
  nor _21117_ (_12744_, _12743_, _12711_);
  nor _21118_ (_12745_, _12744_, _08439_);
  or _21119_ (\oc8051_symbolic_cxrom1.cxrom_data_out [8], _12745_, _12701_);
  and _21120_ (_12746_, _08439_, word_in[9]);
  or _21121_ (_12747_, _08389_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  or _21122_ (_12748_, _08234_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  and _21123_ (_12749_, _12748_, _12747_);
  and _21124_ (_12750_, _12749_, _08441_);
  or _21125_ (_12751_, _08389_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  or _21126_ (_12752_, _08234_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  and _21127_ (_12753_, _12752_, _12751_);
  and _21128_ (_12754_, _12753_, _08440_);
  or _21129_ (_12755_, _12754_, _12750_);
  and _21130_ (_12756_, _12755_, _08402_);
  or _21131_ (_12757_, _08389_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  or _21132_ (_12758_, _08234_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  and _21133_ (_12759_, _12758_, _12757_);
  and _21134_ (_12760_, _12759_, _08441_);
  or _21135_ (_12761_, _08389_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  or _21136_ (_12762_, _08234_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  and _21137_ (_12763_, _12762_, _12761_);
  and _21138_ (_12764_, _12763_, _08440_);
  nor _21139_ (_12765_, _12764_, _12760_);
  nor _21140_ (_12766_, _12765_, _08406_);
  or _21141_ (_12767_, _08389_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  or _21142_ (_12768_, _08234_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  and _21143_ (_12769_, _12768_, _12767_);
  and _21144_ (_12770_, _12769_, _08441_);
  or _21145_ (_12771_, _08389_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  or _21146_ (_12773_, _08234_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  and _21147_ (_12774_, _12773_, _12771_);
  and _21148_ (_12775_, _12774_, _08440_);
  or _21149_ (_12776_, _12775_, _12770_);
  and _21150_ (_12777_, _12776_, _08467_);
  or _21151_ (_12778_, _08389_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  or _21152_ (_12779_, _08234_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  and _21153_ (_12780_, _12779_, _12778_);
  and _21154_ (_12781_, _12780_, _08441_);
  or _21155_ (_12782_, _08389_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  or _21156_ (_12783_, _08234_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  and _21157_ (_12784_, _12783_, _12782_);
  and _21158_ (_12785_, _12784_, _08440_);
  or _21159_ (_12786_, _12785_, _12781_);
  and _21160_ (_12787_, _12786_, _08480_);
  or _21161_ (_12788_, _12787_, _12777_);
  or _21162_ (_12789_, _12788_, _12766_);
  nor _21163_ (_12790_, _12789_, _12756_);
  nor _21164_ (_12791_, _12790_, _08439_);
  or _21165_ (\oc8051_symbolic_cxrom1.cxrom_data_out [9], _12791_, _12746_);
  and _21166_ (_12792_, _08439_, word_in[10]);
  or _21167_ (_12793_, _08389_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  or _21168_ (_12794_, _08234_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  and _21169_ (_12795_, _12794_, _12793_);
  and _21170_ (_12796_, _12795_, _08441_);
  or _21171_ (_12797_, _08389_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  or _21172_ (_12798_, _08234_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  and _21173_ (_12799_, _12798_, _12797_);
  and _21174_ (_12800_, _12799_, _08440_);
  or _21175_ (_12801_, _12800_, _12796_);
  and _21176_ (_12802_, _12801_, _08402_);
  or _21177_ (_12803_, _08389_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  or _21178_ (_12804_, _08234_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  and _21179_ (_12805_, _12804_, _12803_);
  and _21180_ (_12806_, _12805_, _08441_);
  or _21181_ (_12808_, _08389_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  or _21182_ (_12809_, _08234_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  and _21183_ (_12810_, _12809_, _12808_);
  and _21184_ (_12811_, _12810_, _08440_);
  nor _21185_ (_12812_, _12811_, _12806_);
  nor _21186_ (_12813_, _12812_, _08406_);
  or _21187_ (_12814_, _08389_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  or _21188_ (_12815_, _08234_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  and _21189_ (_12816_, _12815_, _12814_);
  and _21190_ (_12817_, _12816_, _08441_);
  or _21191_ (_12818_, _08389_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  or _21192_ (_12819_, _08234_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  and _21193_ (_12820_, _12819_, _12818_);
  and _21194_ (_12821_, _12820_, _08440_);
  or _21195_ (_12822_, _12821_, _12817_);
  and _21196_ (_12823_, _12822_, _08467_);
  or _21197_ (_12824_, _08389_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  or _21198_ (_12825_, _08234_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  and _21199_ (_12826_, _12825_, _12824_);
  and _21200_ (_12827_, _12826_, _08441_);
  or _21201_ (_12828_, _08389_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  or _21202_ (_12829_, _08234_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  and _21203_ (_12830_, _12829_, _12828_);
  and _21204_ (_12831_, _12830_, _08440_);
  or _21205_ (_12832_, _12831_, _12827_);
  and _21206_ (_12833_, _12832_, _08480_);
  or _21207_ (_12834_, _12833_, _12823_);
  or _21208_ (_12835_, _12834_, _12813_);
  nor _21209_ (_12836_, _12835_, _12802_);
  nor _21210_ (_12837_, _12836_, _08439_);
  or _21211_ (\oc8051_symbolic_cxrom1.cxrom_data_out [10], _12837_, _12792_);
  and _21212_ (_12838_, _08439_, word_in[11]);
  or _21213_ (_12839_, _08389_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  or _21214_ (_12840_, _08234_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  and _21215_ (_12841_, _12840_, _12839_);
  and _21216_ (_12842_, _12841_, _08441_);
  or _21217_ (_12843_, _08389_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  or _21218_ (_12844_, _08234_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  and _21219_ (_12845_, _12844_, _12843_);
  and _21220_ (_12846_, _12845_, _08440_);
  or _21221_ (_12847_, _12846_, _12842_);
  and _21222_ (_12848_, _12847_, _08402_);
  or _21223_ (_12849_, _08389_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  or _21224_ (_12850_, _08234_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  and _21225_ (_12851_, _12850_, _12849_);
  and _21226_ (_12852_, _12851_, _08441_);
  or _21227_ (_12853_, _08389_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  or _21228_ (_12854_, _08234_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  and _21229_ (_12855_, _12854_, _12853_);
  and _21230_ (_12856_, _12855_, _08440_);
  nor _21231_ (_12857_, _12856_, _12852_);
  nor _21232_ (_12858_, _12857_, _08406_);
  or _21233_ (_12859_, _08389_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  or _21234_ (_12860_, _08234_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  and _21235_ (_12861_, _12860_, _12859_);
  and _21236_ (_12862_, _12861_, _08441_);
  or _21237_ (_12863_, _08389_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  or _21238_ (_12864_, _08234_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  and _21239_ (_12865_, _12864_, _12863_);
  and _21240_ (_12866_, _12865_, _08440_);
  or _21241_ (_12867_, _12866_, _12862_);
  and _21242_ (_12868_, _12867_, _08467_);
  or _21243_ (_12869_, _08389_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  or _21244_ (_12870_, _08234_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  and _21245_ (_12871_, _12870_, _12869_);
  and _21246_ (_12872_, _12871_, _08441_);
  or _21247_ (_12873_, _08389_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  or _21248_ (_12874_, _08234_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  and _21249_ (_12875_, _12874_, _12873_);
  and _21250_ (_12876_, _12875_, _08440_);
  or _21251_ (_12877_, _12876_, _12872_);
  and _21252_ (_12878_, _12877_, _08480_);
  or _21253_ (_12879_, _12878_, _12868_);
  or _21254_ (_12880_, _12879_, _12858_);
  nor _21255_ (_12881_, _12880_, _12848_);
  nor _21256_ (_12882_, _12881_, _08439_);
  or _21257_ (\oc8051_symbolic_cxrom1.cxrom_data_out [11], _12882_, _12838_);
  and _21258_ (_12883_, _08439_, word_in[12]);
  or _21259_ (_12884_, _08389_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  or _21260_ (_12885_, _08234_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  and _21261_ (_12886_, _12885_, _12884_);
  and _21262_ (_12887_, _12886_, _08441_);
  or _21263_ (_12888_, _08389_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  or _21264_ (_12889_, _08234_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  and _21265_ (_12890_, _12889_, _12888_);
  and _21266_ (_12891_, _12890_, _08440_);
  or _21267_ (_12892_, _12891_, _12887_);
  and _21268_ (_12893_, _12892_, _08402_);
  or _21269_ (_12894_, _08389_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  or _21270_ (_12895_, _08234_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  and _21271_ (_12896_, _12895_, _12894_);
  and _21272_ (_12897_, _12896_, _08441_);
  or _21273_ (_12898_, _08389_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  or _21274_ (_12899_, _08234_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  and _21275_ (_12900_, _12899_, _12898_);
  and _21276_ (_12901_, _12900_, _08440_);
  nor _21277_ (_12902_, _12901_, _12897_);
  nor _21278_ (_12903_, _12902_, _08406_);
  or _21279_ (_12904_, _08389_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  or _21280_ (_12905_, _08234_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  and _21281_ (_12906_, _12905_, _12904_);
  and _21282_ (_12907_, _12906_, _08441_);
  or _21283_ (_12908_, _08389_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  or _21284_ (_12909_, _08234_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  and _21285_ (_12910_, _12909_, _12908_);
  and _21286_ (_12911_, _12910_, _08440_);
  or _21287_ (_12912_, _12911_, _12907_);
  and _21288_ (_12913_, _12912_, _08467_);
  or _21289_ (_12914_, _08389_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  or _21290_ (_12915_, _08234_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  and _21291_ (_12916_, _12915_, _12914_);
  and _21292_ (_12917_, _12916_, _08441_);
  or _21293_ (_12918_, _08389_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  or _21294_ (_12919_, _08234_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  and _21295_ (_12920_, _12919_, _12918_);
  and _21296_ (_12921_, _12920_, _08440_);
  or _21297_ (_12922_, _12921_, _12917_);
  and _21298_ (_12923_, _12922_, _08480_);
  or _21299_ (_12924_, _12923_, _12913_);
  or _21300_ (_12925_, _12924_, _12903_);
  nor _21301_ (_12926_, _12925_, _12893_);
  nor _21302_ (_12927_, _12926_, _08439_);
  or _21303_ (\oc8051_symbolic_cxrom1.cxrom_data_out [12], _12927_, _12883_);
  and _21304_ (_12928_, _08439_, word_in[13]);
  or _21305_ (_12929_, _08389_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  or _21306_ (_12930_, _08234_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  and _21307_ (_12931_, _12930_, _12929_);
  and _21308_ (_12932_, _12931_, _08441_);
  or _21309_ (_12933_, _08389_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  or _21310_ (_12934_, _08234_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  and _21311_ (_12935_, _12934_, _12933_);
  and _21312_ (_12936_, _12935_, _08440_);
  or _21313_ (_12937_, _12936_, _12932_);
  and _21314_ (_12938_, _12937_, _08402_);
  or _21315_ (_12939_, _08389_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  or _21316_ (_12940_, _08234_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  and _21317_ (_12941_, _12940_, _12939_);
  and _21318_ (_12942_, _12941_, _08441_);
  or _21319_ (_12943_, _08389_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  or _21320_ (_12944_, _08234_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  and _21321_ (_12945_, _12944_, _12943_);
  and _21322_ (_12946_, _12945_, _08440_);
  nor _21323_ (_12947_, _12946_, _12942_);
  nor _21324_ (_12948_, _12947_, _08406_);
  or _21325_ (_12949_, _08389_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  or _21326_ (_12950_, _08234_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  and _21327_ (_12951_, _12950_, _12949_);
  and _21328_ (_12952_, _12951_, _08441_);
  or _21329_ (_12953_, _08389_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  or _21330_ (_12954_, _08234_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  and _21331_ (_12955_, _12954_, _12953_);
  and _21332_ (_12956_, _12955_, _08440_);
  or _21333_ (_12957_, _12956_, _12952_);
  and _21334_ (_12958_, _12957_, _08467_);
  or _21335_ (_12959_, _08389_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  or _21336_ (_12960_, _08234_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  and _21337_ (_12961_, _12960_, _12959_);
  and _21338_ (_12962_, _12961_, _08441_);
  or _21339_ (_12963_, _08389_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  or _21340_ (_12964_, _08234_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  and _21341_ (_12965_, _12964_, _12963_);
  and _21342_ (_12966_, _12965_, _08440_);
  or _21343_ (_12967_, _12966_, _12962_);
  and _21344_ (_12968_, _12967_, _08480_);
  or _21345_ (_12969_, _12968_, _12958_);
  or _21346_ (_12970_, _12969_, _12948_);
  nor _21347_ (_12971_, _12970_, _12938_);
  nor _21348_ (_12972_, _12971_, _08439_);
  or _21349_ (\oc8051_symbolic_cxrom1.cxrom_data_out [13], _12972_, _12928_);
  and _21350_ (_12973_, _08439_, word_in[14]);
  or _21351_ (_12974_, _08389_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  or _21352_ (_12975_, _08234_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  and _21353_ (_12976_, _12975_, _12974_);
  and _21354_ (_12977_, _12976_, _08441_);
  or _21355_ (_12978_, _08389_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  or _21356_ (_12979_, _08234_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  and _21357_ (_12980_, _12979_, _12978_);
  and _21358_ (_12981_, _12980_, _08440_);
  or _21359_ (_12982_, _12981_, _12977_);
  and _21360_ (_12983_, _12982_, _08402_);
  or _21361_ (_12984_, _08389_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  or _21362_ (_12985_, _08234_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  and _21363_ (_12986_, _12985_, _12984_);
  and _21364_ (_12987_, _12986_, _08441_);
  or _21365_ (_12988_, _08389_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  or _21366_ (_12989_, _08234_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  and _21367_ (_12990_, _12989_, _12988_);
  and _21368_ (_12991_, _12990_, _08440_);
  nor _21369_ (_12992_, _12991_, _12987_);
  nor _21370_ (_12993_, _12992_, _08406_);
  or _21371_ (_12994_, _08389_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  or _21372_ (_12995_, _08234_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  and _21373_ (_12996_, _12995_, _12994_);
  and _21374_ (_12997_, _12996_, _08441_);
  or _21375_ (_12998_, _08389_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  or _21376_ (_12999_, _08234_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  and _21377_ (_13000_, _12999_, _12998_);
  and _21378_ (_13001_, _13000_, _08440_);
  or _21379_ (_13002_, _13001_, _12997_);
  and _21380_ (_13003_, _13002_, _08467_);
  or _21381_ (_13004_, _08389_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  or _21382_ (_13005_, _08234_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  and _21383_ (_13006_, _13005_, _13004_);
  and _21384_ (_13007_, _13006_, _08441_);
  or _21385_ (_13008_, _08389_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  or _21386_ (_13009_, _08234_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  and _21387_ (_13010_, _13009_, _13008_);
  and _21388_ (_13011_, _13010_, _08440_);
  or _21389_ (_13012_, _13011_, _13007_);
  and _21390_ (_13013_, _13012_, _08480_);
  or _21391_ (_13014_, _13013_, _13003_);
  or _21392_ (_13015_, _13014_, _12993_);
  nor _21393_ (_13016_, _13015_, _12983_);
  nor _21394_ (_13017_, _13016_, _08439_);
  or _21395_ (\oc8051_symbolic_cxrom1.cxrom_data_out [14], _13017_, _12973_);
  and _21396_ (_13018_, _08533_, word_in[16]);
  and _21397_ (_13019_, _12395_, _08257_);
  and _21398_ (_13020_, _12389_, _08260_);
  or _21399_ (_13021_, _13020_, _13019_);
  and _21400_ (_13022_, _12384_, _08279_);
  and _21401_ (_13023_, _12379_, _08267_);
  or _21402_ (_13024_, _13023_, _13022_);
  or _21403_ (_13025_, _13024_, _13021_);
  or _21404_ (_13026_, _13025_, _08502_);
  and _21405_ (_13027_, _12409_, _08260_);
  and _21406_ (_13028_, _12401_, _08267_);
  or _21407_ (_13029_, _13028_, _13027_);
  and _21408_ (_13030_, _12415_, _08257_);
  and _21409_ (_13031_, _12405_, _08279_);
  or _21410_ (_13032_, _13031_, _13030_);
  nor _21411_ (_13033_, _13032_, _13029_);
  nand _21412_ (_13034_, _13033_, _08502_);
  nand _21413_ (_13035_, _13034_, _13026_);
  nor _21414_ (_13036_, _13035_, _08533_);
  or _21415_ (\oc8051_symbolic_cxrom1.cxrom_data_out [16], _13036_, _13018_);
  and _21416_ (_13037_, _08533_, word_in[17]);
  and _21417_ (_13038_, _12428_, _08279_);
  and _21418_ (_13039_, _12424_, _08267_);
  or _21419_ (_13040_, _13039_, _13038_);
  and _21420_ (_13041_, _12438_, _08257_);
  and _21421_ (_13042_, _12432_, _08260_);
  or _21422_ (_13043_, _13042_, _13041_);
  or _21423_ (_13044_, _13043_, _13040_);
  or _21424_ (_13045_, _13044_, _08502_);
  and _21425_ (_13046_, _12460_, _08257_);
  and _21426_ (_13047_, _12449_, _08279_);
  or _21427_ (_13048_, _13047_, _13046_);
  and _21428_ (_13049_, _12453_, _08260_);
  and _21429_ (_13050_, _12445_, _08267_);
  or _21430_ (_13051_, _13050_, _13049_);
  nor _21431_ (_13052_, _13051_, _13048_);
  nand _21432_ (_13053_, _13052_, _08502_);
  nand _21433_ (_13054_, _13053_, _13045_);
  nor _21434_ (_13055_, _13054_, _08533_);
  or _21435_ (\oc8051_symbolic_cxrom1.cxrom_data_out [17], _13055_, _13037_);
  and _21436_ (_13056_, _08533_, word_in[18]);
  and _21437_ (_13057_, _12484_, _08257_);
  and _21438_ (_13058_, _12478_, _08260_);
  or _21439_ (_13059_, _13058_, _13057_);
  and _21440_ (_13060_, _12474_, _08279_);
  and _21441_ (_13061_, _12470_, _08267_);
  or _21442_ (_13062_, _13061_, _13060_);
  nor _21443_ (_13063_, _13062_, _13059_);
  nor _21444_ (_13064_, _13063_, _08502_);
  and _21445_ (_13065_, _12504_, _08257_);
  and _21446_ (_13066_, _12498_, _08260_);
  or _21447_ (_13067_, _13066_, _13065_);
  and _21448_ (_13068_, _12494_, _08279_);
  and _21449_ (_13069_, _12490_, _08267_);
  or _21450_ (_13070_, _13069_, _13068_);
  or _21451_ (_13071_, _13070_, _13067_);
  and _21452_ (_13072_, _13071_, _08502_);
  nor _21453_ (_13073_, _13072_, _13064_);
  nor _21454_ (_13074_, _13073_, _08533_);
  or _21455_ (\oc8051_symbolic_cxrom1.cxrom_data_out [18], _13074_, _13056_);
  and _21456_ (_13075_, _08533_, word_in[19]);
  and _21457_ (_13076_, _12524_, _08257_);
  and _21458_ (_13077_, _12517_, _08279_);
  or _21459_ (_13078_, _13077_, _13076_);
  and _21460_ (_13079_, _12528_, _08260_);
  and _21461_ (_13080_, _12513_, _08267_);
  or _21462_ (_13081_, _13080_, _13079_);
  or _21463_ (_13082_, _13081_, _13078_);
  or _21464_ (_13083_, _13082_, _08502_);
  and _21465_ (_13084_, _12535_, _08279_);
  and _21466_ (_13085_, _12539_, _08267_);
  or _21467_ (_13086_, _13085_, _13084_);
  and _21468_ (_13087_, _12544_, _08257_);
  and _21469_ (_13088_, _12548_, _08260_);
  or _21470_ (_13089_, _13088_, _13087_);
  nor _21471_ (_13090_, _13089_, _13086_);
  nand _21472_ (_13091_, _13090_, _08502_);
  nand _21473_ (_13092_, _13091_, _13083_);
  nor _21474_ (_13093_, _13092_, _08533_);
  or _21475_ (\oc8051_symbolic_cxrom1.cxrom_data_out [19], _13093_, _13075_);
  and _21476_ (_13094_, _08533_, word_in[20]);
  and _21477_ (_13095_, _12572_, _08257_);
  and _21478_ (_13096_, _12566_, _08279_);
  or _21479_ (_13097_, _13096_, _13095_);
  and _21480_ (_13098_, _12562_, _08260_);
  and _21481_ (_13099_, _12558_, _08267_);
  or _21482_ (_13100_, _13099_, _13098_);
  or _21483_ (_13101_, _13100_, _13097_);
  or _21484_ (_13102_, _13101_, _08502_);
  and _21485_ (_13103_, _12582_, _08279_);
  and _21486_ (_13104_, _12578_, _08267_);
  or _21487_ (_13105_, _13104_, _13103_);
  and _21488_ (_13107_, _12592_, _08257_);
  and _21489_ (_13108_, _12586_, _08260_);
  or _21490_ (_13110_, _13108_, _13107_);
  nor _21491_ (_13111_, _13110_, _13105_);
  nand _21492_ (_13112_, _13111_, _08502_);
  nand _21493_ (_13113_, _13112_, _13102_);
  nor _21494_ (_13114_, _13113_, _08533_);
  or _21495_ (\oc8051_symbolic_cxrom1.cxrom_data_out [20], _13114_, _13094_);
  and _21496_ (_13115_, _08533_, word_in[21]);
  and _21497_ (_13116_, _12610_, _08260_);
  and _21498_ (_13117_, _12616_, _08257_);
  or _21499_ (_13118_, _13117_, _13116_);
  and _21500_ (_13119_, _12606_, _08279_);
  and _21501_ (_13120_, _12602_, _08286_);
  or _21502_ (_13121_, _13120_, _13119_);
  or _21503_ (_13122_, _13121_, _13118_);
  or _21504_ (_13123_, _13122_, _08502_);
  and _21505_ (_13124_, _12626_, _08279_);
  and _21506_ (_13125_, _12622_, _08267_);
  or _21507_ (_13126_, _13125_, _13124_);
  and _21508_ (_13127_, _12636_, _08257_);
  and _21509_ (_13128_, _12630_, _08260_);
  or _21510_ (_13130_, _13128_, _13127_);
  nor _21511_ (_13131_, _13130_, _13126_);
  nand _21512_ (_13133_, _13131_, _08502_);
  nand _21513_ (_13134_, _13133_, _13123_);
  nor _21514_ (_13136_, _13134_, _08533_);
  or _21515_ (\oc8051_symbolic_cxrom1.cxrom_data_out [21], _13136_, _13115_);
  and _21516_ (_13137_, _08533_, word_in[22]);
  and _21517_ (_13138_, _12659_, _08257_);
  and _21518_ (_13140_, _12645_, _08279_);
  or _21519_ (_13141_, _13140_, _13138_);
  and _21520_ (_13143_, _12649_, _08260_);
  and _21521_ (_13144_, _12653_, _08267_);
  or _21522_ (_13145_, _13144_, _13143_);
  or _21523_ (_13146_, _13145_, _13141_);
  or _21524_ (_13147_, _13146_, _08502_);
  and _21525_ (_13148_, _12679_, _08257_);
  and _21526_ (_13149_, _12665_, _08279_);
  or _21527_ (_13151_, _13149_, _13148_);
  and _21528_ (_13152_, _12673_, _08260_);
  and _21529_ (_13153_, _12669_, _08267_);
  or _21530_ (_13155_, _13153_, _13152_);
  nor _21531_ (_13156_, _13155_, _13151_);
  nand _21532_ (_13158_, _13156_, _08502_);
  nand _21533_ (_13159_, _13158_, _13147_);
  nor _21534_ (_13160_, _13159_, _08533_);
  or _21535_ (\oc8051_symbolic_cxrom1.cxrom_data_out [22], _13160_, _13137_);
  and _21536_ (_13161_, _08595_, word_in[24]);
  and _21537_ (_13162_, _12708_, _08441_);
  and _21538_ (_13164_, _12704_, _08440_);
  or _21539_ (_13165_, _13164_, _13162_);
  and _21540_ (_13166_, _13165_, _08567_);
  and _21541_ (_13168_, _12718_, _08441_);
  and _21542_ (_13169_, _12714_, _08440_);
  or _21543_ (_13170_, _13169_, _13168_);
  and _21544_ (_13171_, _13170_, _08572_);
  and _21545_ (_13172_, _12728_, _08441_);
  and _21546_ (_13173_, _12724_, _08440_);
  or _21547_ (_13174_, _13173_, _13172_);
  and _21548_ (_13176_, _13174_, _08607_);
  and _21549_ (_13177_, _12738_, _08441_);
  and _21550_ (_13178_, _12734_, _08440_);
  or _21551_ (_13179_, _13178_, _13177_);
  and _21552_ (_13180_, _13179_, _08613_);
  or _21553_ (_13181_, _13180_, _13176_);
  or _21554_ (_13182_, _13181_, _13171_);
  nor _21555_ (_13183_, _13182_, _13166_);
  nor _21556_ (_13184_, _13183_, _08595_);
  or _21557_ (\oc8051_symbolic_cxrom1.cxrom_data_out [24], _13184_, _13161_);
  and _21558_ (_13185_, _08595_, word_in[25]);
  and _21559_ (_13186_, _12753_, _08441_);
  and _21560_ (_13187_, _12749_, _08440_);
  or _21561_ (_13188_, _13187_, _13186_);
  and _21562_ (_13189_, _13188_, _08567_);
  and _21563_ (_13190_, _12763_, _08441_);
  and _21564_ (_13192_, _12759_, _08440_);
  or _21565_ (_13193_, _13192_, _13190_);
  and _21566_ (_13195_, _13193_, _08572_);
  and _21567_ (_13196_, _12774_, _08441_);
  and _21568_ (_13198_, _12769_, _08440_);
  or _21569_ (_13199_, _13198_, _13196_);
  and _21570_ (_13200_, _13199_, _08607_);
  and _21571_ (_13201_, _12784_, _08441_);
  and _21572_ (_13202_, _12780_, _08440_);
  or _21573_ (_13204_, _13202_, _13201_);
  and _21574_ (_13205_, _13204_, _08613_);
  or _21575_ (_13207_, _13205_, _13200_);
  or _21576_ (_13208_, _13207_, _13195_);
  nor _21577_ (_13210_, _13208_, _13189_);
  nor _21578_ (_13211_, _13210_, _08595_);
  or _21579_ (\oc8051_symbolic_cxrom1.cxrom_data_out [25], _13211_, _13185_);
  and _21580_ (_13213_, _08595_, word_in[26]);
  and _21581_ (_13214_, _12799_, _08441_);
  and _21582_ (_13216_, _12795_, _08440_);
  or _21583_ (_13217_, _13216_, _13214_);
  and _21584_ (_13218_, _13217_, _08567_);
  and _21585_ (_13220_, _12810_, _08441_);
  and _21586_ (_13221_, _12805_, _08440_);
  or _21587_ (_13223_, _13221_, _13220_);
  and _21588_ (_13224_, _13223_, _08572_);
  and _21589_ (_13225_, _12820_, _08441_);
  and _21590_ (_13226_, _12816_, _08440_);
  or _21591_ (_13227_, _13226_, _13225_);
  and _21592_ (_13228_, _13227_, _08607_);
  and _21593_ (_13229_, _12830_, _08441_);
  and _21594_ (_13230_, _12826_, _08440_);
  or _21595_ (_13231_, _13230_, _13229_);
  and _21596_ (_13232_, _13231_, _08613_);
  or _21597_ (_13233_, _13232_, _13228_);
  or _21598_ (_13234_, _13233_, _13224_);
  nor _21599_ (_13235_, _13234_, _13218_);
  nor _21600_ (_13236_, _13235_, _08595_);
  or _21601_ (\oc8051_symbolic_cxrom1.cxrom_data_out [26], _13236_, _13213_);
  and _21602_ (_13238_, _08595_, word_in[27]);
  and _21603_ (_13239_, _12855_, _08441_);
  and _21604_ (_13240_, _12851_, _08440_);
  or _21605_ (_13241_, _13240_, _13239_);
  and _21606_ (_13243_, _13241_, _08572_);
  and _21607_ (_13244_, _12845_, _08441_);
  and _21608_ (_13246_, _12841_, _08440_);
  or _21609_ (_13247_, _13246_, _13244_);
  and _21610_ (_13248_, _13247_, _08567_);
  and _21611_ (_13249_, _12865_, _08441_);
  and _21612_ (_13251_, _12861_, _08440_);
  or _21613_ (_13252_, _13251_, _13249_);
  and _21614_ (_13253_, _13252_, _08607_);
  and _21615_ (_13254_, _12875_, _08441_);
  and _21616_ (_13255_, _12871_, _08440_);
  or _21617_ (_13256_, _13255_, _13254_);
  and _21618_ (_13257_, _13256_, _08613_);
  or _21619_ (_13258_, _13257_, _13253_);
  or _21620_ (_13259_, _13258_, _13248_);
  nor _21621_ (_13260_, _13259_, _13243_);
  nor _21622_ (_13261_, _13260_, _08595_);
  or _21623_ (\oc8051_symbolic_cxrom1.cxrom_data_out [27], _13261_, _13238_);
  and _21624_ (_13263_, _08595_, word_in[28]);
  and _21625_ (_13264_, _12890_, _08441_);
  and _21626_ (_13265_, _12886_, _08440_);
  or _21627_ (_13266_, _13265_, _13264_);
  and _21628_ (_13267_, _13266_, _08567_);
  and _21629_ (_13268_, _12900_, _08441_);
  and _21630_ (_13269_, _12896_, _08440_);
  or _21631_ (_13270_, _13269_, _13268_);
  and _21632_ (_13272_, _13270_, _08572_);
  and _21633_ (_13273_, _12910_, _08441_);
  and _21634_ (_13274_, _12906_, _08440_);
  or _21635_ (_13275_, _13274_, _13273_);
  and _21636_ (_13277_, _13275_, _08607_);
  and _21637_ (_13278_, _12920_, _08441_);
  and _21638_ (_13280_, _12916_, _08440_);
  or _21639_ (_13281_, _13280_, _13278_);
  and _21640_ (_13283_, _13281_, _08613_);
  or _21641_ (_13284_, _13283_, _13277_);
  or _21642_ (_13285_, _13284_, _13272_);
  nor _21643_ (_13286_, _13285_, _13267_);
  nor _21644_ (_13287_, _13286_, _08595_);
  or _21645_ (\oc8051_symbolic_cxrom1.cxrom_data_out [28], _13287_, _13263_);
  and _21646_ (_13288_, _08595_, word_in[29]);
  and _21647_ (_13289_, _12945_, _08441_);
  and _21648_ (_13290_, _12941_, _08440_);
  or _21649_ (_13291_, _13290_, _13289_);
  and _21650_ (_13292_, _13291_, _08572_);
  and _21651_ (_13294_, _12935_, _08441_);
  and _21652_ (_13295_, _12931_, _08440_);
  or _21653_ (_13297_, _13295_, _13294_);
  and _21654_ (_13298_, _13297_, _08567_);
  and _21655_ (_13299_, _12955_, _08441_);
  and _21656_ (_13300_, _12951_, _08440_);
  or _21657_ (_13302_, _13300_, _13299_);
  and _21658_ (_13303_, _13302_, _08607_);
  and _21659_ (_13304_, _12965_, _08441_);
  and _21660_ (_13305_, _12961_, _08440_);
  or _21661_ (_13306_, _13305_, _13304_);
  and _21662_ (_13307_, _13306_, _08613_);
  or _21663_ (_13308_, _13307_, _13303_);
  or _21664_ (_13309_, _13308_, _13298_);
  nor _21665_ (_13310_, _13309_, _13292_);
  nor _21666_ (_13311_, _13310_, _08595_);
  or _21667_ (\oc8051_symbolic_cxrom1.cxrom_data_out [29], _13311_, _13288_);
  and _21668_ (_13312_, _08595_, word_in[30]);
  and _21669_ (_13313_, _12980_, _08441_);
  and _21670_ (_13314_, _12976_, _08440_);
  or _21671_ (_13315_, _13314_, _13313_);
  and _21672_ (_13316_, _13315_, _08567_);
  and _21673_ (_13317_, _12990_, _08441_);
  and _21674_ (_13318_, _12986_, _08440_);
  or _21675_ (_13319_, _13318_, _13317_);
  and _21676_ (_13320_, _13319_, _08572_);
  and _21677_ (_13321_, _13000_, _08441_);
  and _21678_ (_13322_, _12996_, _08440_);
  or _21679_ (_13323_, _13322_, _13321_);
  and _21680_ (_13324_, _13323_, _08607_);
  and _21681_ (_13325_, _13010_, _08441_);
  and _21682_ (_13326_, _13006_, _08440_);
  or _21683_ (_13327_, _13326_, _13325_);
  and _21684_ (_13328_, _13327_, _08613_);
  or _21685_ (_13329_, _13328_, _13324_);
  or _21686_ (_13331_, _13329_, _13320_);
  nor _21687_ (_13332_, _13331_, _13316_);
  nor _21688_ (_13333_, _13332_, _08595_);
  or _21689_ (\oc8051_symbolic_cxrom1.cxrom_data_out [30], _13333_, _13312_);
  and _21690_ (_13334_, _05552_, \oc8051_top_1.oc8051_memory_interface1.int_ack_buff );
  and _21691_ (_11498_, _13334_, _05671_);
  and _21692_ (_11504_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , _05552_);
  nor _21693_ (_11517_, _11469_, rst);
  or _21694_ (_13335_, _05550_, \oc8051_top_1.oc8051_rom1.data_o [9]);
  nand _21695_ (_13336_, _05550_, _11609_);
  and _21696_ (_13337_, _13336_, _05552_);
  and _21697_ (_11551_, _13337_, _13335_);
  or _21698_ (_13339_, _09144_, _09105_);
  nor _21699_ (_13341_, _09039_, _09145_);
  and _21700_ (_13342_, _13341_, _13339_);
  nor _21701_ (_13343_, _09038_, _06489_);
  or _21702_ (_13344_, _13343_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _21703_ (_13345_, _13344_, _13342_);
  or _21704_ (_13346_, _05605_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and _21705_ (_13347_, _13346_, _05552_);
  and _21706_ (_11554_, _13347_, _13345_);
  nor _21707_ (_13349_, _09142_, _09139_);
  nor _21708_ (_13350_, _13349_, _09143_);
  or _21709_ (_13352_, _13350_, _09039_);
  or _21710_ (_13353_, _09038_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _21711_ (_13354_, _13353_, _07933_);
  and _21712_ (_13355_, _13354_, _13352_);
  and _21713_ (_13356_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and _21714_ (_13357_, _13356_, _05552_);
  or _21715_ (_11588_, _13357_, _13355_);
  nand _21716_ (_13358_, _07711_, _06973_);
  and _21717_ (_13359_, _08048_, _06060_);
  nor _21718_ (_13360_, _06060_, _06201_);
  nor _21719_ (_13361_, _13360_, _13359_);
  or _21720_ (_13362_, _13361_, _08924_);
  and _21721_ (_13363_, _08935_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor _21722_ (_13365_, _13363_, _07260_);
  and _21723_ (_13366_, _13365_, _13362_);
  nand _21724_ (_13367_, _13366_, _13358_);
  or _21725_ (_13368_, _08228_, _07261_);
  and _21726_ (_13369_, _13368_, _13367_);
  and _21727_ (_11659_, _13369_, _05552_);
  nand _21728_ (_13371_, _06949_, _06560_);
  or _21729_ (_13372_, _06949_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  and _21730_ (_13373_, _13372_, _05552_);
  and _21731_ (_11681_, _13373_, _13371_);
  nor _21732_ (_13374_, _07211_, _06330_);
  and _21733_ (_13375_, _07211_, _06330_);
  or _21734_ (_13377_, _13375_, _13374_);
  and _21735_ (_11685_, _13377_, _05552_);
  and _21736_ (_13379_, _12299_, \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  or _21737_ (_13380_, _10898_, _05820_);
  and _21738_ (_13381_, _13380_, _10905_);
  or _21739_ (_13382_, _13381_, _10941_);
  or _21740_ (_13383_, _10943_, _10899_);
  or _21741_ (_13384_, _13383_, _13382_);
  or _21742_ (_13385_, _11174_, _12282_);
  and _21743_ (_13386_, _06567_, _05830_);
  or _21744_ (_13387_, _13386_, _12307_);
  or _21745_ (_13389_, _13387_, _13385_);
  or _21746_ (_13390_, _13389_, _10927_);
  or _21747_ (_13391_, _13390_, _13384_);
  or _21748_ (_13392_, _11160_, _11151_);
  and _21749_ (_13394_, _06567_, _05846_);
  or _21750_ (_13395_, _13394_, _12272_);
  or _21751_ (_13397_, _13395_, _13392_);
  or _21752_ (_13398_, _12328_, _11155_);
  or _21753_ (_13399_, _13398_, _12291_);
  or _21754_ (_13400_, _13399_, _13397_);
  or _21755_ (_13401_, _13400_, _13391_);
  and _21756_ (_13402_, _13401_, _06576_);
  or _21757_ (_11720_, _13402_, _13379_);
  and _21758_ (_11741_, _07646_, _05552_);
  nor _21759_ (_13404_, _07939_, _07388_);
  and _21760_ (_13405_, _07939_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  or _21761_ (_13407_, _13405_, _13404_);
  and _21762_ (_11748_, _13407_, _05552_);
  and _21763_ (_13408_, _07939_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  and _21764_ (_13409_, _07976_, _07937_);
  or _21765_ (_13410_, _13409_, _13408_);
  and _21766_ (_11755_, _13410_, _05552_);
  and _21767_ (_13411_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9], _05556_);
  and _21768_ (_13412_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _21769_ (_13413_, _13412_, _13411_);
  and _21770_ (_11758_, _13413_, _05552_);
  not _21771_ (_13414_, _11774_);
  or _21772_ (_13415_, _12037_, _11828_);
  or _21773_ (_13416_, _12029_, _12032_);
  and _21774_ (_13417_, _13416_, _13415_);
  nor _21775_ (_13418_, _13417_, _06487_);
  and _21776_ (_13419_, _13417_, _06487_);
  or _21777_ (_13420_, _13419_, _13418_);
  and _21778_ (_13421_, _13420_, _12161_);
  and _21779_ (_13422_, _11811_, _07574_);
  and _21780_ (_13423_, _11784_, _07600_);
  nor _21781_ (_13424_, _11805_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor _21782_ (_13425_, _13424_, _11806_);
  and _21783_ (_13426_, _13425_, _11792_);
  and _21784_ (_13427_, _11780_, _11391_);
  and _21785_ (_13428_, _11817_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or _21786_ (_13429_, _13428_, _13427_);
  or _21787_ (_13430_, _13429_, _13426_);
  or _21788_ (_13431_, _13430_, _13423_);
  or _21789_ (_13432_, _13431_, _13422_);
  or _21790_ (_13433_, _13432_, _13421_);
  or _21791_ (_13434_, _13433_, _13414_);
  nor _21792_ (_13435_, _12071_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor _21793_ (_13436_, _13435_, _12072_);
  or _21794_ (_13437_, _13436_, _11774_);
  and _21795_ (_13438_, _13437_, _05552_);
  and _21796_ (_11798_, _13438_, _13434_);
  nand _21797_ (_13439_, _12028_, _11828_);
  or _21798_ (_13440_, _12036_, _11828_);
  and _21799_ (_13441_, _13440_, _13439_);
  nand _21800_ (_13442_, _13441_, _06085_);
  or _21801_ (_13443_, _13441_, _06085_);
  and _21802_ (_13444_, _13443_, _12161_);
  and _21803_ (_13445_, _13444_, _13442_);
  and _21804_ (_13446_, _11811_, _07635_);
  and _21805_ (_13447_, _11784_, _07663_);
  nor _21806_ (_13448_, _11804_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor _21807_ (_13449_, _13448_, _11805_);
  and _21808_ (_13450_, _13449_, _11792_);
  and _21809_ (_13451_, _11780_, _11449_);
  and _21810_ (_13452_, _11817_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or _21811_ (_13453_, _13452_, _13451_);
  or _21812_ (_13454_, _13453_, _13450_);
  nor _21813_ (_13455_, _13454_, _13447_);
  nand _21814_ (_13456_, _13455_, _11774_);
  or _21815_ (_13457_, _13456_, _13446_);
  or _21816_ (_13458_, _13457_, _13445_);
  nor _21817_ (_13459_, _12069_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor _21818_ (_13460_, _13459_, _12071_);
  or _21819_ (_13461_, _13460_, _11774_);
  and _21820_ (_13462_, _13461_, _05552_);
  and _21821_ (_11826_, _13462_, _13458_);
  not _21822_ (_13463_, _11650_);
  and _21823_ (_13464_, _11704_, _13463_);
  not _21824_ (_13465_, _11509_);
  not _21825_ (_13466_, _11452_);
  not _21826_ (_13467_, _11335_);
  nand _21827_ (_13468_, _11395_, _13467_);
  or _21828_ (_13469_, _13468_, _13466_);
  or _21829_ (_13471_, _13469_, _13465_);
  not _21830_ (_13472_, _13471_);
  and _21831_ (_13473_, _11763_, _11279_);
  and _21832_ (_13474_, _13473_, _13472_);
  and _21833_ (_13475_, _13474_, _13464_);
  and _21834_ (_13476_, _13475_, _07485_);
  nor _21835_ (_13477_, _13476_, rst);
  and _21836_ (_13478_, _07711_, _05552_);
  or _21837_ (_13479_, _13478_, _13477_);
  and _21838_ (_13480_, _11704_, _11650_);
  not _21839_ (_13481_, _11763_);
  nor _21840_ (_13482_, _13481_, _11279_);
  and _21841_ (_13484_, _13482_, _13480_);
  nor _21842_ (_13485_, _11395_, _13466_);
  and _21843_ (_13486_, _11509_, _13467_);
  and _21844_ (_13487_, _13486_, _13485_);
  and _21845_ (_13488_, _13487_, _13484_);
  nand _21846_ (_13489_, _13488_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  nor _21847_ (_13491_, _11763_, _11279_);
  and _21848_ (_13492_, _13491_, _13480_);
  and _21849_ (_13494_, _13487_, _13492_);
  nand _21850_ (_13495_, _13494_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and _21851_ (_13496_, _13495_, _13489_);
  nor _21852_ (_13497_, _11704_, _13463_);
  and _21853_ (_13498_, _13491_, _13497_);
  and _21854_ (_13499_, _13487_, _13498_);
  nand _21855_ (_13500_, _13499_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and _21856_ (_13501_, _13482_, _13464_);
  and _21857_ (_13502_, _13487_, _13501_);
  nand _21858_ (_13503_, _13502_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  and _21859_ (_13504_, _13503_, _13500_);
  and _21860_ (_13505_, _13504_, _13496_);
  and _21861_ (_13507_, _13484_, _13472_);
  nand _21862_ (_13508_, _13507_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  nor _21863_ (_13509_, _11704_, _11650_);
  and _21864_ (_13510_, _13482_, _13509_);
  and _21865_ (_13511_, _13487_, _13510_);
  nand _21866_ (_13512_, _13511_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  and _21867_ (_13513_, _13512_, _13508_);
  nor _21868_ (_13514_, _13468_, _11452_);
  and _21869_ (_13515_, _13514_, _11509_);
  and _21870_ (_13516_, _13515_, _13484_);
  nand _21871_ (_13517_, _13516_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and _21872_ (_13518_, _13514_, _13465_);
  and _21873_ (_13519_, _13509_, _13481_);
  and _21874_ (_13520_, _13519_, _11279_);
  and _21875_ (_13521_, _13520_, _13518_);
  nand _21876_ (_13522_, _13521_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and _21877_ (_13523_, _13522_, _13517_);
  and _21878_ (_13524_, _13523_, _13513_);
  and _21879_ (_13525_, _13524_, _13505_);
  not _21880_ (_13526_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and _21881_ (_13527_, _13497_, _13482_);
  nand _21882_ (_13528_, _13527_, _13472_);
  or _21883_ (_13529_, _13528_, _13526_);
  not _21884_ (_13530_, _13510_);
  nor _21885_ (_13531_, _13530_, _13471_);
  nand _21886_ (_13532_, _13531_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and _21887_ (_13533_, _13532_, _13529_);
  and _21888_ (_13534_, _13501_, _13472_);
  nand _21889_ (_13535_, _13534_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and _21890_ (_13536_, _13498_, _13472_);
  nand _21891_ (_13537_, _13536_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and _21892_ (_13538_, _13537_, _13535_);
  and _21893_ (_13539_, _13538_, _13533_);
  nor _21894_ (_13540_, _13469_, _11509_);
  and _21895_ (_13541_, _13540_, _13527_);
  nand _21896_ (_13542_, _13541_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  and _21897_ (_13544_, _13484_, _13540_);
  nand _21898_ (_13545_, _13544_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  and _21899_ (_13546_, _13545_, _13542_);
  and _21900_ (_13547_, _13492_, _13472_);
  nand _21901_ (_13548_, _13547_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and _21902_ (_13549_, _13520_, _13472_);
  nand _21903_ (_13550_, _13549_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  and _21904_ (_13551_, _13550_, _13548_);
  and _21905_ (_13552_, _13551_, _13546_);
  and _21906_ (_13553_, _13552_, _13539_);
  and _21907_ (_13554_, _13553_, _13525_);
  and _21908_ (_13555_, _13497_, _13474_);
  nand _21909_ (_13556_, _13555_, _11700_);
  and _21910_ (_13557_, _13480_, _13473_);
  and _21911_ (_13559_, _13557_, _13465_);
  nor _21912_ (_13560_, _11395_, _11452_);
  and _21913_ (_13561_, _13560_, _13467_);
  and _21914_ (_13562_, _13561_, _13559_);
  nand _21915_ (_13563_, _13562_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  and _21916_ (_13565_, _13563_, _13556_);
  nand _21917_ (_13566_, _13475_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  nand _21918_ (_13567_, _13509_, _13473_);
  nor _21919_ (_13568_, _13567_, _13471_);
  nand _21920_ (_13570_, _13568_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and _21921_ (_13571_, _13570_, _13566_);
  and _21922_ (_13572_, _13571_, _13565_);
  not _21923_ (_13573_, _13557_);
  nor _21924_ (_13574_, _13573_, _13471_);
  and _21925_ (_13575_, _12283_, _05852_);
  or _21926_ (_13576_, _13575_, _05855_);
  nor _21927_ (_13577_, _13576_, _11169_);
  and _21928_ (_13578_, _10898_, _05854_);
  and _21929_ (_13579_, _13578_, _05669_);
  nor _21930_ (_13581_, _12331_, _13579_);
  and _21931_ (_13582_, _13581_, _13577_);
  and _21932_ (_13583_, _10909_, _10843_);
  or _21933_ (_13584_, _12330_, _05811_);
  nor _21934_ (_13585_, _13584_, _13583_);
  and _21935_ (_13586_, _13585_, _12315_);
  and _21936_ (_13588_, _13586_, _13582_);
  and _21937_ (_13589_, _13588_, _12319_);
  and _21938_ (_13591_, _13589_, _11159_);
  nor _21939_ (_13592_, _13591_, _11085_);
  nor _21940_ (_13593_, _13592_, p0_in[0]);
  not _21941_ (_13594_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  and _21942_ (_13595_, _13592_, _13594_);
  nor _21943_ (_13596_, _13595_, _13593_);
  nand _21944_ (_13597_, _13596_, _13574_);
  and _21945_ (_13598_, _13540_, _13557_);
  nor _21946_ (_13599_, _13592_, p1_in[0]);
  not _21947_ (_13600_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and _21948_ (_13601_, _13592_, _13600_);
  nor _21949_ (_13602_, _13601_, _13599_);
  nand _21950_ (_13603_, _13602_, _13598_);
  and _21951_ (_13604_, _13603_, _13597_);
  and _21952_ (_13605_, _13518_, _13557_);
  nor _21953_ (_13606_, _13592_, p3_in[0]);
  not _21954_ (_13607_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and _21955_ (_13608_, _13592_, _13607_);
  nor _21956_ (_13609_, _13608_, _13606_);
  nand _21957_ (_13610_, _13609_, _13605_);
  and _21958_ (_13611_, _13515_, _13557_);
  nor _21959_ (_13612_, _13592_, p2_in[0]);
  not _21960_ (_13613_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and _21961_ (_13614_, _13592_, _13613_);
  nor _21962_ (_13615_, _13614_, _13612_);
  nand _21963_ (_13616_, _13615_, _13611_);
  and _21964_ (_13617_, _13616_, _13610_);
  and _21965_ (_13618_, _13617_, _13604_);
  and _21966_ (_13619_, _13618_, _13572_);
  nor _21967_ (_13620_, _11509_, _11335_);
  and _21968_ (_13621_, _13620_, _13485_);
  and _21969_ (_13622_, _13621_, _13557_);
  nand _21970_ (_13623_, _07362_, _07275_);
  nand _21971_ (_13624_, _08920_, _13623_);
  or _21972_ (_13625_, _08920_, _13623_);
  nand _21973_ (_13626_, _13625_, _13624_);
  and _21974_ (_13627_, _12189_, _06973_);
  nor _21975_ (_13628_, _08057_, _06157_);
  or _21976_ (_13629_, _13628_, _08062_);
  and _21977_ (_13630_, _13629_, _08923_);
  and _21978_ (_13631_, _08935_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or _21979_ (_13632_, _13631_, _07260_);
  or _21980_ (_13633_, _13632_, _13630_);
  or _21981_ (_13634_, _13633_, _13627_);
  or _21982_ (_13635_, _12215_, _07261_);
  and _21983_ (_13636_, _13635_, _13634_);
  and _21984_ (_13637_, _07635_, _06973_);
  nand _21985_ (_13638_, _08635_, _06763_);
  or _21986_ (_13639_, _08635_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and _21987_ (_13640_, _13639_, _08923_);
  and _21988_ (_13641_, _13640_, _13638_);
  and _21989_ (_13642_, _08935_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or _21990_ (_13643_, _13642_, _07260_);
  or _21991_ (_13644_, _13643_, _13641_);
  or _21992_ (_13645_, _13644_, _13637_);
  or _21993_ (_13646_, _07663_, _07261_);
  and _21994_ (_13647_, _13646_, _13645_);
  or _21995_ (_13648_, _13647_, _13636_);
  nand _21996_ (_13649_, _13647_, _13636_);
  and _21997_ (_13650_, _13649_, _13648_);
  nand _21998_ (_13651_, _13650_, _13626_);
  or _21999_ (_13652_, _13650_, _13626_);
  nand _22000_ (_13653_, _13652_, _13651_);
  nand _22001_ (_13654_, _13368_, _13367_);
  nand _22002_ (_13655_, _13654_, _08942_);
  or _22003_ (_13656_, _13654_, _08942_);
  nand _22004_ (_13657_, _13656_, _13655_);
  or _22005_ (_13658_, _12137_, _12136_);
  nand _22006_ (_13659_, _08144_, _06973_);
  and _22007_ (_13660_, _08935_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor _22008_ (_13661_, _08013_, _06213_);
  nor _22009_ (_13662_, _13661_, _08015_);
  nor _22010_ (_13663_, _13662_, _08924_);
  nor _22011_ (_13664_, _13663_, _13660_);
  and _22012_ (_13665_, _13664_, _07261_);
  and _22013_ (_13666_, _13665_, _13659_);
  and _22014_ (_13667_, _08200_, _07260_);
  nor _22015_ (_13668_, _13667_, _13666_);
  nand _22016_ (_13669_, _13668_, _13658_);
  or _22017_ (_13670_, _13668_, _13658_);
  and _22018_ (_13671_, _13670_, _13669_);
  nand _22019_ (_13672_, _13671_, _13657_);
  or _22020_ (_13673_, _13671_, _13657_);
  nand _22021_ (_13674_, _13673_, _13672_);
  nand _22022_ (_13675_, _13674_, _13653_);
  or _22023_ (_13676_, _13674_, _13653_);
  nand _22024_ (_13677_, _13676_, _13675_);
  nand _22025_ (_13678_, _13677_, _13622_);
  and _22026_ (_13679_, _13557_, _11509_);
  and _22027_ (_13681_, _13561_, _13679_);
  nand _22028_ (_13683_, _13681_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and _22029_ (_13684_, _13683_, _13678_);
  and _22030_ (_13685_, _13684_, _13619_);
  and _22031_ (_13686_, _13685_, _13554_);
  and _22032_ (_13687_, _13622_, _11591_);
  and _22033_ (_13688_, _13509_, _13474_);
  and _22034_ (_13689_, _13688_, _07485_);
  nor _22035_ (_13690_, _13689_, _13687_);
  nor _22036_ (_13691_, _13690_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not _22037_ (_13692_, _13691_);
  nor _22038_ (_13693_, _10859_, _05971_);
  not _22039_ (_13694_, _13519_);
  and _22040_ (_13695_, _13694_, _13693_);
  and _22041_ (_13696_, _13695_, _11515_);
  or _22042_ (_13697_, _07260_, _06965_);
  and _22043_ (_13698_, _13681_, _13697_);
  nor _22044_ (_13699_, _13698_, _13696_);
  and _22045_ (_13700_, _13699_, _11772_);
  and _22046_ (_13701_, _13700_, _13692_);
  not _22047_ (_13702_, _13701_);
  nor _22048_ (_13703_, _13702_, _13686_);
  not _22049_ (_13704_, _13476_);
  nor _22050_ (_13705_, _13494_, _13488_);
  nor _22051_ (_13706_, _13502_, _13499_);
  and _22052_ (_13707_, _13706_, _13705_);
  nor _22053_ (_13708_, _13511_, _13507_);
  nor _22054_ (_13710_, _13521_, _13516_);
  and _22055_ (_13711_, _13710_, _13708_);
  and _22056_ (_13712_, _13711_, _13707_);
  not _22057_ (_13713_, _13528_);
  nor _22058_ (_13715_, _13531_, _13713_);
  nor _22059_ (_13716_, _13536_, _13534_);
  and _22060_ (_13718_, _13716_, _13715_);
  nor _22061_ (_13719_, _13544_, _13541_);
  nor _22062_ (_13721_, _13549_, _13547_);
  and _22063_ (_13722_, _13721_, _13719_);
  and _22064_ (_13723_, _13722_, _13718_);
  and _22065_ (_13724_, _13723_, _13712_);
  nor _22066_ (_13725_, _13681_, _13622_);
  not _22067_ (_13727_, _13468_);
  nand _22068_ (_13728_, _13557_, _13727_);
  nor _22069_ (_13729_, _13568_, _13475_);
  nor _22070_ (_13730_, _13562_, _13555_);
  and _22071_ (_13731_, _13730_, _13729_);
  and _22072_ (_13732_, _13731_, _13728_);
  and _22073_ (_13733_, _13732_, _13725_);
  nand _22074_ (_13734_, _13733_, _13724_);
  nand _22075_ (_13735_, _13734_, _13701_);
  nand _22076_ (_13736_, _13735_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  nand _22077_ (_13737_, _13736_, _13704_);
  or _22078_ (_13738_, _13737_, _13703_);
  and _22079_ (_11841_, _13738_, _13479_);
  or _22080_ (_13739_, _06948_, _06063_);
  or _22081_ (_13740_, _09508_, _13739_);
  not _22082_ (_13741_, _09503_);
  or _22083_ (_13742_, _13741_, _06309_);
  and _22084_ (_13743_, _13742_, _06068_);
  or _22085_ (_13744_, _13743_, _13740_);
  and _22086_ (_13745_, _13744_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  and _22087_ (_13746_, _12264_, _06307_);
  or _22088_ (_13747_, _13746_, _13745_);
  and _22089_ (_11869_, _13747_, _05552_);
  and _22090_ (_13748_, _09505_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  nor _22091_ (_13749_, _09505_, _06560_);
  or _22092_ (_13750_, _13749_, _13748_);
  or _22093_ (_13751_, _13750_, _06955_);
  or _22094_ (_13752_, _06068_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  and _22095_ (_13753_, _13752_, _05552_);
  and _22096_ (_11880_, _13753_, _13751_);
  and _22097_ (_13754_, _07951_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  and _22098_ (_13755_, _07946_, _07949_);
  or _22099_ (_13756_, _13755_, _13754_);
  and _22100_ (_11882_, _13756_, _05552_);
  nand _22101_ (_13757_, _13735_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  nand _22102_ (_13758_, _13488_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  nand _22103_ (_13759_, _13494_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and _22104_ (_13760_, _13759_, _13758_);
  nand _22105_ (_13762_, _13502_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  nand _22106_ (_13763_, _13499_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and _22107_ (_13764_, _13763_, _13762_);
  and _22108_ (_13765_, _13764_, _13760_);
  nand _22109_ (_13766_, _13507_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  nand _22110_ (_13767_, _13511_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and _22111_ (_13768_, _13767_, _13766_);
  nand _22112_ (_13769_, _13516_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  nand _22113_ (_13770_, _13521_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and _22114_ (_13771_, _13770_, _13769_);
  and _22115_ (_13772_, _13771_, _13768_);
  and _22116_ (_13773_, _13772_, _13765_);
  nand _22117_ (_13774_, _13531_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  not _22118_ (_13775_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  or _22119_ (_13776_, _13528_, _13775_);
  and _22120_ (_13777_, _13776_, _13774_);
  nand _22121_ (_13778_, _13536_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nand _22122_ (_13779_, _13534_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and _22123_ (_13780_, _13779_, _13778_);
  and _22124_ (_13781_, _13780_, _13777_);
  nand _22125_ (_13782_, _13541_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  nand _22126_ (_13783_, _13544_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and _22127_ (_13784_, _13783_, _13782_);
  nand _22128_ (_13785_, _13547_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nand _22129_ (_13786_, _13549_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  and _22130_ (_13787_, _13786_, _13785_);
  and _22131_ (_13788_, _13787_, _13784_);
  and _22132_ (_13789_, _13788_, _13781_);
  and _22133_ (_13790_, _13789_, _13773_);
  nand _22134_ (_13791_, _13555_, _11503_);
  nand _22135_ (_13792_, _13562_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and _22136_ (_13793_, _13792_, _13791_);
  nand _22137_ (_13794_, _13475_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  nand _22138_ (_13795_, _13568_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  and _22139_ (_13796_, _13795_, _13794_);
  and _22140_ (_13797_, _13796_, _13793_);
  nor _22141_ (_13798_, _13592_, p2_in[4]);
  not _22142_ (_13799_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and _22143_ (_13800_, _13592_, _13799_);
  nor _22144_ (_13801_, _13800_, _13798_);
  nand _22145_ (_13802_, _13801_, _13611_);
  nor _22146_ (_13803_, _13592_, p3_in[4]);
  not _22147_ (_13804_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and _22148_ (_13805_, _13592_, _13804_);
  nor _22149_ (_13806_, _13805_, _13803_);
  nand _22150_ (_13807_, _13806_, _13605_);
  and _22151_ (_13808_, _13807_, _13802_);
  nor _22152_ (_13809_, _13592_, p0_in[4]);
  not _22153_ (_13810_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and _22154_ (_13811_, _13592_, _13810_);
  nor _22155_ (_13812_, _13811_, _13809_);
  nand _22156_ (_13813_, _13812_, _13574_);
  nor _22157_ (_13814_, _13592_, p1_in[4]);
  not _22158_ (_13815_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and _22159_ (_13816_, _13592_, _13815_);
  nor _22160_ (_13817_, _13816_, _13814_);
  nand _22161_ (_13818_, _13817_, _13598_);
  and _22162_ (_13819_, _13818_, _13813_);
  and _22163_ (_13820_, _13819_, _13808_);
  and _22164_ (_13821_, _13820_, _13797_);
  nand _22165_ (_13822_, _13681_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nand _22166_ (_13823_, _13622_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and _22167_ (_13824_, _13823_, _13822_);
  and _22168_ (_13825_, _13824_, _13821_);
  and _22169_ (_13826_, _13825_, _13790_);
  or _22170_ (_13827_, _13826_, _13702_);
  and _22171_ (_13828_, _13827_, _13757_);
  nand _22172_ (_13829_, _13828_, _13704_);
  or _22173_ (_13830_, _13704_, _12189_);
  and _22174_ (_13831_, _13830_, _05552_);
  and _22175_ (_11885_, _13831_, _13829_);
  nand _22176_ (_13832_, _13735_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  nand _22177_ (_13833_, _13494_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  nand _22178_ (_13834_, _13488_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and _22179_ (_13835_, _13834_, _13833_);
  nand _22180_ (_13836_, _13499_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  nand _22181_ (_13837_, _13502_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and _22182_ (_13838_, _13837_, _13836_);
  and _22183_ (_13839_, _13838_, _13835_);
  nand _22184_ (_13840_, _13507_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  nand _22185_ (_13841_, _13511_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and _22186_ (_13842_, _13841_, _13840_);
  nand _22187_ (_13843_, _13516_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  nand _22188_ (_13844_, _13521_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and _22189_ (_13845_, _13844_, _13843_);
  and _22190_ (_13846_, _13845_, _13842_);
  and _22191_ (_13847_, _13846_, _13839_);
  nand _22192_ (_13848_, _13531_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nand _22193_ (_13849_, _13713_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  and _22194_ (_13850_, _13849_, _13848_);
  nand _22195_ (_13851_, _13534_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  nand _22196_ (_13852_, _13536_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and _22197_ (_00002_, _13852_, _13851_);
  and _22198_ (_00003_, _00002_, _13850_);
  nand _22199_ (_00004_, _13541_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  nand _22200_ (_00005_, _13544_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  and _22201_ (_00006_, _00005_, _00004_);
  nand _22202_ (_00007_, _13547_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  nand _22203_ (_00008_, _13549_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  and _22204_ (_00009_, _00008_, _00007_);
  and _22205_ (_00010_, _00009_, _00006_);
  and _22206_ (_00011_, _00010_, _00003_);
  and _22207_ (_00012_, _00011_, _13847_);
  nand _22208_ (_00013_, _13475_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  nand _22209_ (_00014_, _13568_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  and _22210_ (_00015_, _00014_, _00013_);
  nand _22211_ (_00016_, _13555_, _11251_);
  nand _22212_ (_00017_, _13562_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and _22213_ (_00018_, _00017_, _00016_);
  and _22214_ (_00019_, _00018_, _00015_);
  nor _22215_ (_00020_, _13592_, p0_in[3]);
  not _22216_ (_00021_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and _22217_ (_00022_, _13592_, _00021_);
  nor _22218_ (_00023_, _00022_, _00020_);
  nand _22219_ (_00024_, _00023_, _13574_);
  nor _22220_ (_00026_, _13592_, p1_in[3]);
  not _22221_ (_00027_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and _22222_ (_00028_, _13592_, _00027_);
  nor _22223_ (_00029_, _00028_, _00026_);
  nand _22224_ (_00030_, _00029_, _13598_);
  and _22225_ (_00031_, _00030_, _00024_);
  nor _22226_ (_00032_, _13592_, p3_in[3]);
  not _22227_ (_00033_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and _22228_ (_00034_, _13592_, _00033_);
  nor _22229_ (_00035_, _00034_, _00032_);
  nand _22230_ (_00036_, _00035_, _13605_);
  nor _22231_ (_00037_, _13592_, p2_in[3]);
  not _22232_ (_00038_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and _22233_ (_00039_, _13592_, _00038_);
  nor _22234_ (_00040_, _00039_, _00037_);
  nand _22235_ (_00041_, _00040_, _13611_);
  and _22236_ (_00042_, _00041_, _00036_);
  and _22237_ (_00043_, _00042_, _00031_);
  and _22238_ (_00044_, _00043_, _00019_);
  nand _22239_ (_00045_, _13681_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nand _22240_ (_00046_, _13622_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and _22241_ (_00047_, _00046_, _00045_);
  and _22242_ (_00048_, _00047_, _00044_);
  and _22243_ (_00049_, _00048_, _00012_);
  or _22244_ (_00050_, _00049_, _13702_);
  and _22245_ (_00051_, _00050_, _13832_);
  nand _22246_ (_00052_, _00051_, _13704_);
  or _22247_ (_00053_, _13704_, _07483_);
  and _22248_ (_00054_, _00053_, _05552_);
  and _22249_ (_11888_, _00054_, _00052_);
  and _22250_ (_00055_, _13499_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and _22251_ (_00056_, _13502_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  or _22252_ (_00057_, _00056_, _00055_);
  and _22253_ (_00058_, _13494_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and _22254_ (_00059_, _13488_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or _22255_ (_00061_, _00059_, _00058_);
  or _22256_ (_00062_, _00061_, _00057_);
  and _22257_ (_00063_, _13507_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and _22258_ (_00064_, _13511_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  or _22259_ (_00065_, _00064_, _00063_);
  and _22260_ (_00066_, _13516_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and _22261_ (_00067_, _13521_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or _22262_ (_00068_, _00067_, _00066_);
  or _22263_ (_00069_, _00068_, _00065_);
  or _22264_ (_00070_, _00069_, _00062_);
  and _22265_ (_00072_, _13531_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  not _22266_ (_00073_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  nor _22267_ (_00074_, _13528_, _00073_);
  or _22268_ (_00075_, _00074_, _00072_);
  and _22269_ (_00077_, _13534_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  and _22270_ (_00078_, _13536_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  or _22271_ (_00079_, _00078_, _00077_);
  or _22272_ (_00080_, _00079_, _00075_);
  and _22273_ (_00081_, _13541_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  and _22274_ (_00082_, _13544_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  or _22275_ (_00083_, _00082_, _00081_);
  and _22276_ (_00084_, _13547_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _22277_ (_00086_, _13549_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  or _22278_ (_00087_, _00086_, _00084_);
  or _22279_ (_00088_, _00087_, _00083_);
  or _22280_ (_00089_, _00088_, _00080_);
  or _22281_ (_00090_, _00089_, _00070_);
  and _22282_ (_00091_, _13475_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and _22283_ (_00092_, _13568_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or _22284_ (_00093_, _00092_, _00091_);
  and _22285_ (_00094_, _13555_, _11759_);
  and _22286_ (_00095_, _13562_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or _22287_ (_00096_, _00095_, _00094_);
  or _22288_ (_00097_, _00096_, _00093_);
  or _22289_ (_00098_, _13592_, p3_in[2]);
  not _22290_ (_00099_, _13592_);
  or _22291_ (_00100_, _00099_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and _22292_ (_00101_, _00100_, _00098_);
  and _22293_ (_00102_, _00101_, _13605_);
  or _22294_ (_00103_, _13592_, p2_in[2]);
  or _22295_ (_00104_, _00099_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and _22296_ (_00105_, _00104_, _00103_);
  and _22297_ (_00106_, _00105_, _13611_);
  or _22298_ (_00107_, _00106_, _00102_);
  or _22299_ (_00108_, _13592_, p1_in[2]);
  or _22300_ (_00109_, _00099_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and _22301_ (_00110_, _00109_, _00108_);
  and _22302_ (_00111_, _00110_, _13598_);
  or _22303_ (_00112_, _13592_, p0_in[2]);
  or _22304_ (_00113_, _00099_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and _22305_ (_00114_, _00113_, _00112_);
  and _22306_ (_00115_, _00114_, _13574_);
  or _22307_ (_00116_, _00115_, _00111_);
  or _22308_ (_00117_, _00116_, _00107_);
  or _22309_ (_00118_, _00117_, _00097_);
  and _22310_ (_00119_, _13622_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  and _22311_ (_00120_, _13681_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or _22312_ (_00121_, _00120_, _00119_);
  or _22313_ (_00123_, _00121_, _00118_);
  or _22314_ (_00124_, _00123_, _00090_);
  and _22315_ (_00125_, _00124_, _13701_);
  and _22316_ (_00126_, _13735_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  or _22317_ (_00127_, _00126_, _00125_);
  or _22318_ (_00128_, _00127_, _13476_);
  or _22319_ (_00129_, _13704_, _08144_);
  and _22320_ (_00130_, _00129_, _05552_);
  and _22321_ (_11894_, _00130_, _00128_);
  and _22322_ (_00131_, _13502_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and _22323_ (_00132_, _13499_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  or _22324_ (_00133_, _00132_, _00131_);
  and _22325_ (_00134_, _13494_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and _22326_ (_00135_, _13488_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or _22327_ (_00136_, _00135_, _00134_);
  or _22328_ (_00137_, _00136_, _00133_);
  and _22329_ (_00138_, _13507_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  and _22330_ (_00139_, _13511_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  or _22331_ (_00140_, _00139_, _00138_);
  and _22332_ (_00141_, _13516_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and _22333_ (_00142_, _13521_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  or _22334_ (_00143_, _00142_, _00141_);
  or _22335_ (_00144_, _00143_, _00140_);
  or _22336_ (_00145_, _00144_, _00137_);
  not _22337_ (_00146_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  nor _22338_ (_00147_, _13528_, _00146_);
  and _22339_ (_00148_, _13531_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  or _22340_ (_00149_, _00148_, _00147_);
  and _22341_ (_00150_, _13536_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and _22342_ (_00151_, _13534_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  or _22343_ (_00152_, _00151_, _00150_);
  or _22344_ (_00154_, _00152_, _00149_);
  and _22345_ (_00155_, _13544_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  and _22346_ (_00156_, _13541_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  or _22347_ (_00157_, _00156_, _00155_);
  and _22348_ (_00158_, _13547_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and _22349_ (_00160_, _13549_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  or _22350_ (_00161_, _00160_, _00158_);
  or _22351_ (_00162_, _00161_, _00157_);
  or _22352_ (_00163_, _00162_, _00154_);
  or _22353_ (_00164_, _00163_, _00145_);
  and _22354_ (_00165_, _13475_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and _22355_ (_00166_, _13568_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or _22356_ (_00167_, _00166_, _00165_);
  and _22357_ (_00168_, _13555_, _11627_);
  and _22358_ (_00169_, _13562_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  or _22359_ (_00170_, _00169_, _00168_);
  or _22360_ (_00171_, _00170_, _00167_);
  or _22361_ (_00172_, _13592_, p2_in[1]);
  not _22362_ (_00173_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  nand _22363_ (_00174_, _13592_, _00173_);
  and _22364_ (_00175_, _00174_, _00172_);
  and _22365_ (_00176_, _00175_, _13611_);
  or _22366_ (_00177_, _13592_, p3_in[1]);
  or _22367_ (_00178_, _00099_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and _22368_ (_00179_, _00178_, _00177_);
  and _22369_ (_00180_, _00179_, _13605_);
  or _22370_ (_00181_, _00180_, _00176_);
  or _22371_ (_00182_, _13592_, p0_in[1]);
  or _22372_ (_00183_, _00099_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and _22373_ (_00184_, _00183_, _00182_);
  and _22374_ (_00185_, _00184_, _13574_);
  or _22375_ (_00186_, _13592_, p1_in[1]);
  or _22376_ (_00187_, _00099_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and _22377_ (_00188_, _00187_, _00186_);
  and _22378_ (_00189_, _00188_, _13598_);
  or _22379_ (_00190_, _00189_, _00185_);
  or _22380_ (_00191_, _00190_, _00181_);
  or _22381_ (_00192_, _00191_, _00171_);
  and _22382_ (_00193_, _13622_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and _22383_ (_00194_, _13681_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or _22384_ (_00195_, _00194_, _00193_);
  or _22385_ (_00196_, _00195_, _00192_);
  or _22386_ (_00197_, _00196_, _00164_);
  and _22387_ (_00198_, _00197_, _13701_);
  and _22388_ (_00199_, _13735_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  or _22389_ (_00200_, _00199_, _00198_);
  or _22390_ (_00202_, _00200_, _13476_);
  or _22391_ (_00203_, _13704_, _08102_);
  and _22392_ (_00204_, _00203_, _05552_);
  and _22393_ (_11897_, _00204_, _00202_);
  nor _22394_ (_11963_, _05646_, rst);
  or _22395_ (_00207_, _05550_, \oc8051_top_1.oc8051_rom1.data_o [6]);
  nand _22396_ (_00208_, _05550_, _05786_);
  and _22397_ (_00209_, _00208_, _05552_);
  and _22398_ (_11974_, _00209_, _00207_);
  and _22399_ (_00210_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and _22400_ (_00211_, _12140_, \oc8051_top_1.oc8051_rom1.data_o [23]);
  or _22401_ (_00212_, _00211_, _00210_);
  and _22402_ (_11981_, _00212_, _05552_);
  and _22403_ (_00213_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and _22404_ (_00214_, _12140_, \oc8051_top_1.oc8051_rom1.data_o [16]);
  or _22405_ (_00215_, _00214_, _00213_);
  and _22406_ (_11984_, _00215_, _05552_);
  or _22407_ (_00216_, _05550_, \oc8051_top_1.oc8051_rom1.data_o [28]);
  nand _22408_ (_00217_, _05550_, _11052_);
  and _22409_ (_00218_, _00217_, _05552_);
  and _22410_ (_11992_, _00218_, _00216_);
  nor _22411_ (_12003_, _11646_, rst);
  and _22412_ (_00220_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and _22413_ (_00221_, _12140_, \oc8051_top_1.oc8051_rom1.data_o [25]);
  or _22414_ (_00222_, _00221_, _00220_);
  and _22415_ (_12011_, _00222_, _05552_);
  nand _22416_ (_00223_, _10860_, _06527_);
  nor _22417_ (_00224_, _00223_, _05971_);
  and _22418_ (_00225_, _00224_, _06910_);
  or _22419_ (_00226_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  or _22420_ (_00227_, _00226_, _00225_);
  nand _22421_ (_00228_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  nand _22422_ (_00229_, _00228_, _00225_);
  or _22423_ (_00230_, _00229_, _08926_);
  and _22424_ (_00231_, _00230_, _00227_);
  and _22425_ (_00232_, _08990_, _06927_);
  or _22426_ (_00233_, _00232_, _00231_);
  nand _22427_ (_00234_, _00232_, _07975_);
  and _22428_ (_00236_, _00234_, _05552_);
  and _22429_ (_12023_, _00236_, _00233_);
  or _22430_ (_00237_, _07668_, _07255_);
  or _22431_ (_00238_, _07670_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and _22432_ (_00239_, _00238_, _05552_);
  and _22433_ (_12026_, _00239_, _00237_);
  nor _22434_ (_12033_, _11872_, rst);
  and _22435_ (_00240_, _06771_, _06525_);
  and _22436_ (_00241_, _00240_, _07443_);
  nand _22437_ (_00242_, _00241_, _08041_);
  or _22438_ (_00243_, _00241_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  and _22439_ (_00244_, _00243_, _05552_);
  and _22440_ (_12042_, _00244_, _00242_);
  and _22441_ (_00245_, _08989_, _06056_);
  and _22442_ (_00246_, _00245_, _06927_);
  and _22443_ (_00248_, _00246_, _05560_);
  and _22444_ (_00249_, _00248_, _11490_);
  and _22445_ (_00250_, \oc8051_top_1.oc8051_sfr1.pres_ow , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  and _22446_ (_00252_, _00250_, _05560_);
  and _22447_ (_00253_, _05573_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr );
  and _22448_ (_00254_, _00253_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  nor _22449_ (_00255_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  nor _22450_ (_00256_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  and _22451_ (_00257_, _00256_, _00255_);
  and _22452_ (_00258_, _00257_, _00254_);
  nor _22453_ (_00259_, _00258_, _00252_);
  not _22454_ (_00260_, _00259_);
  and _22455_ (_00261_, _00260_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  and _22456_ (_00262_, _00259_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  nor _22457_ (_00263_, _00262_, _00261_);
  and _22458_ (_00264_, _06524_, _06308_);
  and _22459_ (_00265_, _00264_, _06927_);
  nor _22460_ (_00266_, _00265_, _00263_);
  and _22461_ (_00267_, _00246_, _05573_);
  not _22462_ (_00268_, _00267_);
  nor _22463_ (_00270_, _00268_, _06560_);
  or _22464_ (_00272_, _00270_, _00266_);
  or _22465_ (_00273_, _00272_, _00249_);
  and _22466_ (_12049_, _00273_, _05552_);
  and _22467_ (_00275_, _00248_, _11234_);
  and _22468_ (_00276_, _00260_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  and _22469_ (_00277_, _00259_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  nor _22470_ (_00278_, _00277_, _00276_);
  nor _22471_ (_00279_, _00278_, _00265_);
  and _22472_ (_00280_, _00267_, _11238_);
  or _22473_ (_00281_, _00280_, _00279_);
  or _22474_ (_00282_, _00281_, _00275_);
  and _22475_ (_12055_, _00282_, _05552_);
  nor _22476_ (_00283_, _11802_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor _22477_ (_00284_, _00283_, _11803_);
  and _22478_ (_00285_, _00284_, _11792_);
  and _22479_ (_00286_, _11811_, _07483_);
  not _22480_ (_00287_, _11784_);
  nor _22481_ (_00288_, _00287_, _07515_);
  and _22482_ (_00289_, _11780_, _11275_);
  and _22483_ (_00290_, _11817_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  or _22484_ (_00292_, _00290_, _00289_);
  or _22485_ (_00293_, _00292_, _00288_);
  or _22486_ (_00294_, _00293_, _00286_);
  nor _22487_ (_00295_, _00294_, _00285_);
  nand _22488_ (_00296_, _00295_, _11774_);
  and _22489_ (_00297_, _12025_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  or _22490_ (_00298_, _00297_, _12155_);
  or _22491_ (_00299_, _12034_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _22492_ (_00300_, _00299_, _12035_);
  or _22493_ (_00301_, _00300_, _11828_);
  and _22494_ (_00302_, _00301_, _12054_);
  and _22495_ (_00303_, _00302_, _00298_);
  or _22496_ (_00304_, _00303_, _00296_);
  nor _22497_ (_00305_, _12066_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor _22498_ (_00306_, _00305_, _12068_);
  or _22499_ (_00307_, _00306_, _11774_);
  and _22500_ (_00308_, _00307_, _05552_);
  and _22501_ (_12058_, _00308_, _00304_);
  nor _22502_ (_00309_, _12017_, _11854_);
  nor _22503_ (_00310_, _00309_, _12018_);
  and _22504_ (_00311_, _00310_, _12054_);
  or _22505_ (_00312_, _11817_, _11784_);
  and _22506_ (_00313_, _00312_, _07574_);
  nor _22507_ (_00314_, _11102_, _09047_);
  not _22508_ (_00315_, _11848_);
  and _22509_ (_00316_, _00315_, _11780_);
  and _22510_ (_00317_, _11792_, _11391_);
  or _22511_ (_00318_, _00317_, _00316_);
  or _22512_ (_00319_, _00318_, _00314_);
  or _22513_ (_00320_, _00319_, _00313_);
  or _22514_ (_00321_, _00320_, _00311_);
  and _22515_ (_00322_, _00321_, _11774_);
  nor _22516_ (_00323_, _12060_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and _22517_ (_00324_, _12060_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or _22518_ (_00325_, _00324_, _00323_);
  nor _22519_ (_00326_, _00325_, _11774_);
  or _22520_ (_00327_, _00326_, _00322_);
  and _22521_ (_12065_, _00327_, _05552_);
  and _22522_ (_00329_, _00254_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  and _22523_ (_00330_, _00329_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  nor _22524_ (_00332_, _00330_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  and _22525_ (_00333_, _00330_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  nor _22526_ (_00334_, _00333_, _00332_);
  nor _22527_ (_00335_, _00246_, rst);
  and _22528_ (_12067_, _00335_, _00334_);
  and _22529_ (_00337_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  nor _22530_ (_00338_, _05550_, _05786_);
  or _22531_ (_00339_, _00338_, _00337_);
  and _22532_ (_12070_, _00339_, _05552_);
  nor _22533_ (_00340_, _09150_, _09094_);
  nor _22534_ (_00341_, _00340_, _09151_);
  or _22535_ (_00343_, _00341_, _09039_);
  or _22536_ (_00344_, _09038_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and _22537_ (_00345_, _00344_, _07933_);
  and _22538_ (_00346_, _00345_, _00343_);
  and _22539_ (_00347_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and _22540_ (_00348_, _00347_, _05552_);
  or _22541_ (_12078_, _00348_, _00346_);
  and _22542_ (_00349_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  nor _22543_ (_00350_, _05550_, _11739_);
  or _22544_ (_00351_, _00350_, _00349_);
  and _22545_ (_12079_, _00351_, _05552_);
  nor _22546_ (_12084_, \oc8051_top_1.oc8051_sfr1.prescaler [0], rst);
  nor _22547_ (_00352_, _09137_, _09116_);
  nor _22548_ (_00353_, _00352_, _09139_);
  or _22549_ (_00354_, _00353_, _09039_);
  or _22550_ (_00355_, _09038_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and _22551_ (_00356_, _00355_, _05605_);
  and _22552_ (_00357_, _00356_, _00354_);
  and _22553_ (_00358_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3], \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _22554_ (_00359_, _00358_, _00357_);
  and _22555_ (_12087_, _00359_, _05552_);
  and _22556_ (_00360_, _09123_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  or _22557_ (_00361_, _07919_, _05622_);
  nand _22558_ (_00362_, _07919_, _05622_);
  and _22559_ (_00363_, _00362_, _00361_);
  nand _22560_ (_00364_, _00363_, _00360_);
  or _22561_ (_00365_, _00363_, _00360_);
  and _22562_ (_00366_, _00365_, _00364_);
  or _22563_ (_00367_, _00366_, _05548_);
  or _22564_ (_00368_, _05547_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and _22565_ (_00369_, _00368_, _07933_);
  and _22566_ (_12102_, _00369_, _00367_);
  and _22567_ (_00370_, _05916_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  or _22568_ (_00371_, _00370_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and _22569_ (_12105_, _00371_, _05552_);
  nor _22570_ (_12110_, _11943_, rst);
  not _22571_ (_00372_, \oc8051_top_1.oc8051_sfr1.prescaler [2]);
  and _22572_ (_00373_, \oc8051_top_1.oc8051_sfr1.prescaler [1], \oc8051_top_1.oc8051_sfr1.prescaler [0]);
  and _22573_ (_00374_, _00373_, _00372_);
  and _22574_ (_00375_, _00374_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  nor _22575_ (_00376_, _00373_, _00372_);
  or _22576_ (_00377_, _00376_, _00374_);
  nand _22577_ (_00378_, _00377_, _05552_);
  nor _22578_ (_12113_, _00378_, _00375_);
  or _22579_ (_00379_, \oc8051_top_1.oc8051_sfr1.prescaler [1], \oc8051_top_1.oc8051_sfr1.prescaler [0]);
  nor _22580_ (_00380_, _00373_, rst);
  and _22581_ (_12115_, _00380_, _00379_);
  and _22582_ (_00381_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], _07768_);
  and _22583_ (_00382_, \oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or _22584_ (_00383_, _00382_, _00381_);
  and _22585_ (_12135_, _00383_, _05552_);
  nor _22586_ (_00384_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and _22587_ (_00385_, _00384_, _05573_);
  and _22588_ (_00386_, _00385_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  not _22589_ (_00387_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  nor _22590_ (_00388_, _00385_, _00387_);
  or _22591_ (_00389_, _00388_, _00386_);
  or _22592_ (_00390_, _00389_, _00225_);
  or _22593_ (_00391_, _08013_, _00387_);
  nand _22594_ (_00392_, _00391_, _00225_);
  or _22595_ (_00393_, _00392_, _08015_);
  and _22596_ (_00394_, _00393_, _00390_);
  or _22597_ (_00396_, _00394_, _00232_);
  nand _22598_ (_00397_, _00232_, _08041_);
  and _22599_ (_00398_, _00397_, _05552_);
  and _22600_ (_12151_, _00398_, _00396_);
  nand _22601_ (_00399_, _00241_, _06560_);
  or _22602_ (_00400_, _00241_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  and _22603_ (_00401_, _00400_, _05552_);
  and _22604_ (_12158_, _00401_, _00399_);
  and _22605_ (_00402_, _00248_, _06307_);
  and _22606_ (_00403_, _00260_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  and _22607_ (_00404_, _00259_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  nor _22608_ (_00405_, _00404_, _00403_);
  nor _22609_ (_00406_, _00405_, _00265_);
  nor _22610_ (_00407_, _00268_, _07388_);
  or _22611_ (_00408_, _00407_, _00406_);
  or _22612_ (_00409_, _00408_, _00402_);
  and _22613_ (_12191_, _00409_, _05552_);
  nor _22614_ (_00410_, _12059_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor _22615_ (_00411_, _00410_, _12060_);
  or _22616_ (_00412_, _00411_, _11774_);
  and _22617_ (_00413_, _00412_, _05552_);
  and _22618_ (_00414_, _00312_, _07635_);
  nor _22619_ (_00415_, _11102_, _09106_);
  not _22620_ (_00416_, _11872_);
  and _22621_ (_00417_, _00416_, _11780_);
  and _22622_ (_00418_, _11792_, _11449_);
  or _22623_ (_00419_, _00418_, _00417_);
  or _22624_ (_00420_, _00419_, _00415_);
  or _22625_ (_00421_, _00420_, _00414_);
  or _22626_ (_00422_, _11876_, _11877_);
  and _22627_ (_00423_, _00422_, _12015_);
  nor _22628_ (_00424_, _00422_, _12015_);
  or _22629_ (_00425_, _00424_, _00423_);
  nand _22630_ (_00426_, _00425_, _12054_);
  nand _22631_ (_00427_, _00426_, _11774_);
  or _22632_ (_00428_, _00427_, _00421_);
  and _22633_ (_12275_, _00428_, _00413_);
  nand _22634_ (_00429_, _08386_, _06949_);
  or _22635_ (_00430_, _06949_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  and _22636_ (_00431_, _00430_, _05552_);
  and _22637_ (_12281_, _00431_, _00429_);
  and _22638_ (_00432_, _00312_, _12189_);
  and _22639_ (_00433_, _11792_, _11470_);
  not _22640_ (_00434_, _11900_);
  and _22641_ (_00435_, _00434_, _11780_);
  or _22642_ (_00436_, _00435_, _00433_);
  or _22643_ (_00437_, _12013_, _12010_);
  and _22644_ (_00438_, _12054_, _12014_);
  and _22645_ (_00439_, _00438_, _00437_);
  or _22646_ (_00440_, _00439_, _00436_);
  or _22647_ (_00441_, _00440_, _00432_);
  or _22648_ (_00442_, _11102_, _09107_);
  nand _22649_ (_00443_, _00442_, _11774_);
  or _22650_ (_00444_, _00443_, _00441_);
  nor _22651_ (_00445_, _08238_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor _22652_ (_00446_, _00445_, _12059_);
  or _22653_ (_00447_, _00446_, _11774_);
  and _22654_ (_00448_, _00447_, _05552_);
  and _22655_ (_12286_, _00448_, _00444_);
  and _22656_ (_00449_, _00225_, _10632_);
  nand _22657_ (_00450_, _00449_, _06763_);
  not _22658_ (_00451_, _00232_);
  or _22659_ (_00452_, _00449_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  and _22660_ (_00453_, _00452_, _00451_);
  and _22661_ (_00454_, _00453_, _00450_);
  nor _22662_ (_00455_, _00451_, _06560_);
  or _22663_ (_00456_, _00455_, _00454_);
  and _22664_ (_12294_, _00456_, _05552_);
  nand _22665_ (_00457_, _00241_, _07388_);
  or _22666_ (_00458_, _00241_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  and _22667_ (_00459_, _00458_, _05552_);
  and _22668_ (_12323_, _00459_, _00457_);
  and _22669_ (_00460_, _00248_, _11367_);
  and _22670_ (_00461_, _00260_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  and _22671_ (_00462_, _00259_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  nor _22672_ (_00463_, _00462_, _00461_);
  nor _22673_ (_00464_, _00463_, _00265_);
  nor _22674_ (_00465_, _00268_, _06306_);
  or _22675_ (_00466_, _00465_, _00464_);
  or _22676_ (_00467_, _00466_, _00460_);
  and _22677_ (_12326_, _00467_, _05552_);
  or _22678_ (_00468_, _11774_, _08240_);
  and _22679_ (_00469_, _00468_, _05552_);
  and _22680_ (_00470_, _00312_, _07483_);
  nor _22681_ (_00471_, _11102_, _09048_);
  not _22682_ (_00472_, _11921_);
  and _22683_ (_00473_, _00472_, _11780_);
  and _22684_ (_00474_, _11792_, _11275_);
  or _22685_ (_00476_, _00474_, _00473_);
  or _22686_ (_00477_, _00476_, _00471_);
  or _22687_ (_00478_, _00477_, _00470_);
  or _22688_ (_00479_, _11925_, _11926_);
  nor _22689_ (_00480_, _00479_, _12008_);
  and _22690_ (_00481_, _00479_, _12008_);
  or _22691_ (_00482_, _00481_, _00480_);
  nand _22692_ (_00483_, _00482_, _12054_);
  nand _22693_ (_00484_, _00483_, _11774_);
  or _22694_ (_00485_, _00484_, _00478_);
  and _22695_ (_12343_, _00485_, _00469_);
  or _22696_ (_00486_, _11774_, _08253_);
  and _22697_ (_00487_, _00486_, _05552_);
  and _22698_ (_00488_, _00312_, _08144_);
  nor _22699_ (_00489_, _11102_, _08236_);
  and _22700_ (_00490_, _11944_, _11780_);
  and _22701_ (_00491_, _11792_, _11747_);
  or _22702_ (_00492_, _00491_, _00490_);
  or _22703_ (_00493_, _00492_, _00489_);
  or _22704_ (_00494_, _00493_, _00488_);
  nor _22705_ (_00495_, _12006_, _12004_);
  nor _22706_ (_00496_, _00495_, _12007_);
  nand _22707_ (_00497_, _00496_, _12054_);
  nand _22708_ (_00498_, _00497_, _11774_);
  or _22709_ (_00499_, _00498_, _00494_);
  and _22710_ (_12346_, _00499_, _00487_);
  and _22711_ (_00500_, _08058_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  or _22712_ (_00501_, _00500_, _08062_);
  and _22713_ (_00502_, _00501_, _00225_);
  not _22714_ (_00503_, _00225_);
  or _22715_ (_00504_, _00503_, _08059_);
  and _22716_ (_00505_, _00504_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  or _22717_ (_00506_, _00505_, _00232_);
  or _22718_ (_00507_, _00506_, _00502_);
  nand _22719_ (_00508_, _00232_, _07388_);
  and _22720_ (_00509_, _00508_, _05552_);
  and _22721_ (_12356_, _00509_, _00507_);
  and _22722_ (_00510_, _00248_, _07439_);
  not _22723_ (_00511_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  nor _22724_ (_00512_, _00259_, _00511_);
  and _22725_ (_00513_, _00259_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  nor _22726_ (_00515_, _00513_, _00512_);
  nor _22727_ (_00516_, _00515_, _00265_);
  nor _22728_ (_00517_, _00268_, _08386_);
  or _22729_ (_00518_, _00517_, _00516_);
  or _22730_ (_00519_, _00518_, _00510_);
  and _22731_ (_12358_, _00519_, _05552_);
  and _22732_ (_00520_, _00312_, _08102_);
  and _22733_ (_00521_, _11811_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  and _22734_ (_00522_, _11968_, _11780_);
  and _22735_ (_00523_, _11792_, _11617_);
  or _22736_ (_00524_, _00523_, _00522_);
  or _22737_ (_00525_, _00524_, _00521_);
  nor _22738_ (_00526_, _12000_, _11998_);
  nor _22739_ (_00527_, _00526_, _12001_);
  and _22740_ (_00528_, _00527_, _12054_);
  or _22741_ (_00529_, _00528_, _00525_);
  nor _22742_ (_00531_, _00529_, _00520_);
  nand _22743_ (_00532_, _00531_, _11774_);
  or _22744_ (_00534_, _11774_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  and _22745_ (_00535_, _00534_, _05552_);
  and _22746_ (_12361_, _00535_, _00532_);
  and _22747_ (_00536_, _00312_, _07711_);
  or _22748_ (_00537_, _11997_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  not _22749_ (_00538_, _11998_);
  and _22750_ (_00539_, _12161_, _00538_);
  and _22751_ (_00540_, _00539_, _00537_);
  and _22752_ (_00541_, _11994_, _11780_);
  and _22753_ (_00542_, _11792_, _11691_);
  and _22754_ (_00543_, _11811_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  or _22755_ (_00544_, _00543_, _00542_);
  or _22756_ (_00545_, _00544_, _00541_);
  or _22757_ (_00546_, _00545_, _00540_);
  nor _22758_ (_00547_, _00546_, _00536_);
  nand _22759_ (_00548_, _00547_, _11774_);
  or _22760_ (_00550_, _11774_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and _22761_ (_00551_, _00550_, _05552_);
  and _22762_ (_12370_, _00551_, _00548_);
  and _22763_ (_00552_, _00225_, _08635_);
  nand _22764_ (_00553_, _00552_, _06763_);
  or _22765_ (_00554_, _00552_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  and _22766_ (_00555_, _00554_, _00451_);
  and _22767_ (_00556_, _00555_, _00553_);
  nor _22768_ (_00557_, _00451_, _06306_);
  or _22769_ (_00558_, _00557_, _00556_);
  and _22770_ (_12383_, _00558_, _05552_);
  and _22771_ (_00559_, _00312_, _07255_);
  and _22772_ (_00560_, _11792_, _11328_);
  not _22773_ (_00561_, _07758_);
  and _22774_ (_00562_, _11780_, _00561_);
  or _22775_ (_00563_, _00562_, _00560_);
  or _22776_ (_00564_, _11830_, _11829_);
  not _22777_ (_00565_, _00564_);
  nand _22778_ (_00566_, _00565_, _12019_);
  or _22779_ (_00567_, _00565_, _12019_);
  and _22780_ (_00568_, _00567_, _12054_);
  and _22781_ (_00569_, _00568_, _00566_);
  or _22782_ (_00570_, _00569_, _00563_);
  or _22783_ (_00571_, _00570_, _00559_);
  or _22784_ (_00572_, _11102_, _09046_);
  nand _22785_ (_00573_, _00572_, _11774_);
  or _22786_ (_00574_, _00573_, _00571_);
  nor _22787_ (_00575_, _00324_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and _22788_ (_00576_, _12061_, _12060_);
  nor _22789_ (_00577_, _00576_, _00575_);
  or _22790_ (_00578_, _00577_, _11774_);
  and _22791_ (_00579_, _00578_, _05552_);
  and _22792_ (_12440_, _00579_, _00574_);
  and _22793_ (_00580_, \oc8051_top_1.oc8051_memory_interface1.reti , \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  nor _22794_ (_00581_, _00580_, _08998_);
  and _22795_ (_00582_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _08998_);
  and _22796_ (_00583_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _22797_ (_00584_, _00583_, _00582_);
  and _22798_ (_00585_, _00584_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  nor _22799_ (_00586_, _00585_, _08996_);
  not _22800_ (_00587_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  nor _22801_ (_00588_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  nor _22802_ (_00589_, _00588_, _00587_);
  and _22803_ (_00590_, _00589_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  not _22804_ (_00591_, _00590_);
  not _22805_ (_00592_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  nor _22806_ (_00593_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  nor _22807_ (_00594_, _00593_, _00592_);
  nand _22808_ (_00595_, _00594_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and _22809_ (_00596_, _00595_, _00591_);
  and _22810_ (_00597_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and _22811_ (_00598_, _00597_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  not _22812_ (_00599_, _00598_);
  and _22813_ (_00600_, _00599_, _00596_);
  and _22814_ (_00601_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and _22815_ (_00602_, _00601_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  not _22816_ (_00603_, _00602_);
  and _22817_ (_00605_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and _22818_ (_00607_, _00605_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and _22819_ (_00608_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and _22820_ (_00609_, _00608_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  nor _22821_ (_00610_, _00609_, _00607_);
  and _22822_ (_00611_, _00610_, _00603_);
  and _22823_ (_00612_, _00611_, _00600_);
  nor _22824_ (_00613_, _00612_, _00586_);
  and _22825_ (_00614_, _08996_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  not _22826_ (_00615_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and _22827_ (_00616_, _00589_, _00615_);
  not _22828_ (_00617_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and _22829_ (_00618_, _00594_, _00617_);
  nor _22830_ (_00619_, _00618_, _00616_);
  not _22831_ (_00620_, _00619_);
  and _22832_ (_00621_, _00620_, _00614_);
  not _22833_ (_00622_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and _22834_ (_00623_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and _22835_ (_00624_, _00623_, _00622_);
  and _22836_ (_00625_, _00624_, _00614_);
  or _22837_ (_00626_, _00625_, _00621_);
  or _22838_ (_00627_, _00626_, _00613_);
  nand _22839_ (_00628_, _00613_, _00600_);
  and _22840_ (_00629_, _00628_, _00627_);
  and _22841_ (_00630_, _00629_, _00581_);
  or _22842_ (_00631_, _00630_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  not _22843_ (_00632_, _00581_);
  not _22844_ (_00633_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and _22845_ (_00634_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  and _22846_ (_00635_, _00634_, _00633_);
  not _22847_ (_00636_, _00635_);
  not _22848_ (_00637_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and _22849_ (_00638_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and _22850_ (_00639_, _00638_, _00637_);
  not _22851_ (_00640_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and _22852_ (_00641_, _00608_, _00640_);
  nor _22853_ (_00642_, _00641_, _00639_);
  and _22854_ (_00643_, _00642_, _00636_);
  not _22855_ (_00644_, _00624_);
  and _22856_ (_00645_, _00643_, _00644_);
  nand _22857_ (_00646_, _00645_, _00619_);
  nand _22858_ (_00647_, _00646_, _00614_);
  nor _22859_ (_00648_, _00647_, _00613_);
  not _22860_ (_00649_, _00648_);
  or _22861_ (_00650_, _00649_, _00643_);
  or _22862_ (_00651_, _00611_, _00586_);
  and _22863_ (_00652_, _00651_, _00650_);
  or _22864_ (_00653_, _00652_, _00632_);
  and _22865_ (_00654_, _00653_, _05552_);
  and _22866_ (_12455_, _00654_, _00631_);
  and _22867_ (_00655_, _12024_, _11828_);
  and _22868_ (_00656_, _12021_, _11796_);
  nor _22869_ (_00657_, _00656_, _11828_);
  or _22870_ (_00658_, _00657_, _00655_);
  nand _22871_ (_00659_, _00658_, _06219_);
  or _22872_ (_00660_, _00658_, _06219_);
  and _22873_ (_00661_, _00660_, _12161_);
  and _22874_ (_00662_, _00661_, _00659_);
  and _22875_ (_00663_, _11811_, _08144_);
  nor _22876_ (_00664_, _00287_, _08200_);
  and _22877_ (_00665_, _11780_, _11747_);
  and _22878_ (_00666_, _11792_, _05781_);
  and _22879_ (_00667_, _11817_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  or _22880_ (_00668_, _00667_, _00666_);
  or _22881_ (_00669_, _00668_, _00665_);
  nor _22882_ (_00670_, _00669_, _00664_);
  nand _22883_ (_00671_, _00670_, _11774_);
  or _22884_ (_00672_, _00671_, _00663_);
  or _22885_ (_00673_, _00672_, _00662_);
  and _22886_ (_00674_, _00324_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and _22887_ (_00675_, _00674_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and _22888_ (_00676_, _00675_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  nand _22889_ (_00677_, _00676_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  or _22890_ (_00678_, _00676_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and _22891_ (_00679_, _00678_, _00677_);
  or _22892_ (_00680_, _00679_, _11774_);
  and _22893_ (_00681_, _00680_, _05552_);
  and _22894_ (_12467_, _00681_, _00673_);
  and _22895_ (_00683_, _12021_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  or _22896_ (_00685_, _00683_, _11828_);
  nand _22897_ (_00686_, _12022_, _11828_);
  and _22898_ (_00687_, _00686_, _00685_);
  and _22899_ (_00688_, _00687_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  or _22900_ (_00689_, _00687_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nand _22901_ (_00690_, _00689_, _12161_);
  nor _22902_ (_00691_, _00690_, _00688_);
  and _22903_ (_00692_, _11811_, _08102_);
  nor _22904_ (_00693_, _00287_, _08173_);
  and _22905_ (_00694_, _11792_, _05803_);
  and _22906_ (_00695_, _11780_, _11617_);
  and _22907_ (_00696_, _11817_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  or _22908_ (_00697_, _00696_, _00695_);
  or _22909_ (_00698_, _00697_, _00694_);
  nor _22910_ (_00699_, _00698_, _00693_);
  nand _22911_ (_00700_, _00699_, _11774_);
  or _22912_ (_00701_, _00700_, _00692_);
  or _22913_ (_00702_, _00701_, _00691_);
  nor _22914_ (_00703_, _00675_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  nor _22915_ (_00704_, _00703_, _00676_);
  or _22916_ (_00705_, _00704_, _11774_);
  and _22917_ (_00706_, _00705_, _05552_);
  and _22918_ (_12520_, _00706_, _00702_);
  and _22919_ (_00707_, _11811_, _07711_);
  and _22920_ (_00708_, _11784_, _08228_);
  and _22921_ (_00709_, _11792_, _07781_);
  and _22922_ (_00710_, _11780_, _11691_);
  or _22923_ (_00711_, _00710_, _00709_);
  and _22924_ (_00712_, _11817_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  or _22925_ (_00713_, _00712_, _00711_);
  or _22926_ (_00714_, _00713_, _00708_);
  or _22927_ (_00715_, _00686_, _00683_);
  and _22928_ (_00716_, _12021_, _06192_);
  nor _22929_ (_00717_, _12021_, _06192_);
  or _22930_ (_00718_, _00717_, _00716_);
  or _22931_ (_00719_, _00718_, _11828_);
  and _22932_ (_00720_, _00719_, _00715_);
  and _22933_ (_00721_, _00720_, _12054_);
  or _22934_ (_00722_, _00721_, _00714_);
  or _22935_ (_00723_, _00722_, _00707_);
  or _22936_ (_00724_, _00723_, _13414_);
  nor _22937_ (_00725_, _00576_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor _22938_ (_00726_, _00725_, _00675_);
  or _22939_ (_00727_, _00726_, _11774_);
  and _22940_ (_00728_, _00727_, _05552_);
  and _22941_ (_12523_, _00728_, _00724_);
  nor _22942_ (_12598_, _11193_, rst);
  nor _22943_ (_00729_, _08041_, _07939_);
  and _22944_ (_00730_, _07939_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  or _22945_ (_00731_, _00730_, _00729_);
  and _22946_ (_12772_, _00731_, _05552_);
  and _22947_ (_12807_, _05552_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  and _22948_ (pc_log_change, _05608_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  and _22949_ (_00732_, _10861_, _08013_);
  or _22950_ (_00733_, _00732_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and _22951_ (_00734_, _00733_, _08992_);
  nand _22952_ (_00735_, _00732_, _06763_);
  and _22953_ (_00736_, _00735_, _00734_);
  nor _22954_ (_00737_, _08992_, _08041_);
  or _22955_ (_00738_, _00737_, _00736_);
  and _22956_ (_13106_, _00738_, _05552_);
  and _22957_ (_00739_, _10861_, _06060_);
  or _22958_ (_00740_, _00739_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and _22959_ (_00741_, _00740_, _08992_);
  nand _22960_ (_00742_, _00739_, _06763_);
  and _22961_ (_00743_, _00742_, _00741_);
  and _22962_ (_00744_, _08991_, _11238_);
  or _22963_ (_00745_, _00744_, _00743_);
  and _22964_ (_13109_, _00745_, _05552_);
  and _22965_ (_00746_, _10633_, _07443_);
  nand _22966_ (_00747_, _00746_, _06306_);
  and _22967_ (_00748_, _13775_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  not _22968_ (_00749_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and _22969_ (_00750_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _00749_);
  nor _22970_ (_00751_, _00750_, _00748_);
  and _22971_ (_00752_, _08989_, _08635_);
  and _22972_ (_00753_, _00752_, _07443_);
  nor _22973_ (_00754_, _00753_, _00751_);
  not _22974_ (_00755_, _00754_);
  and _22975_ (_00756_, _00755_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  not _22976_ (_00757_, _00751_);
  not _22977_ (_00758_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and _22978_ (_00759_, _00758_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  not _22979_ (_00760_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and _22980_ (_00761_, \oc8051_top_1.oc8051_sfr1.pres_ow , _00760_);
  not _22981_ (_00762_, t1_i);
  and _22982_ (_00763_, _00762_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and _22983_ (_00764_, _00763_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff );
  or _22984_ (_00765_, _00764_, _00761_);
  and _22985_ (_00766_, _00765_, _00759_);
  and _22986_ (_00767_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and _22987_ (_00768_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  and _22988_ (_00769_, _00768_, _00767_);
  and _22989_ (_00770_, _00769_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and _22990_ (_00772_, _00770_, _00766_);
  nor _22991_ (_00773_, _00772_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and _22992_ (_00774_, _00772_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  nor _22993_ (_00775_, _00774_, _00773_);
  and _22994_ (_00776_, _00775_, _00757_);
  and _22995_ (_00777_, _00774_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and _22996_ (_00778_, _00777_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and _22997_ (_00779_, _00778_, _00748_);
  and _22998_ (_00780_, _00779_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  nor _22999_ (_00781_, _00780_, _00776_);
  nor _23000_ (_00782_, _00781_, _00753_);
  or _23001_ (_00783_, _00782_, _00756_);
  or _23002_ (_00784_, _00783_, _00746_);
  and _23003_ (_00785_, _00784_, _05552_);
  and _23004_ (_13129_, _00785_, _00747_);
  nand _23005_ (_00786_, _00746_, _07388_);
  and _23006_ (_00787_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  nor _23007_ (_00788_, _00787_, _00753_);
  not _23008_ (_00789_, _00788_);
  and _23009_ (_00790_, _00789_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and _23010_ (_00791_, _00779_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  not _23011_ (_00792_, _00787_);
  and _23012_ (_00794_, _00769_, _00766_);
  and _23013_ (_00795_, _00794_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  nor _23014_ (_00796_, _00794_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  nor _23015_ (_00797_, _00796_, _00795_);
  and _23016_ (_00798_, _00797_, _00792_);
  nor _23017_ (_00799_, _00798_, _00791_);
  nor _23018_ (_00800_, _00799_, _00753_);
  or _23019_ (_00801_, _00800_, _00790_);
  or _23020_ (_00802_, _00801_, _00746_);
  and _23021_ (_00803_, _00802_, _05552_);
  and _23022_ (_13132_, _00803_, _00786_);
  nand _23023_ (_00804_, _00779_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nor _23024_ (_00805_, _00804_, _00753_);
  and _23025_ (_00806_, _00766_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and _23026_ (_00808_, _00806_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  and _23027_ (_00809_, _00808_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  nor _23028_ (_00810_, _00809_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nor _23029_ (_00811_, _00810_, _00794_);
  and _23030_ (_00812_, _00811_, _00788_);
  and _23031_ (_00813_, _00789_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  or _23032_ (_00814_, _00813_, _00812_);
  or _23033_ (_00816_, _00814_, _00805_);
  or _23034_ (_00817_, _00816_, _00746_);
  nand _23035_ (_00818_, _00746_, _06560_);
  and _23036_ (_00819_, _00818_, _05552_);
  and _23037_ (_13135_, _00819_, _00817_);
  nand _23038_ (_00820_, _00746_, _08386_);
  nand _23039_ (_00821_, _00779_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nor _23040_ (_00822_, _00821_, _00753_);
  and _23041_ (_00823_, _00755_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and _23042_ (_00824_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and _23043_ (_00825_, _00824_, _00795_);
  nor _23044_ (_00826_, _00774_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nor _23045_ (_00827_, _00826_, _00825_);
  and _23046_ (_00828_, _00827_, _00754_);
  or _23047_ (_00829_, _00828_, _00823_);
  or _23048_ (_00830_, _00829_, _00822_);
  or _23049_ (_00831_, _00830_, _00746_);
  and _23050_ (_00832_, _00831_, _05552_);
  and _23051_ (_13139_, _00832_, _00820_);
  nor _23052_ (_00833_, _00580_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nand _23053_ (_00834_, _00833_, _00648_);
  and _23054_ (_00835_, _00833_, _00613_);
  or _23055_ (_00836_, _00835_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0]);
  and _23056_ (_00837_, _00836_, _05552_);
  and _23057_ (_13142_, _00837_, _00834_);
  not _23058_ (_00838_, _00580_);
  or _23059_ (_00839_, _00838_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and _23060_ (_00840_, _00839_, _05552_);
  not _23061_ (_00841_, _00610_);
  or _23062_ (_00842_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and _23063_ (_00843_, _00842_, _00841_);
  nor _23064_ (_00844_, _00595_, _08998_);
  nor _23065_ (_00845_, _00844_, _00598_);
  and _23066_ (_00846_, _00590_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or _23067_ (_00847_, _00846_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and _23068_ (_00848_, _00847_, _00610_);
  and _23069_ (_00849_, _00848_, _00845_);
  or _23070_ (_00850_, _00849_, _00843_);
  and _23071_ (_00851_, _00850_, _00603_);
  and _23072_ (_00852_, _00610_, _00598_);
  or _23073_ (_00853_, _00852_, _00602_);
  and _23074_ (_00854_, _00853_, _09009_);
  or _23075_ (_00855_, _00854_, _00851_);
  and _23076_ (_00856_, _00855_, _00613_);
  not _23077_ (_00857_, _00613_);
  and _23078_ (_00858_, _00842_, _00636_);
  or _23079_ (_00859_, _00858_, _00643_);
  and _23080_ (_00860_, _00624_, _09009_);
  not _23081_ (_00861_, _00642_);
  and _23082_ (_00862_, _00618_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _23083_ (_00863_, _00862_, _00624_);
  and _23084_ (_00864_, _00616_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or _23085_ (_00865_, _00864_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and _23086_ (_00866_, _00865_, _00863_);
  or _23087_ (_00867_, _00866_, _00861_);
  or _23088_ (_00868_, _00867_, _00860_);
  and _23089_ (_00869_, _00868_, _00859_);
  and _23090_ (_00870_, _00635_, _09009_);
  or _23091_ (_00871_, _00870_, _00647_);
  or _23092_ (_00872_, _00871_, _00869_);
  not _23093_ (_00873_, _00647_);
  or _23094_ (_00874_, _00873_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and _23095_ (_00875_, _00874_, _00872_);
  and _23096_ (_00876_, _00875_, _00857_);
  or _23097_ (_00877_, _00876_, _00856_);
  or _23098_ (_00878_, _00877_, _00580_);
  and _23099_ (_13150_, _00878_, _00840_);
  and _23100_ (_00879_, _00789_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and _23101_ (_00880_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and _23102_ (_00881_, _00824_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and _23103_ (_00882_, _00881_, _00880_);
  and _23104_ (_00883_, _00882_, _00769_);
  and _23105_ (_00884_, _00883_, _00748_);
  nor _23106_ (_00885_, _00766_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nor _23107_ (_00886_, _00885_, _00806_);
  and _23108_ (_00887_, _00886_, _00792_);
  nor _23109_ (_00888_, _00887_, _00884_);
  nor _23110_ (_00889_, _00888_, _00753_);
  or _23111_ (_00890_, _00889_, _00746_);
  or _23112_ (_00891_, _00890_, _00879_);
  nand _23113_ (_00892_, _00746_, _07945_);
  and _23114_ (_00893_, _00892_, _05552_);
  and _23115_ (_13154_, _00893_, _00891_);
  nor _23116_ (_00895_, _08386_, _07939_);
  and _23117_ (_00896_, _07939_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  or _23118_ (_00897_, _00896_, _00895_);
  and _23119_ (_13157_, _00897_, _05552_);
  nand _23120_ (_00898_, _00779_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nor _23121_ (_00899_, _00898_, _00753_);
  nor _23122_ (_00900_, _00806_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nor _23123_ (_00901_, _00900_, _00808_);
  and _23124_ (_00902_, _00901_, _00788_);
  or _23125_ (_00903_, _00902_, _00899_);
  and _23126_ (_00904_, _00789_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  or _23127_ (_00905_, _00904_, _00746_);
  or _23128_ (_00906_, _00905_, _00903_);
  nand _23129_ (_00907_, _00746_, _07975_);
  and _23130_ (_00908_, _00907_, _05552_);
  and _23131_ (_13163_, _00908_, _00906_);
  nor _23132_ (_00909_, _00808_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  or _23133_ (_00911_, _00909_, _00809_);
  nand _23134_ (_00912_, _00911_, _00788_);
  or _23135_ (_00913_, _00788_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  and _23136_ (_00914_, _00913_, _00912_);
  nand _23137_ (_00915_, _00779_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nor _23138_ (_00916_, _00915_, _00753_);
  or _23139_ (_00918_, _00916_, _00746_);
  or _23140_ (_00919_, _00918_, _00914_);
  nand _23141_ (_00920_, _00746_, _08041_);
  and _23142_ (_00921_, _00920_, _05552_);
  and _23143_ (_13167_, _00921_, _00919_);
  nand _23144_ (_00923_, _00648_, _00581_);
  and _23145_ (_00924_, _00613_, _00581_);
  or _23146_ (_00926_, _00924_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0]);
  and _23147_ (_00927_, _00926_, _05552_);
  and _23148_ (_13175_, _00927_, _00923_);
  not _23149_ (_00929_, _00746_);
  and _23150_ (_00931_, _00883_, _00766_);
  or _23151_ (_00932_, _00931_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  not _23152_ (_00934_, _00750_);
  and _23153_ (_00935_, _00931_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nor _23154_ (_00936_, _00935_, _00934_);
  and _23155_ (_00937_, _00936_, _00932_);
  nor _23156_ (_00939_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  not _23157_ (_00940_, _00939_);
  and _23158_ (_00942_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and _23159_ (_00943_, _00942_, _00772_);
  nor _23160_ (_00944_, _00943_, _00940_);
  or _23161_ (_00945_, _00944_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and _23162_ (_00946_, _00880_, _00794_);
  and _23163_ (_00947_, _00944_, _00946_);
  or _23164_ (_00948_, _00947_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and _23165_ (_00949_, _00948_, _00945_);
  nor _23166_ (_00950_, _00949_, _00937_);
  nor _23167_ (_00951_, _00950_, _00753_);
  not _23168_ (_00952_, _00753_);
  nor _23169_ (_00953_, _00952_, _07975_);
  or _23170_ (_00954_, _00953_, _00951_);
  and _23171_ (_00955_, _00954_, _00929_);
  and _23172_ (_00956_, _00746_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  or _23173_ (_00957_, _00956_, _00955_);
  and _23174_ (_13191_, _00957_, _05552_);
  nand _23175_ (_00958_, _00753_, _08041_);
  nand _23176_ (_00959_, _00943_, _00939_);
  nor _23177_ (_00960_, _00959_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and _23178_ (_00961_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and _23179_ (_00963_, _00961_, _00931_);
  or _23180_ (_00964_, _00935_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nand _23181_ (_00965_, _00964_, _00750_);
  nor _23182_ (_00967_, _00965_, _00963_);
  and _23183_ (_00968_, _00945_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  or _23184_ (_00969_, _00968_, _00967_);
  or _23185_ (_00971_, _00969_, _00960_);
  or _23186_ (_00972_, _00971_, _00753_);
  and _23187_ (_00973_, _00972_, _00929_);
  and _23188_ (_00974_, _00973_, _00958_);
  and _23189_ (_00975_, _00746_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  or _23190_ (_00976_, _00975_, _00974_);
  and _23191_ (_13194_, _00976_, _05552_);
  and _23192_ (_00977_, _00753_, _11238_);
  not _23193_ (_00978_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and _23194_ (_00979_, _00939_, _00795_);
  and _23195_ (_00980_, _00825_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and _23196_ (_00981_, _00980_, _00750_);
  nor _23197_ (_00982_, _00981_, _00979_);
  nand _23198_ (_00983_, _00982_, _00978_);
  or _23199_ (_00984_, _00982_, _00978_);
  nand _23200_ (_00985_, _00984_, _00983_);
  nor _23201_ (_00986_, _00985_, _00753_);
  or _23202_ (_00987_, _00986_, _00746_);
  or _23203_ (_00988_, _00987_, _00977_);
  nand _23204_ (_00989_, _00746_, _00978_);
  and _23205_ (_00991_, _00989_, _05552_);
  and _23206_ (_13197_, _00991_, _00988_);
  nand _23207_ (_00993_, _00753_, _07388_);
  or _23208_ (_00994_, _00963_, _00934_);
  and _23209_ (_00995_, _00961_, _00749_);
  and _23210_ (_00997_, _00995_, _00946_);
  or _23211_ (_00998_, _00997_, _00750_);
  and _23212_ (_01000_, _00998_, _00994_);
  nand _23213_ (_01001_, _01000_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and _23214_ (_01002_, _01001_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nor _23215_ (_01003_, _01001_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  or _23216_ (_01004_, _01003_, _01002_);
  or _23217_ (_01005_, _01004_, _00753_);
  and _23218_ (_01006_, _01005_, _00929_);
  and _23219_ (_01007_, _01006_, _00993_);
  and _23220_ (_01008_, _00746_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  or _23221_ (_01009_, _01008_, _01007_);
  and _23222_ (_13203_, _01009_, _05552_);
  nand _23223_ (_01010_, _00753_, _08386_);
  and _23224_ (_01011_, _00961_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and _23225_ (_01012_, _01011_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and _23226_ (_01013_, _01012_, _00931_);
  nor _23227_ (_01014_, _01013_, _00934_);
  and _23228_ (_01015_, _01012_, _00749_);
  and _23229_ (_01016_, _01015_, _00946_);
  nor _23230_ (_01017_, _01016_, _00750_);
  nor _23231_ (_01018_, _01017_, _01014_);
  nand _23232_ (_01019_, _01018_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and _23233_ (_01020_, _01019_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nor _23234_ (_01021_, _01019_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  or _23235_ (_01022_, _01021_, _01020_);
  or _23236_ (_01023_, _01022_, _00753_);
  and _23237_ (_01024_, _01023_, _00929_);
  and _23238_ (_01025_, _01024_, _01010_);
  and _23239_ (_01026_, _00746_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  or _23240_ (_01027_, _01026_, _01025_);
  and _23241_ (_13206_, _01027_, _05552_);
  nand _23242_ (_01029_, _00753_, _06306_);
  or _23243_ (_01030_, _01018_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and _23244_ (_01031_, _01030_, _01019_);
  or _23245_ (_01032_, _01031_, _00753_);
  and _23246_ (_01033_, _01032_, _00929_);
  and _23247_ (_01035_, _01033_, _01029_);
  and _23248_ (_01036_, _00746_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  or _23249_ (_01038_, _01036_, _01035_);
  and _23250_ (_13209_, _01038_, _05552_);
  nand _23251_ (_01039_, _00753_, _06560_);
  or _23252_ (_01040_, _01000_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and _23253_ (_01041_, _01040_, _01001_);
  or _23254_ (_01043_, _01041_, _00753_);
  and _23255_ (_01045_, _01043_, _00929_);
  and _23256_ (_01047_, _01045_, _01039_);
  and _23257_ (_01048_, _00746_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or _23258_ (_01049_, _01048_, _01047_);
  and _23259_ (_13212_, _01049_, _05552_);
  not _23260_ (_01050_, t0_i);
  and _23261_ (_01051_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , _01050_);
  nor _23262_ (_01052_, _01051_, _00073_);
  not _23263_ (_01053_, _01052_);
  not _23264_ (_01054_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  nor _23265_ (_01055_, \oc8051_top_1.oc8051_sfr1.pres_ow , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  nor _23266_ (_01056_, _01055_, _01054_);
  and _23267_ (_01058_, _01056_, _01053_);
  and _23268_ (_01059_, _01058_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  nor _23269_ (_01060_, _01059_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and _23270_ (_01061_, _01059_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  or _23271_ (_01063_, _01061_, _01060_);
  not _23272_ (_01064_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and _23273_ (_01066_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  and _23274_ (_01067_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  and _23275_ (_01068_, _01067_, _01066_);
  and _23276_ (_01069_, _01068_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and _23277_ (_01070_, _01069_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and _23278_ (_01071_, _01070_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and _23279_ (_01072_, _01071_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and _23280_ (_01074_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], _13526_);
  and _23281_ (_01075_, _01074_, _01058_);
  nand _23282_ (_01076_, _01075_, _01072_);
  or _23283_ (_01078_, _01076_, _01064_);
  and _23284_ (_01079_, _01078_, _01063_);
  and _23285_ (_01081_, _08989_, _08057_);
  and _23286_ (_01082_, _01081_, _07443_);
  nor _23287_ (_01084_, _01082_, _01079_);
  and _23288_ (_01085_, _01082_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  or _23289_ (_01087_, _01085_, _01084_);
  and _23290_ (_01089_, _10627_, _07443_);
  not _23291_ (_01091_, _01089_);
  and _23292_ (_01093_, _01091_, _01087_);
  nor _23293_ (_01095_, _01091_, _07975_);
  or _23294_ (_01096_, _01095_, _01093_);
  and _23295_ (_13215_, _01096_, _05552_);
  not _23296_ (_01098_, _01058_);
  nor _23297_ (_01100_, _01082_, _01098_);
  or _23298_ (_01101_, _01100_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and _23299_ (_01102_, _01074_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand _23300_ (_01104_, _01102_, _01072_);
  nand _23301_ (_01105_, _01104_, _01059_);
  or _23302_ (_01106_, _01105_, _01082_);
  and _23303_ (_01107_, _01106_, _01101_);
  or _23304_ (_01108_, _01107_, _01089_);
  nand _23305_ (_01109_, _01089_, _07945_);
  and _23306_ (_01110_, _01109_, _05552_);
  and _23307_ (_13219_, _01110_, _01108_);
  not _23308_ (_01111_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  nand _23309_ (_01112_, _01082_, _01111_);
  and _23310_ (_01113_, _01061_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  nor _23311_ (_01114_, _01061_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  nor _23312_ (_01115_, _01114_, _01113_);
  and _23313_ (_01116_, _01071_, _01058_);
  and _23314_ (_01117_, _01116_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and _23315_ (_01118_, _01074_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _23316_ (_01119_, _01118_, _01117_);
  or _23317_ (_01120_, _01119_, _01115_);
  or _23318_ (_01121_, _01120_, _01082_);
  and _23319_ (_01122_, _01121_, _01112_);
  or _23320_ (_01123_, _01122_, _01089_);
  nand _23321_ (_01124_, _01089_, _08041_);
  and _23322_ (_01126_, _01124_, _05552_);
  and _23323_ (_13237_, _01126_, _01123_);
  and _23324_ (_01127_, _01068_, _01058_);
  nor _23325_ (_01128_, _01127_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and _23326_ (_01129_, _01127_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  nor _23327_ (_01131_, _01129_, _01128_);
  and _23328_ (_01132_, _01072_, _01058_);
  and _23329_ (_01133_, _01074_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _23330_ (_01134_, _01133_, _01132_);
  nor _23331_ (_01136_, _01134_, _01131_);
  nor _23332_ (_01137_, _01136_, _01082_);
  and _23333_ (_01138_, _01082_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  or _23334_ (_01139_, _01138_, _01137_);
  and _23335_ (_01140_, _01139_, _01091_);
  nor _23336_ (_01141_, _01091_, _07388_);
  or _23337_ (_01142_, _01141_, _01140_);
  and _23338_ (_13242_, _01142_, _05552_);
  nor _23339_ (_01144_, _01113_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  nor _23340_ (_01145_, _01144_, _01127_);
  and _23341_ (_01146_, _01074_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and _23342_ (_01147_, _01146_, _01117_);
  or _23343_ (_01148_, _01147_, _01145_);
  or _23344_ (_01149_, _01148_, _01082_);
  not _23345_ (_01151_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  nand _23346_ (_01152_, _01082_, _01151_);
  and _23347_ (_01153_, _01152_, _01091_);
  and _23348_ (_01154_, _01153_, _01149_);
  nor _23349_ (_01155_, _01091_, _06560_);
  or _23350_ (_01156_, _01155_, _01154_);
  and _23351_ (_13245_, _01156_, _05552_);
  or _23352_ (_01157_, _00838_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and _23353_ (_01158_, _01157_, _05552_);
  and _23354_ (_01159_, _00853_, _09008_);
  or _23355_ (_01160_, _08998_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  or _23356_ (_01161_, _01160_, _00610_);
  and _23357_ (_01162_, _01161_, _00603_);
  and _23358_ (_01163_, _00590_, _08998_);
  or _23359_ (_01164_, _01163_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  nor _23360_ (_01165_, _00595_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _23361_ (_01166_, _01165_, _00598_);
  and _23362_ (_01167_, _01166_, _01164_);
  or _23363_ (_01168_, _01167_, _00841_);
  and _23364_ (_01170_, _01168_, _01162_);
  or _23365_ (_01171_, _01170_, _01159_);
  and _23366_ (_01172_, _01171_, _00613_);
  and _23367_ (_01173_, _01160_, _00636_);
  or _23368_ (_01174_, _01173_, _00643_);
  and _23369_ (_01175_, _00624_, _09008_);
  and _23370_ (_01176_, _00618_, _08998_);
  nor _23371_ (_01177_, _01176_, _00624_);
  and _23372_ (_01178_, _00616_, _08998_);
  or _23373_ (_01179_, _01178_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and _23374_ (_01180_, _01179_, _01177_);
  or _23375_ (_01181_, _01180_, _00861_);
  or _23376_ (_01183_, _01181_, _01175_);
  and _23377_ (_01184_, _01183_, _01174_);
  and _23378_ (_01185_, _00635_, _09008_);
  or _23379_ (_01186_, _01185_, _00647_);
  or _23380_ (_01187_, _01186_, _01184_);
  or _23381_ (_01188_, _00873_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and _23382_ (_01189_, _01188_, _01187_);
  and _23383_ (_01190_, _01189_, _00857_);
  or _23384_ (_01191_, _01190_, _01172_);
  or _23385_ (_01192_, _01191_, _00580_);
  and _23386_ (_13250_, _01192_, _01158_);
  or _23387_ (_01194_, _08998_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  or _23388_ (_01195_, _01194_, _00603_);
  not _23389_ (_01196_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  or _23390_ (_01197_, _01163_, _01196_);
  nand _23391_ (_01198_, _01197_, _01166_);
  or _23392_ (_01199_, _00599_, _08997_);
  and _23393_ (_01200_, _01199_, _01198_);
  or _23394_ (_01202_, _01200_, _00609_);
  not _23395_ (_01203_, _00607_);
  not _23396_ (_01204_, _00609_);
  or _23397_ (_01205_, _01194_, _01204_);
  and _23398_ (_01206_, _01205_, _01203_);
  and _23399_ (_01208_, _01206_, _01202_);
  and _23400_ (_01209_, _00607_, _08997_);
  or _23401_ (_01210_, _01209_, _00602_);
  or _23402_ (_01212_, _01210_, _01208_);
  and _23403_ (_01213_, _01212_, _01195_);
  or _23404_ (_01214_, _01213_, _00857_);
  or _23405_ (_01215_, _01194_, _00636_);
  or _23406_ (_01217_, _01178_, _01196_);
  nand _23407_ (_01218_, _01217_, _01177_);
  or _23408_ (_01219_, _00644_, _08997_);
  and _23409_ (_01220_, _01219_, _01218_);
  or _23410_ (_01221_, _01220_, _00641_);
  not _23411_ (_01222_, _00639_);
  not _23412_ (_01223_, _00641_);
  or _23413_ (_01224_, _01194_, _01223_);
  and _23414_ (_01225_, _01224_, _01222_);
  and _23415_ (_01226_, _01225_, _01221_);
  and _23416_ (_01227_, _00639_, _08997_);
  or _23417_ (_01228_, _01227_, _00635_);
  or _23418_ (_01229_, _01228_, _01226_);
  and _23419_ (_01230_, _01229_, _01215_);
  or _23420_ (_01231_, _01230_, _00649_);
  and _23421_ (_01232_, _01231_, _01214_);
  or _23422_ (_01233_, _01232_, _00580_);
  nor _23423_ (_01234_, _00873_, _00613_);
  nor _23424_ (_01235_, _01234_, _00580_);
  or _23425_ (_01236_, _01235_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  and _23426_ (_01237_, _01236_, _05552_);
  and _23427_ (_13262_, _01237_, _01233_);
  and _23428_ (_01238_, _05552_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  and _23429_ (_13271_, _01238_, _00580_);
  or _23430_ (_01239_, _00641_, _00624_);
  and _23431_ (_01240_, _00619_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or _23432_ (_01241_, _01240_, _01239_);
  and _23433_ (_01242_, _01241_, _01222_);
  and _23434_ (_01243_, _00648_, _00636_);
  and _23435_ (_01244_, _01243_, _01242_);
  or _23436_ (_01245_, _00609_, _00598_);
  and _23437_ (_01246_, _00596_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or _23438_ (_01247_, _01246_, _01245_);
  and _23439_ (_01248_, _01247_, _01203_);
  and _23440_ (_01249_, _00613_, _00603_);
  and _23441_ (_01250_, _01249_, _01248_);
  or _23442_ (_01251_, _01250_, _00580_);
  or _23443_ (_01252_, _01251_, _01244_);
  nand _23444_ (_01253_, _00580_, _05910_);
  and _23445_ (_01254_, _01253_, _05552_);
  and _23446_ (_13276_, _01254_, _01252_);
  nor _23447_ (_01255_, _00616_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nor _23448_ (_01256_, _01255_, _00618_);
  or _23449_ (_01257_, _01256_, _00624_);
  and _23450_ (_01258_, _01257_, _01223_);
  or _23451_ (_01259_, _01258_, _00639_);
  and _23452_ (_01260_, _01259_, _01243_);
  or _23453_ (_01261_, _00590_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and _23454_ (_01262_, _01261_, _00595_);
  or _23455_ (_01263_, _01262_, _00598_);
  and _23456_ (_01264_, _01263_, _01204_);
  or _23457_ (_01266_, _01264_, _00607_);
  and _23458_ (_01267_, _01266_, _01249_);
  or _23459_ (_01268_, _01267_, _00580_);
  or _23460_ (_01269_, _01268_, _01260_);
  or _23461_ (_01270_, _00838_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and _23462_ (_01271_, _01270_, _05552_);
  and _23463_ (_13279_, _01271_, _01269_);
  and _23464_ (_01272_, _00580_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  or _23465_ (_01273_, _01272_, _01235_);
  and _23466_ (_13282_, _01273_, _05552_);
  not _23467_ (_01274_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  nor _23468_ (_01275_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  not _23469_ (_01276_, _01275_);
  and _23470_ (_01277_, _01276_, _01058_);
  nand _23471_ (_01278_, _01277_, _01071_);
  nor _23472_ (_01279_, _01278_, _01082_);
  nor _23473_ (_01280_, _01279_, _01274_);
  not _23474_ (_01281_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or _23475_ (_01282_, _01076_, _01281_);
  not _23476_ (_01283_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  nor _23477_ (_01284_, _01275_, _01283_);
  and _23478_ (_01285_, _01284_, _01129_);
  nand _23479_ (_01286_, _01285_, _01278_);
  and _23480_ (_01287_, _01286_, _01282_);
  nor _23481_ (_01288_, _01287_, _01082_);
  or _23482_ (_01289_, _01288_, _01280_);
  and _23483_ (_01290_, _01289_, _01091_);
  nor _23484_ (_01291_, _01091_, _08386_);
  or _23485_ (_01292_, _01291_, _01290_);
  and _23486_ (_13293_, _01292_, _05552_);
  and _23487_ (_13296_, _00580_, _07727_);
  and _23488_ (_01293_, _01129_, _01276_);
  and _23489_ (_01294_, _01293_, _01283_);
  not _23490_ (_01295_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nor _23491_ (_01296_, _01076_, _01295_);
  nor _23492_ (_01297_, _01296_, _01294_);
  nor _23493_ (_01298_, _01297_, _01082_);
  not _23494_ (_01299_, _01293_);
  or _23495_ (_01300_, _01299_, _01082_);
  and _23496_ (_01301_, _01300_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  or _23497_ (_01302_, _01301_, _01298_);
  and _23498_ (_01303_, _01302_, _01091_);
  nor _23499_ (_01304_, _01091_, _06306_);
  or _23500_ (_01305_, _01304_, _01303_);
  and _23501_ (_13301_, _01305_, _05552_);
  nand _23502_ (_01306_, _01082_, _08386_);
  and _23503_ (_01307_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and _23504_ (_01308_, _01307_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _23505_ (_01309_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and _23506_ (_01310_, _01309_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _23507_ (_01311_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], \oc8051_top_1.oc8051_sfr1.pres_ow );
  and _23508_ (_01312_, _01311_, _01310_);
  and _23509_ (_01313_, _01312_, _01308_);
  and _23510_ (_01314_, _01313_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or _23511_ (_01315_, _01314_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and _23512_ (_01316_, _01312_, _01307_);
  and _23513_ (_01317_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and _23514_ (_01318_, _01317_, _01316_);
  nand _23515_ (_01319_, _01318_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and _23516_ (_01320_, _01319_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _23517_ (_01321_, _01320_, _01315_);
  and _23518_ (_01322_, _01308_, _01310_);
  and _23519_ (_01323_, _01322_, _01129_);
  nor _23520_ (_01324_, _01323_, _01281_);
  and _23521_ (_01325_, _01323_, _01281_);
  or _23522_ (_01326_, _01325_, _01324_);
  and _23523_ (_01327_, _01326_, _01275_);
  and _23524_ (_01328_, _01310_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and _23525_ (_01329_, _01328_, _01117_);
  nand _23526_ (_01330_, _01329_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or _23527_ (_01331_, _01330_, _01295_);
  nand _23528_ (_01332_, _01331_, _01281_);
  and _23529_ (_01333_, _00146_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or _23530_ (_01334_, _01331_, _01281_);
  and _23531_ (_01335_, _01334_, _01333_);
  and _23532_ (_01336_, _01335_, _01332_);
  or _23533_ (_01337_, _01336_, _01327_);
  or _23534_ (_01338_, _01337_, _01321_);
  or _23535_ (_01339_, _01338_, _01082_);
  and _23536_ (_01340_, _01339_, _01091_);
  and _23537_ (_01341_, _01340_, _01306_);
  and _23538_ (_01342_, _01089_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or _23539_ (_01343_, _01342_, _01341_);
  and _23540_ (_13330_, _01343_, _05552_);
  nand _23541_ (_01344_, _01082_, _08041_);
  and _23542_ (_01345_, _01309_, _01129_);
  or _23543_ (_01346_, _01345_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _23544_ (_01347_, _01345_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nor _23545_ (_01348_, _01347_, _01276_);
  and _23546_ (_01349_, _01348_, _01346_);
  and _23547_ (_01350_, _01309_, _01132_);
  or _23548_ (_01351_, _01350_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nand _23549_ (_01353_, _01310_, _01132_);
  and _23550_ (_01354_, _01353_, _01333_);
  and _23551_ (_01356_, _01354_, _01351_);
  and _23552_ (_01357_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and _23553_ (_01358_, _01311_, _01309_);
  or _23554_ (_01359_, _01358_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nand _23555_ (_01360_, _01359_, _01357_);
  nor _23556_ (_01361_, _01360_, _01312_);
  or _23557_ (_01362_, _01361_, _01118_);
  or _23558_ (_01364_, _01362_, _01356_);
  or _23559_ (_01365_, _01364_, _01349_);
  or _23560_ (_01367_, _01365_, _01082_);
  and _23561_ (_01368_, _01367_, _01091_);
  and _23562_ (_01369_, _01368_, _01344_);
  and _23563_ (_01370_, _01089_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  or _23564_ (_01371_, _01370_, _01369_);
  and _23565_ (_13338_, _01371_, _05552_);
  nand _23566_ (_01372_, _01082_, _06560_);
  or _23567_ (_01373_, _01347_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and _23568_ (_01374_, _01347_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  nor _23569_ (_01375_, _01374_, _01276_);
  and _23570_ (_01376_, _01375_, _01373_);
  or _23571_ (_01377_, _01312_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and _23572_ (_01378_, _01312_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  not _23573_ (_01379_, _01378_);
  and _23574_ (_01380_, _01379_, _01357_);
  and _23575_ (_01381_, _01380_, _01377_);
  and _23576_ (_01382_, _01132_, _00146_);
  and _23577_ (_01383_, _01382_, _01310_);
  or _23578_ (_01384_, _01383_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  or _23579_ (_01385_, _01333_, _01074_);
  nand _23580_ (_01386_, _01383_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and _23581_ (_01388_, _01386_, _01385_);
  and _23582_ (_01389_, _01388_, _01384_);
  or _23583_ (_01390_, _01389_, _01381_);
  or _23584_ (_01392_, _01390_, _01376_);
  or _23585_ (_01393_, _01392_, _01082_);
  and _23586_ (_01394_, _01393_, _01091_);
  and _23587_ (_01396_, _01394_, _01372_);
  and _23588_ (_01397_, _01089_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  or _23589_ (_01398_, _01397_, _01396_);
  and _23590_ (_13340_, _01398_, _05552_);
  nand _23591_ (_01399_, _01082_, _07388_);
  or _23592_ (_01400_, _01374_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _23593_ (_01401_, _01374_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nor _23594_ (_01402_, _01401_, _01276_);
  and _23595_ (_01404_, _01402_, _01400_);
  and _23596_ (_01405_, _01328_, _01132_);
  or _23597_ (_01406_, _01405_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _23598_ (_01407_, _01330_, _01333_);
  and _23599_ (_01408_, _01407_, _01406_);
  or _23600_ (_01409_, _01378_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nand _23601_ (_01410_, _01409_, _01357_);
  nor _23602_ (_01411_, _01410_, _01316_);
  or _23603_ (_01412_, _01411_, _01133_);
  or _23604_ (_01413_, _01412_, _01408_);
  or _23605_ (_01414_, _01413_, _01404_);
  or _23606_ (_01415_, _01414_, _01082_);
  and _23607_ (_01416_, _01415_, _01091_);
  and _23608_ (_01417_, _01416_, _01399_);
  and _23609_ (_01418_, _01089_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or _23610_ (_01419_, _01418_, _01417_);
  and _23611_ (_13348_, _01419_, _05552_);
  nand _23612_ (_01420_, _01082_, _06306_);
  or _23613_ (_01422_, _01401_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nand _23614_ (_01423_, _01401_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _23615_ (_01424_, _01423_, _01275_);
  and _23616_ (_01425_, _01424_, _01422_);
  or _23617_ (_01426_, _01316_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  not _23618_ (_01427_, _01313_);
  and _23619_ (_01428_, _01427_, _01357_);
  and _23620_ (_01429_, _01428_, _01426_);
  and _23621_ (_01430_, _01405_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _23622_ (_01431_, _01430_, _00146_);
  nor _23623_ (_01432_, _01431_, _01295_);
  and _23624_ (_01433_, _01431_, _01295_);
  or _23625_ (_01434_, _01433_, _01432_);
  and _23626_ (_01435_, _01434_, _01385_);
  or _23627_ (_01438_, _01435_, _01429_);
  or _23628_ (_01439_, _01438_, _01425_);
  or _23629_ (_01440_, _01439_, _01082_);
  and _23630_ (_01441_, _01440_, _01091_);
  and _23631_ (_01442_, _01441_, _01420_);
  and _23632_ (_01443_, _01089_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  or _23633_ (_01445_, _01443_, _01442_);
  and _23634_ (_13351_, _01445_, _05552_);
  nand _23635_ (_01446_, _01082_, _07975_);
  nand _23636_ (_01448_, _01382_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand _23637_ (_01450_, _01448_, _01064_);
  not _23638_ (_01451_, _01350_);
  and _23639_ (_01452_, _01451_, _01333_);
  or _23640_ (_01454_, _01452_, _01074_);
  and _23641_ (_01455_, _01454_, _01450_);
  and _23642_ (_01456_, _01311_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or _23643_ (_01457_, _01456_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  not _23644_ (_01458_, _01358_);
  and _23645_ (_01460_, _01458_, _01357_);
  and _23646_ (_01461_, _01460_, _01457_);
  and _23647_ (_01462_, _01129_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or _23648_ (_01463_, _01462_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nor _23649_ (_01464_, _01345_, _01276_);
  and _23650_ (_01465_, _01464_, _01463_);
  or _23651_ (_01466_, _01465_, _01461_);
  or _23652_ (_01467_, _01466_, _01455_);
  or _23653_ (_01468_, _01467_, _01082_);
  and _23654_ (_01469_, _01468_, _01446_);
  or _23655_ (_01470_, _01469_, _01089_);
  nand _23656_ (_01471_, _01089_, _01064_);
  and _23657_ (_01472_, _01471_, _05552_);
  and _23658_ (_13364_, _01472_, _01470_);
  or _23659_ (_01473_, _01382_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and _23660_ (_01474_, _01448_, _01385_);
  and _23661_ (_01475_, _01474_, _01473_);
  nor _23662_ (_01476_, _01311_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nor _23663_ (_01477_, _01476_, _01456_);
  and _23664_ (_01478_, _01477_, _01357_);
  or _23665_ (_01479_, _01129_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nor _23666_ (_01481_, _01462_, _01276_);
  and _23667_ (_01482_, _01481_, _01479_);
  or _23668_ (_01483_, _01482_, _01478_);
  or _23669_ (_01484_, _01483_, _01475_);
  or _23670_ (_01485_, _01484_, _01082_);
  nand _23671_ (_01486_, _01082_, _07945_);
  and _23672_ (_01487_, _01486_, _01485_);
  or _23673_ (_01488_, _01487_, _01089_);
  or _23674_ (_01489_, _01091_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and _23675_ (_01491_, _01489_, _05552_);
  and _23676_ (_13370_, _01491_, _01488_);
  and _23677_ (_01492_, _00245_, _07443_);
  nor _23678_ (_01494_, _01492_, _13526_);
  and _23679_ (_01495_, _01492_, _11238_);
  or _23680_ (_01496_, _01495_, _01494_);
  and _23681_ (_13376_, _01496_, _05552_);
  nor _23682_ (_01497_, _01492_, _00146_);
  and _23683_ (_01498_, _01492_, _11234_);
  or _23684_ (_01499_, _01498_, _01497_);
  and _23685_ (_13378_, _01499_, _05552_);
  or _23686_ (_01500_, _01492_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  and _23687_ (_01501_, _01500_, _05552_);
  nand _23688_ (_01502_, _01492_, _06560_);
  and _23689_ (_13388_, _01502_, _01501_);
  or _23690_ (_01503_, _01492_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and _23691_ (_01504_, _01503_, _05552_);
  nand _23692_ (_01505_, _01492_, _07388_);
  and _23693_ (_13393_, _01505_, _01504_);
  or _23694_ (_01506_, _01492_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and _23695_ (_01507_, _01506_, _05552_);
  nand _23696_ (_01508_, _01492_, _08041_);
  and _23697_ (_13396_, _01508_, _01507_);
  or _23698_ (_01509_, _01492_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and _23699_ (_01510_, _01509_, _05552_);
  nand _23700_ (_01511_, _01492_, _08386_);
  and _23701_ (_13403_, _01511_, _01510_);
  or _23702_ (_01512_, _01492_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and _23703_ (_01513_, _01512_, _05552_);
  nand _23704_ (_01514_, _01492_, _06306_);
  and _23705_ (_13406_, _01514_, _01513_);
  and _23706_ (_13470_, _08073_, _05552_);
  and _23707_ (_01515_, _00224_, _06765_);
  and _23708_ (_01516_, _01515_, _08635_);
  nand _23709_ (_01517_, _01516_, _06763_);
  nor _23710_ (_01518_, _06001_, _05989_);
  and _23711_ (_01519_, _01518_, _06926_);
  and _23712_ (_01520_, _01519_, _00240_);
  not _23713_ (_01521_, _01520_);
  or _23714_ (_01522_, _01516_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and _23715_ (_01523_, _01522_, _01521_);
  and _23716_ (_01524_, _01523_, _01517_);
  nor _23717_ (_01525_, _01521_, _06306_);
  or _23718_ (_01526_, _01525_, _01524_);
  and _23719_ (_13483_, _01526_, _05552_);
  and _23720_ (_01527_, _06054_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  or _23721_ (_01528_, _01527_, _08062_);
  and _23722_ (_01529_, _01528_, _01515_);
  nor _23723_ (_01530_, _06059_, _06054_);
  not _23724_ (_01531_, _01515_);
  or _23725_ (_01532_, _01531_, _01530_);
  and _23726_ (_01533_, _01532_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  or _23727_ (_01534_, _01533_, _01520_);
  or _23728_ (_01535_, _01534_, _01529_);
  nand _23729_ (_01536_, _01520_, _07388_);
  and _23730_ (_01537_, _01536_, _05552_);
  and _23731_ (_13490_, _01537_, _01535_);
  and _23732_ (_01538_, _01515_, _10632_);
  nand _23733_ (_01540_, _01538_, _06763_);
  or _23734_ (_01541_, _01538_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and _23735_ (_01543_, _01541_, _01521_);
  and _23736_ (_01544_, _01543_, _01540_);
  nor _23737_ (_01546_, _01521_, _06560_);
  or _23738_ (_01548_, _01546_, _01544_);
  and _23739_ (_13493_, _01548_, _05552_);
  and _23740_ (_13506_, _07677_, _05552_);
  and _23741_ (_01550_, _01515_, _06060_);
  nand _23742_ (_01551_, _01550_, _06763_);
  or _23743_ (_01552_, _01550_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and _23744_ (_01553_, _01552_, _01521_);
  and _23745_ (_01554_, _01553_, _01551_);
  and _23746_ (_01555_, _01520_, _11238_);
  or _23747_ (_01556_, _01555_, _01554_);
  and _23748_ (_13543_, _01556_, _05552_);
  and _23749_ (_01557_, _08990_, _06779_);
  or _23750_ (_01558_, _06770_, _06769_);
  not _23751_ (_01559_, _01558_);
  and _23752_ (_01560_, _10860_, _06779_);
  nand _23753_ (_01561_, _01560_, _01559_);
  and _23754_ (_01562_, _01561_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or _23755_ (_01563_, _01562_, _01557_);
  and _23756_ (_01564_, _06055_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or _23757_ (_01565_, _01564_, _08015_);
  and _23758_ (_01567_, _01565_, _01560_);
  or _23759_ (_01568_, _01567_, _01563_);
  nand _23760_ (_01570_, _01557_, _08041_);
  and _23761_ (_01572_, _01570_, _05552_);
  and _23762_ (_13558_, _01572_, _01568_);
  not _23763_ (_01573_, _01557_);
  and _23764_ (_01574_, _06064_, _05989_);
  and _23765_ (_01575_, _13693_, _01574_);
  and _23766_ (_01576_, _01575_, _06765_);
  and _23767_ (_01577_, _01576_, _06056_);
  or _23768_ (_01578_, _01577_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and _23769_ (_01579_, _01578_, _01573_);
  nand _23770_ (_01580_, _01577_, _06763_);
  and _23771_ (_01581_, _01580_, _01579_);
  nor _23772_ (_01582_, _01573_, _07975_);
  or _23773_ (_01583_, _01582_, _01581_);
  and _23774_ (_13564_, _01583_, _05552_);
  and _23775_ (_01585_, _01560_, _06060_);
  or _23776_ (_01586_, _01585_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and _23777_ (_01588_, _01586_, _01573_);
  nand _23778_ (_01589_, _01585_, _06763_);
  and _23779_ (_01590_, _01589_, _01588_);
  and _23780_ (_01591_, _01557_, _11238_);
  or _23781_ (_01592_, _01591_, _01590_);
  and _23782_ (_13569_, _01592_, _05552_);
  and _23783_ (_01595_, _01560_, _08365_);
  or _23784_ (_01597_, _01595_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and _23785_ (_01598_, _01597_, _01573_);
  nand _23786_ (_01599_, _01595_, _06763_);
  and _23787_ (_01600_, _01599_, _01598_);
  nor _23788_ (_01601_, _01573_, _08386_);
  or _23789_ (_01602_, _01601_, _01600_);
  and _23790_ (_13580_, _01602_, _05552_);
  and _23791_ (_01603_, _01560_, _08635_);
  or _23792_ (_01604_, _01603_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and _23793_ (_01605_, _01604_, _01573_);
  nand _23794_ (_01606_, _01603_, _06763_);
  and _23795_ (_01607_, _01606_, _01605_);
  nor _23796_ (_01608_, _01573_, _06306_);
  or _23797_ (_01609_, _01608_, _01607_);
  and _23798_ (_13587_, _01609_, _05552_);
  not _23799_ (_01610_, _01560_);
  or _23800_ (_01611_, _01610_, _08059_);
  and _23801_ (_01612_, _01611_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  or _23802_ (_01613_, _01612_, _01557_);
  and _23803_ (_01614_, _08058_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  or _23804_ (_01615_, _01614_, _08062_);
  and _23805_ (_01616_, _01615_, _01560_);
  or _23806_ (_01617_, _01616_, _01613_);
  nand _23807_ (_01618_, _01557_, _07388_);
  and _23808_ (_01619_, _01618_, _05552_);
  and _23809_ (_13590_, _01619_, _01617_);
  nand _23810_ (_13680_, _11699_, _05552_);
  nor _23811_ (_01620_, _07951_, _07388_);
  and _23812_ (_01621_, _07951_, _06070_);
  or _23813_ (_01622_, _01621_, _06062_);
  and _23814_ (_01623_, _01622_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  or _23815_ (_01624_, _06948_, _06309_);
  or _23816_ (_01625_, _01624_, _06058_);
  and _23817_ (_01626_, _06068_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  and _23818_ (_01627_, _01626_, _01625_);
  or _23819_ (_01628_, _01627_, _01623_);
  or _23820_ (_01629_, _01628_, _01620_);
  and _23821_ (_13682_, _01629_, _05552_);
  nor _23822_ (_13709_, _11250_, rst);
  nor _23823_ (_13714_, _11344_, rst);
  nor _23824_ (_13717_, _11429_, rst);
  nor _23825_ (_13720_, _11502_, rst);
  nand _23826_ (_13726_, _11757_, _05552_);
  and _23827_ (_01632_, _06068_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  and _23828_ (_01633_, _01632_, _13739_);
  and _23829_ (_01634_, _06070_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  and _23830_ (_01635_, _07976_, _06309_);
  or _23831_ (_01636_, _01635_, _01634_);
  or _23832_ (_01637_, _01636_, _01633_);
  and _23833_ (_13761_, _01637_, _05552_);
  and _23834_ (_01638_, _13740_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  and _23835_ (_01639_, _06068_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  and _23836_ (_01640_, _01639_, _13742_);
  and _23837_ (_01641_, _09504_, _07946_);
  or _23838_ (_01642_, _01641_, _01640_);
  or _23839_ (_01643_, _01642_, _01638_);
  and _23840_ (_00025_, _01643_, _05552_);
  and _23841_ (_01644_, _06072_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  and _23842_ (_01645_, _11490_, _06310_);
  or _23843_ (_01646_, _01645_, _01644_);
  and _23844_ (_00060_, _01646_, _05552_);
  and _23845_ (_01647_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor _23846_ (_01648_, _05550_, _11609_);
  or _23847_ (_01649_, _01648_, _01647_);
  and _23848_ (_00071_, _01649_, _05552_);
  and _23849_ (_01650_, _06072_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  and _23850_ (_01651_, _07439_, _06310_);
  or _23851_ (_01652_, _01651_, _01650_);
  and _23852_ (_00076_, _01652_, _05552_);
  and _23853_ (_00085_, _07522_, _05552_);
  nor _23854_ (_01653_, _09030_, _06811_);
  and _23855_ (_01654_, _09030_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  or _23856_ (_01655_, _01654_, _01653_);
  and _23857_ (_00122_, _01655_, _05552_);
  and _23858_ (_00153_, _07610_, _05552_);
  and _23859_ (_01656_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and _23860_ (_01657_, _12140_, \oc8051_top_1.oc8051_rom1.data_o [30]);
  or _23861_ (_01658_, _01657_, _01656_);
  and _23862_ (_00159_, _01658_, _05552_);
  or _23863_ (_01659_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  nand _23864_ (_01660_, _05550_, _05652_);
  and _23865_ (_01661_, _01660_, _05552_);
  and _23866_ (_00201_, _01661_, _01659_);
  and _23867_ (_00205_, _12169_, _05552_);
  and _23868_ (_01662_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  nor _23869_ (_01663_, _05550_, _07743_);
  or _23870_ (_01665_, _01663_, _01662_);
  and _23871_ (_00206_, _01665_, _05552_);
  and _23872_ (_01667_, _06068_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  and _23873_ (_01668_, _01667_, _13739_);
  and _23874_ (_01669_, _06070_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  and _23875_ (_01670_, _11726_, _06310_);
  or _23876_ (_01671_, _01670_, _01669_);
  or _23877_ (_01672_, _01671_, _01668_);
  and _23878_ (_00219_, _01672_, _05552_);
  and _23879_ (_00235_, _07454_, _05552_);
  nor _23880_ (_01673_, _09505_, _06811_);
  and _23881_ (_01674_, _09505_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  or _23882_ (_01675_, _01674_, _06955_);
  or _23883_ (_01676_, _01675_, _01673_);
  or _23884_ (_01677_, _06068_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  and _23885_ (_01678_, _01677_, _05552_);
  and _23886_ (_00247_, _01678_, _01676_);
  and _23887_ (_01679_, _11076_, _05886_);
  or _23888_ (_01681_, _11174_, _05833_);
  or _23889_ (_01682_, _11155_, _11078_);
  not _23890_ (_01683_, _11170_);
  or _23891_ (_01684_, _13392_, _01683_);
  or _23892_ (_01685_, _01684_, _01682_);
  or _23893_ (_01687_, _01685_, _01681_);
  and _23894_ (_01688_, _01687_, _11084_);
  or _23895_ (_01689_, _01688_, _01679_);
  and _23896_ (_00251_, _01689_, _05552_);
  nand _23897_ (_01690_, _10861_, _06056_);
  nor _23898_ (_01691_, _01690_, _06763_);
  nand _23899_ (_01692_, _09001_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  or _23900_ (_01693_, _09012_, _09006_);
  or _23901_ (_01694_, _01693_, _01692_);
  nand _23902_ (_01695_, _01694_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  nand _23903_ (_01696_, _01695_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and _23904_ (_01697_, _01696_, _01690_);
  or _23905_ (_01698_, _01697_, _08991_);
  or _23906_ (_01699_, _01698_, _01691_);
  nand _23907_ (_01700_, _08991_, _07975_);
  and _23908_ (_01701_, _01700_, _05552_);
  and _23909_ (_00269_, _01701_, _01699_);
  nand _23910_ (_01702_, _11098_, _05552_);
  nor _23911_ (_02255_, _01702_, _11141_);
  and _23912_ (_00271_, _02255_, _11258_);
  nand _23913_ (_01703_, _10861_, _10632_);
  nor _23914_ (_01704_, _01703_, _06763_);
  and _23915_ (_01705_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or _23916_ (_01706_, _01692_, _09013_);
  and _23917_ (_01707_, _01706_, _01705_);
  and _23918_ (_01708_, _01707_, _01703_);
  or _23919_ (_01709_, _01708_, _08991_);
  or _23920_ (_01710_, _01709_, _01704_);
  nand _23921_ (_01711_, _08991_, _06560_);
  and _23922_ (_01712_, _01711_, _05552_);
  and _23923_ (_00274_, _01712_, _01710_);
  or _23924_ (_01714_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  nand _23925_ (_01715_, _05550_, _05695_);
  and _23926_ (_01716_, _01715_, _05552_);
  and _23927_ (_00291_, _01716_, _01714_);
  and _23928_ (_01717_, _06068_, _06062_);
  nand _23929_ (_01718_, _01717_, _07945_);
  or _23930_ (_01719_, _01717_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  and _23931_ (_01720_, _01719_, _01718_);
  and _23932_ (_00328_, _01720_, _05552_);
  and _23933_ (_00331_, _08113_, _05552_);
  and _23934_ (_01721_, _01560_, _06771_);
  or _23935_ (_01722_, _01721_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and _23936_ (_01723_, _01722_, _01573_);
  nand _23937_ (_01724_, _01721_, _06763_);
  and _23938_ (_01725_, _01724_, _01723_);
  nor _23939_ (_01726_, _01573_, _06811_);
  or _23940_ (_01727_, _01726_, _01725_);
  and _23941_ (_00336_, _01727_, _05552_);
  and _23942_ (_01728_, _05567_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  and _23943_ (_01729_, _01728_, _05576_);
  or _23944_ (_01730_, _01729_, _06320_);
  and _23945_ (_01731_, _01730_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  nand _23946_ (_01732_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor _23947_ (_01733_, _01732_, _05586_);
  or _23948_ (_01734_, _01733_, _13411_);
  or _23949_ (_01735_, _01734_, _01731_);
  and _23950_ (_00342_, _01735_, _05552_);
  and _23951_ (_00475_, _07698_, _05552_);
  or _23952_ (_01736_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  and _23953_ (_01738_, _10626_, _10860_);
  or _23954_ (_01739_, _01738_, _01736_);
  not _23955_ (_01740_, _06771_);
  nor _23956_ (_01741_, _01740_, _06763_);
  nand _23957_ (_01742_, _01740_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  nand _23958_ (_01743_, _01742_, _01738_);
  or _23959_ (_01744_, _01743_, _01741_);
  and _23960_ (_01745_, _01744_, _01739_);
  and _23961_ (_01746_, _10626_, _08990_);
  or _23962_ (_01747_, _01746_, _01745_);
  nand _23963_ (_01748_, _01746_, _06811_);
  and _23964_ (_01749_, _01748_, _05552_);
  and _23965_ (_00514_, _01749_, _01747_);
  and _23966_ (_01750_, _07262_, _06915_);
  nand _23967_ (_01751_, _01750_, _06060_);
  or _23968_ (_01752_, _01751_, _07635_);
  not _23969_ (_01753_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nand _23970_ (_01754_, _01751_, _01753_);
  and _23971_ (_01755_, _01754_, _06524_);
  and _23972_ (_01756_, _01755_, _01752_);
  nor _23973_ (_01757_, _06774_, _01753_);
  and _23974_ (_01758_, _01750_, _08635_);
  nand _23975_ (_01759_, _01758_, _06763_);
  or _23976_ (_01760_, _01758_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and _23977_ (_01762_, _01760_, _06775_);
  and _23978_ (_01763_, _01762_, _01759_);
  or _23979_ (_01764_, _01763_, _01757_);
  or _23980_ (_01765_, _01764_, _01756_);
  and _23981_ (_00530_, _01765_, _05552_);
  or _23982_ (_01766_, _01751_, _12189_);
  not _23983_ (_01767_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nand _23984_ (_01768_, _01751_, _01767_);
  and _23985_ (_01769_, _01768_, _06524_);
  and _23986_ (_01770_, _01769_, _01766_);
  nor _23987_ (_01771_, _06774_, _01767_);
  not _23988_ (_01772_, _01750_);
  or _23989_ (_01773_, _01772_, _01530_);
  and _23990_ (_01774_, _01773_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and _23991_ (_01775_, _06054_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  or _23992_ (_01776_, _01775_, _08062_);
  and _23993_ (_01777_, _01776_, _01750_);
  or _23994_ (_01778_, _01777_, _01774_);
  and _23995_ (_01779_, _01778_, _06775_);
  or _23996_ (_01780_, _01779_, _01771_);
  or _23997_ (_01781_, _01780_, _01770_);
  and _23998_ (_00533_, _01781_, _05552_);
  or _23999_ (_01782_, _05550_, \oc8051_top_1.oc8051_rom1.data_o [10]);
  nand _24000_ (_01783_, _05550_, _11739_);
  and _24001_ (_01784_, _01783_, _05552_);
  and _24002_ (_00549_, _01784_, _01782_);
  not _24003_ (_01785_, _06321_);
  and _24004_ (_01786_, _09817_, _01785_);
  or _24005_ (_01787_, _01729_, _06319_);
  and _24006_ (_01788_, _05585_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  and _24007_ (_01789_, _01788_, _01787_);
  or _24008_ (_00604_, _01789_, _01786_);
  and _24009_ (_01790_, _05917_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  or _24010_ (_01791_, _01790_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  and _24011_ (_00606_, _01791_, _05552_);
  nor _24012_ (_01792_, _00329_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  nor _24013_ (_01793_, _01792_, _00330_);
  and _24014_ (_00682_, _01793_, _00335_);
  nor _24015_ (_01795_, _00254_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  nor _24016_ (_01796_, _01795_, _00329_);
  and _24017_ (_00684_, _01796_, _00335_);
  and _24018_ (_01798_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor _24019_ (_01799_, _05550_, _08689_);
  or _24020_ (_01800_, _01799_, _01798_);
  and _24021_ (_00771_, _01800_, _05552_);
  and _24022_ (_01801_, _01081_, _10626_);
  and _24023_ (_01802_, _00752_, _10626_);
  nor _24024_ (_01803_, _01802_, _01801_);
  and _24025_ (_01804_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and _24026_ (_01805_, _01804_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and _24027_ (_01806_, _01805_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and _24028_ (_01807_, _01806_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and _24029_ (_01808_, _01807_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and _24030_ (_01809_, _01808_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and _24031_ (_01810_, _01809_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and _24032_ (_01811_, _01810_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and _24033_ (_01812_, _01811_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and _24034_ (_01813_, _01812_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and _24035_ (_01814_, _01813_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and _24036_ (_01815_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  and _24037_ (_01816_, _01815_, _01814_);
  and _24038_ (_01818_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  and _24039_ (_01819_, _01818_, _01816_);
  or _24040_ (_01820_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1], \oc8051_top_1.oc8051_sfr1.pres_ow );
  not _24041_ (_01821_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or _24042_ (_01822_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _01821_);
  and _24043_ (_01823_, _01822_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and _24044_ (_01824_, _01823_, _01820_);
  not _24045_ (_01825_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and _24046_ (_01826_, _10638_, _01825_);
  and _24047_ (_01827_, _01826_, _10639_);
  not _24048_ (_01828_, _01827_);
  and _24049_ (_01829_, _01828_, _01824_);
  and _24050_ (_01830_, _01829_, _01819_);
  nand _24051_ (_01831_, _01830_, _10639_);
  nand _24052_ (_01832_, _01831_, _01803_);
  or _24053_ (_01833_, _01803_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and _24054_ (_01834_, _01833_, _05552_);
  and _24055_ (_00793_, _01834_, _01832_);
  or _24056_ (_01835_, _01751_, _08144_);
  not _24057_ (_01836_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  nand _24058_ (_01837_, _01751_, _01836_);
  and _24059_ (_01838_, _01837_, _06524_);
  and _24060_ (_01839_, _01838_, _01835_);
  nor _24061_ (_01840_, _06774_, _01836_);
  nand _24062_ (_01841_, _01750_, _01559_);
  and _24063_ (_01842_, _01841_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and _24064_ (_01843_, _06055_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or _24065_ (_01844_, _01843_, _08015_);
  and _24066_ (_01845_, _01844_, _01750_);
  or _24067_ (_01846_, _01845_, _01842_);
  and _24068_ (_01847_, _01846_, _06775_);
  or _24069_ (_01848_, _01847_, _01840_);
  or _24070_ (_01849_, _01848_, _01839_);
  and _24071_ (_00807_, _01849_, _05552_);
  or _24072_ (_01850_, _01751_, _08102_);
  not _24073_ (_01851_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  nand _24074_ (_01852_, _01751_, _01851_);
  and _24075_ (_01853_, _01852_, _06524_);
  and _24076_ (_01854_, _01853_, _01850_);
  nor _24077_ (_01855_, _06774_, _01851_);
  and _24078_ (_01856_, _01750_, _06056_);
  nand _24079_ (_01857_, _01856_, _06763_);
  or _24080_ (_01858_, _01856_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and _24081_ (_01859_, _01858_, _06775_);
  and _24082_ (_01860_, _01859_, _01857_);
  or _24083_ (_01861_, _01860_, _01855_);
  or _24084_ (_01862_, _01861_, _01854_);
  and _24085_ (_00815_, _01862_, _05552_);
  and _24086_ (_00894_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _05552_);
  and _24087_ (_00910_, _07995_, _05552_);
  not _24088_ (_01865_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and _24089_ (_01866_, _10638_, _01865_);
  or _24090_ (_01867_, _01866_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or _24091_ (_01868_, _01867_, _01738_);
  nand _24092_ (_01869_, _08366_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  nand _24093_ (_01870_, _01869_, _01738_);
  or _24094_ (_01871_, _01870_, _08367_);
  and _24095_ (_01872_, _01871_, _01868_);
  or _24096_ (_01873_, _01872_, _01746_);
  nand _24097_ (_01874_, _01746_, _08386_);
  and _24098_ (_01875_, _01874_, _05552_);
  and _24099_ (_00917_, _01875_, _01873_);
  not _24100_ (_01876_, _01746_);
  and _24101_ (_01877_, _01738_, _08635_);
  or _24102_ (_01878_, _01877_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and _24103_ (_01879_, _01878_, _01876_);
  nand _24104_ (_01880_, _01877_, _06763_);
  and _24105_ (_01881_, _01880_, _01879_);
  nor _24106_ (_01882_, _01876_, _06306_);
  or _24107_ (_01883_, _01882_, _01881_);
  and _24108_ (_00922_, _01883_, _05552_);
  or _24109_ (_01885_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  not _24110_ (_01886_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nand _24111_ (_01888_, pc_log_change, _01886_);
  and _24112_ (_01889_, _01888_, _05552_);
  and _24113_ (_00925_, _01889_, _01885_);
  not _24114_ (_01890_, _01738_);
  or _24115_ (_01891_, _01890_, _08059_);
  and _24116_ (_01892_, _01891_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  or _24117_ (_01893_, _01892_, _01746_);
  and _24118_ (_01894_, _08058_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  or _24119_ (_01896_, _01894_, _08062_);
  and _24120_ (_01897_, _01896_, _01738_);
  or _24121_ (_01898_, _01897_, _01893_);
  nand _24122_ (_01900_, _01746_, _07388_);
  and _24123_ (_01901_, _01900_, _05552_);
  and _24124_ (_00928_, _01901_, _01898_);
  and _24125_ (_01902_, _01738_, _10632_);
  or _24126_ (_01903_, _01902_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and _24127_ (_01905_, _01903_, _01876_);
  nand _24128_ (_01906_, _01902_, _06763_);
  and _24129_ (_01907_, _01906_, _01905_);
  nor _24130_ (_01908_, _01876_, _06560_);
  or _24131_ (_01909_, _01908_, _01907_);
  and _24132_ (_00930_, _01909_, _05552_);
  or _24133_ (_01910_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  not _24134_ (_01911_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nand _24135_ (_01912_, pc_log_change, _01911_);
  and _24136_ (_01913_, _01912_, _05552_);
  and _24137_ (_00933_, _01913_, _01910_);
  or _24138_ (_01914_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  not _24139_ (_01915_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nand _24140_ (_01916_, pc_log_change, _01915_);
  and _24141_ (_01917_, _01916_, _05552_);
  and _24142_ (_00938_, _01917_, _01914_);
  and _24143_ (_01919_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  not _24144_ (_01920_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor _24145_ (_01921_, pc_log_change, _01920_);
  or _24146_ (_01922_, _01921_, _01919_);
  and _24147_ (_00941_, _01922_, _05552_);
  and _24148_ (_01923_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  not _24149_ (_01924_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nor _24150_ (_01925_, pc_log_change, _01924_);
  or _24151_ (_01926_, _01925_, _01923_);
  and _24152_ (_00962_, _01926_, _05552_);
  nand _24153_ (_01927_, _01738_, _01559_);
  and _24154_ (_01928_, _01927_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or _24155_ (_01929_, _01928_, _01746_);
  and _24156_ (_01930_, _06055_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or _24157_ (_01931_, _01930_, _08015_);
  and _24158_ (_01933_, _01931_, _01738_);
  or _24159_ (_01934_, _01933_, _01929_);
  nand _24160_ (_01935_, _01746_, _08041_);
  and _24161_ (_01936_, _01935_, _05552_);
  and _24162_ (_00966_, _01936_, _01934_);
  and _24163_ (_01937_, _01575_, _08007_);
  and _24164_ (_01938_, _01937_, _06056_);
  or _24165_ (_01939_, _01938_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  and _24166_ (_01940_, _01939_, _01876_);
  nand _24167_ (_01941_, _01938_, _06763_);
  and _24168_ (_01942_, _01941_, _01940_);
  nor _24169_ (_01943_, _01876_, _07975_);
  or _24170_ (_01944_, _01943_, _01942_);
  and _24171_ (_00970_, _01944_, _05552_);
  and _24172_ (_01945_, _01738_, _06060_);
  or _24173_ (_01946_, _01945_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and _24174_ (_01947_, _01946_, _01876_);
  nand _24175_ (_01948_, _01945_, _06763_);
  and _24176_ (_01949_, _01948_, _01947_);
  and _24177_ (_01950_, _01746_, _11238_);
  or _24178_ (_01951_, _01950_, _01949_);
  and _24179_ (_00990_, _01951_, _05552_);
  or _24180_ (_01952_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nand _24181_ (_01953_, pc_log_change, _06192_);
  and _24182_ (_01954_, _01953_, _05552_);
  and _24183_ (_00992_, _01954_, _01952_);
  and _24184_ (_01955_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  not _24185_ (_01956_, pc_log_change);
  and _24186_ (_01957_, _01956_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  or _24187_ (_01958_, _01957_, _01955_);
  and _24188_ (_00996_, _01958_, _05552_);
  and _24189_ (_01959_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  not _24190_ (_01960_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor _24191_ (_01961_, pc_log_change, _01960_);
  or _24192_ (_01962_, _01961_, _01959_);
  and _24193_ (_00999_, _01962_, _05552_);
  and _24194_ (_01963_, _01824_, _01816_);
  and _24195_ (_01964_, _01963_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  nor _24196_ (_01965_, _01963_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  nor _24197_ (_01966_, _01965_, _01964_);
  not _24198_ (_01967_, _10641_);
  and _24199_ (_01968_, _01967_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and _24200_ (_01969_, _01968_, _01824_);
  and _24201_ (_01970_, _01969_, _01819_);
  or _24202_ (_01971_, _01970_, _01827_);
  or _24203_ (_01972_, _01971_, _01966_);
  or _24204_ (_01973_, _01828_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and _24205_ (_01974_, _01973_, _01803_);
  and _24206_ (_01975_, _01974_, _01972_);
  and _24207_ (_01976_, _01801_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or _24208_ (_01977_, _01976_, _01975_);
  not _24209_ (_01978_, _01802_);
  nor _24210_ (_01979_, _01978_, _08386_);
  or _24211_ (_01980_, _01979_, _01977_);
  and _24212_ (_01028_, _01980_, _05552_);
  and _24213_ (_01981_, _01801_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  and _24214_ (_01982_, _01824_, _01814_);
  and _24215_ (_01983_, _01982_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  nor _24216_ (_01984_, _01983_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  nor _24217_ (_01985_, _01984_, _01963_);
  and _24218_ (_01986_, _01967_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and _24219_ (_01987_, _01986_, _01824_);
  and _24220_ (_01988_, _01987_, _01819_);
  or _24221_ (_01989_, _01988_, _01827_);
  or _24222_ (_01990_, _01989_, _01985_);
  or _24223_ (_01991_, _01828_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and _24224_ (_01992_, _01991_, _01803_);
  and _24225_ (_01993_, _01992_, _01990_);
  nor _24226_ (_01994_, _01978_, _06306_);
  or _24227_ (_01995_, _01994_, _01993_);
  or _24228_ (_01996_, _01995_, _01981_);
  and _24229_ (_01034_, _01996_, _05552_);
  not _24230_ (_01997_, _01801_);
  or _24231_ (_01998_, _01997_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or _24232_ (_01999_, _01982_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  nor _24233_ (_02000_, _01983_, _01827_);
  or _24234_ (_02001_, _02000_, _01801_);
  and _24235_ (_02002_, _02001_, _01999_);
  and _24236_ (_02003_, _01827_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and _24237_ (_02005_, _01967_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and _24238_ (_02006_, _02005_, _01830_);
  or _24239_ (_02007_, _02006_, _02003_);
  or _24240_ (_02008_, _02007_, _02002_);
  and _24241_ (_02009_, _02008_, _01998_);
  or _24242_ (_02011_, _02009_, _01802_);
  nand _24243_ (_02013_, _01802_, _07388_);
  and _24244_ (_02014_, _02013_, _05552_);
  and _24245_ (_01037_, _02014_, _02011_);
  or _24246_ (_02015_, _01279_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  not _24247_ (_02016_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and _24248_ (_02017_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], _02016_);
  or _24249_ (_02018_, _02017_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  nand _24250_ (_02019_, _02018_, _01132_);
  or _24251_ (_02020_, _02019_, _01082_);
  and _24252_ (_02021_, _02020_, _01091_);
  and _24253_ (_02022_, _02021_, _02015_);
  nor _24254_ (_02023_, _01091_, _06811_);
  or _24255_ (_02024_, _02023_, _02022_);
  and _24256_ (_01042_, _02024_, _05552_);
  nor _24257_ (_02025_, _01082_, rst);
  not _24258_ (_02026_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 );
  nor _24259_ (_02027_, _01311_, _02026_);
  and _24260_ (_02028_, _01322_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and _24261_ (_02029_, _02028_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and _24262_ (_02030_, _02029_, _01311_);
  or _24263_ (_02031_, _02030_, _02027_);
  nand _24264_ (_02032_, _02031_, _01357_);
  nor _24265_ (_02033_, _02032_, _01089_);
  and _24266_ (_01044_, _02033_, _02025_);
  nand _24267_ (_02034_, _01082_, _06811_);
  and _24268_ (_02035_, _01431_, _01317_);
  or _24269_ (_02036_, _02035_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand _24270_ (_02037_, _02035_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and _24271_ (_02038_, _02037_, _01385_);
  and _24272_ (_02039_, _02038_, _02036_);
  nor _24273_ (_02040_, _01318_, _02016_);
  and _24274_ (_02041_, _01318_, _02016_);
  or _24275_ (_02042_, _02041_, _02040_);
  and _24276_ (_02043_, _02042_, _01357_);
  and _24277_ (_02044_, _01069_, _01058_);
  and _24278_ (_02045_, _02044_, _02028_);
  or _24279_ (_02046_, _02045_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and _24280_ (_02047_, _02044_, _02029_);
  nor _24281_ (_02048_, _02047_, _01276_);
  and _24282_ (_02049_, _02048_, _02046_);
  or _24283_ (_02050_, _02049_, _02043_);
  or _24284_ (_02051_, _02050_, _02039_);
  or _24285_ (_02052_, _02051_, _01082_);
  and _24286_ (_02053_, _02052_, _01091_);
  and _24287_ (_02054_, _02053_, _02034_);
  and _24288_ (_02055_, _01089_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or _24289_ (_02056_, _02055_, _02054_);
  and _24290_ (_01046_, _02056_, _05552_);
  or _24291_ (_02057_, _01492_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and _24292_ (_02058_, _02057_, _05552_);
  nand _24293_ (_02059_, _01492_, _06811_);
  and _24294_ (_01057_, _02059_, _02058_);
  and _24295_ (_02060_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  not _24296_ (_02061_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  nor _24297_ (_02062_, pc_log_change, _02061_);
  or _24298_ (_02063_, _02062_, _02060_);
  and _24299_ (_01062_, _02063_, _05552_);
  or _24300_ (_02064_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  not _24301_ (_02065_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  nand _24302_ (_02066_, pc_log_change, _02065_);
  and _24303_ (_02067_, _02066_, _05552_);
  and _24304_ (_01065_, _02067_, _02064_);
  and _24305_ (_02068_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor _24306_ (_02069_, pc_log_change, _01886_);
  or _24307_ (_02070_, _02069_, _02068_);
  and _24308_ (_01073_, _02070_, _05552_);
  and _24309_ (_02071_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nor _24310_ (_02072_, pc_log_change, _01915_);
  or _24311_ (_02073_, _02072_, _02071_);
  and _24312_ (_01077_, _02073_, _05552_);
  and _24313_ (_01080_, t0_i, _05552_);
  and _24314_ (_01083_, t1_i, _05552_);
  and _24315_ (_02075_, _01967_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and _24316_ (_02076_, _01824_, _01819_);
  and _24317_ (_02077_, _02076_, _02075_);
  not _24318_ (_02078_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  nand _24319_ (_02079_, _01824_, _01813_);
  and _24320_ (_02080_, _02079_, _02078_);
  nor _24321_ (_02081_, _02080_, _01982_);
  or _24322_ (_02082_, _02081_, _01827_);
  or _24323_ (_02083_, _02082_, _02077_);
  nor _24324_ (_02084_, _01828_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  nor _24325_ (_02085_, _02084_, _01801_);
  and _24326_ (_02086_, _02085_, _02083_);
  and _24327_ (_02087_, _01801_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or _24328_ (_02088_, _02087_, _01802_);
  or _24329_ (_02090_, _02088_, _02086_);
  nand _24330_ (_02091_, _01802_, _06560_);
  and _24331_ (_02092_, _02091_, _05552_);
  and _24332_ (_01086_, _02092_, _02090_);
  nand _24333_ (_02093_, _00753_, _06811_);
  and _24334_ (_02094_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and _24335_ (_02095_, _02094_, _01011_);
  and _24336_ (_02096_, _02095_, _00931_);
  and _24337_ (_02097_, _02096_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  or _24338_ (_02098_, _02097_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and _24339_ (_02099_, _02097_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor _24340_ (_02100_, _02099_, _00934_);
  and _24341_ (_02101_, _02100_, _02098_);
  and _24342_ (_02102_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and _24343_ (_02103_, _02102_, _01012_);
  and _24344_ (_02104_, _02103_, _00946_);
  or _24345_ (_02105_, _02104_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and _24346_ (_02106_, _02104_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor _24347_ (_02107_, _02106_, _00940_);
  and _24348_ (_02108_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  or _24349_ (_02109_, _02108_, _02107_);
  and _24350_ (_02110_, _02109_, _02105_);
  or _24351_ (_02111_, _02110_, _02101_);
  or _24352_ (_02112_, _02111_, _00753_);
  and _24353_ (_02113_, _02112_, _00929_);
  and _24354_ (_02114_, _02113_, _02093_);
  and _24355_ (_02115_, _00746_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  or _24356_ (_02116_, _02115_, _02114_);
  and _24357_ (_01088_, _02116_, _05552_);
  and _24358_ (_02118_, _01098_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  or _24359_ (_02119_, _02118_, _02047_);
  and _24360_ (_02120_, _02119_, _01275_);
  or _24361_ (_02121_, _02118_, _01132_);
  or _24362_ (_02122_, _02118_, _02029_);
  and _24363_ (_02123_, _02122_, _01333_);
  or _24364_ (_02124_, _02123_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _24365_ (_02125_, _02124_, _02121_);
  nor _24366_ (_02126_, _02125_, _02120_);
  nor _24367_ (_02127_, _02126_, _01089_);
  and _24368_ (_01090_, _02127_, _02025_);
  not _24369_ (_02128_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  nor _24370_ (_02129_, _00766_, _02128_);
  or _24371_ (_02130_, _02129_, _02106_);
  and _24372_ (_02131_, _02130_, _00939_);
  or _24373_ (_02132_, _02129_, _02099_);
  and _24374_ (_02133_, _02132_, _00750_);
  and _24375_ (_02134_, _00787_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  and _24376_ (_02135_, _02129_, _00748_);
  or _24377_ (_02136_, _02135_, _00779_);
  or _24378_ (_02137_, _02136_, _02134_);
  or _24379_ (_02138_, _02137_, _02133_);
  or _24380_ (_02139_, _02138_, _02131_);
  nor _24381_ (_02140_, _00746_, rst);
  and _24382_ (_02141_, _02140_, _00952_);
  and _24383_ (_01092_, _02141_, _02139_);
  nand _24384_ (_02142_, _00746_, _06811_);
  and _24385_ (_02143_, _00755_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and _24386_ (_02144_, _00779_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor _24387_ (_02145_, _00825_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  nor _24388_ (_02146_, _02145_, _00980_);
  and _24389_ (_02147_, _02146_, _00757_);
  nor _24390_ (_02148_, _02147_, _02144_);
  nor _24391_ (_02149_, _02148_, _00753_);
  or _24392_ (_02150_, _02149_, _02143_);
  or _24393_ (_02151_, _02150_, _00746_);
  and _24394_ (_02152_, _02151_, _05552_);
  and _24395_ (_01094_, _02152_, _02142_);
  and _24396_ (_02154_, _01967_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and _24397_ (_02155_, _02154_, _02076_);
  and _24398_ (_02156_, _01824_, _01812_);
  or _24399_ (_02157_, _02156_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and _24400_ (_02158_, _02157_, _02079_);
  or _24401_ (_02159_, _02158_, _01827_);
  or _24402_ (_02160_, _02159_, _02155_);
  nor _24403_ (_02161_, _01828_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  nor _24404_ (_02162_, _02161_, _01801_);
  and _24405_ (_02163_, _02162_, _02160_);
  and _24406_ (_02164_, _01801_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or _24407_ (_02166_, _02164_, _01802_);
  or _24408_ (_02167_, _02166_, _02163_);
  nand _24409_ (_02169_, _01802_, _08041_);
  and _24410_ (_02170_, _02169_, _05552_);
  and _24411_ (_01097_, _02170_, _02167_);
  and _24412_ (_02171_, _01967_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  and _24413_ (_02172_, _02171_, _02076_);
  and _24414_ (_02173_, _01824_, _01811_);
  nor _24415_ (_02174_, _02173_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  nor _24416_ (_02175_, _02174_, _02156_);
  or _24417_ (_02176_, _02175_, _01827_);
  or _24418_ (_02177_, _02176_, _02172_);
  nor _24419_ (_02178_, _01828_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  nor _24420_ (_02179_, _02178_, _01801_);
  and _24421_ (_02180_, _02179_, _02177_);
  and _24422_ (_02181_, _01801_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  or _24423_ (_02182_, _02181_, _01802_);
  or _24424_ (_02183_, _02182_, _02180_);
  nand _24425_ (_02184_, _01802_, _07975_);
  and _24426_ (_02185_, _02184_, _05552_);
  and _24427_ (_01103_, _02185_, _02183_);
  nor _24428_ (_01125_, _11139_, rst);
  or _24429_ (_02186_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  not _24430_ (_02187_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nand _24431_ (_02188_, pc_log_change, _02187_);
  and _24432_ (_02189_, _02188_, _05552_);
  and _24433_ (_01130_, _02189_, _02186_);
  or _24434_ (_02191_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nand _24435_ (_02192_, pc_log_change, _06085_);
  and _24436_ (_02193_, _02192_, _05552_);
  and _24437_ (_01135_, _02193_, _02191_);
  and _24438_ (_02194_, _01967_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  and _24439_ (_02195_, _02194_, _02076_);
  and _24440_ (_02196_, _01824_, _01810_);
  nor _24441_ (_02197_, _02196_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nor _24442_ (_02198_, _02197_, _02173_);
  or _24443_ (_02199_, _02198_, _01827_);
  or _24444_ (_02200_, _02199_, _02195_);
  nor _24445_ (_02201_, _01828_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  nor _24446_ (_02202_, _02201_, _01801_);
  and _24447_ (_02203_, _02202_, _02200_);
  and _24448_ (_02204_, _01801_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  or _24449_ (_02205_, _02204_, _01802_);
  or _24450_ (_02206_, _02205_, _02203_);
  nand _24451_ (_02207_, _01802_, _07945_);
  and _24452_ (_02208_, _02207_, _05552_);
  and _24453_ (_01143_, _02208_, _02206_);
  and _24454_ (_02209_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor _24455_ (_02210_, pc_log_change, _02187_);
  or _24456_ (_02211_, _02210_, _02209_);
  and _24457_ (_01150_, _02211_, _05552_);
  nor _24458_ (_02212_, _01997_, _08386_);
  and _24459_ (_02213_, _01967_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and _24460_ (_02214_, _02213_, _02076_);
  and _24461_ (_02215_, _01824_, _01808_);
  or _24462_ (_02216_, _02215_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  nand _24463_ (_02217_, _01824_, _01809_);
  and _24464_ (_02218_, _02217_, _02216_);
  or _24465_ (_02219_, _02218_, _01827_);
  or _24466_ (_02220_, _02219_, _02214_);
  nor _24467_ (_02221_, _01828_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  nor _24468_ (_02222_, _02221_, _01801_);
  and _24469_ (_02223_, _02222_, _02220_);
  or _24470_ (_02224_, _02223_, _01802_);
  or _24471_ (_02225_, _02224_, _02212_);
  or _24472_ (_02226_, _01978_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and _24473_ (_02227_, _02226_, _05552_);
  and _24474_ (_01169_, _02227_, _02225_);
  and _24475_ (_02228_, _01967_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and _24476_ (_02229_, _02228_, _02076_);
  and _24477_ (_02230_, _01824_, _01807_);
  nor _24478_ (_02231_, _02230_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  nor _24479_ (_02232_, _02231_, _02215_);
  or _24480_ (_02233_, _02232_, _01827_);
  or _24481_ (_02234_, _02233_, _02229_);
  nor _24482_ (_02235_, _01828_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  nor _24483_ (_02236_, _02235_, _01801_);
  and _24484_ (_02237_, _02236_, _02234_);
  and _24485_ (_02239_, _09018_, _06059_);
  and _24486_ (_02240_, _02239_, _10626_);
  and _24487_ (_02241_, _02240_, _06524_);
  not _24488_ (_02242_, _02241_);
  nor _24489_ (_02243_, _02242_, _06306_);
  or _24490_ (_02244_, _02243_, _02237_);
  or _24491_ (_02245_, _02244_, _01802_);
  or _24492_ (_02246_, _01978_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and _24493_ (_02247_, _02246_, _05552_);
  and _24494_ (_01182_, _02247_, _02245_);
  and _24495_ (_02248_, _01967_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and _24496_ (_02249_, _02248_, _02076_);
  nand _24497_ (_02250_, _01824_, _01804_);
  and _24498_ (_02251_, _02250_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  nor _24499_ (_02252_, _02250_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or _24500_ (_02254_, _02252_, _01827_);
  or _24501_ (_02256_, _02254_, _02251_);
  or _24502_ (_02257_, _02256_, _02249_);
  nor _24503_ (_02258_, _01828_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  nor _24504_ (_02259_, _02258_, _01801_);
  and _24505_ (_02260_, _02259_, _02257_);
  nor _24506_ (_02261_, _01997_, _08041_);
  or _24507_ (_02262_, _02261_, _01802_);
  or _24508_ (_02263_, _02262_, _02260_);
  or _24509_ (_02264_, _01978_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and _24510_ (_02265_, _02264_, _05552_);
  and _24511_ (_01201_, _02265_, _02263_);
  and _24512_ (_02266_, _01967_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and _24513_ (_02267_, _02266_, _02076_);
  and _24514_ (_02268_, _01824_, _01806_);
  nor _24515_ (_02269_, _02268_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  nor _24516_ (_02270_, _02269_, _02230_);
  or _24517_ (_02271_, _02270_, _01827_);
  or _24518_ (_02272_, _02271_, _02267_);
  nor _24519_ (_02273_, _01828_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  nor _24520_ (_02274_, _02273_, _01801_);
  and _24521_ (_02275_, _02274_, _02272_);
  nor _24522_ (_02276_, _02242_, _07388_);
  or _24523_ (_02277_, _02276_, _02275_);
  or _24524_ (_02278_, _02277_, _01802_);
  or _24525_ (_02279_, _01978_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and _24526_ (_02280_, _02279_, _05552_);
  and _24527_ (_01207_, _02280_, _02278_);
  and _24528_ (_02281_, _01967_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and _24529_ (_02282_, _02281_, _02076_);
  and _24530_ (_02283_, _01824_, _01805_);
  nor _24531_ (_02284_, _02283_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  nor _24532_ (_02285_, _02284_, _02268_);
  or _24533_ (_02287_, _02285_, _01827_);
  or _24534_ (_02288_, _02287_, _02282_);
  nor _24535_ (_02289_, _01828_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  nor _24536_ (_02290_, _02289_, _01801_);
  and _24537_ (_02291_, _02290_, _02288_);
  nor _24538_ (_02292_, _01997_, _06560_);
  or _24539_ (_02293_, _02292_, _01802_);
  or _24540_ (_02294_, _02293_, _02291_);
  or _24541_ (_02295_, _01978_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and _24542_ (_02296_, _02295_, _05552_);
  and _24543_ (_01211_, _02296_, _02294_);
  and _24544_ (_02297_, _01827_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and _24545_ (_02298_, _01824_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  or _24546_ (_02299_, _02298_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and _24547_ (_02300_, _02250_, _01828_);
  and _24548_ (_02301_, _02300_, _02299_);
  or _24549_ (_02302_, _02301_, _02297_);
  or _24550_ (_02303_, _02302_, _01801_);
  and _24551_ (_02304_, _01967_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and _24552_ (_02305_, _02304_, _01830_);
  or _24553_ (_02306_, _02305_, _02303_);
  nand _24554_ (_02307_, _01801_, _07975_);
  and _24555_ (_02308_, _02307_, _02306_);
  or _24556_ (_02309_, _02308_, _01802_);
  or _24557_ (_02310_, _01978_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and _24558_ (_02311_, _02310_, _05552_);
  and _24559_ (_01216_, _02311_, _02309_);
  or _24560_ (_02312_, _01824_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and _24561_ (_02313_, _01967_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  nand _24562_ (_02314_, _02313_, _01819_);
  nand _24563_ (_02315_, _02314_, _02298_);
  and _24564_ (_02316_, _02315_, _02312_);
  or _24565_ (_02317_, _02316_, _01827_);
  nor _24566_ (_02318_, _01828_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  nor _24567_ (_02319_, _02318_, _01801_);
  and _24568_ (_02320_, _02319_, _02317_);
  and _24569_ (_02321_, _01801_, _11238_);
  or _24570_ (_02322_, _02321_, _01802_);
  or _24571_ (_02323_, _02322_, _02320_);
  or _24572_ (_02324_, _01978_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and _24573_ (_02325_, _02324_, _05552_);
  and _24574_ (_01265_, _02325_, _02323_);
  or _24575_ (_02326_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  nand _24576_ (_02327_, _05550_, _05770_);
  and _24577_ (_02329_, _02327_, _05552_);
  and _24578_ (_01352_, _02329_, _02326_);
  not _24579_ (_02331_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  and _24580_ (_02332_, _00258_, _02331_);
  nor _24581_ (_02333_, _00258_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  or _24582_ (_02334_, _02333_, _00252_);
  or _24583_ (_02335_, _02334_, _02332_);
  nor _24584_ (_02336_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  nor _24585_ (_02337_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  nor _24586_ (_02338_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  nor _24587_ (_02339_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  and _24588_ (_02340_, _02339_, _02338_);
  and _24589_ (_02341_, _02340_, _02337_);
  nor _24590_ (_02342_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  and _24591_ (_02343_, _02342_, _00511_);
  and _24592_ (_02344_, _02343_, _02331_);
  and _24593_ (_02345_, _02344_, _02341_);
  nor _24594_ (_02346_, _02345_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  nor _24595_ (_02347_, _02346_, _02336_);
  nand _24596_ (_02348_, _02347_, _00252_);
  and _24597_ (_02349_, _02348_, _02335_);
  nor _24598_ (_02350_, _02349_, _00265_);
  and _24599_ (_02351_, _00248_, _11238_);
  or _24600_ (_02352_, _02351_, _02350_);
  and _24601_ (_01355_, _02352_, _05552_);
  nor _24602_ (_02354_, _10629_, _10643_);
  and _24603_ (_02355_, _02354_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  not _24604_ (_02356_, _02354_);
  and _24605_ (_02357_, _02356_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  or _24606_ (_02358_, _02357_, _02355_);
  or _24607_ (_02359_, _02358_, _10635_);
  nand _24608_ (_02360_, _10635_, _08041_);
  and _24609_ (_02361_, _02360_, _05552_);
  and _24610_ (_01363_, _02361_, _02359_);
  nand _24611_ (_02362_, _10635_, _08386_);
  and _24612_ (_02363_, _02356_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and _24613_ (_02364_, _02354_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or _24614_ (_02365_, _02364_, _02363_);
  or _24615_ (_02366_, _02365_, _10635_);
  and _24616_ (_02367_, _02366_, _05552_);
  and _24617_ (_01366_, _02367_, _02362_);
  nand _24618_ (_02368_, _10635_, _06306_);
  and _24619_ (_02369_, _02356_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and _24620_ (_02370_, _02354_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or _24621_ (_02371_, _02370_, _02369_);
  or _24622_ (_02372_, _02371_, _10635_);
  and _24623_ (_02373_, _02372_, _05552_);
  and _24624_ (_01387_, _02373_, _02368_);
  nand _24625_ (_02374_, _10635_, _07388_);
  and _24626_ (_02375_, _02354_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and _24627_ (_02377_, _02356_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  or _24628_ (_02379_, _02377_, _02375_);
  or _24629_ (_02380_, _02379_, _10635_);
  and _24630_ (_02381_, _02380_, _05552_);
  and _24631_ (_01391_, _02381_, _02374_);
  nand _24632_ (_02383_, _10635_, _06560_);
  or _24633_ (_02384_, _02354_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  nand _24634_ (_02385_, _02354_, _02078_);
  and _24635_ (_02386_, _02385_, _02384_);
  or _24636_ (_02387_, _02386_, _10635_);
  and _24637_ (_02388_, _02387_, _05552_);
  and _24638_ (_01395_, _02388_, _02383_);
  or _24639_ (_02389_, _02354_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  or _24640_ (_02390_, _02356_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and _24641_ (_02391_, _02390_, _02389_);
  or _24642_ (_02392_, _02391_, _10635_);
  nand _24643_ (_02393_, _10635_, _07975_);
  and _24644_ (_02394_, _02393_, _05552_);
  and _24645_ (_01403_, _02394_, _02392_);
  or _24646_ (_02395_, _02354_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  or _24647_ (_02396_, _02356_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and _24648_ (_02397_, _02396_, _02395_);
  or _24649_ (_02398_, _02397_, _10635_);
  nand _24650_ (_02399_, _10635_, _07945_);
  and _24651_ (_02400_, _02399_, _05552_);
  and _24652_ (_01421_, _02400_, _02398_);
  and _24653_ (_02401_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  not _24654_ (_02402_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _24655_ (_02403_, pc_log_change, _02402_);
  or _24656_ (_02404_, _02403_, _02401_);
  and _24657_ (_01437_, _02404_, _05552_);
  and _24658_ (_02405_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  not _24659_ (_02406_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor _24660_ (_02407_, pc_log_change, _02406_);
  or _24661_ (_02408_, _02407_, _02405_);
  and _24662_ (_01444_, _02408_, _05552_);
  and _24663_ (_02409_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  not _24664_ (_02410_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor _24665_ (_02411_, pc_log_change, _02410_);
  or _24666_ (_02412_, _02411_, _02409_);
  and _24667_ (_01447_, _02412_, _05552_);
  and _24668_ (_02414_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  not _24669_ (_02415_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  nor _24670_ (_02416_, pc_log_change, _02415_);
  or _24671_ (_02417_, _02416_, _02414_);
  and _24672_ (_01449_, _02417_, _05552_);
  and _24673_ (_02418_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor _24674_ (_02419_, pc_log_change, _02065_);
  or _24675_ (_02420_, _02419_, _02418_);
  and _24676_ (_01453_, _02420_, _05552_);
  or _24677_ (_02421_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nand _24678_ (_02422_, pc_log_change, _06219_);
  and _24679_ (_02423_, _02422_, _05552_);
  and _24680_ (_01459_, _02423_, _02421_);
  nand _24681_ (_02424_, _10629_, _08386_);
  and _24682_ (_02425_, _10643_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and _24683_ (_02426_, _10642_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  or _24684_ (_02427_, _02426_, _02425_);
  or _24685_ (_02428_, _02427_, _10629_);
  and _24686_ (_02429_, _02428_, _10636_);
  and _24687_ (_02430_, _02429_, _02424_);
  and _24688_ (_02431_, _10635_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  or _24689_ (_02432_, _02431_, _02430_);
  and _24690_ (_01480_, _02432_, _05552_);
  nand _24691_ (_02433_, _10629_, _06306_);
  and _24692_ (_02434_, _10643_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and _24693_ (_02436_, _10642_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or _24694_ (_02437_, _02436_, _02434_);
  or _24695_ (_02438_, _02437_, _10629_);
  and _24696_ (_02439_, _02438_, _10636_);
  and _24697_ (_02440_, _02439_, _02433_);
  and _24698_ (_02441_, _10635_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  or _24699_ (_02442_, _02441_, _02440_);
  and _24700_ (_01490_, _02442_, _05552_);
  and _24701_ (_02443_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor _24702_ (_02444_, pc_log_change, _01911_);
  or _24703_ (_02445_, _02444_, _02443_);
  and _24704_ (_01493_, _02445_, _05552_);
  nand _24705_ (_02446_, _10629_, _07388_);
  and _24706_ (_02447_, _10643_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and _24707_ (_02448_, _10642_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or _24708_ (_02449_, _02448_, _02447_);
  or _24709_ (_02451_, _02449_, _10629_);
  and _24710_ (_02452_, _02451_, _10636_);
  and _24711_ (_02453_, _02452_, _02446_);
  and _24712_ (_02454_, _10635_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  or _24713_ (_02455_, _02454_, _02453_);
  and _24714_ (_01539_, _02455_, _05552_);
  nand _24715_ (_02457_, _10629_, _06560_);
  and _24716_ (_02459_, _10643_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and _24717_ (_02460_, _10642_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or _24718_ (_02461_, _02460_, _02459_);
  or _24719_ (_02462_, _02461_, _10629_);
  and _24720_ (_02463_, _02462_, _10636_);
  and _24721_ (_02464_, _02463_, _02457_);
  and _24722_ (_02466_, _10635_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  or _24723_ (_02467_, _02466_, _02464_);
  and _24724_ (_01542_, _02467_, _05552_);
  nand _24725_ (_02469_, _10629_, _08041_);
  and _24726_ (_02470_, _10643_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and _24727_ (_02472_, _10642_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or _24728_ (_02473_, _02472_, _02470_);
  or _24729_ (_02475_, _02473_, _10629_);
  and _24730_ (_02476_, _02475_, _10636_);
  and _24731_ (_02477_, _02476_, _02469_);
  and _24732_ (_02478_, _10635_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  or _24733_ (_02479_, _02478_, _02477_);
  and _24734_ (_01545_, _02479_, _05552_);
  nand _24735_ (_02480_, _10629_, _07975_);
  or _24736_ (_02481_, _10642_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  or _24737_ (_02482_, _10643_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and _24738_ (_02483_, _02482_, _02481_);
  or _24739_ (_02484_, _02483_, _10629_);
  and _24740_ (_02485_, _02484_, _10636_);
  and _24741_ (_02486_, _02485_, _02480_);
  and _24742_ (_02487_, _10635_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  or _24743_ (_02488_, _02487_, _02486_);
  and _24744_ (_01547_, _02488_, _05552_);
  or _24745_ (_02489_, _10642_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  or _24746_ (_02490_, _10643_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and _24747_ (_02491_, _02490_, _02489_);
  or _24748_ (_02492_, _02491_, _10629_);
  nand _24749_ (_02493_, _10629_, _07945_);
  and _24750_ (_02494_, _02493_, _02492_);
  or _24751_ (_02495_, _02494_, _10635_);
  or _24752_ (_02496_, _10636_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  and _24753_ (_02497_, _02496_, _05552_);
  and _24754_ (_01549_, _02497_, _02495_);
  and _24755_ (_02499_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  not _24756_ (_02500_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nor _24757_ (_02501_, pc_log_change, _02500_);
  or _24758_ (_02502_, _02501_, _02499_);
  and _24759_ (_01566_, _02502_, _05552_);
  and _24760_ (_02504_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  not _24761_ (_02505_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _24762_ (_02506_, pc_log_change, _02505_);
  or _24763_ (_02507_, _02506_, _02504_);
  and _24764_ (_01569_, _02507_, _05552_);
  and _24765_ (_02508_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  and _24766_ (_02509_, _01956_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  or _24767_ (_02510_, _02509_, _02508_);
  and _24768_ (_01571_, _02510_, _05552_);
  and _24769_ (_02511_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  not _24770_ (_02512_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _24771_ (_02513_, pc_log_change, _02512_);
  or _24772_ (_02514_, _02513_, _02511_);
  and _24773_ (_01584_, _02514_, _05552_);
  and _24774_ (_02515_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  and _24775_ (_02516_, _01956_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  or _24776_ (_02517_, _02516_, _02515_);
  and _24777_ (_01587_, _02517_, _05552_);
  or _24778_ (_02518_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  nand _24779_ (_02520_, pc_log_change, _02415_);
  and _24780_ (_02521_, _02520_, _05552_);
  and _24781_ (_01593_, _02521_, _02518_);
  and _24782_ (_02522_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  not _24783_ (_02523_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  nor _24784_ (_02524_, pc_log_change, _02523_);
  or _24785_ (_02525_, _02524_, _02522_);
  and _24786_ (_01594_, _02525_, _05552_);
  and _24787_ (_02526_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  and _24788_ (_02527_, _01956_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  or _24789_ (_02528_, _02527_, _02526_);
  and _24790_ (_01596_, _02528_, _05552_);
  and _24791_ (_01630_, _13647_, _05552_);
  nor _24792_ (_02529_, _07388_, _06953_);
  and _24793_ (_02530_, _06953_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  or _24794_ (_02531_, _02530_, _06955_);
  or _24795_ (_02532_, _02531_, _02529_);
  or _24796_ (_02533_, _06068_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  and _24797_ (_02534_, _02533_, _05552_);
  and _24798_ (_01631_, _02534_, _02532_);
  and _24799_ (_01761_, _10981_, _05552_);
  and _24800_ (_02535_, _06691_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or _24801_ (_01664_, _02535_, _01761_);
  or _24802_ (_02538_, _05550_, \oc8051_top_1.oc8051_rom1.data_o [20]);
  nand _24803_ (_02539_, _05550_, _10995_);
  and _24804_ (_02541_, _02539_, _05552_);
  and _24805_ (_01666_, _02541_, _02538_);
  not _24806_ (_02542_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r );
  not _24807_ (_02543_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re );
  and _24808_ (_02544_, _02543_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  not _24809_ (_02546_, _02544_);
  nor _24810_ (_02547_, _05560_, _05556_);
  and _24811_ (_02548_, _02547_, _02546_);
  and _24812_ (_02549_, _02548_, _05593_);
  nor _24813_ (_02550_, _02549_, _02542_);
  and _24814_ (_02551_, _02549_, rxd_i);
  or _24815_ (_02552_, _02551_, rst);
  or _24816_ (_01680_, _02552_, _02550_);
  and _24817_ (_01686_, _12106_, _05552_);
  and _24818_ (_02553_, _05917_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  or _24819_ (_02554_, _02553_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  and _24820_ (_01713_, _02554_, _05552_);
  and _24821_ (_01737_, _07998_, _05552_);
  nand _24822_ (_02555_, _10635_, _06811_);
  and _24823_ (_02556_, _02356_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  and _24824_ (_02557_, _02354_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  or _24825_ (_02558_, _02557_, _02556_);
  or _24826_ (_02559_, _02558_, _10635_);
  and _24827_ (_02560_, _02559_, _05552_);
  and _24828_ (_01794_, _02560_, _02555_);
  and _24829_ (_02561_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor _24830_ (_02562_, _05550_, _05907_);
  or _24831_ (_02563_, _02562_, _02561_);
  and _24832_ (_01797_, _02563_, _05552_);
  and _24833_ (_02564_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor _24834_ (_02565_, _05550_, _06564_);
  or _24835_ (_02566_, _02565_, _02564_);
  and _24836_ (_01817_, _02566_, _05552_);
  and _24837_ (_01863_, t2ex_i, _05552_);
  nand _24838_ (_02567_, _05547_, _05605_);
  nand _24839_ (_02568_, _02567_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nand _24840_ (_02569_, _02568_, _05917_);
  and _24841_ (_01864_, _02569_, _05552_);
  and _24842_ (_02570_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _05552_);
  and _24843_ (_02572_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _05552_);
  and _24844_ (_02573_, _02572_, _05917_);
  or _24845_ (_01884_, _02573_, _02570_);
  nor _24846_ (_02574_, _05550_, _05548_);
  and _24847_ (_02575_, _00364_, _00361_);
  nor _24848_ (_02576_, _02575_, _05548_);
  and _24849_ (_02577_, _02576_, _05542_);
  nor _24850_ (_02578_, _02576_, _05542_);
  nor _24851_ (_02579_, _02578_, _02577_);
  nor _24852_ (_02580_, _02579_, _02574_);
  and _24853_ (_02581_, _05623_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and _24854_ (_02582_, _02581_, _02574_);
  and _24855_ (_02583_, _02582_, _07929_);
  or _24856_ (_02584_, _02583_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _24857_ (_02585_, _02584_, _02580_);
  and _24858_ (_01887_, _02585_, _05552_);
  and _24859_ (_02586_, _13744_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  and _24860_ (_02587_, _12264_, _11367_);
  or _24861_ (_02588_, _02587_, _02586_);
  and _24862_ (_01895_, _02588_, _05552_);
  nor _24863_ (_01899_, _11993_, rst);
  and _24864_ (_02589_, _11102_, _05552_);
  and _24865_ (_01918_, _02589_, _11774_);
  nand _24866_ (_02590_, _01717_, _06560_);
  or _24867_ (_02591_, _01717_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  and _24868_ (_02592_, _02591_, _05552_);
  and _24869_ (_01932_, _02592_, _02590_);
  nor _24870_ (_02593_, _09030_, _07388_);
  and _24871_ (_02594_, _09030_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  or _24872_ (_02595_, _02594_, _02593_);
  and _24873_ (_02010_, _02595_, _05552_);
  and _24874_ (_02596_, _09030_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  nor _24875_ (_02598_, _09030_, _06560_);
  or _24876_ (_02599_, _02598_, _02596_);
  and _24877_ (_02012_, _02599_, _05552_);
  nor _24878_ (_02600_, t2ex_i, rst);
  and _24879_ (_02074_, _02600_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r );
  nor _24880_ (_02089_, _11967_, rst);
  or _24881_ (_02601_, _12189_, _07668_);
  or _24882_ (_02602_, _07670_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and _24883_ (_02603_, _02602_, _05552_);
  and _24884_ (_02153_, _02603_, _02601_);
  and _24885_ (_02605_, _11367_, _06310_);
  or _24886_ (_02606_, _13739_, _06070_);
  and _24887_ (_02607_, _02606_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  or _24888_ (_02608_, _02607_, _02605_);
  and _24889_ (_02165_, _02608_, _05552_);
  and _24890_ (_02610_, _12189_, _07445_);
  and _24891_ (_02611_, _07486_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or _24892_ (_02613_, _02611_, _07485_);
  or _24893_ (_02614_, _02613_, _02610_);
  or _24894_ (_02615_, _12215_, _07579_);
  and _24895_ (_02616_, _02615_, _05552_);
  and _24896_ (_02168_, _02616_, _02614_);
  nor _24897_ (_02617_, _08386_, _06953_);
  and _24898_ (_02618_, _06953_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  or _24899_ (_02619_, _02618_, _06955_);
  or _24900_ (_02620_, _02619_, _02617_);
  or _24901_ (_02621_, _06068_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  and _24902_ (_02622_, _02621_, _05552_);
  and _24903_ (_02190_, _02622_, _02620_);
  and _24904_ (_02238_, _08982_, _05552_);
  not _24905_ (_02623_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _24906_ (_02624_, _02623_, \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and _24907_ (_02253_, _02624_, _05552_);
  and _24908_ (_02625_, _13744_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  and _24909_ (_02626_, _12264_, _11490_);
  or _24910_ (_02627_, _02626_, _02625_);
  and _24911_ (_02286_, _02627_, _05552_);
  nand _24912_ (_02628_, _01717_, _07388_);
  or _24913_ (_02629_, _01717_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  and _24914_ (_02630_, _02629_, _05552_);
  and _24915_ (_02330_, _02630_, _02628_);
  and _24916_ (_02631_, _01622_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  and _24917_ (_02632_, _06068_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  and _24918_ (_02633_, _02632_, _01625_);
  nor _24919_ (_02634_, _08041_, _07951_);
  or _24920_ (_02635_, _02634_, _02633_);
  or _24921_ (_02637_, _02635_, _02631_);
  and _24922_ (_02353_, _02637_, _05552_);
  nor _24923_ (_02376_, _11448_, rst);
  and _24924_ (_02638_, _05607_, _05545_);
  and _24925_ (_02639_, _02638_, _05884_);
  and _24926_ (_02640_, _07865_, _07784_);
  or _24927_ (_02641_, _02640_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and _24928_ (_02642_, _07788_, _05756_);
  and _24929_ (_02643_, _07898_, _02642_);
  not _24930_ (_02644_, _05733_);
  and _24931_ (_02645_, _07805_, _07788_);
  and _24932_ (_02646_, _07865_, _07810_);
  or _24933_ (_02647_, _02646_, _02645_);
  and _24934_ (_02648_, _02647_, _02644_);
  or _24935_ (_02649_, _02648_, _02643_);
  or _24936_ (_02650_, _02649_, _02641_);
  and _24937_ (_02651_, _02650_, _02639_);
  nor _24938_ (_02652_, _02638_, _05884_);
  or _24939_ (_02653_, _02652_, rst);
  or _24940_ (_02378_, _02653_, _02651_);
  nor _24941_ (_02382_, _11390_, rst);
  nand _24942_ (_02655_, _07945_, _06949_);
  or _24943_ (_02656_, _06949_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  and _24944_ (_02657_, _02656_, _02655_);
  and _24945_ (_02413_, _02657_, _05552_);
  nor _24946_ (_02658_, t2_i, rst);
  and _24947_ (_02435_, _02658_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r );
  and _24948_ (_02659_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and _24949_ (_02660_, _12140_, \oc8051_top_1.oc8051_rom1.data_o [29]);
  or _24950_ (_02661_, _02660_, _02659_);
  and _24951_ (_02450_, _02661_, _05552_);
  and _24952_ (_02456_, _13668_, _05552_);
  and _24953_ (_02458_, _13636_, _05552_);
  and _24954_ (_02662_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _05556_);
  and _24955_ (_02663_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _24956_ (_02664_, _02663_, _02662_);
  and _24957_ (_02465_, _02664_, _05552_);
  and _24958_ (_02665_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _05556_);
  and _24959_ (_02666_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _24960_ (_02667_, _02666_, _02665_);
  and _24961_ (_02468_, _02667_, _05552_);
  and _24962_ (_02669_, _11214_, _06310_);
  and _24963_ (_02670_, _06068_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  and _24964_ (_02671_, _02670_, _13739_);
  and _24965_ (_02672_, _06070_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  or _24966_ (_02673_, _02672_, _02671_);
  or _24967_ (_02674_, _02673_, _02669_);
  and _24968_ (_02471_, _02674_, _05552_);
  and _24969_ (_02675_, _05585_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  or _24970_ (_02474_, _02675_, _05591_);
  and _24971_ (_02498_, _02570_, _00580_);
  nand _24972_ (_02676_, _01717_, _08386_);
  or _24973_ (_02678_, _01717_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  and _24974_ (_02679_, _02678_, _05552_);
  and _24975_ (_02503_, _02679_, _02676_);
  nor _24976_ (_02519_, _08986_, rst);
  and _24977_ (_02680_, _06068_, _06058_);
  not _24978_ (_02681_, _02680_);
  and _24979_ (_02682_, _02681_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  and _24980_ (_02683_, _02680_, _11234_);
  or _24981_ (_02684_, _02683_, _02682_);
  and _24982_ (_02536_, _02684_, _05552_);
  and _24983_ (_02685_, _05917_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  or _24984_ (_02686_, _02685_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and _24985_ (_02537_, _02686_, _05552_);
  and _24986_ (_02687_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _05556_);
  and _24987_ (_02688_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _24988_ (_02689_, _02688_, _02687_);
  and _24989_ (_02540_, _02689_, _05552_);
  nand _24990_ (_02690_, _01717_, _06306_);
  or _24991_ (_02691_, _01717_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  and _24992_ (_02692_, _02691_, _05552_);
  and _24993_ (_02545_, _02692_, _02690_);
  or _24994_ (_02693_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  nand _24995_ (_02694_, _05550_, _05615_);
  and _24996_ (_02695_, _02694_, _05552_);
  and _24997_ (_02571_, _02695_, _02693_);
  and _24998_ (_02597_, _05669_, _05552_);
  and _24999_ (_02696_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  not _25000_ (_02697_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nor _25001_ (_02698_, pc_log_change, _02697_);
  or _25002_ (_02699_, _02698_, _02696_);
  and _25003_ (_02604_, _02699_, _05552_);
  nand _25004_ (_02700_, _01717_, _07975_);
  or _25005_ (_02701_, _01717_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  and _25006_ (_02702_, _02701_, _02700_);
  and _25007_ (_02609_, _02702_, _05552_);
  nand _25008_ (_02703_, _01717_, _08041_);
  or _25009_ (_02704_, _01717_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  and _25010_ (_02705_, _02704_, _05552_);
  and _25011_ (_02612_, _02705_, _02703_);
  nor _25012_ (_02707_, _00613_, _00580_);
  or _25013_ (_02709_, _02707_, _08998_);
  nand _25014_ (_02710_, _01234_, _00833_);
  and _25015_ (_02711_, _02710_, _05552_);
  and _25016_ (_02636_, _02711_, _02709_);
  and _25017_ (_02712_, _06055_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or _25018_ (_02713_, _02712_, _08015_);
  and _25019_ (_02714_, _02713_, _01515_);
  nand _25020_ (_02715_, _01515_, _01559_);
  and _25021_ (_02716_, _02715_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or _25022_ (_02717_, _02716_, _01520_);
  or _25023_ (_02718_, _02717_, _02714_);
  nand _25024_ (_02719_, _01520_, _08041_);
  and _25025_ (_02720_, _02719_, _05552_);
  and _25026_ (_02654_, _02720_, _02718_);
  or _25027_ (_02721_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or _25028_ (_02722_, _02721_, _00636_);
  not _25029_ (_02723_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  or _25030_ (_02724_, _00864_, _02723_);
  nand _25031_ (_02725_, _02724_, _00863_);
  or _25032_ (_02727_, _00644_, _08999_);
  and _25033_ (_02728_, _02727_, _02725_);
  or _25034_ (_02729_, _02728_, _00641_);
  or _25035_ (_02730_, _02721_, _01223_);
  and _25036_ (_02731_, _02730_, _01222_);
  and _25037_ (_02732_, _02731_, _02729_);
  and _25038_ (_02733_, _00639_, _08999_);
  or _25039_ (_02734_, _02733_, _00635_);
  or _25040_ (_02735_, _02734_, _02732_);
  and _25041_ (_02737_, _02735_, _02722_);
  or _25042_ (_02738_, _02737_, _00649_);
  or _25043_ (_02740_, _02721_, _00603_);
  or _25044_ (_02741_, _00846_, _02723_);
  nand _25045_ (_02742_, _02741_, _00845_);
  or _25046_ (_02743_, _00599_, _08999_);
  and _25047_ (_02744_, _02743_, _02742_);
  or _25048_ (_02745_, _02744_, _00609_);
  or _25049_ (_02746_, _02721_, _01204_);
  and _25050_ (_02747_, _02746_, _01203_);
  and _25051_ (_02748_, _02747_, _02745_);
  and _25052_ (_02749_, _00607_, _08999_);
  or _25053_ (_02750_, _02749_, _00602_);
  or _25054_ (_02751_, _02750_, _02748_);
  and _25055_ (_02752_, _02751_, _02740_);
  or _25056_ (_02753_, _02752_, _00857_);
  and _25057_ (_02754_, _02753_, _02738_);
  or _25058_ (_02755_, _02754_, _00580_);
  or _25059_ (_02756_, _01235_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  and _25060_ (_02757_, _02756_, _05552_);
  and _25061_ (_02668_, _02757_, _02755_);
  and _25062_ (_02758_, _00580_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  or _25063_ (_02759_, _02758_, _01235_);
  and _25064_ (_02677_, _02759_, _05552_);
  and _25065_ (_02706_, _08976_, _05552_);
  or _25066_ (_02760_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  nand _25067_ (_02761_, _05550_, _05791_);
  and _25068_ (_02762_, _02761_, _05552_);
  and _25069_ (_02708_, _02762_, _02760_);
  and _25070_ (_02763_, _00225_, _06771_);
  nand _25071_ (_02764_, _02763_, _06763_);
  or _25072_ (_02765_, _02763_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  and _25073_ (_02767_, _02765_, _00451_);
  and _25074_ (_02768_, _02767_, _02764_);
  nor _25075_ (_02769_, _00451_, _06811_);
  or _25076_ (_02770_, _02769_, _02768_);
  and _25077_ (_02726_, _02770_, _05552_);
  and _25078_ (_02771_, _02336_, _00257_);
  and _25079_ (_02772_, _02771_, _02343_);
  and _25080_ (_02773_, _02772_, _02341_);
  not _25081_ (_02774_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  nor _25082_ (_02775_, _00257_, _02774_);
  or _25083_ (_02776_, _02775_, _02773_);
  and _25084_ (_02777_, _02776_, _00254_);
  nand _25085_ (_02778_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  nor _25086_ (_02780_, _02778_, _00253_);
  nor _25087_ (_02781_, _02780_, _02777_);
  nor _25088_ (_02782_, _02781_, _00252_);
  and _25089_ (_02783_, _02345_, _00252_);
  or _25090_ (_02784_, _02783_, _02782_);
  and _25091_ (_02736_, _02784_, _00335_);
  not _25092_ (_02785_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  and _25093_ (_02786_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  not _25094_ (_02787_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and _25095_ (_02788_, _10874_, _02787_);
  or _25096_ (_02789_, _02788_, _12099_);
  nor _25097_ (_02790_, _02789_, _02786_);
  nand _25098_ (_02791_, _02790_, _02785_);
  nor _25099_ (_02792_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  nor _25100_ (_02793_, _02792_, _02790_);
  nand _25101_ (_02794_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  nand _25102_ (_02795_, _02794_, _02793_);
  and _25103_ (_02796_, _02795_, _05552_);
  and _25104_ (_02739_, _02796_, _02791_);
  or _25105_ (_02797_, _00333_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  nand _25106_ (_02798_, _00333_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  and _25107_ (_02799_, _02798_, _02797_);
  and _25108_ (_02766_, _02799_, _00335_);
  or _25109_ (_02800_, _02542_, rxd_i);
  nand _25110_ (_02801_, _02800_, _05574_);
  or _25111_ (_02802_, _05575_, _05561_);
  and _25112_ (_02803_, _02802_, _02801_);
  or _25113_ (_02804_, _05580_, _05572_);
  or _25114_ (_02806_, _02804_, _05562_);
  or _25115_ (_02807_, _02806_, _02803_);
  and _25116_ (_02779_, _02807_, _05585_);
  and _25117_ (_02808_, _01560_, _10632_);
  or _25118_ (_02809_, _02808_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and _25119_ (_02810_, _02809_, _01573_);
  nand _25120_ (_02811_, _02808_, _06763_);
  and _25121_ (_02812_, _02811_, _02810_);
  nor _25122_ (_02813_, _01573_, _06560_);
  or _25123_ (_02814_, _02813_, _02812_);
  and _25124_ (_02805_, _02814_, _05552_);
  and _25125_ (_02816_, _01515_, _06056_);
  nand _25126_ (_02817_, _02816_, _06763_);
  or _25127_ (_02819_, _02816_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and _25128_ (_02820_, _02819_, _01521_);
  and _25129_ (_02822_, _02820_, _02817_);
  nor _25130_ (_02823_, _01521_, _07975_);
  or _25131_ (_02824_, _02823_, _02822_);
  and _25132_ (_02815_, _02824_, _05552_);
  and _25133_ (_02825_, _13744_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  and _25134_ (_02826_, _12264_, _11726_);
  or _25135_ (_02827_, _02826_, _02825_);
  and _25136_ (_02818_, _02827_, _05552_);
  and _25137_ (_02828_, _01515_, _08365_);
  nand _25138_ (_02829_, _02828_, _06763_);
  or _25139_ (_02830_, _02828_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and _25140_ (_02832_, _02830_, _01521_);
  and _25141_ (_02833_, _02832_, _02829_);
  nor _25142_ (_02835_, _01521_, _08386_);
  or _25143_ (_02837_, _02835_, _02833_);
  and _25144_ (_02821_, _02837_, _05552_);
  and _25145_ (_02831_, _02793_, _05552_);
  or _25146_ (_02839_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and _25147_ (_02840_, _02839_, _05552_);
  or _25148_ (_02841_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0]);
  and _25149_ (_02842_, _02841_, _05568_);
  or _25150_ (_02843_, _02842_, _05582_);
  nand _25151_ (_02844_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0]);
  nor _25152_ (_02845_, _02844_, _05582_);
  or _25153_ (_02846_, _02845_, rxd_i);
  and _25154_ (_02847_, _02846_, _02843_);
  and _25155_ (_02848_, _01785_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  or _25156_ (_02849_, _02848_, _02847_);
  and _25157_ (_02834_, _02849_, _02840_);
  nand _25158_ (_02852_, _02773_, _00253_);
  nand _25159_ (_02854_, _02852_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  nor _25160_ (_02855_, _02854_, _02783_);
  or _25161_ (_02856_, _02855_, _00265_);
  and _25162_ (_02836_, _02856_, _05552_);
  or _25163_ (_02857_, _05803_, _08675_);
  or _25164_ (_02858_, _05546_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and _25165_ (_02859_, _02858_, _05552_);
  and _25166_ (_02838_, _02859_, _02857_);
  nand _25167_ (_02860_, _05756_, _05546_);
  or _25168_ (_02861_, _05546_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and _25169_ (_02862_, _02861_, _05552_);
  and _25170_ (_02850_, _02862_, _02860_);
  nand _25171_ (_02863_, _00241_, _06811_);
  or _25172_ (_02864_, _00241_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  and _25173_ (_02865_, _02864_, _05552_);
  and _25174_ (_02851_, _02865_, _02863_);
  and _25175_ (_02866_, _00259_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  and _25176_ (_02868_, _02866_, _00335_);
  and _25177_ (_02869_, _00246_, _05552_);
  and _25178_ (_02870_, _02869_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  or _25179_ (_02853_, _02870_, _02868_);
  nand _25180_ (_02871_, _00645_, _00621_);
  nor _25181_ (_02872_, _02871_, _00613_);
  and _25182_ (_02873_, _00580_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  or _25183_ (_02874_, _00598_, _00580_);
  nor _25184_ (_02875_, _02874_, _00586_);
  not _25185_ (_02876_, _00611_);
  nor _25186_ (_02877_, _02876_, _00596_);
  and _25187_ (_02878_, _02877_, _02875_);
  or _25188_ (_02879_, _02878_, _02873_);
  or _25189_ (_02880_, _02879_, _02872_);
  and _25190_ (_02867_, _02880_, _05552_);
  and _25191_ (_02881_, _10861_, _08057_);
  or _25192_ (_02882_, _02881_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and _25193_ (_02883_, _02882_, _08992_);
  nand _25194_ (_02884_, _02881_, _06763_);
  and _25195_ (_02885_, _02884_, _02883_);
  nor _25196_ (_02886_, _08992_, _07388_);
  or _25197_ (_02887_, _02886_, _02885_);
  and _25198_ (_02889_, _02887_, _05552_);
  and _25199_ (_02888_, _00260_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  and _25200_ (_02890_, _00259_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  or _25201_ (_02891_, _02890_, _02888_);
  and _25202_ (_02892_, _02891_, _00335_);
  nand _25203_ (_02893_, _06560_, _05560_);
  nand _25204_ (_02894_, _08041_, _05573_);
  and _25205_ (_02895_, _02894_, _02869_);
  and _25206_ (_02896_, _02895_, _02893_);
  or _25207_ (_03014_, _02896_, _02892_);
  and _25208_ (_02897_, _00260_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  and _25209_ (_02898_, _00259_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  or _25210_ (_02899_, _02898_, _02897_);
  and _25211_ (_02900_, _02899_, _00335_);
  nand _25212_ (_02901_, _08041_, _05560_);
  nand _25213_ (_02902_, _07975_, _05573_);
  and _25214_ (_02903_, _02902_, _02869_);
  and _25215_ (_02904_, _02903_, _02901_);
  or _25216_ (_03048_, _02904_, _02900_);
  and _25217_ (_02905_, _00260_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  and _25218_ (_02906_, _00259_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  or _25219_ (_02907_, _02906_, _02905_);
  and _25220_ (_02908_, _02907_, _00335_);
  or _25221_ (_02909_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3], _12098_);
  and _25222_ (_02910_, _02909_, _05552_);
  and _25223_ (_02911_, _02910_, _00267_);
  or _25224_ (_03075_, _02911_, _02908_);
  nand _25225_ (_02912_, _01802_, _06811_);
  or _25226_ (_02913_, _01964_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  nand _25227_ (_02914_, _01967_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  and _25228_ (_02915_, _02914_, _01824_);
  nand _25229_ (_02916_, _02915_, _01819_);
  and _25230_ (_02917_, _02916_, _02913_);
  or _25231_ (_02918_, _02917_, _01827_);
  nor _25232_ (_02919_, _01828_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  nor _25233_ (_02920_, _02919_, _01801_);
  and _25234_ (_02921_, _02920_, _02918_);
  nor _25235_ (_02922_, _01802_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  nor _25236_ (_02923_, _02922_, _01803_);
  or _25237_ (_02924_, _02923_, _02921_);
  and _25238_ (_02925_, _02924_, _05552_);
  and _25239_ (_03078_, _02925_, _02912_);
  and _25240_ (_02926_, _01519_, _06061_);
  nand _25241_ (_02927_, _02926_, _06763_);
  or _25242_ (_02928_, _02926_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and _25243_ (_02929_, _02928_, _06775_);
  and _25244_ (_02930_, _02929_, _02927_);
  and _25245_ (_02931_, _02926_, _11238_);
  nor _25246_ (_02932_, _02926_, _13607_);
  or _25247_ (_02933_, _02932_, _02931_);
  and _25248_ (_02934_, _02933_, _06524_);
  nor _25249_ (_02935_, _06774_, _13607_);
  or _25250_ (_02936_, _02935_, rst);
  or _25251_ (_02937_, _02936_, _02934_);
  or _25252_ (_03126_, _02937_, _02930_);
  and _25253_ (_02938_, _08365_, _06768_);
  nand _25254_ (_02939_, _02938_, _06763_);
  or _25255_ (_02940_, _02938_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and _25256_ (_02941_, _02940_, _06775_);
  and _25257_ (_02942_, _02941_, _02939_);
  nor _25258_ (_02943_, _08386_, _06782_);
  and _25259_ (_02944_, _06782_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or _25260_ (_02945_, _02944_, _02943_);
  and _25261_ (_02946_, _02945_, _06524_);
  and _25262_ (_02947_, _06816_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or _25263_ (_02948_, _02947_, rst);
  or _25264_ (_02949_, _02948_, _02946_);
  or _25265_ (_03128_, _02949_, _02942_);
  and _25266_ (_02950_, _06916_, _08013_);
  nand _25267_ (_02951_, _02950_, _06763_);
  or _25268_ (_02952_, _02950_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and _25269_ (_02953_, _02952_, _06775_);
  and _25270_ (_02954_, _02953_, _02951_);
  nand _25271_ (_02955_, _08041_, _06928_);
  or _25272_ (_02956_, _06928_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and _25273_ (_02957_, _02956_, _06524_);
  and _25274_ (_02958_, _02957_, _02955_);
  and _25275_ (_02959_, _06816_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  or _25276_ (_02960_, _02959_, rst);
  or _25277_ (_02961_, _02960_, _02958_);
  or _25278_ (_03132_, _02961_, _02954_);
  or _25279_ (_02962_, _06781_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and _25280_ (_02963_, _02962_, _06775_);
  nand _25281_ (_02964_, _06781_, _06763_);
  and _25282_ (_02965_, _02964_, _02963_);
  and _25283_ (_02966_, _11238_, _06781_);
  nor _25284_ (_02967_, _06781_, _13613_);
  or _25285_ (_02968_, _02967_, _02966_);
  and _25286_ (_02969_, _02968_, _06524_);
  nor _25287_ (_02970_, _06774_, _13613_);
  or _25288_ (_02971_, _02970_, rst);
  or _25289_ (_02972_, _02971_, _02969_);
  or _25290_ (_03134_, _02972_, _02965_);
  and _25291_ (_02973_, _06910_, _06767_);
  nand _25292_ (_02974_, _02973_, _06054_);
  and _25293_ (_02975_, _02974_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  nor _25294_ (_02976_, _01558_, _00021_);
  or _25295_ (_02977_, _02976_, _12129_);
  and _25296_ (_02978_, _02977_, _02973_);
  or _25297_ (_02979_, _02978_, _02975_);
  and _25298_ (_02980_, _02979_, _06775_);
  and _25299_ (_02981_, _07443_, _06061_);
  nand _25300_ (_02982_, _02981_, _06560_);
  or _25301_ (_02983_, _02981_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and _25302_ (_02984_, _02983_, _06524_);
  and _25303_ (_02985_, _02984_, _02982_);
  nor _25304_ (_02986_, _06774_, _00021_);
  or _25305_ (_02987_, _02986_, rst);
  or _25306_ (_02988_, _02987_, _02985_);
  or _25307_ (_03136_, _02988_, _02980_);
  or _25308_ (_02989_, _02981_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  and _25309_ (_02990_, _02989_, _06775_);
  nand _25310_ (_02991_, _02981_, _06763_);
  and _25311_ (_02992_, _02991_, _02990_);
  nand _25312_ (_02993_, _07945_, _02981_);
  and _25313_ (_02994_, _02989_, _06524_);
  and _25314_ (_02995_, _02994_, _02993_);
  nor _25315_ (_02996_, _06774_, _13594_);
  or _25316_ (_02997_, _02996_, rst);
  or _25317_ (_02998_, _02997_, _02995_);
  or _25318_ (_03138_, _02998_, _02992_);
  and _25319_ (_02999_, _00259_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  and _25320_ (_03000_, _00260_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  or _25321_ (_03001_, _03000_, _02999_);
  or _25322_ (_03002_, _03001_, _00265_);
  and _25323_ (_03003_, _03002_, _05552_);
  nand _25324_ (_03004_, _00267_, _06811_);
  and _25325_ (_03153_, _03004_, _03003_);
  and _25326_ (_03005_, _06915_, _06765_);
  and _25327_ (_03006_, _03005_, _08635_);
  nand _25328_ (_03007_, _03006_, _06763_);
  or _25329_ (_03008_, _03006_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and _25330_ (_03009_, _03008_, _06775_);
  and _25331_ (_03010_, _03009_, _03007_);
  not _25332_ (_03011_, _02926_);
  nor _25333_ (_03012_, _03011_, _06306_);
  and _25334_ (_03013_, _03011_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or _25335_ (_03015_, _03013_, _03012_);
  and _25336_ (_03016_, _03015_, _06524_);
  and _25337_ (_03017_, _06816_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or _25338_ (_03018_, _03017_, rst);
  or _25339_ (_03019_, _03018_, _03016_);
  or _25340_ (_03158_, _03019_, _03010_);
  and _25341_ (_03020_, _08635_, _06768_);
  nand _25342_ (_03021_, _03020_, _06763_);
  or _25343_ (_03022_, _03020_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and _25344_ (_03023_, _03022_, _06775_);
  and _25345_ (_03024_, _03023_, _03021_);
  nor _25346_ (_03025_, _06782_, _06306_);
  and _25347_ (_03026_, _06782_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or _25348_ (_03027_, _03026_, _03025_);
  and _25349_ (_03028_, _03027_, _06524_);
  and _25350_ (_03029_, _06816_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or _25351_ (_03030_, _03029_, rst);
  or _25352_ (_03031_, _03030_, _03028_);
  or _25353_ (_03160_, _03031_, _03024_);
  and _25354_ (_03032_, _06916_, _08365_);
  nand _25355_ (_03033_, _03032_, _06763_);
  or _25356_ (_03034_, _03032_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and _25357_ (_03035_, _03034_, _06775_);
  and _25358_ (_03036_, _03035_, _03033_);
  nand _25359_ (_03037_, _08386_, _06928_);
  or _25360_ (_03038_, _06928_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and _25361_ (_03039_, _03038_, _06524_);
  and _25362_ (_03040_, _03039_, _03037_);
  and _25363_ (_03041_, _06816_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  or _25364_ (_03042_, _03041_, rst);
  or _25365_ (_03043_, _03042_, _03040_);
  or _25366_ (_03162_, _03043_, _03036_);
  and _25367_ (_03044_, _06916_, _06056_);
  nand _25368_ (_03045_, _03044_, _06763_);
  or _25369_ (_03046_, _03044_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and _25370_ (_03047_, _03046_, _06775_);
  and _25371_ (_03049_, _03047_, _03045_);
  nand _25372_ (_03050_, _07975_, _06928_);
  or _25373_ (_03051_, _06928_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and _25374_ (_03052_, _03051_, _06524_);
  and _25375_ (_03053_, _03052_, _03050_);
  and _25376_ (_03054_, _06816_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  or _25377_ (_03055_, _03054_, rst);
  or _25378_ (_03056_, _03055_, _03053_);
  or _25379_ (_03164_, _03056_, _03049_);
  and _25380_ (_03057_, _06916_, _08057_);
  nand _25381_ (_03058_, _03057_, _06763_);
  or _25382_ (_03059_, _03057_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and _25383_ (_03060_, _03059_, _06775_);
  and _25384_ (_03061_, _03060_, _03058_);
  nand _25385_ (_03062_, _07388_, _06928_);
  or _25386_ (_03063_, _06928_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and _25387_ (_03064_, _03063_, _06524_);
  and _25388_ (_03065_, _03064_, _03062_);
  nor _25389_ (_03066_, _06774_, _13815_);
  or _25390_ (_03067_, _03066_, rst);
  or _25391_ (_03068_, _03067_, _03065_);
  or _25392_ (_03167_, _03068_, _03061_);
  nand _25393_ (_03069_, _02973_, _01559_);
  and _25394_ (_03070_, _03069_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and _25395_ (_03071_, _06055_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or _25396_ (_03072_, _03071_, _08015_);
  and _25397_ (_03073_, _03072_, _02973_);
  or _25398_ (_03074_, _03073_, _03070_);
  and _25399_ (_03076_, _03074_, _06775_);
  nand _25400_ (_03077_, _08041_, _02981_);
  or _25401_ (_03079_, _02981_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and _25402_ (_03080_, _03079_, _06524_);
  and _25403_ (_03081_, _03080_, _03077_);
  and _25404_ (_03082_, _06816_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or _25405_ (_03083_, _03082_, rst);
  or _25406_ (_03084_, _03083_, _03081_);
  or _25407_ (_03170_, _03084_, _03076_);
  and _25408_ (_03085_, _02973_, _08635_);
  nand _25409_ (_03086_, _03085_, _06763_);
  or _25410_ (_03087_, _03085_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and _25411_ (_03088_, _03087_, _06775_);
  and _25412_ (_03089_, _03088_, _03086_);
  nand _25413_ (_03090_, _02981_, _06306_);
  or _25414_ (_03091_, _02981_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and _25415_ (_03092_, _03091_, _06524_);
  and _25416_ (_03093_, _03092_, _03090_);
  and _25417_ (_03094_, _06816_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  or _25418_ (_03095_, _03094_, rst);
  or _25419_ (_03096_, _03095_, _03093_);
  or _25420_ (_03172_, _03096_, _03089_);
  and _25421_ (_03097_, _08057_, _06768_);
  nand _25422_ (_03098_, _03097_, _06763_);
  or _25423_ (_03099_, _03097_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and _25424_ (_03100_, _03099_, _06775_);
  and _25425_ (_03101_, _03100_, _03098_);
  nor _25426_ (_03102_, _07388_, _06782_);
  nor _25427_ (_03103_, _06781_, _13799_);
  or _25428_ (_03104_, _03103_, _03102_);
  and _25429_ (_03105_, _03104_, _06524_);
  nor _25430_ (_03106_, _06774_, _13799_);
  or _25431_ (_03107_, _03106_, rst);
  or _25432_ (_03108_, _03107_, _03105_);
  or _25433_ (_03256_, _03108_, _03101_);
  and _25434_ (_03109_, _10632_, _06768_);
  nand _25435_ (_03110_, _03109_, _06763_);
  or _25436_ (_03111_, _03109_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and _25437_ (_03112_, _03111_, _06775_);
  and _25438_ (_03113_, _03112_, _03110_);
  nor _25439_ (_03114_, _06782_, _06560_);
  nor _25440_ (_03115_, _06781_, _00038_);
  or _25441_ (_03116_, _03115_, _03114_);
  and _25442_ (_03117_, _03116_, _06524_);
  nor _25443_ (_03118_, _06774_, _00038_);
  or _25444_ (_03119_, _03118_, rst);
  or _25445_ (_03120_, _03119_, _03117_);
  or _25446_ (_03257_, _03120_, _03113_);
  nor _25447_ (_03121_, _09030_, _08041_);
  and _25448_ (_03122_, _09030_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  or _25449_ (_03123_, _03122_, _03121_);
  and _25450_ (_03270_, _03123_, _05552_);
  and _25451_ (_03124_, _08013_, _06768_);
  nand _25452_ (_03125_, _03124_, _06763_);
  or _25453_ (_03127_, _03124_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and _25454_ (_03129_, _03127_, _06775_);
  and _25455_ (_03130_, _03129_, _03125_);
  nor _25456_ (_03131_, _08041_, _06782_);
  and _25457_ (_03133_, _06782_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or _25458_ (_03135_, _03133_, _03131_);
  and _25459_ (_03137_, _03135_, _06524_);
  and _25460_ (_03139_, _06816_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or _25461_ (_03140_, _03139_, rst);
  or _25462_ (_03141_, _03140_, _03137_);
  or _25463_ (_03281_, _03141_, _03130_);
  and _25464_ (_03142_, _06916_, _06060_);
  nand _25465_ (_03143_, _03142_, _06763_);
  or _25466_ (_03144_, _06928_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and _25467_ (_03145_, _03144_, _06775_);
  and _25468_ (_03146_, _03145_, _03143_);
  nand _25469_ (_03147_, _07945_, _06928_);
  and _25470_ (_03148_, _03147_, _06524_);
  and _25471_ (_03149_, _03148_, _03144_);
  nor _25472_ (_03150_, _06774_, _13600_);
  or _25473_ (_03151_, _03150_, rst);
  or _25474_ (_03152_, _03151_, _03149_);
  or _25475_ (_03283_, _03152_, _03146_);
  and _25476_ (_03154_, _03005_, _10632_);
  nand _25477_ (_03155_, _03154_, _06763_);
  or _25478_ (_03156_, _03154_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and _25479_ (_03157_, _03156_, _06775_);
  and _25480_ (_03159_, _03157_, _03155_);
  nor _25481_ (_03161_, _03011_, _06560_);
  nor _25482_ (_03163_, _02926_, _00033_);
  or _25483_ (_03165_, _03163_, _03161_);
  and _25484_ (_03166_, _03165_, _06524_);
  nor _25485_ (_03168_, _06774_, _00033_);
  or _25486_ (_03169_, _03168_, rst);
  or _25487_ (_03171_, _03169_, _03166_);
  or _25488_ (_03286_, _03171_, _03159_);
  and _25489_ (_03173_, _03005_, _08013_);
  nand _25490_ (_03174_, _03173_, _06763_);
  or _25491_ (_03175_, _03173_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and _25492_ (_03176_, _03175_, _06775_);
  and _25493_ (_03177_, _03176_, _03174_);
  nor _25494_ (_03178_, _03011_, _08041_);
  and _25495_ (_03179_, _03011_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or _25496_ (_03180_, _03179_, _03178_);
  and _25497_ (_03181_, _03180_, _06524_);
  and _25498_ (_03182_, _06816_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or _25499_ (_03183_, _03182_, rst);
  or _25500_ (_03184_, _03183_, _03181_);
  or _25501_ (_03287_, _03184_, _03177_);
  nand _25502_ (_03185_, _11223_, _06763_);
  or _25503_ (_03186_, _11223_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and _25504_ (_03187_, _03186_, _06775_);
  and _25505_ (_03188_, _03187_, _03185_);
  nand _25506_ (_03189_, _07975_, _02981_);
  or _25507_ (_03190_, _02981_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and _25508_ (_03191_, _03190_, _06524_);
  and _25509_ (_03192_, _03191_, _03189_);
  and _25510_ (_03193_, _06816_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  or _25511_ (_03194_, _03193_, rst);
  or _25512_ (_03195_, _03194_, _03192_);
  or _25513_ (_03305_, _03195_, _03188_);
  and _25514_ (_03196_, _02973_, _08365_);
  nand _25515_ (_03197_, _03196_, _06763_);
  or _25516_ (_03198_, _03196_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and _25517_ (_03199_, _03198_, _06775_);
  and _25518_ (_03200_, _03199_, _03197_);
  nand _25519_ (_03201_, _08386_, _02981_);
  or _25520_ (_03202_, _02981_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and _25521_ (_03203_, _03202_, _06524_);
  and _25522_ (_03204_, _03203_, _03201_);
  and _25523_ (_03205_, _06816_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  or _25524_ (_03206_, _03205_, rst);
  or _25525_ (_03207_, _03206_, _03204_);
  or _25526_ (_03307_, _03207_, _03200_);
  and _25527_ (_03208_, _02973_, _08057_);
  nand _25528_ (_03209_, _03208_, _06763_);
  or _25529_ (_03210_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and _25530_ (_03211_, _03210_, _06775_);
  and _25531_ (_03212_, _03211_, _03209_);
  nand _25532_ (_03213_, _07388_, _02981_);
  or _25533_ (_03214_, _02981_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and _25534_ (_03215_, _03214_, _06524_);
  and _25535_ (_03216_, _03215_, _03213_);
  nor _25536_ (_03217_, _06774_, _13810_);
  or _25537_ (_03218_, _03217_, rst);
  or _25538_ (_03219_, _03218_, _03216_);
  or _25539_ (_03309_, _03219_, _03212_);
  nand _25540_ (_03220_, _06768_, _06056_);
  nand _25541_ (_03221_, _03220_, _00173_);
  and _25542_ (_03222_, _03221_, _06775_);
  or _25543_ (_03223_, _03220_, _08048_);
  and _25544_ (_03224_, _03223_, _03222_);
  nor _25545_ (_03225_, _07975_, _06782_);
  nor _25546_ (_03226_, _06781_, _00173_);
  or _25547_ (_03227_, _03226_, _03225_);
  and _25548_ (_03228_, _03227_, _06524_);
  nor _25549_ (_03229_, _06774_, _00173_);
  or _25550_ (_03230_, _03229_, rst);
  or _25551_ (_03231_, _03230_, _03228_);
  or _25552_ (_03311_, _03231_, _03224_);
  and _25553_ (_03232_, _06916_, _08635_);
  nand _25554_ (_03233_, _03232_, _06763_);
  or _25555_ (_03234_, _03232_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and _25556_ (_03235_, _03234_, _06775_);
  and _25557_ (_03236_, _03235_, _03233_);
  nand _25558_ (_03237_, _06928_, _06306_);
  or _25559_ (_03238_, _06928_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and _25560_ (_03239_, _03238_, _06524_);
  and _25561_ (_03240_, _03239_, _03237_);
  and _25562_ (_03241_, _06816_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  or _25563_ (_03242_, _03241_, rst);
  or _25564_ (_03243_, _03242_, _03240_);
  or _25565_ (_03312_, _03243_, _03236_);
  and _25566_ (_03244_, _06916_, _10632_);
  nand _25567_ (_03245_, _03244_, _06763_);
  or _25568_ (_03246_, _03244_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and _25569_ (_03247_, _03246_, _06775_);
  and _25570_ (_03248_, _03247_, _03245_);
  nand _25571_ (_03249_, _06928_, _06560_);
  or _25572_ (_03250_, _06928_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and _25573_ (_03251_, _03250_, _06524_);
  and _25574_ (_03252_, _03251_, _03249_);
  nor _25575_ (_03253_, _06774_, _00027_);
  or _25576_ (_03254_, _03253_, rst);
  or _25577_ (_03255_, _03254_, _03252_);
  or _25578_ (_03314_, _03255_, _03248_);
  and _25579_ (_03258_, _03005_, _06056_);
  nand _25580_ (_03259_, _03258_, _06763_);
  or _25581_ (_03260_, _03258_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and _25582_ (_03261_, _03260_, _06775_);
  and _25583_ (_03262_, _03261_, _03259_);
  nor _25584_ (_03263_, _03011_, _07975_);
  and _25585_ (_03264_, _03011_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or _25586_ (_03265_, _03264_, _03263_);
  and _25587_ (_03266_, _03265_, _06524_);
  and _25588_ (_03267_, _06816_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or _25589_ (_03268_, _03267_, rst);
  or _25590_ (_03269_, _03268_, _03266_);
  or _25591_ (_03317_, _03269_, _03262_);
  and _25592_ (_03271_, _03005_, _08365_);
  nand _25593_ (_03272_, _03271_, _06763_);
  or _25594_ (_03273_, _03271_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and _25595_ (_03274_, _03273_, _06775_);
  and _25596_ (_03275_, _03274_, _03272_);
  nor _25597_ (_03277_, _03011_, _08386_);
  and _25598_ (_03278_, _03011_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or _25599_ (_03279_, _03278_, _03277_);
  and _25600_ (_03280_, _03279_, _06524_);
  and _25601_ (_03282_, _06816_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or _25602_ (_03284_, _03282_, rst);
  or _25603_ (_03285_, _03284_, _03280_);
  or _25604_ (_03320_, _03285_, _03275_);
  and _25605_ (_03288_, _03005_, _08057_);
  nand _25606_ (_03289_, _03288_, _06763_);
  or _25607_ (_03290_, _03288_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and _25608_ (_03291_, _03290_, _06775_);
  and _25609_ (_03292_, _03291_, _03289_);
  nor _25610_ (_03293_, _03011_, _07388_);
  nor _25611_ (_03294_, _02926_, _13804_);
  or _25612_ (_03295_, _03294_, _03293_);
  and _25613_ (_03296_, _03295_, _06524_);
  nor _25614_ (_03297_, _06774_, _13804_);
  or _25615_ (_03298_, _03297_, rst);
  or _25616_ (_03299_, _03298_, _03296_);
  or _25617_ (_03322_, _03299_, _03292_);
  nand _25618_ (_03300_, _01717_, _06811_);
  or _25619_ (_03301_, _01717_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  and _25620_ (_03302_, _03301_, _05552_);
  and _25621_ (_03324_, _03302_, _03300_);
  not _25622_ (_03303_, _00833_);
  or _25623_ (_03304_, _03303_, _00652_);
  and _25624_ (_03306_, _00833_, _00629_);
  or _25625_ (_03308_, _03306_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  and _25626_ (_03310_, _03308_, _05552_);
  and _25627_ (_03329_, _03310_, _03304_);
  nor _25628_ (_03313_, _06811_, _06953_);
  and _25629_ (_03315_, _06953_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  or _25630_ (_03316_, _03315_, _06955_);
  or _25631_ (_03318_, _03316_, _03313_);
  or _25632_ (_03319_, _06068_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  and _25633_ (_03321_, _03319_, _05552_);
  and _25634_ (_03332_, _03321_, _03318_);
  or _25635_ (_03323_, _05586_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  or _25636_ (_03325_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _25637_ (_03326_, _03325_, _05560_);
  or _25638_ (_03327_, _03326_, _05562_);
  nand _25639_ (_03328_, _03327_, _03323_);
  nand _25640_ (_03346_, _03328_, _05585_);
  or _25641_ (_03330_, _05710_, _08675_);
  or _25642_ (_03331_, _05546_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and _25643_ (_03333_, _03331_, _05552_);
  and _25644_ (_03347_, _03333_, _03330_);
  and _25645_ (_03334_, _07485_, _07360_);
  or _25646_ (_03335_, _07445_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  and _25647_ (_03336_, _03335_, _07579_);
  or _25648_ (_03337_, _07486_, _07255_);
  and _25649_ (_03338_, _03337_, _03336_);
  or _25650_ (_03339_, _03338_, _03334_);
  and _25651_ (_03398_, _03339_, _05552_);
  or _25652_ (_03340_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  nand _25653_ (_03341_, _05550_, _05768_);
  and _25654_ (_03342_, _03341_, _05552_);
  and _25655_ (_03415_, _03342_, _03340_);
  nor _25656_ (_03424_, _11327_, rst);
  and _25657_ (_03343_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and _25658_ (_03344_, _12140_, \oc8051_top_1.oc8051_rom1.data_o [31]);
  or _25659_ (_03345_, _03344_, _03343_);
  and _25660_ (_03428_, _03345_, _05552_);
  nor _25661_ (_03433_, _11370_, rst);
  nor _25662_ (_03436_, _11418_, rst);
  nor _25663_ (_03439_, _11492_, rst);
  nor _25664_ (_03441_, _11217_, rst);
  nand _25665_ (_03348_, _06949_, _06811_);
  or _25666_ (_03349_, _06949_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  and _25667_ (_03350_, _03349_, _05552_);
  and _25668_ (_03446_, _03350_, _03348_);
  or _25669_ (_03351_, _05550_, \oc8051_top_1.oc8051_rom1.data_o [0]);
  nand _25670_ (_03352_, _05550_, _05656_);
  and _25671_ (_03353_, _03352_, _05552_);
  and _25672_ (_03454_, _03353_, _03351_);
  nor _25673_ (_03467_, _11848_, rst);
  nor _25674_ (_03354_, _01997_, _06811_);
  and _25675_ (_03355_, _01967_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and _25676_ (_03356_, _03355_, _02076_);
  not _25677_ (_03357_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and _25678_ (_03358_, _02217_, _03357_);
  nor _25679_ (_03359_, _03358_, _02196_);
  or _25680_ (_03360_, _03359_, _01827_);
  or _25681_ (_03361_, _03360_, _03356_);
  nor _25682_ (_03362_, _01828_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  nor _25683_ (_03363_, _03362_, _01801_);
  and _25684_ (_03364_, _03363_, _03361_);
  or _25685_ (_03365_, _03364_, _01802_);
  or _25686_ (_03366_, _03365_, _03354_);
  nand _25687_ (_03367_, _01802_, _03357_);
  and _25688_ (_03368_, _03367_, _05552_);
  and _25689_ (_03493_, _03368_, _03366_);
  and _25690_ (_03495_, t2_i, _05552_);
  nand _25691_ (_03369_, _00241_, _07975_);
  or _25692_ (_03370_, _00241_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  and _25693_ (_03371_, _03370_, _05552_);
  and _25694_ (_03522_, _03371_, _03369_);
  and _25695_ (_03372_, _13499_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  and _25696_ (_03373_, _13502_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  or _25697_ (_03374_, _03373_, _03372_);
  and _25698_ (_03375_, _13494_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and _25699_ (_03376_, _13488_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or _25700_ (_03377_, _03376_, _03375_);
  or _25701_ (_03378_, _03377_, _03374_);
  and _25702_ (_03379_, _13507_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and _25703_ (_03380_, _13511_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  or _25704_ (_03381_, _03380_, _03379_);
  and _25705_ (_03382_, _13516_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and _25706_ (_03383_, _13521_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  or _25707_ (_03384_, _03383_, _03382_);
  or _25708_ (_03385_, _03384_, _03381_);
  or _25709_ (_03386_, _03385_, _03378_);
  nor _25710_ (_03387_, _13528_, _00760_);
  and _25711_ (_03388_, _13531_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  or _25712_ (_03389_, _03388_, _03387_);
  and _25713_ (_03390_, _13534_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and _25714_ (_03391_, _13536_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  or _25715_ (_03392_, _03391_, _03390_);
  or _25716_ (_03393_, _03392_, _03389_);
  and _25717_ (_03394_, _13541_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  and _25718_ (_03395_, _13544_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  or _25719_ (_03396_, _03395_, _03394_);
  and _25720_ (_03397_, _13547_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and _25721_ (_03399_, _13549_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  or _25722_ (_03400_, _03399_, _03397_);
  or _25723_ (_03401_, _03400_, _03396_);
  or _25724_ (_03402_, _03401_, _03393_);
  or _25725_ (_03403_, _03402_, _03386_);
  and _25726_ (_03404_, _13555_, _11345_);
  and _25727_ (_03405_, _13562_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  or _25728_ (_03406_, _03405_, _03404_);
  and _25729_ (_03407_, _13475_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and _25730_ (_03408_, _13568_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or _25731_ (_03409_, _03408_, _03407_);
  or _25732_ (_03410_, _03409_, _03406_);
  or _25733_ (_03411_, _13592_, p0_in[6]);
  or _25734_ (_03412_, _00099_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and _25735_ (_03413_, _03412_, _03411_);
  and _25736_ (_03414_, _03413_, _13574_);
  or _25737_ (_03416_, _13592_, p1_in[6]);
  or _25738_ (_03417_, _00099_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and _25739_ (_03418_, _03417_, _03416_);
  and _25740_ (_03419_, _03418_, _13598_);
  or _25741_ (_03420_, _03419_, _03414_);
  or _25742_ (_03421_, _13592_, p3_in[6]);
  or _25743_ (_03422_, _00099_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and _25744_ (_03423_, _03422_, _03421_);
  and _25745_ (_03425_, _03423_, _13605_);
  or _25746_ (_03426_, _13592_, p2_in[6]);
  or _25747_ (_03427_, _00099_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and _25748_ (_03429_, _03427_, _03426_);
  and _25749_ (_03430_, _03429_, _13611_);
  or _25750_ (_03431_, _03430_, _03425_);
  or _25751_ (_03432_, _03431_, _03420_);
  or _25752_ (_03434_, _03432_, _03410_);
  and _25753_ (_03435_, _13622_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and _25754_ (_03437_, _13681_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or _25755_ (_03438_, _03437_, _03435_);
  or _25756_ (_03440_, _03438_, _03434_);
  or _25757_ (_03442_, _03440_, _03403_);
  and _25758_ (_03443_, _03442_, _13701_);
  and _25759_ (_03444_, _13735_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  or _25760_ (_03445_, _03444_, _13476_);
  or _25761_ (_03447_, _03445_, _03443_);
  or _25762_ (_03448_, _13704_, _07574_);
  and _25763_ (_03449_, _03448_, _05552_);
  and _25764_ (_03526_, _03449_, _03447_);
  and _25765_ (_03450_, _05894_, _10917_);
  or _25766_ (_03451_, _13578_, _10937_);
  or _25767_ (_03452_, _03451_, _03450_);
  or _25768_ (_03453_, _03452_, _10901_);
  or _25769_ (_03455_, _03453_, _10934_);
  or _25770_ (_03456_, _11149_, _10913_);
  or _25771_ (_03457_, _03456_, _10941_);
  or _25772_ (_03458_, _11115_, _11088_);
  or _25773_ (_03459_, _03458_, _03457_);
  or _25774_ (_03460_, _11022_, _10943_);
  or _25775_ (_03461_, _11178_, _11015_);
  or _25776_ (_03462_, _03461_, _03460_);
  and _25777_ (_03463_, _12283_, _05837_);
  or _25778_ (_03464_, _03463_, _13575_);
  or _25779_ (_03465_, _03464_, _10929_);
  or _25780_ (_03466_, _03465_, _10908_);
  or _25781_ (_03468_, _03466_, _03462_);
  or _25782_ (_03469_, _03468_, _03459_);
  or _25783_ (_03470_, _03469_, _03455_);
  and _25784_ (_03471_, _03470_, _05547_);
  and _25785_ (_03472_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _25786_ (_03473_, _03472_, _10956_);
  or _25787_ (_03474_, _03473_, _03471_);
  and _25788_ (_03548_, _03474_, _05552_);
  or _25789_ (_03475_, _12332_, _12329_);
  or _25790_ (_03476_, _10933_, _05842_);
  or _25791_ (_03477_, _03476_, _13392_);
  or _25792_ (_03478_, _03477_, _03475_);
  or _25793_ (_03479_, _10851_, _05878_);
  and _25794_ (_03480_, _10929_, _05737_);
  or _25795_ (_03481_, _03480_, _12271_);
  or _25796_ (_03482_, _03481_, _03479_);
  or _25797_ (_03483_, _12308_, _05845_);
  nor _25798_ (_03484_, _03483_, _11022_);
  nand _25799_ (_03485_, _03484_, _12315_);
  or _25800_ (_03486_, _03485_, _03482_);
  or _25801_ (_03487_, _03486_, _12325_);
  or _25802_ (_03488_, _03487_, _03478_);
  and _25803_ (_03489_, _03488_, _05547_);
  and _25804_ (_03490_, \oc8051_top_1.oc8051_decoder1.alu_op [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _25805_ (_03491_, _03490_, _10958_);
  or _25806_ (_03492_, _03491_, _03489_);
  and _25807_ (_03558_, _03492_, _05552_);
  nor _25808_ (_03494_, _09030_, _08386_);
  and _25809_ (_03496_, _09030_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  or _25810_ (_03497_, _03496_, _03494_);
  and _25811_ (_03566_, _03497_, _05552_);
  or _25812_ (_03498_, _01751_, _07483_);
  not _25813_ (_03499_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nand _25814_ (_03500_, _01751_, _03499_);
  and _25815_ (_03501_, _03500_, _06524_);
  and _25816_ (_03502_, _03501_, _03498_);
  nor _25817_ (_03503_, _06774_, _03499_);
  and _25818_ (_03504_, _01750_, _10632_);
  nand _25819_ (_03505_, _03504_, _06763_);
  or _25820_ (_03506_, _03504_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and _25821_ (_03507_, _03506_, _06775_);
  and _25822_ (_03508_, _03507_, _03505_);
  or _25823_ (_03509_, _03508_, _03503_);
  or _25824_ (_03510_, _03509_, _03502_);
  and _25825_ (_03593_, _03510_, _05552_);
  or _25826_ (_03511_, _05689_, _08675_);
  or _25827_ (_03512_, _05546_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and _25828_ (_03513_, _03512_, _05552_);
  and _25829_ (_03600_, _03513_, _03511_);
  or _25830_ (_03514_, _01751_, _07711_);
  not _25831_ (_03515_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nand _25832_ (_03516_, _01751_, _03515_);
  and _25833_ (_03517_, _03516_, _06524_);
  and _25834_ (_03518_, _03517_, _03514_);
  nor _25835_ (_03519_, _06774_, _03515_);
  or _25836_ (_03520_, _01751_, _08048_);
  and _25837_ (_03521_, _03516_, _06775_);
  and _25838_ (_03523_, _03521_, _03520_);
  or _25839_ (_03524_, _03523_, _03519_);
  or _25840_ (_03525_, _03524_, _03518_);
  and _25841_ (_03603_, _03525_, _05552_);
  or _25842_ (_03527_, _06314_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _25843_ (_03528_, _06315_, rst);
  and _25844_ (_03614_, _03528_, _03527_);
  and _25845_ (_03529_, _02973_, _06771_);
  nand _25846_ (_03530_, _03529_, _06763_);
  or _25847_ (_03531_, _03529_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and _25848_ (_03532_, _03531_, _06775_);
  and _25849_ (_03533_, _03532_, _03530_);
  nand _25850_ (_03534_, _02981_, _06811_);
  or _25851_ (_03535_, _02981_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and _25852_ (_03536_, _03535_, _06524_);
  and _25853_ (_03537_, _03536_, _03534_);
  and _25854_ (_03538_, _06816_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  or _25855_ (_03539_, _03538_, rst);
  or _25856_ (_03540_, _03539_, _03537_);
  or _25857_ (_03623_, _03540_, _03533_);
  and _25858_ (_03541_, _07951_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  nor _25859_ (_03542_, _08386_, _07951_);
  or _25860_ (_03543_, _03542_, _03541_);
  and _25861_ (_03636_, _03543_, _05552_);
  or _25862_ (_03544_, _01751_, _07574_);
  not _25863_ (_03545_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  nand _25864_ (_03546_, _01751_, _03545_);
  and _25865_ (_03547_, _03546_, _06524_);
  and _25866_ (_03549_, _03547_, _03544_);
  nor _25867_ (_03550_, _06774_, _03545_);
  and _25868_ (_03551_, _01750_, _08365_);
  nand _25869_ (_03552_, _03551_, _06763_);
  or _25870_ (_03553_, _03551_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and _25871_ (_03554_, _03553_, _06775_);
  and _25872_ (_03555_, _03554_, _03552_);
  or _25873_ (_03556_, _03555_, _03550_);
  or _25874_ (_03557_, _03556_, _03549_);
  and _25875_ (_03638_, _03557_, _05552_);
  and _25876_ (_03651_, _11308_, _05552_);
  and _25877_ (_03559_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], _07768_);
  and _25878_ (_03560_, \oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or _25879_ (_03561_, _03560_, _03559_);
  and _25880_ (_03660_, _03561_, _05552_);
  and _25881_ (_03562_, _07635_, _05552_);
  or _25882_ (_03563_, _03562_, _13477_);
  and _25883_ (_03564_, _13494_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and _25884_ (_03565_, _13488_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  or _25885_ (_03567_, _03565_, _03564_);
  and _25886_ (_03568_, _13502_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and _25887_ (_03569_, _13499_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or _25888_ (_03570_, _03569_, _03568_);
  or _25889_ (_03571_, _03570_, _03567_);
  and _25890_ (_03572_, _13507_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and _25891_ (_03573_, _13511_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  or _25892_ (_03574_, _03573_, _03572_);
  and _25893_ (_03575_, _13516_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and _25894_ (_03576_, _13521_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  or _25895_ (_03577_, _03576_, _03575_);
  or _25896_ (_03578_, _03577_, _03574_);
  or _25897_ (_03579_, _03578_, _03571_);
  nor _25898_ (_03580_, _13528_, _00749_);
  and _25899_ (_03581_, _13531_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  or _25900_ (_03582_, _03581_, _03580_);
  and _25901_ (_03583_, _13536_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and _25902_ (_03584_, _13534_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  or _25903_ (_03585_, _03584_, _03583_);
  or _25904_ (_03586_, _03585_, _03582_);
  and _25905_ (_03587_, _13541_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  and _25906_ (_03588_, _13544_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  or _25907_ (_03589_, _03588_, _03587_);
  and _25908_ (_03590_, _13547_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _25909_ (_03591_, _13549_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  or _25910_ (_03592_, _03591_, _03590_);
  or _25911_ (_03594_, _03592_, _03589_);
  or _25912_ (_03595_, _03594_, _03586_);
  or _25913_ (_03596_, _03595_, _03579_);
  and _25914_ (_03597_, _13555_, _11430_);
  and _25915_ (_03598_, _13562_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  or _25916_ (_03599_, _03598_, _03597_);
  and _25917_ (_03601_, _13475_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and _25918_ (_03602_, _13568_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or _25919_ (_03604_, _03602_, _03601_);
  or _25920_ (_03605_, _03604_, _03599_);
  or _25921_ (_03606_, _13592_, p0_in[5]);
  or _25922_ (_03607_, _00099_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and _25923_ (_03608_, _03607_, _03606_);
  and _25924_ (_03609_, _03608_, _13574_);
  or _25925_ (_03610_, _13592_, p1_in[5]);
  or _25926_ (_03611_, _00099_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and _25927_ (_03612_, _03611_, _03610_);
  and _25928_ (_03613_, _03612_, _13598_);
  or _25929_ (_03615_, _03613_, _03609_);
  or _25930_ (_03616_, _13592_, p2_in[5]);
  or _25931_ (_03617_, _00099_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and _25932_ (_03618_, _03617_, _03616_);
  and _25933_ (_03619_, _03618_, _13611_);
  or _25934_ (_03620_, _13592_, p3_in[5]);
  or _25935_ (_03621_, _00099_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and _25936_ (_03622_, _03621_, _03620_);
  and _25937_ (_03624_, _03622_, _13605_);
  or _25938_ (_03625_, _03624_, _03619_);
  or _25939_ (_03626_, _03625_, _03615_);
  or _25940_ (_03627_, _03626_, _03605_);
  and _25941_ (_03628_, _13681_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and _25942_ (_03629_, _13622_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  or _25943_ (_03630_, _03629_, _03628_);
  or _25944_ (_03631_, _03630_, _03627_);
  or _25945_ (_03632_, _03631_, _03596_);
  and _25946_ (_03633_, _03632_, _13701_);
  and _25947_ (_03634_, _13735_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  or _25948_ (_03635_, _03634_, _13476_);
  or _25949_ (_03637_, _03635_, _03633_);
  and _25950_ (_03665_, _03637_, _03563_);
  and _25951_ (_03639_, _12299_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  and _25952_ (_03640_, _10945_, _10905_);
  or _25953_ (_03641_, _11088_, _05816_);
  or _25954_ (_03642_, _03641_, _03476_);
  or _25955_ (_03643_, _03642_, _03640_);
  or _25956_ (_03644_, _12331_, _12309_);
  or _25957_ (_03646_, _05830_, _05824_);
  and _25958_ (_03647_, _03646_, _10843_);
  or _25959_ (_03648_, _03647_, _13383_);
  or _25960_ (_03649_, _03648_, _03644_);
  or _25961_ (_03650_, _11020_, _05841_);
  or _25962_ (_03652_, _03650_, _05848_);
  or _25963_ (_03653_, _03652_, _03649_);
  or _25964_ (_03654_, _03653_, _03643_);
  or _25965_ (_03655_, _03654_, _13400_);
  and _25966_ (_03656_, _03655_, _06576_);
  or _25967_ (_03671_, _03656_, _03639_);
  nand _25968_ (_03657_, _08041_, _06949_);
  or _25969_ (_03658_, _06949_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  and _25970_ (_03659_, _03658_, _05552_);
  and _25971_ (_03673_, _03659_, _03657_);
  nand _25972_ (_03675_, _11626_, _05552_);
  and _25973_ (_03661_, \oc8051_top_1.oc8051_memory_interface1.cdata [5], _07768_);
  and _25974_ (_03662_, \oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or _25975_ (_03663_, _03662_, _03661_);
  and _25976_ (_03679_, _03663_, _05552_);
  nand _25977_ (_03664_, _00647_, _08996_);
  or _25978_ (_03666_, _03664_, _00613_);
  nor _25979_ (_03667_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _08998_);
  nand _25980_ (_03668_, _03667_, _00580_);
  and _25981_ (_03669_, _03668_, _05552_);
  and _25982_ (_03681_, _03669_, _03666_);
  or _25983_ (_03670_, _05550_, \oc8051_top_1.oc8051_rom1.data_o [21]);
  nand _25984_ (_03672_, _05550_, _11057_);
  and _25985_ (_03674_, _03672_, _05552_);
  and _25986_ (_03688_, _03674_, _03670_);
  nor _25987_ (_03705_, _11900_, rst);
  and _25988_ (_03676_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], _07768_);
  and _25989_ (_03677_, \oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or _25990_ (_03678_, _03677_, _03676_);
  and _25991_ (_03712_, _03678_, _05552_);
  nand _25992_ (_03680_, _00241_, _07945_);
  or _25993_ (_03682_, _00241_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  and _25994_ (_03683_, _03682_, _05552_);
  and _25995_ (_03714_, _03683_, _03680_);
  nand _25996_ (_03684_, _00241_, _08386_);
  or _25997_ (_03685_, _00241_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  and _25998_ (_03686_, _03685_, _05552_);
  and _25999_ (_03718_, _03686_, _03684_);
  nor _26000_ (_03687_, _08041_, _06953_);
  and _26001_ (_03689_, _06953_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  or _26002_ (_03690_, _03689_, _06955_);
  or _26003_ (_03691_, _03690_, _03687_);
  or _26004_ (_03692_, _06068_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  and _26005_ (_03693_, _03692_, _05552_);
  and _26006_ (_03720_, _03693_, _03691_);
  nor _26007_ (_03750_, _11672_, rst);
  and _26008_ (_03694_, _03005_, _06771_);
  nand _26009_ (_03695_, _03694_, _06763_);
  or _26010_ (_03696_, _03694_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and _26011_ (_03697_, _03696_, _06775_);
  and _26012_ (_03698_, _03697_, _03695_);
  nor _26013_ (_03699_, _03011_, _06811_);
  and _26014_ (_03700_, _03011_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or _26015_ (_03701_, _03700_, _03699_);
  and _26016_ (_03702_, _03701_, _06524_);
  and _26017_ (_03703_, _06816_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or _26018_ (_03704_, _03703_, rst);
  or _26019_ (_03706_, _03704_, _03702_);
  or _26020_ (_03760_, _03706_, _03698_);
  and _26021_ (_03707_, _01622_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  nor _26022_ (_03708_, _07951_, _06560_);
  and _26023_ (_03709_, _06068_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  and _26024_ (_03710_, _03709_, _01625_);
  or _26025_ (_03711_, _03710_, _03708_);
  or _26026_ (_03713_, _03711_, _03707_);
  and _26027_ (_03769_, _03713_, _05552_);
  and _26028_ (_03715_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], _07768_);
  and _26029_ (_03716_, \oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or _26030_ (_03717_, _03716_, _03715_);
  and _26031_ (_03771_, _03717_, _05552_);
  or _26032_ (_03719_, _10982_, _08102_);
  or _26033_ (_03721_, _10981_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1]);
  and _26034_ (_03722_, _03721_, _05552_);
  and _26035_ (_03775_, _03722_, _03719_);
  and _26036_ (_03723_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and _26037_ (_03724_, _12140_, \oc8051_top_1.oc8051_rom1.data_o [19]);
  or _26038_ (_03725_, _03724_, _03723_);
  and _26039_ (_03784_, _03725_, _05552_);
  or _26040_ (_03726_, _10982_, _07711_);
  or _26041_ (_03727_, _10981_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  and _26042_ (_03728_, _03727_, _05552_);
  and _26043_ (_03814_, _03728_, _03726_);
  and _26044_ (_03729_, _12299_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  nand _26045_ (_03730_, _06568_, _05738_);
  nor _26046_ (_03731_, _05854_, _05840_);
  nand _26047_ (_03732_, _03731_, _10906_);
  nand _26048_ (_03733_, _03732_, _05894_);
  and _26049_ (_03734_, _03733_, _11166_);
  and _26050_ (_03735_, _03734_, _03730_);
  nand _26051_ (_03736_, _05861_, _05818_);
  or _26052_ (_03737_, _13583_, _10851_);
  and _26053_ (_03738_, _05855_, _05818_);
  nor _26054_ (_03739_, _03738_, _03737_);
  and _26055_ (_03740_, _03739_, _03736_);
  nand _26056_ (_03741_, _10929_, _05738_);
  or _26057_ (_03743_, _13575_, _12284_);
  nor _26058_ (_03744_, _03743_, _10924_);
  and _26059_ (_03745_, _03744_, _03741_);
  nor _26060_ (_03746_, _03456_, _12307_);
  and _26061_ (_03747_, _03746_, _03745_);
  and _26062_ (_03748_, _03747_, _03740_);
  nand _26063_ (_03749_, _03748_, _03735_);
  and _26064_ (_03751_, _03749_, _06576_);
  or _26065_ (_03824_, _03751_, _03729_);
  nand _26066_ (_03752_, _00241_, _06306_);
  or _26067_ (_03753_, _00241_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  and _26068_ (_03754_, _03753_, _05552_);
  and _26069_ (_03844_, _03754_, _03752_);
  and _26070_ (_03846_, _05552_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  nor _26071_ (_03755_, _07951_, _06811_);
  and _26072_ (_03756_, _01622_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  and _26073_ (_03757_, _06068_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  and _26074_ (_03758_, _03757_, _01625_);
  or _26075_ (_03759_, _03758_, _03756_);
  or _26076_ (_03761_, _03759_, _03755_);
  and _26077_ (_03850_, _03761_, _05552_);
  or _26078_ (_03762_, _05550_, \oc8051_top_1.oc8051_rom1.data_o [5]);
  nand _26079_ (_03763_, _05550_, _05748_);
  and _26080_ (_03764_, _03763_, _05552_);
  and _26081_ (_03873_, _03764_, _03762_);
  and _26082_ (_03765_, _08874_, rxd_i);
  not _26083_ (_03766_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0]);
  nor _26084_ (_03767_, _08874_, _03766_);
  or _26085_ (_03768_, _03767_, _03765_);
  and _26086_ (_03881_, _03768_, _05552_);
  and _26087_ (_03883_, _07209_, _05552_);
  and _26088_ (_03770_, _07939_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  nor _26089_ (_03772_, _07939_, _06811_);
  or _26090_ (_03773_, _03772_, _03770_);
  and _26091_ (_03888_, _03773_, _05552_);
  or _26092_ (_03774_, _01751_, _07255_);
  not _26093_ (_03776_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  nand _26094_ (_03777_, _01751_, _03776_);
  and _26095_ (_03778_, _03777_, _06524_);
  and _26096_ (_03779_, _03778_, _03774_);
  nor _26097_ (_03780_, _06774_, _03776_);
  and _26098_ (_03781_, _01750_, _06771_);
  nand _26099_ (_03782_, _03781_, _06763_);
  or _26100_ (_03783_, _03781_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and _26101_ (_03785_, _03783_, _06775_);
  and _26102_ (_03786_, _03785_, _03782_);
  or _26103_ (_03787_, _03786_, _03780_);
  or _26104_ (_03788_, _03787_, _03779_);
  and _26105_ (_03895_, _03788_, _05552_);
  and _26106_ (_03789_, _05550_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and _26107_ (_03790_, _12140_, \oc8051_top_1.oc8051_rom1.data_o [4]);
  or _26108_ (_03791_, _03790_, _03789_);
  and _26109_ (_03902_, _03791_, _05552_);
  and _26110_ (_03792_, _06068_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  and _26111_ (_03793_, _03792_, _13739_);
  and _26112_ (_03794_, _07946_, _06309_);
  and _26113_ (_03795_, _06070_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  or _26114_ (_03796_, _03795_, _03794_);
  or _26115_ (_03797_, _03796_, _03793_);
  and _26116_ (_03914_, _03797_, _05552_);
  or _26117_ (_03798_, _05550_, \oc8051_top_1.oc8051_rom1.data_o [3]);
  nand _26118_ (_03799_, _05550_, _05699_);
  and _26119_ (_03800_, _03799_, _05552_);
  and _26120_ (_03936_, _03800_, _03798_);
  not _26121_ (_03801_, _01819_);
  not _26122_ (_03802_, _10639_);
  and _26123_ (_03803_, _01824_, _03802_);
  and _26124_ (_03804_, _03803_, _01803_);
  nand _26125_ (_03805_, _03804_, _03801_);
  or _26126_ (_03806_, _03804_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  and _26127_ (_03807_, _03806_, _05552_);
  and _26128_ (_03966_, _03807_, _03805_);
  not _26129_ (_03808_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  or _26130_ (_03809_, _03808_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  or _26131_ (_03810_, _03809_, _05560_);
  and _26132_ (_03811_, _03810_, _00384_);
  or _26133_ (_03812_, _03811_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or _26134_ (_03813_, _03812_, _00225_);
  or _26135_ (_03815_, _06060_, _05570_);
  nand _26136_ (_03816_, _03815_, _00225_);
  or _26137_ (_03817_, _03816_, _13359_);
  and _26138_ (_03818_, _03817_, _03813_);
  or _26139_ (_03819_, _03818_, _00232_);
  nand _26140_ (_03820_, _00232_, _07945_);
  and _26141_ (_03821_, _03820_, _05552_);
  and _26142_ (_03974_, _03821_, _03819_);
  or _26143_ (_03822_, _05550_, \oc8051_top_1.oc8051_rom1.data_o [11]);
  nand _26144_ (_03823_, _05550_, _11002_);
  and _26145_ (_03825_, _03823_, _05552_);
  and _26146_ (_04015_, _03825_, _03822_);
  or _26147_ (_03826_, _05550_, \oc8051_top_1.oc8051_rom1.data_o [15]);
  nand _26148_ (_03827_, _05550_, _07743_);
  and _26149_ (_03828_, _03827_, _05552_);
  and _26150_ (_04017_, _03828_, _03826_);
  and _26151_ (_03829_, _00225_, _08365_);
  nand _26152_ (_03830_, _03829_, _06763_);
  or _26153_ (_03831_, _03829_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  and _26154_ (_03832_, _03831_, _00451_);
  and _26155_ (_03833_, _03832_, _03830_);
  nor _26156_ (_03834_, _00451_, _08386_);
  or _26157_ (_03835_, _03834_, _03833_);
  and _26158_ (_04020_, _03835_, _05552_);
  or _26159_ (_03836_, _13701_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  and _26160_ (_03837_, _13488_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  and _26161_ (_03838_, _13494_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or _26162_ (_03839_, _03838_, _03837_);
  and _26163_ (_03840_, _13502_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and _26164_ (_03841_, _13499_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  or _26165_ (_03842_, _03841_, _03840_);
  or _26166_ (_03843_, _03842_, _03839_);
  and _26167_ (_03845_, _13507_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and _26168_ (_03847_, _13511_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  or _26169_ (_03848_, _03847_, _03845_);
  and _26170_ (_03849_, _13516_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and _26171_ (_03851_, _13521_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  or _26172_ (_03852_, _03851_, _03849_);
  or _26173_ (_03853_, _03852_, _03848_);
  or _26174_ (_03854_, _03853_, _03843_);
  and _26175_ (_03855_, _13531_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  nor _26176_ (_03856_, _13528_, _00758_);
  or _26177_ (_03857_, _03856_, _03855_);
  and _26178_ (_03858_, _13534_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and _26179_ (_03859_, _13536_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  or _26180_ (_03860_, _03859_, _03858_);
  or _26181_ (_03861_, _03860_, _03857_);
  and _26182_ (_03862_, _13541_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  and _26183_ (_03863_, _13544_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  or _26184_ (_03864_, _03863_, _03862_);
  and _26185_ (_03865_, _13547_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and _26186_ (_03866_, _13549_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or _26187_ (_03867_, _03866_, _03865_);
  or _26188_ (_03868_, _03867_, _03864_);
  or _26189_ (_03869_, _03868_, _03861_);
  or _26190_ (_03870_, _03869_, _03854_);
  and _26191_ (_03871_, _13475_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and _26192_ (_03872_, _13568_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or _26193_ (_03874_, _03872_, _03871_);
  and _26194_ (_03875_, _13555_, _11308_);
  and _26195_ (_03876_, _13562_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  or _26196_ (_03877_, _03876_, _03875_);
  or _26197_ (_03878_, _03877_, _03874_);
  or _26198_ (_03879_, _13592_, p3_in[7]);
  or _26199_ (_03880_, _00099_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and _26200_ (_03882_, _03880_, _03879_);
  and _26201_ (_03884_, _03882_, _13605_);
  or _26202_ (_03885_, _13592_, p2_in[7]);
  or _26203_ (_03886_, _00099_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and _26204_ (_03887_, _03886_, _03885_);
  and _26205_ (_03889_, _03887_, _13611_);
  or _26206_ (_03890_, _03889_, _03884_);
  or _26207_ (_03891_, _13592_, p1_in[7]);
  or _26208_ (_03892_, _00099_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and _26209_ (_03893_, _03892_, _03891_);
  and _26210_ (_03894_, _03893_, _13598_);
  or _26211_ (_03896_, _13592_, p0_in[7]);
  or _26212_ (_03897_, _00099_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and _26213_ (_03898_, _03897_, _03896_);
  and _26214_ (_03899_, _03898_, _13574_);
  or _26215_ (_03900_, _03899_, _03894_);
  or _26216_ (_03901_, _03900_, _03890_);
  or _26217_ (_03903_, _03901_, _03878_);
  and _26218_ (_03904_, _13622_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  and _26219_ (_03905_, _13681_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or _26220_ (_03906_, _03905_, _03904_);
  or _26221_ (_03907_, _03906_, _03903_);
  or _26222_ (_03908_, _03907_, _03870_);
  and _26223_ (_03909_, _13735_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  or _26224_ (_03910_, _03909_, _03908_);
  and _26225_ (_03911_, _03910_, _03836_);
  or _26226_ (_03912_, _03911_, _13476_);
  or _26227_ (_03913_, _13704_, _07255_);
  and _26228_ (_03915_, _03913_, _05552_);
  and _26229_ (_04036_, _03915_, _03912_);
  nor _26230_ (_03916_, _00374_, rst);
  or _26231_ (_03917_, _00373_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  nand _26232_ (_03918_, _00373_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  and _26233_ (_03919_, _03918_, _03917_);
  and _26234_ (_04039_, _03919_, _03916_);
  or _26235_ (_03920_, _05550_, \oc8051_top_1.oc8051_rom1.data_o [2]);
  nand _26236_ (_03921_, _05550_, _05677_);
  and _26237_ (_03922_, _03921_, _05552_);
  and _26238_ (_04044_, _03922_, _03920_);
  and _26239_ (_04050_, _05552_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  nor _26240_ (_03923_, _07951_, _06306_);
  and _26241_ (_03924_, _01622_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  and _26242_ (_03925_, _06068_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  and _26243_ (_03926_, _03925_, _01625_);
  or _26244_ (_03927_, _03926_, _03924_);
  or _26245_ (_03928_, _03927_, _03923_);
  and _26246_ (_04052_, _03928_, _05552_);
  and _26247_ (_04054_, _05552_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  or _26248_ (_03929_, _12308_, _10851_);
  or _26249_ (_03930_, _12280_, _10913_);
  or _26250_ (_03931_, _03930_, _03929_);
  or _26251_ (_03932_, _03931_, _11088_);
  and _26252_ (_03933_, _03932_, _05547_);
  and _26253_ (_03934_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _26254_ (_03935_, _03934_, _05901_);
  or _26255_ (_03937_, _03935_, _03933_);
  and _26256_ (_04062_, _03937_, _05552_);
  and _26257_ (_03938_, _01740_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or _26258_ (_03939_, _03938_, _01741_);
  and _26259_ (_03940_, _03939_, _08009_);
  nand _26260_ (_03941_, _11591_, _06763_);
  nor _26261_ (_03942_, _11591_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor _26262_ (_03943_, _03942_, _08009_);
  and _26263_ (_03944_, _03943_, _03941_);
  or _26264_ (_03945_, _03944_, _06531_);
  or _26265_ (_03946_, _03945_, _03940_);
  nand _26266_ (_03947_, _06811_, _06531_);
  and _26267_ (_03948_, _03947_, _05552_);
  and _26268_ (_04069_, _03948_, _03946_);
  and _26269_ (_04074_, _07117_, _05552_);
  and _26270_ (_03949_, _01234_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  and _26271_ (_03950_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _08998_);
  nor _26272_ (_03951_, _03950_, _03667_);
  nor _26273_ (_03952_, _03951_, _00857_);
  or _26274_ (_03953_, _03952_, _00580_);
  or _26275_ (_03954_, _03953_, _03949_);
  or _26276_ (_03955_, _03951_, _00838_);
  and _26277_ (_03956_, _03955_, _05552_);
  and _26278_ (_04077_, _03956_, _03954_);
  nor _26279_ (_04080_, _11095_, rst);
  or _26280_ (_03957_, _05550_, \oc8051_top_1.oc8051_rom1.data_o [1]);
  nand _26281_ (_03958_, _05550_, _05611_);
  and _26282_ (_03959_, _03958_, _05552_);
  and _26283_ (_04082_, _03959_, _03957_);
  and _26284_ (_03960_, _12299_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and _26285_ (_03961_, _06567_, _05857_);
  or _26286_ (_03962_, _03961_, _05831_);
  or _26287_ (_03963_, _03962_, _11133_);
  or _26288_ (_03964_, _11570_, _11124_);
  and _26289_ (_03965_, _06570_, _05894_);
  or _26290_ (_03967_, _13386_, _03965_);
  or _26291_ (_03968_, _03967_, _03964_);
  or _26292_ (_03969_, _11127_, _11167_);
  or _26293_ (_03970_, _03969_, _11573_);
  or _26294_ (_03971_, _03970_, _03968_);
  or _26295_ (_03972_, _03971_, _03963_);
  and _26296_ (_03973_, _03972_, _06576_);
  or _26297_ (_04091_, _03973_, _03960_);
  and _26298_ (_04128_, _07200_, _05552_);
  and _26299_ (_04133_, _00375_, _05552_);
  or _26300_ (_04142_, _08764_, _06568_);
  and _26301_ (_03975_, _05803_, _07781_);
  and _26302_ (_03976_, _03975_, _05781_);
  or _26303_ (_03977_, _07897_, _07775_);
  and _26304_ (_03978_, _03977_, _03976_);
  and _26305_ (_03979_, _07898_, _07807_);
  or _26306_ (_03980_, _03979_, _02640_);
  or _26307_ (_03981_, _03980_, _03978_);
  or _26308_ (_03982_, _07853_, _07840_);
  and _26309_ (_03983_, _07862_, _05710_);
  or _26310_ (_03984_, _07923_, _03983_);
  or _26311_ (_03985_, _03984_, _03982_);
  nand _26312_ (_03986_, _07848_, _07815_);
  nor _26313_ (_03987_, _07798_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and _26314_ (_03988_, _03987_, _03986_);
  nand _26315_ (_03989_, _03988_, _07786_);
  nand _26316_ (_03990_, _07867_, _07864_);
  or _26317_ (_03991_, _03990_, _03989_);
  or _26318_ (_03992_, _03991_, _03985_);
  or _26319_ (_03993_, _03992_, _03981_);
  or _26320_ (_03994_, _03993_, _02649_);
  and _26321_ (_03995_, _03994_, _05608_);
  nor _26322_ (_03996_, _02639_, _05891_);
  or _26323_ (_03997_, _03996_, rst);
  or _26324_ (_04144_, _03997_, _03995_);
  and _26325_ (_04147_, _13702_, _13477_);
  and _26326_ (_03998_, _13621_, _11279_);
  or _26327_ (_03999_, _13677_, _13481_);
  or _26328_ (_04000_, _11763_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and _26329_ (_04001_, _04000_, _13480_);
  and _26330_ (_04002_, _04001_, _03999_);
  and _26331_ (_04003_, _13509_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  and _26332_ (_04004_, _13497_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  or _26333_ (_04005_, _04004_, _04003_);
  and _26334_ (_04006_, _04005_, _13481_);
  and _26335_ (_04007_, _11763_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  nor _26336_ (_04008_, _11763_, _07468_);
  or _26337_ (_04009_, _04008_, _04007_);
  and _26338_ (_04010_, _04009_, _13464_);
  and _26339_ (_04011_, _13509_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and _26340_ (_04012_, _13497_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  or _26341_ (_04013_, _04012_, _04011_);
  and _26342_ (_04014_, _04013_, _11763_);
  or _26343_ (_04016_, _04014_, _04010_);
  or _26344_ (_04018_, _04016_, _04006_);
  or _26345_ (_04019_, _04018_, _04002_);
  and _26346_ (_04021_, _04019_, _03998_);
  not _26347_ (_04022_, _11279_);
  and _26348_ (_04023_, _11763_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and _26349_ (_04024_, _13481_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  or _26350_ (_04025_, _04024_, _04023_);
  and _26351_ (_04026_, _04025_, _13509_);
  and _26352_ (_04027_, _11763_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and _26353_ (_04028_, _13481_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  or _26354_ (_04029_, _04028_, _04027_);
  and _26355_ (_04030_, _04029_, _13464_);
  nor _26356_ (_04031_, _11763_, _00592_);
  and _26357_ (_04032_, _11763_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  or _26358_ (_04033_, _04032_, _04031_);
  and _26359_ (_04034_, _04033_, _13480_);
  or _26360_ (_04035_, _04034_, _04030_);
  nor _26361_ (_04037_, _11763_, _00587_);
  and _26362_ (_04038_, _11763_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  or _26363_ (_04040_, _04038_, _04037_);
  and _26364_ (_04041_, _04040_, _13497_);
  or _26365_ (_04042_, _04041_, _04035_);
  or _26366_ (_04043_, _04042_, _04026_);
  and _26367_ (_04045_, _04043_, _13515_);
  and _26368_ (_04046_, _11763_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and _26369_ (_04047_, _13481_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or _26370_ (_04048_, _04047_, _04046_);
  and _26371_ (_04049_, _04048_, _13509_);
  and _26372_ (_04051_, _11763_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and _26373_ (_04053_, _13481_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or _26374_ (_04055_, _04053_, _04051_);
  and _26375_ (_04056_, _04055_, _13464_);
  nor _26376_ (_04057_, _11763_, _01054_);
  and _26377_ (_04058_, _11763_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  or _26378_ (_04059_, _04058_, _04057_);
  and _26379_ (_04060_, _04059_, _13480_);
  or _26380_ (_04061_, _04060_, _04056_);
  and _26381_ (_04063_, _13481_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and _26382_ (_04064_, _11763_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or _26383_ (_04065_, _04064_, _04063_);
  and _26384_ (_04066_, _04065_, _13497_);
  or _26385_ (_04067_, _04066_, _04061_);
  or _26386_ (_04068_, _04067_, _04049_);
  and _26387_ (_04070_, _04068_, _13472_);
  or _26388_ (_04071_, _04070_, _04045_);
  and _26389_ (_04072_, _11763_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and _26390_ (_04073_, _13481_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or _26391_ (_04075_, _04073_, _04072_);
  and _26392_ (_04076_, _04075_, _13464_);
  nor _26393_ (_04078_, _11763_, _02787_);
  and _26394_ (_04079_, _11763_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  or _26395_ (_04081_, _04079_, _04078_);
  and _26396_ (_04083_, _04081_, _13480_);
  or _26397_ (_04084_, _04083_, _04076_);
  and _26398_ (_04085_, _11763_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and _26399_ (_04086_, _13481_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  or _26400_ (_04087_, _04086_, _04085_);
  and _26401_ (_04088_, _04087_, _13509_);
  nor _26402_ (_04089_, _11763_, _12096_);
  and _26403_ (_04090_, _11763_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or _26404_ (_04092_, _04090_, _04089_);
  and _26405_ (_04093_, _04092_, _13497_);
  or _26406_ (_04094_, _04093_, _04088_);
  or _26407_ (_04095_, _04094_, _04084_);
  and _26408_ (_04096_, _04095_, _13487_);
  or _26409_ (_04097_, _04096_, _04071_);
  and _26410_ (_04098_, _04097_, _04022_);
  and _26411_ (_04099_, _13620_, _11279_);
  and _26412_ (_04100_, _04099_, _13560_);
  nor _26413_ (_04101_, _04100_, _03998_);
  and _26414_ (_04102_, _11509_, _11279_);
  and _26415_ (_04103_, _13561_, _04102_);
  nor _26416_ (_04104_, _13469_, _04022_);
  nor _26417_ (_04105_, _04104_, _04103_);
  and _26418_ (_04106_, _04105_, _04101_);
  nor _26419_ (_04107_, _13487_, _13727_);
  or _26420_ (_04108_, _04107_, _11279_);
  nand _26421_ (_04109_, _13514_, _11279_);
  and _26422_ (_04110_, _04109_, \oc8051_top_1.oc8051_sfr1.bit_out );
  and _26423_ (_04111_, _04110_, _04108_);
  and _26424_ (_04112_, _04111_, _04106_);
  nor _26425_ (_04113_, _13471_, _04022_);
  and _26426_ (_04114_, _00114_, _11763_);
  and _26427_ (_04115_, _03413_, _13481_);
  or _26428_ (_04116_, _04115_, _04114_);
  and _26429_ (_04117_, _04116_, _13464_);
  and _26430_ (_04118_, _13812_, _13481_);
  and _26431_ (_04119_, _13596_, _11763_);
  or _26432_ (_04120_, _04119_, _04118_);
  and _26433_ (_04121_, _04120_, _13480_);
  or _26434_ (_04122_, _04121_, _04117_);
  and _26435_ (_04123_, _00184_, _11763_);
  and _26436_ (_04124_, _03608_, _13481_);
  or _26437_ (_04125_, _04124_, _04123_);
  and _26438_ (_04126_, _04125_, _13497_);
  and _26439_ (_04127_, _03898_, _13481_);
  and _26440_ (_04129_, _00023_, _11763_);
  or _26441_ (_04130_, _04129_, _04127_);
  and _26442_ (_04131_, _04130_, _13509_);
  or _26443_ (_04132_, _04131_, _04126_);
  or _26444_ (_04134_, _04132_, _04122_);
  and _26445_ (_04135_, _04134_, _04113_);
  or _26446_ (_04136_, _04135_, _04112_);
  and _26447_ (_04137_, _11763_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  nor _26448_ (_04138_, _11763_, _03545_);
  or _26449_ (_04139_, _04138_, _04137_);
  and _26450_ (_04140_, _04139_, _13464_);
  nor _26451_ (_04141_, _11763_, _01767_);
  and _26452_ (_04143_, _11763_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  or _26453_ (_04145_, _04143_, _04141_);
  and _26454_ (_04146_, _04145_, _13480_);
  or _26455_ (_04148_, _04146_, _04140_);
  and _26456_ (_04149_, _11763_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nor _26457_ (_04150_, _11763_, _03776_);
  or _26458_ (_04151_, _04150_, _04149_);
  and _26459_ (_04152_, _04151_, _13509_);
  nor _26460_ (_04153_, _11763_, _01753_);
  and _26461_ (_04155_, _11763_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  or _26462_ (_04156_, _04155_, _04153_);
  and _26463_ (_04157_, _04156_, _13497_);
  or _26464_ (_04158_, _04157_, _04152_);
  or _26465_ (_04159_, _04158_, _04148_);
  and _26466_ (_04160_, _04159_, _04100_);
  and _26467_ (_04161_, _11763_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor _26468_ (_04162_, _11763_, _06396_);
  or _26469_ (_04163_, _04162_, _04161_);
  and _26470_ (_04164_, _04163_, _13464_);
  nor _26471_ (_04165_, _11763_, _06157_);
  and _26472_ (_04167_, _11763_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or _26473_ (_04169_, _04167_, _04165_);
  and _26474_ (_04170_, _04169_, _13480_);
  or _26475_ (_04171_, _04170_, _04164_);
  and _26476_ (_04172_, _11763_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor _26477_ (_04173_, _11763_, _06361_);
  or _26478_ (_04174_, _04173_, _04172_);
  and _26479_ (_04175_, _04174_, _13509_);
  nor _26480_ (_04177_, _11763_, _06103_);
  and _26481_ (_04178_, _11763_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or _26482_ (_04180_, _04178_, _04177_);
  and _26483_ (_04182_, _04180_, _13497_);
  or _26484_ (_04183_, _04182_, _04175_);
  or _26485_ (_04185_, _04183_, _04171_);
  and _26486_ (_04187_, _04185_, _04103_);
  or _26487_ (_04189_, _04187_, _04160_);
  or _26488_ (_04190_, _04189_, _04136_);
  nor _26489_ (_04191_, _11763_, _03808_);
  and _26490_ (_04192_, _11763_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  or _26491_ (_04193_, _04192_, _04191_);
  and _26492_ (_04194_, _04193_, _13497_);
  or _26493_ (_04195_, _04194_, _11279_);
  and _26494_ (_04196_, _11763_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  and _26495_ (_04197_, _13481_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  or _26496_ (_04198_, _04197_, _04196_);
  and _26497_ (_04199_, _04198_, _13464_);
  and _26498_ (_04200_, _13481_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and _26499_ (_04201_, _11763_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or _26500_ (_04202_, _04201_, _04200_);
  and _26501_ (_04203_, _04202_, _13480_);
  and _26502_ (_04204_, _11763_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  nor _26503_ (_04205_, _11763_, _12098_);
  or _26504_ (_04206_, _04205_, _04204_);
  and _26505_ (_04207_, _04206_, _13509_);
  or _26506_ (_04208_, _04207_, _04203_);
  or _26507_ (_04209_, _04208_, _04199_);
  or _26508_ (_04210_, _04209_, _04195_);
  and _26509_ (_04211_, _13602_, _11763_);
  and _26510_ (_04212_, _13817_, _13481_);
  or _26511_ (_04213_, _04212_, _04211_);
  and _26512_ (_04214_, _04213_, _13480_);
  and _26513_ (_04215_, _00188_, _11763_);
  and _26514_ (_04216_, _03612_, _13481_);
  or _26515_ (_04217_, _04216_, _04215_);
  and _26516_ (_04218_, _04217_, _13497_);
  or _26517_ (_04219_, _04218_, _04022_);
  or _26518_ (_04220_, _04219_, _04214_);
  and _26519_ (_04222_, _00110_, _13464_);
  and _26520_ (_04223_, _00029_, _13509_);
  or _26521_ (_04224_, _04223_, _04222_);
  and _26522_ (_04225_, _04224_, _11763_);
  and _26523_ (_04226_, _03418_, _13464_);
  and _26524_ (_04227_, _03893_, _13509_);
  or _26525_ (_04228_, _04227_, _04226_);
  and _26526_ (_04229_, _04228_, _13481_);
  or _26527_ (_04230_, _04229_, _04225_);
  or _26528_ (_04231_, _04230_, _04220_);
  and _26529_ (_04232_, _04231_, _13540_);
  and _26530_ (_04233_, _04232_, _04210_);
  and _26531_ (_04234_, _13615_, _11763_);
  and _26532_ (_04235_, _13801_, _13481_);
  or _26533_ (_04236_, _04235_, _04234_);
  and _26534_ (_04237_, _04236_, _13480_);
  and _26535_ (_04238_, _00175_, _11763_);
  and _26536_ (_04239_, _03618_, _13481_);
  or _26537_ (_04240_, _04239_, _04238_);
  and _26538_ (_04241_, _04240_, _13497_);
  or _26539_ (_04242_, _04241_, _13465_);
  or _26540_ (_04243_, _04242_, _04237_);
  and _26541_ (_04244_, _00105_, _13464_);
  and _26542_ (_04245_, _00040_, _13509_);
  or _26543_ (_04246_, _04245_, _04244_);
  and _26544_ (_04247_, _04246_, _11763_);
  and _26545_ (_04248_, _03429_, _13464_);
  and _26546_ (_04249_, _03887_, _13509_);
  or _26547_ (_04250_, _04249_, _04248_);
  and _26548_ (_04251_, _04250_, _13481_);
  or _26549_ (_04252_, _04251_, _04247_);
  or _26550_ (_04253_, _04252_, _04243_);
  and _26551_ (_04254_, _13609_, _11763_);
  and _26552_ (_04255_, _13806_, _13481_);
  or _26553_ (_04256_, _04255_, _04254_);
  and _26554_ (_04257_, _04256_, _13480_);
  and _26555_ (_04258_, _00179_, _11763_);
  and _26556_ (_04259_, _03622_, _13481_);
  or _26557_ (_04260_, _04259_, _04258_);
  and _26558_ (_04261_, _04260_, _13497_);
  or _26559_ (_04262_, _04261_, _11509_);
  nor _26560_ (_04263_, _04262_, _04257_);
  nand _26561_ (_04264_, _00101_, _13464_);
  nand _26562_ (_04265_, _00035_, _13509_);
  and _26563_ (_04266_, _04265_, _04264_);
  or _26564_ (_04267_, _04266_, _13481_);
  nand _26565_ (_04268_, _03423_, _13464_);
  nand _26566_ (_04269_, _03882_, _13509_);
  and _26567_ (_04270_, _04269_, _04268_);
  or _26568_ (_04271_, _04270_, _11763_);
  and _26569_ (_04272_, _04271_, _04267_);
  and _26570_ (_04273_, _04272_, _04263_);
  nor _26571_ (_04274_, _04273_, _04109_);
  and _26572_ (_04276_, _04274_, _04253_);
  and _26573_ (_04277_, _13518_, _04022_);
  nor _26574_ (_04278_, _11763_, _00617_);
  and _26575_ (_04279_, _11763_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  or _26576_ (_04280_, _04279_, _04278_);
  and _26577_ (_04281_, _04280_, _13480_);
  nor _26578_ (_04282_, _11763_, _00615_);
  and _26579_ (_04283_, _11763_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  or _26580_ (_04285_, _04283_, _04282_);
  and _26581_ (_04286_, _04285_, _13497_);
  or _26582_ (_04287_, _04286_, _04281_);
  and _26583_ (_04288_, _11763_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and _26584_ (_04289_, _13481_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  or _26585_ (_04290_, _04289_, _04288_);
  and _26586_ (_04291_, _04290_, _13464_);
  and _26587_ (_04292_, _11763_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and _26588_ (_04293_, _13481_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  or _26589_ (_04294_, _04293_, _04292_);
  and _26590_ (_04296_, _04294_, _13509_);
  or _26591_ (_04297_, _04296_, _04291_);
  or _26592_ (_04298_, _04297_, _04287_);
  and _26593_ (_04299_, _04298_, _04277_);
  and _26594_ (_04300_, _11769_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  or _26595_ (_04301_, _04300_, _04299_);
  or _26596_ (_04302_, _04301_, _04276_);
  or _26597_ (_04303_, _04302_, _04233_);
  or _26598_ (_04304_, _04303_, _04190_);
  or _26599_ (_04305_, _04304_, _04098_);
  or _26600_ (_04306_, _04305_, _04021_);
  and _26601_ (_04307_, _04103_, _06965_);
  nor _26602_ (_04308_, _04307_, _11518_);
  nand _26603_ (_04309_, _04300_, _06763_);
  and _26604_ (_04310_, _04309_, _04308_);
  and _26605_ (_04311_, _04310_, _04306_);
  and _26606_ (_04312_, _11763_, _11214_);
  nor _26607_ (_04313_, _11763_, _06811_);
  or _26608_ (_04314_, _04313_, _04312_);
  and _26609_ (_04315_, _04314_, _13509_);
  nor _26610_ (_04316_, _11763_, _07388_);
  and _26611_ (_04317_, _11763_, _11238_);
  or _26612_ (_04318_, _04317_, _04316_);
  and _26613_ (_04319_, _04318_, _13480_);
  nor _26614_ (_04320_, _11763_, _08386_);
  and _26615_ (_04321_, _11763_, _11726_);
  or _26616_ (_04322_, _04321_, _04320_);
  and _26617_ (_04323_, _04322_, _13464_);
  or _26618_ (_04324_, _04323_, _04319_);
  nor _26619_ (_04325_, _11763_, _06306_);
  and _26620_ (_04326_, _11763_, _11234_);
  or _26621_ (_04327_, _04326_, _04325_);
  and _26622_ (_04328_, _04327_, _13497_);
  or _26623_ (_04329_, _04328_, _04324_);
  nor _26624_ (_04330_, _04329_, _04315_);
  nor _26625_ (_04331_, _04330_, _04308_);
  or _26626_ (_04332_, _04331_, _04311_);
  and _26627_ (_04154_, _04332_, _05552_);
  and _26628_ (_04333_, _02681_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  and _26629_ (_04334_, _02680_, _11238_);
  or _26630_ (_04335_, _04334_, _04333_);
  and _26631_ (_04166_, _04335_, _05552_);
  or _26632_ (_04336_, _05781_, _08675_);
  or _26633_ (_04337_, _05546_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and _26634_ (_04338_, _04337_, _05552_);
  and _26635_ (_04168_, _04338_, _04336_);
  and _26636_ (_04339_, _12299_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  or _26637_ (_04340_, _11559_, _10913_);
  nand _26638_ (_04341_, _05894_, _05840_);
  nand _26639_ (_04342_, _10923_, _04341_);
  or _26640_ (_04343_, _04342_, _04340_);
  not _26641_ (_04344_, _11088_);
  nand _26642_ (_04345_, _11111_, _04344_);
  or _26643_ (_04346_, _04345_, _04343_);
  or _26644_ (_04347_, _04346_, _12332_);
  or _26645_ (_04348_, _04347_, _12327_);
  and _26646_ (_04349_, _04348_, _06576_);
  or _26647_ (_04176_, _04349_, _04339_);
  and _26648_ (_04350_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and _26649_ (_04351_, _05858_, _05547_);
  or _26650_ (_04353_, _04351_, _04350_);
  or _26651_ (_04354_, _04353_, _05901_);
  and _26652_ (_04179_, _04354_, _05552_);
  or _26653_ (_04355_, _03961_, _05889_);
  or _26654_ (_04356_, _05890_, _05547_);
  and _26655_ (_04357_, _04356_, _04355_);
  and _26656_ (_04358_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _26657_ (_04359_, _04358_, _10956_);
  or _26658_ (_04360_, _04359_, _04357_);
  and _26659_ (_04181_, _04360_, _05552_);
  and _26660_ (_04361_, _12299_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  or _26661_ (_04362_, _11174_, _05829_);
  or _26662_ (_04363_, _03647_, _12331_);
  or _26663_ (_04364_, _04363_, _04362_);
  or _26664_ (_04365_, _12324_, _11167_);
  or _26665_ (_04366_, _04365_, _03483_);
  or _26666_ (_04367_, _04366_, _03641_);
  or _26667_ (_04368_, _04367_, _04364_);
  and _26668_ (_04369_, _04368_, _06576_);
  or _26669_ (_04184_, _04369_, _04361_);
  and _26670_ (_04370_, _12299_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  or _26671_ (_04371_, _03743_, _05855_);
  or _26672_ (_04372_, _13578_, _10847_);
  or _26673_ (_04373_, _04372_, _04371_);
  or _26674_ (_04374_, _03737_, _10897_);
  or _26675_ (_04375_, _04374_, _04373_);
  or _26676_ (_04376_, _12270_, _11152_);
  or _26677_ (_04377_, _04376_, _12334_);
  or _26678_ (_04378_, _04377_, _04375_);
  or _26679_ (_04379_, _04378_, _12327_);
  and _26680_ (_04380_, _04379_, _06576_);
  or _26681_ (_04186_, _04380_, _04370_);
  and _26682_ (_04381_, _13384_, _05547_);
  nand _26683_ (_04382_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  nand _26684_ (_04383_, _04382_, _10959_);
  or _26685_ (_04384_, _04383_, _04381_);
  and _26686_ (_04188_, _04384_, _05552_);
  or _26687_ (_04385_, _12308_, _11033_);
  or _26688_ (_04386_, _04385_, _05876_);
  or _26689_ (_04387_, _04386_, _11180_);
  or _26690_ (_04388_, _03479_, _05873_);
  or _26691_ (_04389_, _04388_, _04387_);
  or _26692_ (_04390_, _12332_, _10849_);
  or _26693_ (_04391_, _04390_, _04389_);
  or _26694_ (_04392_, _04391_, _05868_);
  and _26695_ (_04393_, _04392_, _05547_);
  and _26696_ (_04394_, \oc8051_top_1.oc8051_decoder1.wr , \oc8051_top_1.oc8051_sfr1.wait_data );
  or _26697_ (_04395_, _04394_, _05903_);
  or _26698_ (_04396_, _04395_, _04393_);
  and _26699_ (_04221_, _04396_, _05552_);
  or _26700_ (_04397_, _05550_, \oc8051_top_1.oc8051_rom1.data_o [14]);
  nand _26701_ (_04398_, _05550_, _11383_);
  and _26702_ (_04399_, _04398_, _05552_);
  and _26703_ (_04275_, _04399_, _04397_);
  or _26704_ (_04400_, _05550_, \oc8051_top_1.oc8051_rom1.data_o [13]);
  nand _26705_ (_04401_, _05550_, _11441_);
  and _26706_ (_04402_, _04401_, _05552_);
  and _26707_ (_04284_, _04402_, _04400_);
  or _26708_ (_04403_, _07668_, _07635_);
  or _26709_ (_04404_, _07670_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and _26710_ (_04405_, _04404_, _05552_);
  and _26711_ (_04295_, _04405_, _04403_);
  or _26712_ (_04406_, _05550_, \oc8051_top_1.oc8051_rom1.data_o [12]);
  nand _26713_ (_04407_, _05550_, _11061_);
  and _26714_ (_04408_, _04407_, _05552_);
  and _26715_ (_04352_, _04408_, _04406_);
  and _26716_ (_04409_, _01515_, _06771_);
  nand _26717_ (_04410_, _04409_, _06763_);
  or _26718_ (_04411_, _04409_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and _26719_ (_04412_, _04411_, _01521_);
  and _26720_ (_04413_, _04412_, _04410_);
  nor _26721_ (_04415_, _01521_, _06811_);
  or _26722_ (_04416_, _04415_, _04413_);
  and _26723_ (_04414_, _04416_, _05552_);
  and _26724_ (_04417_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  not _26725_ (_04418_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  nor _26726_ (_04419_, pc_log_change, _04418_);
  or _26727_ (_04420_, _04419_, _04417_);
  and _26728_ (_04429_, _04420_, _05552_);
  not _26729_ (_04421_, cy_reg);
  and _26730_ (_04422_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and _26731_ (_04423_, _04422_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor _26732_ (_04424_, _04423_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and _26733_ (_04425_, _04423_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _26734_ (_04426_, _04425_, _04424_);
  and _26735_ (_04427_, _04426_, _08302_);
  nor _26736_ (_04428_, _04422_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor _26737_ (_04430_, _04428_, _04423_);
  or _26738_ (_04431_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [4]);
  and _26739_ (_04432_, _04431_, _04422_);
  nand _26740_ (_04433_, _04432_, _04430_);
  nor _26741_ (_04434_, _04433_, _04427_);
  nor _26742_ (_04435_, _04426_, \oc8051_symbolic_cxrom1.regvalid [0]);
  nand _26743_ (_04436_, _04426_, _08796_);
  nand _26744_ (_04437_, _04436_, _04423_);
  nor _26745_ (_04438_, _04437_, _04435_);
  or _26746_ (_04439_, _04438_, _04434_);
  and _26747_ (_04440_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _02500_);
  nand _26748_ (_04441_, _04426_, _08298_);
  or _26749_ (_04442_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [6]);
  and _26750_ (_04443_, _04442_, _04430_);
  and _26751_ (_04444_, _04443_, _04441_);
  not _26752_ (_04445_, _04430_);
  nor _26753_ (_04446_, _04426_, _08424_);
  and _26754_ (_04447_, _04426_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or _26755_ (_04448_, _04447_, _04446_);
  and _26756_ (_04449_, _04448_, _04445_);
  or _26757_ (_04450_, _04449_, _04444_);
  and _26758_ (_04451_, _04450_, _04440_);
  or _26759_ (_04452_, _04451_, _04439_);
  nor _26760_ (_04453_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  or _26761_ (_04454_, _04426_, \oc8051_symbolic_cxrom1.regvalid [5]);
  or _26762_ (_04455_, _02512_, \oc8051_symbolic_cxrom1.regvalid [13]);
  and _26763_ (_04456_, _04455_, _04430_);
  and _26764_ (_04457_, _04456_, _04454_);
  nor _26765_ (_04458_, _04426_, _08276_);
  and _26766_ (_04459_, _04426_, \oc8051_symbolic_cxrom1.regvalid [9]);
  or _26767_ (_04460_, _04459_, _04458_);
  and _26768_ (_04461_, _04460_, _04445_);
  or _26769_ (_04462_, _04461_, _04457_);
  and _26770_ (_04463_, _04462_, _04453_);
  and _26771_ (_04464_, _02505_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  or _26772_ (_04465_, _04426_, \oc8051_symbolic_cxrom1.regvalid [7]);
  or _26773_ (_04466_, _02512_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and _26774_ (_04467_, _04466_, _04430_);
  and _26775_ (_04468_, _04467_, _04465_);
  nor _26776_ (_04469_, _04426_, _08262_);
  and _26777_ (_04470_, _04426_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or _26778_ (_04471_, _04470_, _04469_);
  and _26779_ (_04472_, _04471_, _04445_);
  or _26780_ (_04473_, _04472_, _04468_);
  and _26781_ (_04474_, _04473_, _04464_);
  or _26782_ (_04475_, _04474_, _04463_);
  or _26783_ (_04476_, _04475_, _04452_);
  and _26784_ (_04477_, _04464_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  and _26785_ (_04478_, _04453_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  or _26786_ (_04479_, _04478_, _04477_);
  and _26787_ (_04480_, _04440_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  and _26788_ (_04481_, _04422_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  or _26789_ (_04482_, _04481_, _04480_);
  or _26790_ (_04483_, _04482_, _04479_);
  or _26791_ (_04484_, _04483_, _04445_);
  not _26792_ (_04485_, _04426_);
  and _26793_ (_04486_, _04440_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  and _26794_ (_04487_, _04422_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  or _26795_ (_04488_, _04487_, _04486_);
  and _26796_ (_04489_, _04464_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  and _26797_ (_04491_, _04453_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  or _26798_ (_04492_, _04491_, _04489_);
  or _26799_ (_04493_, _04492_, _04488_);
  or _26800_ (_04494_, _04493_, _04430_);
  and _26801_ (_04495_, _04494_, _04485_);
  and _26802_ (_04496_, _04495_, _04484_);
  and _26803_ (_04497_, _04440_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  and _26804_ (_04498_, _04422_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  or _26805_ (_04499_, _04498_, _04497_);
  and _26806_ (_04500_, _04464_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  and _26807_ (_04501_, _04453_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  or _26808_ (_04502_, _04501_, _04500_);
  or _26809_ (_04503_, _04502_, _04499_);
  or _26810_ (_04504_, _04503_, _04430_);
  and _26811_ (_04505_, _04440_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  and _26812_ (_04506_, _04422_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  or _26813_ (_04507_, _04506_, _04505_);
  and _26814_ (_04508_, _04464_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  and _26815_ (_04509_, _04453_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  or _26816_ (_04510_, _04509_, _04508_);
  or _26817_ (_04511_, _04510_, _04507_);
  or _26818_ (_04512_, _04511_, _04445_);
  and _26819_ (_04513_, _04512_, _04426_);
  and _26820_ (_04514_, _04513_, _04504_);
  or _26821_ (_04515_, _04514_, _04496_);
  and _26822_ (_04516_, _04515_, _04476_);
  and _26823_ (_04517_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and _26824_ (_04518_, _04517_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and _26825_ (_04519_, _04518_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  and _26826_ (_04520_, _04519_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  and _26827_ (_04521_, _04520_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  and _26828_ (_04522_, _04521_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  and _26829_ (_04523_, _04522_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  and _26830_ (_04524_, _04523_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  and _26831_ (_04525_, _04524_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  and _26832_ (_04526_, _04525_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  and _26833_ (_04527_, _04526_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  and _26834_ (_04528_, _04527_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  and _26835_ (_04529_, _04528_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor _26836_ (_04530_, _04528_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor _26837_ (_04531_, _04530_, _04529_);
  and _26838_ (_04532_, _04531_, _04516_);
  nor _26839_ (_04533_, _04526_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor _26840_ (_04534_, _04533_, _04527_);
  and _26841_ (_04535_, _04534_, _04516_);
  and _26842_ (_04536_, _04535_, _02061_);
  nor _26843_ (_04537_, _04527_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  nor _26844_ (_04538_, _04537_, _04528_);
  and _26845_ (_04539_, _04538_, _04516_);
  nor _26846_ (_04540_, _04538_, _04516_);
  nor _26847_ (_04541_, _04540_, _04539_);
  nor _26848_ (_04542_, _04524_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  nor _26849_ (_04543_, _04542_, _04525_);
  and _26850_ (_04544_, _04543_, _04516_);
  and _26851_ (_04545_, _04544_, _02523_);
  nor _26852_ (_04546_, _04525_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  nor _26853_ (_04547_, _04546_, _04526_);
  and _26854_ (_04548_, _04547_, _04516_);
  nor _26855_ (_04549_, _04547_, _04516_);
  nor _26856_ (_04550_, _04549_, _04548_);
  nor _26857_ (_04551_, _04543_, _04516_);
  nor _26858_ (_04552_, _04551_, _04544_);
  not _26859_ (_04553_, _04552_);
  nor _26860_ (_04554_, _04523_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  nor _26861_ (_04555_, _04554_, _04524_);
  and _26862_ (_04556_, _04555_, _04516_);
  nor _26863_ (_04557_, _04522_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor _26864_ (_04558_, _04557_, _04523_);
  and _26865_ (_04559_, _04558_, _04516_);
  nor _26866_ (_04560_, _04555_, _04516_);
  nor _26867_ (_04561_, _04560_, _04556_);
  nor _26868_ (_04562_, _04521_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  nor _26869_ (_04563_, _04562_, _04522_);
  and _26870_ (_04564_, _04563_, _04516_);
  nor _26871_ (_04565_, _04563_, _04516_);
  nor _26872_ (_04566_, _04520_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nor _26873_ (_04567_, _04566_, _04521_);
  and _26874_ (_04568_, _04440_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  and _26875_ (_04569_, _04422_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  or _26876_ (_04570_, _04569_, _04568_);
  and _26877_ (_04572_, _04464_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  and _26878_ (_04573_, _04453_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  or _26879_ (_04574_, _04573_, _04572_);
  or _26880_ (_04575_, _04574_, _04570_);
  or _26881_ (_04576_, _04575_, _04430_);
  and _26882_ (_04577_, _04440_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  and _26883_ (_04578_, _04453_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  or _26884_ (_04579_, _04578_, _04577_);
  and _26885_ (_04580_, _04464_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  and _26886_ (_04581_, _04422_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  or _26887_ (_04582_, _04581_, _04580_);
  or _26888_ (_04583_, _04582_, _04579_);
  or _26889_ (_04584_, _04583_, _04445_);
  and _26890_ (_04585_, _04584_, _04576_);
  or _26891_ (_04586_, _04585_, _04485_);
  and _26892_ (_04587_, _04440_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  and _26893_ (_04588_, _04422_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  or _26894_ (_04589_, _04588_, _04587_);
  and _26895_ (_04590_, _04464_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  and _26896_ (_04591_, _04453_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  or _26897_ (_04592_, _04591_, _04590_);
  or _26898_ (_04593_, _04592_, _04589_);
  or _26899_ (_04594_, _04593_, _04430_);
  and _26900_ (_04595_, _04464_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  and _26901_ (_04596_, _04453_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  or _26902_ (_04597_, _04596_, _04595_);
  and _26903_ (_04598_, _04440_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  and _26904_ (_04599_, _04422_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  or _26905_ (_04600_, _04599_, _04598_);
  or _26906_ (_04601_, _04600_, _04597_);
  or _26907_ (_04602_, _04601_, _04445_);
  and _26908_ (_04603_, _04602_, _04594_);
  or _26909_ (_04604_, _04603_, _04426_);
  and _26910_ (_04605_, _04604_, _04586_);
  and _26911_ (_04606_, _04605_, _04476_);
  and _26912_ (_04607_, _04606_, _04567_);
  nor _26913_ (_04608_, _04606_, _04567_);
  nor _26914_ (_04609_, _04608_, _04607_);
  not _26915_ (_04610_, _04609_);
  and _26916_ (_04611_, _04440_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  and _26917_ (_04612_, _04422_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  or _26918_ (_04613_, _04612_, _04611_);
  and _26919_ (_04614_, _04464_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  and _26920_ (_04615_, _04453_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  or _26921_ (_04616_, _04615_, _04614_);
  or _26922_ (_04617_, _04616_, _04613_);
  or _26923_ (_04618_, _04617_, _04445_);
  and _26924_ (_04619_, _04440_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  and _26925_ (_04620_, _04422_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  or _26926_ (_04621_, _04620_, _04619_);
  and _26927_ (_04622_, _04464_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  and _26928_ (_04623_, _04453_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  or _26929_ (_04624_, _04623_, _04622_);
  or _26930_ (_04625_, _04624_, _04621_);
  or _26931_ (_04626_, _04625_, _04430_);
  and _26932_ (_04627_, _04626_, _04485_);
  and _26933_ (_04628_, _04627_, _04618_);
  and _26934_ (_04629_, _04440_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  and _26935_ (_04630_, _04422_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  or _26936_ (_04631_, _04630_, _04629_);
  and _26937_ (_04632_, _04464_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  and _26938_ (_04633_, _04453_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  or _26939_ (_04634_, _04633_, _04632_);
  or _26940_ (_04635_, _04634_, _04631_);
  or _26941_ (_04636_, _04635_, _04430_);
  and _26942_ (_04637_, _04440_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  and _26943_ (_04638_, _04422_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  or _26944_ (_04639_, _04638_, _04637_);
  and _26945_ (_04640_, _04464_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  and _26946_ (_04641_, _04453_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  or _26947_ (_04642_, _04641_, _04640_);
  or _26948_ (_04643_, _04642_, _04639_);
  or _26949_ (_04644_, _04643_, _04445_);
  and _26950_ (_04645_, _04644_, _04426_);
  and _26951_ (_04646_, _04645_, _04636_);
  or _26952_ (_04647_, _04646_, _04628_);
  and _26953_ (_04648_, _04647_, _04476_);
  nor _26954_ (_04649_, _04519_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  nor _26955_ (_04650_, _04649_, _04520_);
  and _26956_ (_04651_, _04650_, _04648_);
  nor _26957_ (_04652_, _04650_, _04648_);
  nor _26958_ (_04653_, _04652_, _04651_);
  not _26959_ (_04654_, _04653_);
  nor _26960_ (_04655_, _04518_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nor _26961_ (_04656_, _04655_, _04519_);
  and _26962_ (_04657_, _04464_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  and _26963_ (_04658_, _04453_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  or _26964_ (_04659_, _04658_, _04657_);
  and _26965_ (_04660_, _04440_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  and _26966_ (_04661_, _04422_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  or _26967_ (_04662_, _04661_, _04660_);
  or _26968_ (_04663_, _04662_, _04659_);
  or _26969_ (_04664_, _04663_, _04445_);
  and _26970_ (_04665_, _04440_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  and _26971_ (_04666_, _04422_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  or _26972_ (_04667_, _04666_, _04665_);
  and _26973_ (_04668_, _04464_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  and _26974_ (_04669_, _04453_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  or _26975_ (_04670_, _04669_, _04668_);
  or _26976_ (_04671_, _04670_, _04667_);
  or _26977_ (_04672_, _04671_, _04430_);
  and _26978_ (_04673_, _04672_, _04485_);
  and _26979_ (_04674_, _04673_, _04664_);
  and _26980_ (_04675_, _04440_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  and _26981_ (_04676_, _04422_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  or _26982_ (_04677_, _04676_, _04675_);
  and _26983_ (_04678_, _04464_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  and _26984_ (_04679_, _04453_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  or _26985_ (_04680_, _04679_, _04678_);
  or _26986_ (_04681_, _04680_, _04677_);
  or _26987_ (_04682_, _04681_, _04430_);
  and _26988_ (_04683_, _04440_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  and _26989_ (_04684_, _04422_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  or _26990_ (_04685_, _04684_, _04683_);
  and _26991_ (_04686_, _04464_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  and _26992_ (_04687_, _04453_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  or _26993_ (_04688_, _04687_, _04686_);
  or _26994_ (_04689_, _04688_, _04685_);
  or _26995_ (_04690_, _04689_, _04445_);
  and _26996_ (_04691_, _04690_, _04426_);
  and _26997_ (_04692_, _04691_, _04682_);
  or _26998_ (_04693_, _04692_, _04674_);
  and _26999_ (_04694_, _04693_, _04476_);
  and _27000_ (_04695_, _04694_, _04656_);
  nor _27001_ (_04696_, _04517_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _27002_ (_04697_, _04696_, _04518_);
  and _27003_ (_04698_, _04464_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  and _27004_ (_04699_, _04453_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  or _27005_ (_04700_, _04699_, _04698_);
  and _27006_ (_04701_, _04440_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  and _27007_ (_04702_, _04422_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  or _27008_ (_04703_, _04702_, _04701_);
  or _27009_ (_04704_, _04703_, _04700_);
  or _27010_ (_04705_, _04704_, _04445_);
  and _27011_ (_04706_, _04440_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  and _27012_ (_04707_, _04422_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  or _27013_ (_04708_, _04707_, _04706_);
  and _27014_ (_04709_, _04464_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  and _27015_ (_04710_, _04453_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  or _27016_ (_04711_, _04710_, _04709_);
  or _27017_ (_04712_, _04711_, _04708_);
  or _27018_ (_04713_, _04712_, _04430_);
  and _27019_ (_04714_, _04713_, _04485_);
  and _27020_ (_04715_, _04714_, _04705_);
  and _27021_ (_04716_, _04440_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  and _27022_ (_04717_, _04422_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  or _27023_ (_04718_, _04717_, _04716_);
  and _27024_ (_04719_, _04464_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  and _27025_ (_04720_, _04453_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  or _27026_ (_04721_, _04720_, _04719_);
  or _27027_ (_04722_, _04721_, _04718_);
  or _27028_ (_04723_, _04722_, _04430_);
  and _27029_ (_04724_, _04440_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  and _27030_ (_04725_, _04422_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  or _27031_ (_04726_, _04725_, _04724_);
  and _27032_ (_04727_, _04464_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  and _27033_ (_04728_, _04453_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  or _27034_ (_04729_, _04728_, _04727_);
  or _27035_ (_04730_, _04729_, _04726_);
  or _27036_ (_04731_, _04730_, _04445_);
  and _27037_ (_04732_, _04731_, _04426_);
  and _27038_ (_04733_, _04732_, _04723_);
  or _27039_ (_04734_, _04733_, _04715_);
  and _27040_ (_04735_, _04734_, _04476_);
  and _27041_ (_04736_, _04735_, _04697_);
  nor _27042_ (_04737_, _04735_, _04697_);
  and _27043_ (_04738_, _02500_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and _27044_ (_04739_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _01920_);
  nor _27045_ (_04740_, _04739_, _04738_);
  not _27046_ (_04741_, _04740_);
  and _27047_ (_04742_, _04440_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  and _27048_ (_04743_, _04422_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  or _27049_ (_04744_, _04743_, _04742_);
  and _27050_ (_04745_, _04464_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  and _27051_ (_04746_, _04453_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  or _27052_ (_04747_, _04746_, _04745_);
  or _27053_ (_04748_, _04747_, _04744_);
  or _27054_ (_04749_, _04748_, _04430_);
  and _27055_ (_04750_, _04464_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  and _27056_ (_04751_, _04453_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  or _27057_ (_04752_, _04751_, _04750_);
  and _27058_ (_04753_, _04440_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  and _27059_ (_04754_, _04422_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  or _27060_ (_04755_, _04754_, _04753_);
  or _27061_ (_04756_, _04755_, _04752_);
  or _27062_ (_04757_, _04756_, _04445_);
  and _27063_ (_04758_, _04757_, _04749_);
  or _27064_ (_04759_, _04758_, _04485_);
  and _27065_ (_04760_, _04464_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  and _27066_ (_04761_, _04453_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  or _27067_ (_04762_, _04761_, _04760_);
  and _27068_ (_04763_, _04440_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  and _27069_ (_04764_, _04422_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  or _27070_ (_04765_, _04764_, _04763_);
  or _27071_ (_04766_, _04765_, _04762_);
  or _27072_ (_04767_, _04766_, _04430_);
  and _27073_ (_04768_, _04464_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  and _27074_ (_04769_, _04453_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  or _27075_ (_04770_, _04769_, _04768_);
  and _27076_ (_04771_, _04440_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  and _27077_ (_04772_, _04422_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  or _27078_ (_04773_, _04772_, _04771_);
  or _27079_ (_04774_, _04773_, _04770_);
  or _27080_ (_04775_, _04774_, _04445_);
  and _27081_ (_04776_, _04775_, _04767_);
  or _27082_ (_04777_, _04776_, _04426_);
  and _27083_ (_04778_, _04777_, _04759_);
  and _27084_ (_04779_, _04778_, _04476_);
  and _27085_ (_04780_, _04779_, _04741_);
  and _27086_ (_04781_, _04464_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  and _27087_ (_04782_, _04453_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  or _27088_ (_04783_, _04782_, _04781_);
  and _27089_ (_04784_, _04440_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  and _27090_ (_04785_, _04422_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  or _27091_ (_04786_, _04785_, _04784_);
  or _27092_ (_04787_, _04786_, _04783_);
  or _27093_ (_04788_, _04787_, _04445_);
  and _27094_ (_04789_, _04440_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  and _27095_ (_04790_, _04422_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  or _27096_ (_04791_, _04790_, _04789_);
  and _27097_ (_04792_, _04464_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  and _27098_ (_04793_, _04453_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  or _27099_ (_04794_, _04793_, _04792_);
  or _27100_ (_04795_, _04794_, _04791_);
  or _27101_ (_04796_, _04795_, _04430_);
  and _27102_ (_04797_, _04796_, _04485_);
  and _27103_ (_04798_, _04797_, _04788_);
  and _27104_ (_04799_, _04440_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  and _27105_ (_04800_, _04422_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  or _27106_ (_04801_, _04800_, _04799_);
  and _27107_ (_04802_, _04464_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  and _27108_ (_04803_, _04453_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  or _27109_ (_04804_, _04803_, _04802_);
  or _27110_ (_04805_, _04804_, _04801_);
  or _27111_ (_04806_, _04805_, _04430_);
  and _27112_ (_04807_, _04440_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  and _27113_ (_04808_, _04422_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  or _27114_ (_04809_, _04808_, _04807_);
  and _27115_ (_04810_, _04464_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  and _27116_ (_04811_, _04453_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  or _27117_ (_04812_, _04811_, _04810_);
  or _27118_ (_04813_, _04812_, _04809_);
  or _27119_ (_04814_, _04813_, _04445_);
  and _27120_ (_04815_, _04814_, _04426_);
  and _27121_ (_04816_, _04815_, _04806_);
  or _27122_ (_04817_, _04816_, _04798_);
  and _27123_ (_04818_, _04817_, _04476_);
  and _27124_ (_04819_, _04818_, _02500_);
  and _27125_ (_04820_, _04440_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and _27126_ (_04821_, _04422_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  or _27127_ (_04822_, _04821_, _04820_);
  and _27128_ (_04823_, _04464_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and _27129_ (_04824_, _04453_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  or _27130_ (_04825_, _04824_, _04823_);
  or _27131_ (_04826_, _04825_, _04822_);
  or _27132_ (_04827_, _04826_, _04430_);
  and _27133_ (_04828_, _04440_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and _27134_ (_04829_, _04422_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  or _27135_ (_04830_, _04829_, _04828_);
  and _27136_ (_04831_, _04464_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  and _27137_ (_04832_, _04453_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  or _27138_ (_04833_, _04832_, _04831_);
  or _27139_ (_04834_, _04833_, _04830_);
  or _27140_ (_04835_, _04834_, _04445_);
  and _27141_ (_04836_, _04835_, _04827_);
  or _27142_ (_04837_, _04836_, _04485_);
  and _27143_ (_04838_, _04440_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  and _27144_ (_04839_, _04422_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  or _27145_ (_04840_, _04839_, _04838_);
  and _27146_ (_04841_, _04464_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  and _27147_ (_04842_, _04453_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  or _27148_ (_04843_, _04842_, _04841_);
  or _27149_ (_04844_, _04843_, _04840_);
  or _27150_ (_04845_, _04844_, _04445_);
  and _27151_ (_04846_, _04464_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  and _27152_ (_04847_, _04453_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  or _27153_ (_04848_, _04847_, _04846_);
  and _27154_ (_04849_, _04440_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  and _27155_ (_04850_, _04422_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  or _27156_ (_04851_, _04850_, _04849_);
  or _27157_ (_04852_, _04851_, _04848_);
  or _27158_ (_04853_, _04852_, _04430_);
  and _27159_ (_04854_, _04853_, _04845_);
  or _27160_ (_04855_, _04854_, _04426_);
  and _27161_ (_04856_, _04855_, _04837_);
  and _27162_ (_04857_, _04856_, _04476_);
  and _27163_ (_04858_, _04857_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _27164_ (_04859_, _04818_, _02500_);
  nor _27165_ (_04860_, _04859_, _04819_);
  and _27166_ (_04861_, _04860_, _04858_);
  nor _27167_ (_04862_, _04861_, _04819_);
  nor _27168_ (_04863_, _04779_, _04741_);
  nor _27169_ (_04864_, _04863_, _04780_);
  not _27170_ (_04865_, _04864_);
  nor _27171_ (_04866_, _04865_, _04862_);
  nor _27172_ (_04867_, _04866_, _04780_);
  nor _27173_ (_04868_, _04867_, _04737_);
  nor _27174_ (_04869_, _04868_, _04736_);
  nor _27175_ (_04870_, _04694_, _04656_);
  nor _27176_ (_04871_, _04870_, _04695_);
  not _27177_ (_04872_, _04871_);
  nor _27178_ (_04873_, _04872_, _04869_);
  nor _27179_ (_04874_, _04873_, _04695_);
  nor _27180_ (_04875_, _04874_, _04654_);
  nor _27181_ (_04876_, _04875_, _04651_);
  nor _27182_ (_04877_, _04876_, _04610_);
  nor _27183_ (_04878_, _04877_, _04607_);
  nor _27184_ (_04879_, _04878_, _04565_);
  or _27185_ (_04880_, _04879_, _04564_);
  nor _27186_ (_04881_, _04558_, _04516_);
  nor _27187_ (_04882_, _04881_, _04559_);
  and _27188_ (_04883_, _04882_, _04880_);
  and _27189_ (_04884_, _04883_, _04561_);
  or _27190_ (_04885_, _04884_, _04559_);
  nor _27191_ (_04886_, _04885_, _04556_);
  nor _27192_ (_04887_, _04886_, _04553_);
  and _27193_ (_04888_, _04887_, _04550_);
  or _27194_ (_04889_, _04888_, _04548_);
  nor _27195_ (_04890_, _04889_, _04545_);
  nor _27196_ (_04891_, _04534_, _04516_);
  nor _27197_ (_04892_, _04891_, _04535_);
  not _27198_ (_04893_, _04892_);
  nor _27199_ (_04894_, _04893_, _04890_);
  and _27200_ (_04895_, _04894_, _04541_);
  or _27201_ (_04896_, _04895_, _04539_);
  nor _27202_ (_04897_, _04896_, _04536_);
  nor _27203_ (_04898_, _04531_, _04516_);
  nor _27204_ (_04899_, _04898_, _04532_);
  not _27205_ (_04900_, _04899_);
  nor _27206_ (_04901_, _04900_, _04897_);
  nor _27207_ (_04902_, _04901_, _04532_);
  nor _27208_ (_04903_, _04529_, _04418_);
  and _27209_ (_04904_, _04529_, _04418_);
  or _27210_ (_04905_, _04904_, _04903_);
  and _27211_ (_04906_, _04905_, _04516_);
  nor _27212_ (_04907_, _04905_, _04516_);
  nor _27213_ (_04908_, _04907_, _04906_);
  nor _27214_ (_04909_, _04908_, _04902_);
  and _27215_ (_04910_, _04908_, _04902_);
  or _27216_ (_04911_, _04910_, _04909_);
  nor _27217_ (_04912_, _04911_, _04421_);
  nor _27218_ (_04913_, _04905_, cy_reg);
  nor _27219_ (_04914_, _04913_, _04912_);
  nor _27220_ (_04915_, _04914_, _02697_);
  and _27221_ (_04916_, _04914_, _02697_);
  or _27222_ (_04917_, _04916_, _04915_);
  nor _27223_ (_04918_, _04894_, _04535_);
  and _27224_ (_04919_, _04918_, _04541_);
  nor _27225_ (_04920_, _04918_, _04541_);
  nor _27226_ (_04921_, _04920_, _04919_);
  nor _27227_ (_04922_, _04921_, _04421_);
  and _27228_ (_04923_, _04538_, _04421_);
  nor _27229_ (_04924_, _04923_, _04922_);
  nor _27230_ (_04925_, _04924_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and _27231_ (_04926_, _04924_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nor _27232_ (_04927_, _04547_, cy_reg);
  nor _27233_ (_04928_, _04887_, _04544_);
  nor _27234_ (_04929_, _04928_, _04550_);
  and _27235_ (_04930_, _04928_, _04550_);
  or _27236_ (_04931_, _04930_, _04929_);
  nor _27237_ (_04932_, _04931_, _04421_);
  nor _27238_ (_04933_, _04932_, _04927_);
  and _27239_ (_04934_, _04933_, _01924_);
  nor _27240_ (_04935_, _04933_, _01924_);
  and _27241_ (_04936_, _04555_, _04421_);
  nor _27242_ (_04937_, _04883_, _04559_);
  and _27243_ (_04938_, _04937_, _04561_);
  nor _27244_ (_04939_, _04937_, _04561_);
  nor _27245_ (_04940_, _04939_, _04938_);
  nor _27246_ (_04941_, _04940_, _04421_);
  nor _27247_ (_04942_, _04941_, _04936_);
  nor _27248_ (_04943_, _04942_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and _27249_ (_04944_, _04942_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nor _27250_ (_04945_, _04563_, cy_reg);
  nor _27251_ (_04946_, _04564_, _04565_);
  and _27252_ (_04947_, _04946_, _04878_);
  nor _27253_ (_04948_, _04946_, _04878_);
  or _27254_ (_04949_, _04948_, _04947_);
  nor _27255_ (_04950_, _04949_, _04421_);
  nor _27256_ (_04951_, _04950_, _04945_);
  nor _27257_ (_04952_, _04951_, _02415_);
  and _27258_ (_04953_, _04951_, _02415_);
  and _27259_ (_04954_, _04567_, _04421_);
  and _27260_ (_04955_, _04876_, _04610_);
  nor _27261_ (_04956_, _04955_, _04877_);
  and _27262_ (_04957_, _04956_, cy_reg);
  nor _27263_ (_04958_, _04957_, _04954_);
  and _27264_ (_04959_, _04958_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  nor _27265_ (_04960_, _04958_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  and _27266_ (_04961_, _04650_, _04421_);
  and _27267_ (_04962_, _04874_, _04654_);
  nor _27268_ (_04963_, _04962_, _04875_);
  and _27269_ (_04964_, _04963_, cy_reg);
  nor _27270_ (_04965_, _04964_, _04961_);
  and _27271_ (_04966_, _04965_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nor _27272_ (_04967_, _04965_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  and _27273_ (_04968_, _04656_, _04421_);
  and _27274_ (_04969_, _04872_, _04869_);
  nor _27275_ (_04970_, _04969_, _04873_);
  and _27276_ (_04971_, _04970_, cy_reg);
  nor _27277_ (_04972_, _04971_, _04968_);
  and _27278_ (_04973_, _04972_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  nor _27279_ (_04974_, _04697_, cy_reg);
  nor _27280_ (_04975_, _04737_, _04736_);
  nor _27281_ (_04976_, _04975_, _04867_);
  and _27282_ (_04977_, _04975_, _04867_);
  or _27283_ (_04978_, _04977_, _04976_);
  nor _27284_ (_04979_, _04978_, _04421_);
  nor _27285_ (_04980_, _04979_, _04974_);
  nor _27286_ (_04981_, _04980_, _02406_);
  and _27287_ (_04982_, _04980_, _02406_);
  nor _27288_ (_04983_, _04740_, cy_reg);
  and _27289_ (_04984_, _04865_, _04862_);
  nor _27290_ (_04985_, _04984_, _04866_);
  and _27291_ (_04986_, _04985_, cy_reg);
  nor _27292_ (_04987_, _04986_, _04983_);
  and _27293_ (_04988_, _04987_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and _27294_ (_04989_, _04857_, cy_reg);
  not _27295_ (_04990_, _04989_);
  nor _27296_ (_04991_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _27297_ (_04992_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _27298_ (_04993_, _04992_, _04991_);
  nor _27299_ (_04994_, _04993_, _04990_);
  and _27300_ (_04995_, _04993_, _04990_);
  or _27301_ (_04996_, _04995_, _04994_);
  nor _27302_ (_04997_, cy_reg, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nor _27303_ (_04998_, _04860_, _04858_);
  nor _27304_ (_04999_, _04998_, _04861_);
  and _27305_ (_05000_, _04999_, cy_reg);
  nor _27306_ (_05001_, _05000_, _04997_);
  nor _27307_ (_05002_, _05001_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and _27308_ (_05003_, _05001_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  or _27309_ (_05004_, _05003_, _05002_);
  or _27310_ (_05005_, _05004_, _04996_);
  nor _27311_ (_05006_, _04987_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or _27312_ (_05007_, _05006_, _05005_);
  or _27313_ (_05008_, _05007_, _04988_);
  or _27314_ (_05009_, _05008_, _04982_);
  or _27315_ (_05010_, _05009_, _04981_);
  nor _27316_ (_05011_, _04972_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  or _27317_ (_05012_, _05011_, _05010_);
  or _27318_ (_05013_, _05012_, _04973_);
  or _27319_ (_05014_, _05013_, _04967_);
  or _27320_ (_05015_, _05014_, _04966_);
  or _27321_ (_05016_, _05015_, _04960_);
  or _27322_ (_05017_, _05016_, _04959_);
  or _27323_ (_05018_, _05017_, _04953_);
  or _27324_ (_05019_, _05018_, _04952_);
  and _27325_ (_05020_, _04558_, _04421_);
  nor _27326_ (_05021_, _04882_, _04880_);
  nor _27327_ (_05022_, _05021_, _04883_);
  and _27328_ (_05023_, _05022_, cy_reg);
  nor _27329_ (_05024_, _05023_, _05020_);
  nor _27330_ (_05025_, _05024_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  and _27331_ (_05026_, _05024_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  or _27332_ (_05027_, _05026_, _05025_);
  or _27333_ (_05028_, _05027_, _05019_);
  or _27334_ (_05029_, _05028_, _04944_);
  or _27335_ (_05030_, _05029_, _04943_);
  and _27336_ (_05031_, _04543_, _04421_);
  and _27337_ (_05032_, _04886_, _04553_);
  nor _27338_ (_05033_, _05032_, _04887_);
  and _27339_ (_05034_, _05033_, cy_reg);
  nor _27340_ (_05035_, _05034_, _05031_);
  and _27341_ (_05036_, _05035_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nor _27342_ (_05037_, _05035_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  or _27343_ (_05038_, _05037_, _05036_);
  or _27344_ (_05039_, _05038_, _05030_);
  or _27345_ (_05040_, _05039_, _04935_);
  or _27346_ (_05041_, _05040_, _04934_);
  and _27347_ (_05042_, _04534_, _04421_);
  and _27348_ (_05043_, _04893_, _04890_);
  nor _27349_ (_05044_, _05043_, _04894_);
  and _27350_ (_05045_, _05044_, cy_reg);
  nor _27351_ (_05046_, _05045_, _05042_);
  and _27352_ (_05047_, _05046_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nor _27353_ (_05048_, _05046_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  or _27354_ (_05049_, _05048_, _05047_);
  or _27355_ (_05050_, _05049_, _05041_);
  or _27356_ (_05051_, _05050_, _04926_);
  or _27357_ (_05052_, _05051_, _04925_);
  and _27358_ (_05053_, _04531_, _04421_);
  and _27359_ (_05054_, _04900_, _04897_);
  nor _27360_ (_05055_, _05054_, _04901_);
  and _27361_ (_05056_, _05055_, cy_reg);
  nor _27362_ (_05057_, _05056_, _05053_);
  and _27363_ (_05058_, _05057_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nor _27364_ (_05059_, _05057_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  or _27365_ (_05060_, _05059_, _05058_);
  or _27366_ (_05061_, _05060_, _05052_);
  or _27367_ (_05062_, _05061_, _04917_);
  nor _27368_ (_05063_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor _27369_ (_05064_, _05063_, _02410_);
  nor _27370_ (_05065_, _05064_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _27371_ (_05066_, _05064_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor _27372_ (_05067_, _05066_, _05065_);
  or _27373_ (_05068_, _01960_, \oc8051_symbolic_cxrom1.regvalid [2]);
  or _27374_ (_05069_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_symbolic_cxrom1.regvalid [0]);
  and _27375_ (_05070_, _05069_, _05068_);
  or _27376_ (_05071_, _05070_, _05067_);
  and _27377_ (_05072_, _05063_, _02410_);
  nor _27378_ (_05073_, _05072_, _05064_);
  not _27379_ (_05074_, _05073_);
  or _27380_ (_05075_, _01960_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or _27381_ (_05076_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_symbolic_cxrom1.regvalid [8]);
  nand _27382_ (_05077_, _05076_, _05075_);
  nand _27383_ (_05078_, _05077_, _05067_);
  and _27384_ (_05079_, _05078_, _05074_);
  and _27385_ (_05080_, _05079_, _05071_);
  and _27386_ (_05081_, _05067_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and _27387_ (_05082_, _02406_, \oc8051_symbolic_cxrom1.regvalid [4]);
  or _27388_ (_05083_, _05082_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  or _27389_ (_05084_, _05083_, _05081_);
  and _27390_ (_05085_, _05067_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and _27391_ (_05086_, _02406_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or _27392_ (_05087_, _05086_, _01960_);
  or _27393_ (_05088_, _05087_, _05085_);
  and _27394_ (_05089_, _05088_, _05073_);
  and _27395_ (_05090_, _05089_, _05084_);
  or _27396_ (_05091_, _05090_, _05080_);
  and _27397_ (_05092_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and _27398_ (_05093_, _05092_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor _27399_ (_05094_, _05092_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor _27400_ (_05095_, _05094_, _05093_);
  not _27401_ (_05096_, _05095_);
  nor _27402_ (_05097_, _05093_, _02406_);
  and _27403_ (_05098_, _05093_, _02406_);
  nor _27404_ (_05099_, _05098_, _05097_);
  or _27405_ (_05100_, _05099_, \oc8051_symbolic_cxrom1.regvalid [14]);
  or _27406_ (_05101_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [6]);
  and _27407_ (_05102_, _05101_, _05100_);
  or _27408_ (_05103_, _05102_, _05096_);
  nand _27409_ (_05104_, _05099_, _08424_);
  or _27410_ (_05105_, _05099_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and _27411_ (_05106_, _05105_, _05104_);
  or _27412_ (_05107_, _05106_, _05095_);
  and _27413_ (_05108_, _05107_, _05103_);
  or _27414_ (_05109_, _05108_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor _27415_ (_05110_, _05099_, _08796_);
  and _27416_ (_05111_, _05099_, \oc8051_symbolic_cxrom1.regvalid [0]);
  or _27417_ (_05112_, _05111_, _05110_);
  and _27418_ (_05113_, _05112_, _05096_);
  or _27419_ (_05114_, _05099_, \oc8051_symbolic_cxrom1.regvalid [12]);
  or _27420_ (_05115_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [4]);
  and _27421_ (_05116_, _05115_, _05095_);
  and _27422_ (_05117_, _05116_, _05114_);
  or _27423_ (_05118_, _05117_, _01960_);
  or _27424_ (_05119_, _05118_, _05113_);
  and _27425_ (_05120_, _02406_, \oc8051_symbolic_cxrom1.regvalid [7]);
  and _27426_ (_05121_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [15]);
  or _27427_ (_05122_, _05121_, _05120_);
  and _27428_ (_05123_, _05122_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or _27429_ (_05124_, _02406_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or _27430_ (_05125_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [3]);
  and _27431_ (_05126_, _05125_, _02410_);
  and _27432_ (_05127_, _05126_, _05124_);
  or _27433_ (_05128_, _05127_, _05123_);
  and _27434_ (_05129_, _05128_, _05092_);
  and _27435_ (_05130_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0], _01960_);
  or _27436_ (_05131_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [5]);
  or _27437_ (_05132_, _02406_, \oc8051_symbolic_cxrom1.regvalid [13]);
  and _27438_ (_05133_, _05132_, _05131_);
  or _27439_ (_05134_, _05133_, _02410_);
  or _27440_ (_05135_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [1]);
  or _27441_ (_05136_, _02406_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and _27442_ (_05137_, _05136_, _05135_);
  or _27443_ (_05138_, _05137_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and _27444_ (_05139_, _05138_, _05134_);
  and _27445_ (_05140_, _05139_, _05130_);
  or _27446_ (_05141_, _05140_, _05129_);
  and _27447_ (_05143_, _05128_, _01960_);
  or _27448_ (_05144_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [9]);
  and _27449_ (_05145_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or _27450_ (_05146_, _02406_, \oc8051_symbolic_cxrom1.regvalid [1]);
  and _27451_ (_05147_, _05146_, _05145_);
  and _27452_ (_05148_, _05147_, _05144_);
  and _27453_ (_05149_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], _02410_);
  and _27454_ (_05150_, _05149_, _05133_);
  or _27455_ (_05151_, _05150_, _05148_);
  or _27456_ (_05152_, _05151_, _05143_);
  and _27457_ (_05153_, _05152_, _05141_);
  and _27458_ (_05154_, _05153_, _05119_);
  and _27459_ (_05155_, _05154_, _05109_);
  and _27460_ (_05156_, _05155_, _05091_);
  and _27461_ (_05157_, _05067_, \oc8051_symbolic_cxrom1.regvalid [15]);
  or _27462_ (_05158_, _05120_, _05074_);
  or _27463_ (_05159_, _05158_, _05157_);
  and _27464_ (_05160_, _05159_, _01960_);
  nor _27465_ (_05161_, _05067_, _08262_);
  and _27466_ (_05162_, _05067_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or _27467_ (_05163_, _05162_, _05161_);
  or _27468_ (_05164_, _05163_, _05073_);
  and _27469_ (_05165_, _05164_, _05160_);
  or _27470_ (_05166_, _05165_, _05151_);
  and _27471_ (_05167_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [8]);
  and _27472_ (_05168_, _02406_, \oc8051_symbolic_cxrom1.regvalid [0]);
  or _27473_ (_05169_, _05168_, _05167_);
  and _27474_ (_05170_, _05169_, _02410_);
  and _27475_ (_05171_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [12]);
  or _27476_ (_05172_, _05171_, _05082_);
  and _27477_ (_05173_, _05172_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or _27478_ (_05174_, _05173_, _05170_);
  and _27479_ (_05175_, _05174_, _01960_);
  or _27480_ (_05176_, _05099_, \oc8051_symbolic_cxrom1.regvalid [13]);
  and _27481_ (_05177_, _05131_, _05095_);
  and _27482_ (_05178_, _05177_, _05176_);
  or _27483_ (_05179_, _05099_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nand _27484_ (_05180_, _05099_, _08276_);
  and _27485_ (_05181_, _05180_, _05096_);
  and _27486_ (_05182_, _05181_, _05179_);
  or _27487_ (_05183_, _05182_, _05178_);
  and _27488_ (_05184_, _05183_, _05175_);
  or _27489_ (_05185_, _05099_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nand _27490_ (_05186_, _05099_, _08262_);
  and _27491_ (_05187_, _05186_, _05096_);
  and _27492_ (_05188_, _05187_, _05185_);
  or _27493_ (_05189_, _05099_, \oc8051_symbolic_cxrom1.regvalid [15]);
  or _27494_ (_05190_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [7]);
  and _27495_ (_05191_, _05190_, _05095_);
  and _27496_ (_05192_, _05191_, _05189_);
  or _27497_ (_05193_, _05192_, _05188_);
  and _27498_ (_05194_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [14]);
  or _27499_ (_05195_, _05086_, _02410_);
  or _27500_ (_05196_, _05195_, _05194_);
  or _27501_ (_05197_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [2]);
  or _27502_ (_05198_, _02406_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and _27503_ (_05199_, _05198_, _05197_);
  or _27504_ (_05200_, _05199_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and _27505_ (_05201_, _05200_, _05196_);
  and _27506_ (_05202_, _05201_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and _27507_ (_05203_, _05172_, _05149_);
  or _27508_ (_05204_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [8]);
  or _27509_ (_05205_, _02406_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and _27510_ (_05206_, _05205_, _05145_);
  and _27511_ (_05207_, _05206_, _05204_);
  or _27512_ (_05208_, _05207_, _05203_);
  and _27513_ (_05209_, _05208_, _05202_);
  and _27514_ (_05210_, _05209_, _05193_);
  or _27515_ (_05211_, _05210_, _05184_);
  or _27516_ (_05212_, _05208_, _05201_);
  and _27517_ (_05213_, _05212_, _02402_);
  and _27518_ (_05214_, _05213_, _05211_);
  and _27519_ (_05215_, _05214_, _05166_);
  or _27520_ (_05216_, _05215_, _05156_);
  nor _27521_ (_05217_, _04453_, _01920_);
  nor _27522_ (_05218_, _05217_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and _27523_ (_05219_, _05217_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _27524_ (_05220_, _05219_, _05218_);
  nand _27525_ (_05221_, _05220_, _08298_);
  nor _27526_ (_05222_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and _27527_ (_05223_, _05222_, _02505_);
  nor _27528_ (_05224_, _05223_, _05217_);
  and _27529_ (_05225_, _05224_, _04442_);
  and _27530_ (_05226_, _05225_, _05221_);
  not _27531_ (_05227_, _05224_);
  and _27532_ (_05228_, _05220_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor _27533_ (_05229_, _05220_, _08424_);
  or _27534_ (_05230_, _05229_, _05228_);
  and _27535_ (_05231_, _05230_, _05227_);
  or _27536_ (_05232_, _05231_, _05226_);
  and _27537_ (_05233_, _05232_, _04422_);
  nand _27538_ (_05234_, _05220_, _08967_);
  or _27539_ (_05235_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [5]);
  and _27540_ (_05236_, _05235_, _05224_);
  and _27541_ (_05237_, _05236_, _05234_);
  and _27542_ (_05238_, _05220_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor _27543_ (_05239_, _05220_, _08276_);
  or _27544_ (_05240_, _05239_, _05238_);
  and _27545_ (_05241_, _05240_, _05227_);
  or _27546_ (_05242_, _05241_, _05237_);
  and _27547_ (_05243_, _05242_, _04464_);
  or _27548_ (_05244_, _05243_, _05233_);
  nand _27549_ (_05245_, _05220_, _08270_);
  or _27550_ (_05246_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [7]);
  and _27551_ (_05247_, _05246_, _05224_);
  and _27552_ (_05248_, _05247_, _05245_);
  and _27553_ (_05249_, _05220_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor _27554_ (_05250_, _05220_, _08262_);
  or _27555_ (_05251_, _05250_, _05249_);
  and _27556_ (_05252_, _05251_, _05227_);
  or _27557_ (_05253_, _05252_, _05248_);
  and _27558_ (_05254_, _05253_, _04453_);
  nand _27559_ (_05255_, _05220_, _08302_);
  and _27560_ (_05256_, _05224_, _04431_);
  and _27561_ (_05257_, _05256_, _05255_);
  and _27562_ (_05258_, _05220_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor _27563_ (_05259_, _05220_, _08293_);
  or _27564_ (_05260_, _05259_, _05258_);
  and _27565_ (_05261_, _05260_, _05227_);
  or _27566_ (_05262_, _05261_, _05257_);
  and _27567_ (_05263_, _05262_, _04440_);
  or _27568_ (_05264_, _05263_, _05254_);
  or _27569_ (_05265_, _05264_, _05244_);
  not _27570_ (_05266_, _04422_);
  nor _27571_ (_05267_, \oc8051_symbolic_cxrom1.regarray[11] [3], \oc8051_symbolic_cxrom1.regarray[11] [2]);
  nor _27572_ (_05268_, \oc8051_symbolic_cxrom1.regarray[11] [1], \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and _27573_ (_05269_, _05268_, _05267_);
  or _27574_ (_05270_, _05269_, _05266_);
  nor _27575_ (_05271_, \oc8051_symbolic_cxrom1.regarray[9] [1], \oc8051_symbolic_cxrom1.regarray[9] [0]);
  nor _27576_ (_05272_, \oc8051_symbolic_cxrom1.regarray[9] [3], \oc8051_symbolic_cxrom1.regarray[9] [2]);
  nand _27577_ (_05273_, _05272_, _05271_);
  nand _27578_ (_05274_, _05273_, _04440_);
  and _27579_ (_05275_, _05274_, _05270_);
  nor _27580_ (_05276_, \oc8051_symbolic_cxrom1.regarray[10] [1], \oc8051_symbolic_cxrom1.regarray[10] [0]);
  nor _27581_ (_05277_, \oc8051_symbolic_cxrom1.regarray[10] [3], \oc8051_symbolic_cxrom1.regarray[10] [2]);
  nand _27582_ (_05278_, _05277_, _05276_);
  nand _27583_ (_05279_, _05278_, _04464_);
  not _27584_ (_05280_, _04453_);
  nor _27585_ (_05281_, \oc8051_symbolic_cxrom1.regarray[8] [1], \oc8051_symbolic_cxrom1.regarray[8] [0]);
  nor _27586_ (_05282_, \oc8051_symbolic_cxrom1.regarray[8] [3], \oc8051_symbolic_cxrom1.regarray[8] [2]);
  and _27587_ (_05283_, _05282_, _05281_);
  or _27588_ (_05284_, _05283_, _05280_);
  and _27589_ (_05285_, _05284_, _05279_);
  and _27590_ (_05286_, _05285_, _05275_);
  and _27591_ (_05287_, _04422_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  and _27592_ (_05288_, _04464_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  or _27593_ (_05289_, _05288_, _05287_);
  and _27594_ (_05290_, _04453_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  and _27595_ (_05291_, _04440_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  or _27596_ (_05292_, _05291_, _05290_);
  or _27597_ (_05293_, _05292_, _05289_);
  nand _27598_ (_05294_, _04464_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  nand _27599_ (_05295_, _04440_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  and _27600_ (_05296_, _05295_, _05294_);
  nand _27601_ (_05297_, _04422_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  nand _27602_ (_05298_, _04453_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  and _27603_ (_05299_, _05298_, _05297_);
  and _27604_ (_05300_, _05299_, _05296_);
  or _27605_ (_05301_, \oc8051_symbolic_cxrom1.regarray[9] [5], \oc8051_symbolic_cxrom1.regarray[9] [4]);
  nand _27606_ (_05302_, _05301_, _04440_);
  or _27607_ (_05303_, \oc8051_symbolic_cxrom1.regarray[10] [5], \oc8051_symbolic_cxrom1.regarray[10] [4]);
  nand _27608_ (_05304_, _05303_, _04464_);
  and _27609_ (_05305_, _05304_, _05302_);
  or _27610_ (_05306_, \oc8051_symbolic_cxrom1.regarray[11] [5], \oc8051_symbolic_cxrom1.regarray[11] [4]);
  nand _27611_ (_05307_, _05306_, _04422_);
  or _27612_ (_05308_, \oc8051_symbolic_cxrom1.regarray[8] [5], \oc8051_symbolic_cxrom1.regarray[8] [4]);
  nand _27613_ (_05309_, _05308_, _04453_);
  and _27614_ (_05310_, _05309_, _05307_);
  and _27615_ (_05311_, _05310_, _05305_);
  and _27616_ (_05312_, _05311_, _05300_);
  and _27617_ (_05313_, _05312_, _05293_);
  and _27618_ (_05314_, _05313_, _05286_);
  or _27619_ (_05315_, _05314_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor _27620_ (_05316_, \oc8051_symbolic_cxrom1.regarray[12] [1], \oc8051_symbolic_cxrom1.regarray[12] [0]);
  nor _27621_ (_05317_, \oc8051_symbolic_cxrom1.regarray[12] [3], \oc8051_symbolic_cxrom1.regarray[12] [2]);
  and _27622_ (_05318_, _05317_, _05316_);
  or _27623_ (_05319_, _05318_, _05280_);
  nor _27624_ (_05320_, \oc8051_symbolic_cxrom1.regarray[15] [3], \oc8051_symbolic_cxrom1.regarray[15] [2]);
  nor _27625_ (_05321_, \oc8051_symbolic_cxrom1.regarray[15] [1], \oc8051_symbolic_cxrom1.regarray[15] [0]);
  and _27626_ (_05322_, _05321_, _05320_);
  or _27627_ (_05323_, _05322_, _05266_);
  and _27628_ (_05324_, _05323_, _05319_);
  nor _27629_ (_05325_, \oc8051_symbolic_cxrom1.regarray[14] [1], \oc8051_symbolic_cxrom1.regarray[14] [0]);
  nor _27630_ (_05326_, \oc8051_symbolic_cxrom1.regarray[14] [3], \oc8051_symbolic_cxrom1.regarray[14] [2]);
  nand _27631_ (_05327_, _05326_, _05325_);
  nand _27632_ (_05328_, _05327_, _04464_);
  nor _27633_ (_05329_, \oc8051_symbolic_cxrom1.regarray[13] [1], \oc8051_symbolic_cxrom1.regarray[13] [0]);
  nor _27634_ (_05330_, \oc8051_symbolic_cxrom1.regarray[13] [3], \oc8051_symbolic_cxrom1.regarray[13] [2]);
  nand _27635_ (_05331_, _05330_, _05329_);
  nand _27636_ (_05332_, _05331_, _04440_);
  and _27637_ (_05333_, _05332_, _05328_);
  and _27638_ (_05334_, _05333_, _05324_);
  and _27639_ (_05335_, _04422_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  and _27640_ (_05336_, _04464_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  or _27641_ (_05337_, _05336_, _05335_);
  and _27642_ (_05338_, _04440_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  and _27643_ (_05339_, _04453_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  or _27644_ (_05340_, _05339_, _05338_);
  or _27645_ (_05341_, _05340_, _05337_);
  nand _27646_ (_05342_, _04464_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  or _27647_ (_05343_, \oc8051_symbolic_cxrom1.regarray[14] [5], \oc8051_symbolic_cxrom1.regarray[14] [4]);
  nand _27648_ (_05344_, _05343_, _04464_);
  and _27649_ (_05345_, _05344_, _05342_);
  nand _27650_ (_05346_, _04422_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  nand _27651_ (_05347_, _04453_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  and _27652_ (_05348_, _05347_, _05346_);
  and _27653_ (_05349_, _05348_, _05345_);
  nand _27654_ (_05350_, _04440_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  or _27655_ (_05351_, \oc8051_symbolic_cxrom1.regarray[12] [5], \oc8051_symbolic_cxrom1.regarray[12] [4]);
  nand _27656_ (_05352_, _05351_, _04453_);
  and _27657_ (_05353_, _05352_, _05350_);
  or _27658_ (_05354_, \oc8051_symbolic_cxrom1.regarray[15] [5], \oc8051_symbolic_cxrom1.regarray[15] [4]);
  nand _27659_ (_05355_, _05354_, _04422_);
  or _27660_ (_05356_, \oc8051_symbolic_cxrom1.regarray[13] [5], \oc8051_symbolic_cxrom1.regarray[13] [4]);
  nand _27661_ (_05357_, _05356_, _04440_);
  and _27662_ (_05358_, _05357_, _05355_);
  and _27663_ (_05359_, _05358_, _05353_);
  and _27664_ (_05360_, _05359_, _05349_);
  and _27665_ (_05361_, _05360_, _05341_);
  and _27666_ (_05362_, _05361_, _05334_);
  or _27667_ (_05363_, _05362_, _01920_);
  and _27668_ (_05364_, _05363_, _05315_);
  or _27669_ (_05365_, _05364_, _02512_);
  or _27670_ (_05366_, \oc8051_symbolic_cxrom1.regarray[6] [3], \oc8051_symbolic_cxrom1.regarray[6] [2]);
  nand _27671_ (_05367_, _05366_, _04464_);
  and _27672_ (_05368_, _05367_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  or _27673_ (_05369_, \oc8051_symbolic_cxrom1.regarray[7] [3], \oc8051_symbolic_cxrom1.regarray[7] [2]);
  nand _27674_ (_05370_, _05369_, _04422_);
  or _27675_ (_05371_, \oc8051_symbolic_cxrom1.regarray[5] [3], \oc8051_symbolic_cxrom1.regarray[5] [2]);
  nand _27676_ (_05372_, _05371_, _04440_);
  and _27677_ (_05373_, _05372_, _05370_);
  or _27678_ (_05374_, \oc8051_symbolic_cxrom1.regarray[4] [3], \oc8051_symbolic_cxrom1.regarray[4] [2]);
  nand _27679_ (_05375_, _05374_, _04453_);
  or _27680_ (_05376_, \oc8051_symbolic_cxrom1.regarray[4] [5], \oc8051_symbolic_cxrom1.regarray[4] [4]);
  nand _27681_ (_05377_, _05376_, _04453_);
  and _27682_ (_05378_, _05377_, _05375_);
  and _27683_ (_05379_, _05378_, _05373_);
  and _27684_ (_05380_, _05379_, _05368_);
  nand _27685_ (_05381_, _04440_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  or _27686_ (_05382_, \oc8051_symbolic_cxrom1.regarray[5] [5], \oc8051_symbolic_cxrom1.regarray[5] [4]);
  nand _27687_ (_05383_, _05382_, _04440_);
  and _27688_ (_05384_, _05383_, _05381_);
  or _27689_ (_05385_, \oc8051_symbolic_cxrom1.regarray[7] [5], \oc8051_symbolic_cxrom1.regarray[7] [4]);
  nand _27690_ (_05386_, _05385_, _04422_);
  or _27691_ (_05387_, \oc8051_symbolic_cxrom1.regarray[6] [5], \oc8051_symbolic_cxrom1.regarray[6] [4]);
  nand _27692_ (_05388_, _05387_, _04464_);
  and _27693_ (_05389_, _05388_, _05386_);
  and _27694_ (_05390_, _05389_, _05384_);
  nand _27695_ (_05391_, _04464_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  or _27696_ (_05392_, \oc8051_symbolic_cxrom1.regarray[4] [1], \oc8051_symbolic_cxrom1.regarray[4] [0]);
  nand _27697_ (_05393_, _05392_, _04453_);
  and _27698_ (_05394_, _05393_, _05391_);
  nand _27699_ (_05395_, _04422_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  nand _27700_ (_05396_, _04453_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  and _27701_ (_05397_, _05396_, _05395_);
  and _27702_ (_05398_, _05397_, _05394_);
  and _27703_ (_05399_, _05398_, _05390_);
  and _27704_ (_05400_, _04440_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  and _27705_ (_05401_, _04453_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  or _27706_ (_05402_, _05401_, _05400_);
  and _27707_ (_05403_, _04422_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  and _27708_ (_05404_, _04464_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  or _27709_ (_05405_, _05404_, _05403_);
  or _27710_ (_05406_, _05405_, _05402_);
  or _27711_ (_05407_, \oc8051_symbolic_cxrom1.regarray[6] [1], \oc8051_symbolic_cxrom1.regarray[6] [0]);
  nand _27712_ (_05408_, _05407_, _04464_);
  or _27713_ (_05409_, \oc8051_symbolic_cxrom1.regarray[7] [1], \oc8051_symbolic_cxrom1.regarray[7] [0]);
  nand _27714_ (_05410_, _05409_, _04422_);
  or _27715_ (_05411_, \oc8051_symbolic_cxrom1.regarray[5] [1], \oc8051_symbolic_cxrom1.regarray[5] [0]);
  nand _27716_ (_05412_, _05411_, _04440_);
  and _27717_ (_05413_, _05412_, _05410_);
  and _27718_ (_05414_, _05413_, _05408_);
  and _27719_ (_05415_, _05414_, _05406_);
  and _27720_ (_05416_, _05415_, _05399_);
  and _27721_ (_05417_, _05416_, _05380_);
  nand _27722_ (_05418_, _04440_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  and _27723_ (_05419_, _05418_, _01920_);
  or _27724_ (_05420_, \oc8051_symbolic_cxrom1.regarray[0] [5], \oc8051_symbolic_cxrom1.regarray[0] [4]);
  nand _27725_ (_05421_, _05420_, _04453_);
  or _27726_ (_05422_, \oc8051_symbolic_cxrom1.regarray[0] [1], \oc8051_symbolic_cxrom1.regarray[0] [0]);
  nand _27727_ (_05423_, _05422_, _04453_);
  and _27728_ (_05424_, _05423_, _05421_);
  or _27729_ (_05425_, \oc8051_symbolic_cxrom1.regarray[2] [3], \oc8051_symbolic_cxrom1.regarray[2] [2]);
  nand _27730_ (_05426_, _05425_, _04464_);
  or _27731_ (_05427_, \oc8051_symbolic_cxrom1.regarray[1] [3], \oc8051_symbolic_cxrom1.regarray[1] [2]);
  nand _27732_ (_05428_, _05427_, _04440_);
  and _27733_ (_05429_, _05428_, _05426_);
  and _27734_ (_05430_, _05429_, _05424_);
  and _27735_ (_05431_, _05430_, _05419_);
  nand _27736_ (_05432_, _04453_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  or _27737_ (_05433_, \oc8051_symbolic_cxrom1.regarray[1] [5], \oc8051_symbolic_cxrom1.regarray[1] [4]);
  nand _27738_ (_05434_, _05433_, _04440_);
  and _27739_ (_05435_, _05434_, _05432_);
  or _27740_ (_05436_, \oc8051_symbolic_cxrom1.regarray[3] [5], \oc8051_symbolic_cxrom1.regarray[3] [4]);
  nand _27741_ (_05437_, _05436_, _04422_);
  or _27742_ (_05438_, \oc8051_symbolic_cxrom1.regarray[2] [5], \oc8051_symbolic_cxrom1.regarray[2] [4]);
  nand _27743_ (_05439_, _05438_, _04464_);
  and _27744_ (_05440_, _05439_, _05437_);
  and _27745_ (_05441_, _05440_, _05435_);
  nand _27746_ (_05442_, _04464_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  nand _27747_ (_05443_, _04422_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  and _27748_ (_05444_, _05443_, _05442_);
  or _27749_ (_05445_, \oc8051_symbolic_cxrom1.regarray[3] [3], \oc8051_symbolic_cxrom1.regarray[3] [2]);
  nand _27750_ (_05446_, _05445_, _04422_);
  or _27751_ (_05447_, \oc8051_symbolic_cxrom1.regarray[0] [3], \oc8051_symbolic_cxrom1.regarray[0] [2]);
  nand _27752_ (_05448_, _05447_, _04453_);
  and _27753_ (_05449_, _05448_, _05446_);
  and _27754_ (_05450_, _05449_, _05444_);
  and _27755_ (_05451_, _05450_, _05441_);
  and _27756_ (_05452_, _04453_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  and _27757_ (_05453_, _04440_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  or _27758_ (_05454_, _05453_, _05452_);
  and _27759_ (_05455_, _04464_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  and _27760_ (_05456_, _04422_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  or _27761_ (_05457_, _05456_, _05455_);
  or _27762_ (_05458_, _05457_, _05454_);
  or _27763_ (_05459_, \oc8051_symbolic_cxrom1.regarray[2] [1], \oc8051_symbolic_cxrom1.regarray[2] [0]);
  nand _27764_ (_05460_, _05459_, _04464_);
  or _27765_ (_05461_, \oc8051_symbolic_cxrom1.regarray[3] [1], \oc8051_symbolic_cxrom1.regarray[3] [0]);
  nand _27766_ (_05462_, _05461_, _04422_);
  or _27767_ (_05463_, \oc8051_symbolic_cxrom1.regarray[1] [1], \oc8051_symbolic_cxrom1.regarray[1] [0]);
  nand _27768_ (_05464_, _05463_, _04440_);
  and _27769_ (_05465_, _05464_, _05462_);
  and _27770_ (_05466_, _05465_, _05460_);
  and _27771_ (_05467_, _05466_, _05458_);
  and _27772_ (_05468_, _05467_, _05451_);
  and _27773_ (_05469_, _05468_, _05431_);
  or _27774_ (_05470_, _05469_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or _27775_ (_05471_, _05470_, _05417_);
  and _27776_ (_05472_, _05246_, _04466_);
  or _27777_ (_05473_, _05472_, _01920_);
  or _27778_ (_05474_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [3]);
  or _27779_ (_05475_, _02512_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and _27780_ (_05476_, _05475_, _05474_);
  or _27781_ (_05477_, _05476_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and _27782_ (_05478_, _05477_, _05473_);
  and _27783_ (_05479_, _05478_, _04440_);
  and _27784_ (_05480_, _04464_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  or _27785_ (_05481_, _02512_, \oc8051_symbolic_cxrom1.regvalid [0]);
  or _27786_ (_05482_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [8]);
  and _27787_ (_05483_, _05482_, _05481_);
  and _27788_ (_05484_, _05483_, _05480_);
  or _27789_ (_05485_, _02512_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or _27790_ (_05486_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [9]);
  and _27791_ (_05487_, _05486_, _05485_);
  and _27792_ (_05488_, _05487_, _04423_);
  or _27793_ (_05489_, _05488_, _05484_);
  or _27794_ (_05490_, _05489_, _05479_);
  or _27795_ (_05491_, _02512_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and _27796_ (_05492_, _05491_, _04431_);
  or _27797_ (_05493_, _05492_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _27798_ (_05494_, _05235_, _04455_);
  or _27799_ (_05495_, _05494_, _02505_);
  and _27800_ (_05496_, _05495_, _04739_);
  and _27801_ (_05497_, _05496_, _05493_);
  or _27802_ (_05498_, _02512_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and _27803_ (_05499_, _04442_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and _27804_ (_05500_, _05499_, _05498_);
  or _27805_ (_05501_, _02512_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or _27806_ (_05502_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [2]);
  and _27807_ (_05503_, _05502_, _01920_);
  and _27808_ (_05504_, _05503_, _05501_);
  or _27809_ (_05505_, _05504_, _05500_);
  and _27810_ (_05506_, _05505_, _04453_);
  or _27811_ (_05507_, _05506_, _05497_);
  or _27812_ (_05508_, _05507_, _05490_);
  and _27813_ (_05509_, _05505_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and _27814_ (_05510_, _05492_, _04738_);
  or _27815_ (_05511_, _02512_, \oc8051_symbolic_cxrom1.regvalid [8]);
  or _27816_ (_05512_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [0]);
  and _27817_ (_05513_, _05512_, _05222_);
  and _27818_ (_05514_, _05513_, _05511_);
  or _27819_ (_05515_, _05514_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  or _27820_ (_05516_, _05515_, _05510_);
  or _27821_ (_05517_, _05516_, _05509_);
  and _27822_ (_05518_, _05478_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and _27823_ (_05519_, _05494_, _04738_);
  and _27824_ (_05520_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [9]);
  and _27825_ (_05521_, _02512_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or _27826_ (_05522_, _05521_, _05520_);
  and _27827_ (_05523_, _05522_, _05222_);
  or _27828_ (_05524_, _05523_, _02505_);
  or _27829_ (_05525_, _05524_, _05519_);
  or _27830_ (_05526_, _05525_, _05518_);
  nor _27831_ (_05527_, _01956_, first_instr);
  and _27832_ (_05528_, _05527_, _05526_);
  and _27833_ (_05529_, _05528_, _05517_);
  and _27834_ (_05530_, _05529_, _05508_);
  and _27835_ (_05531_, _05530_, _05471_);
  and _27836_ (_05532_, _05531_, _05365_);
  and _27837_ (_05533_, _05532_, _04476_);
  and _27838_ (_05534_, _05533_, _05265_);
  and _27839_ (_05535_, _05534_, _05216_);
  and _27840_ (property_invalid_jc, _05535_, _05062_);
  or _27841_ (_05536_, pc_log_change_r, _04421_);
  nand _27842_ (_05537_, pc_log_change_r, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nand _27843_ (_00000_, _05537_, _05536_);
  and _27844_ (_05538_, _01956_, first_instr);
  or _27845_ (_00001_, _05538_, rst);
  dff _27846_ (cy_reg, _00000_, clk);
  dff _27847_ (pc_log_change_r, pc_log_change, clk);
  dff _27848_ (first_instr, _00001_, clk);
  dff _27849_ (\oc8051_symbolic_cxrom1.regarray[15] [0], _13870_, clk);
  dff _27850_ (\oc8051_symbolic_cxrom1.regarray[15] [1], _13871_, clk);
  dff _27851_ (\oc8051_symbolic_cxrom1.regarray[15] [2], _13872_, clk);
  dff _27852_ (\oc8051_symbolic_cxrom1.regarray[15] [3], _13873_, clk);
  dff _27853_ (\oc8051_symbolic_cxrom1.regarray[15] [4], _13874_, clk);
  dff _27854_ (\oc8051_symbolic_cxrom1.regarray[15] [5], _13875_, clk);
  dff _27855_ (\oc8051_symbolic_cxrom1.regarray[15] [6], _13876_, clk);
  dff _27856_ (\oc8051_symbolic_cxrom1.regarray[15] [7], _13877_, clk);
  dff _27857_ (\oc8051_symbolic_cxrom1.regarray[14] [0], _09923_, clk);
  dff _27858_ (\oc8051_symbolic_cxrom1.regarray[14] [1], _09925_, clk);
  dff _27859_ (\oc8051_symbolic_cxrom1.regarray[14] [2], _09926_, clk);
  dff _27860_ (\oc8051_symbolic_cxrom1.regarray[14] [3], _09929_, clk);
  dff _27861_ (\oc8051_symbolic_cxrom1.regarray[14] [4], _09932_, clk);
  dff _27862_ (\oc8051_symbolic_cxrom1.regarray[14] [5], _09935_, clk);
  dff _27863_ (\oc8051_symbolic_cxrom1.regarray[14] [6], _09939_, clk);
  dff _27864_ (\oc8051_symbolic_cxrom1.regarray[14] [7], _09941_, clk);
  dff _27865_ (\oc8051_symbolic_cxrom1.regarray[13] [0], _13869_, clk);
  dff _27866_ (\oc8051_symbolic_cxrom1.regarray[13] [1], _09832_, clk);
  dff _27867_ (\oc8051_symbolic_cxrom1.regarray[13] [2], _09836_, clk);
  dff _27868_ (\oc8051_symbolic_cxrom1.regarray[13] [3], _09840_, clk);
  dff _27869_ (\oc8051_symbolic_cxrom1.regarray[13] [4], _09842_, clk);
  dff _27870_ (\oc8051_symbolic_cxrom1.regarray[13] [5], _09845_, clk);
  dff _27871_ (\oc8051_symbolic_cxrom1.regarray[13] [6], _09847_, clk);
  dff _27872_ (\oc8051_symbolic_cxrom1.regarray[13] [7], _09850_, clk);
  dff _27873_ (\oc8051_symbolic_cxrom1.regarray[12] [0], _09751_, clk);
  dff _27874_ (\oc8051_symbolic_cxrom1.regarray[12] [1], _09755_, clk);
  dff _27875_ (\oc8051_symbolic_cxrom1.regarray[12] [2], _09758_, clk);
  dff _27876_ (\oc8051_symbolic_cxrom1.regarray[12] [3], _09760_, clk);
  dff _27877_ (\oc8051_symbolic_cxrom1.regarray[12] [4], _09762_, clk);
  dff _27878_ (\oc8051_symbolic_cxrom1.regarray[12] [5], _09765_, clk);
  dff _27879_ (\oc8051_symbolic_cxrom1.regarray[12] [6], _09769_, clk);
  dff _27880_ (\oc8051_symbolic_cxrom1.regarray[12] [7], _09772_, clk);
  dff _27881_ (\oc8051_symbolic_cxrom1.regarray[11] [0], _13861_, clk);
  dff _27882_ (\oc8051_symbolic_cxrom1.regarray[11] [1], _13862_, clk);
  dff _27883_ (\oc8051_symbolic_cxrom1.regarray[11] [2], _13863_, clk);
  dff _27884_ (\oc8051_symbolic_cxrom1.regarray[11] [3], _13864_, clk);
  dff _27885_ (\oc8051_symbolic_cxrom1.regarray[11] [4], _13865_, clk);
  dff _27886_ (\oc8051_symbolic_cxrom1.regarray[11] [5], _13866_, clk);
  dff _27887_ (\oc8051_symbolic_cxrom1.regarray[11] [6], _13867_, clk);
  dff _27888_ (\oc8051_symbolic_cxrom1.regarray[11] [7], _13868_, clk);
  dff _27889_ (\oc8051_symbolic_cxrom1.regarray[10] [0], _13853_, clk);
  dff _27890_ (\oc8051_symbolic_cxrom1.regarray[10] [1], _13854_, clk);
  dff _27891_ (\oc8051_symbolic_cxrom1.regarray[10] [2], _13855_, clk);
  dff _27892_ (\oc8051_symbolic_cxrom1.regarray[10] [3], _13856_, clk);
  dff _27893_ (\oc8051_symbolic_cxrom1.regarray[10] [4], _13857_, clk);
  dff _27894_ (\oc8051_symbolic_cxrom1.regarray[10] [5], _13858_, clk);
  dff _27895_ (\oc8051_symbolic_cxrom1.regarray[10] [6], _13859_, clk);
  dff _27896_ (\oc8051_symbolic_cxrom1.regarray[10] [7], _13860_, clk);
  dff _27897_ (\oc8051_symbolic_cxrom1.regarray[9] [0], _13898_, clk);
  dff _27898_ (\oc8051_symbolic_cxrom1.regarray[9] [1], _13899_, clk);
  dff _27899_ (\oc8051_symbolic_cxrom1.regarray[9] [2], _13900_, clk);
  dff _27900_ (\oc8051_symbolic_cxrom1.regarray[9] [3], _13901_, clk);
  dff _27901_ (\oc8051_symbolic_cxrom1.regarray[9] [4], _13902_, clk);
  dff _27902_ (\oc8051_symbolic_cxrom1.regarray[9] [5], _13903_, clk);
  dff _27903_ (\oc8051_symbolic_cxrom1.regarray[9] [6], _13904_, clk);
  dff _27904_ (\oc8051_symbolic_cxrom1.regarray[9] [7], _13905_, clk);
  dff _27905_ (\oc8051_symbolic_cxrom1.regarray[8] [0], _09403_, clk);
  dff _27906_ (\oc8051_symbolic_cxrom1.regarray[8] [1], _09408_, clk);
  dff _27907_ (\oc8051_symbolic_cxrom1.regarray[8] [2], _13892_, clk);
  dff _27908_ (\oc8051_symbolic_cxrom1.regarray[8] [3], _13893_, clk);
  dff _27909_ (\oc8051_symbolic_cxrom1.regarray[8] [4], _13894_, clk);
  dff _27910_ (\oc8051_symbolic_cxrom1.regarray[8] [5], _13895_, clk);
  dff _27911_ (\oc8051_symbolic_cxrom1.regarray[8] [6], _13896_, clk);
  dff _27912_ (\oc8051_symbolic_cxrom1.regarray[8] [7], _13897_, clk);
  dff _27913_ (\oc8051_symbolic_cxrom1.regarray[7] [0], _13884_, clk);
  dff _27914_ (\oc8051_symbolic_cxrom1.regarray[7] [1], _13885_, clk);
  dff _27915_ (\oc8051_symbolic_cxrom1.regarray[7] [2], _13886_, clk);
  dff _27916_ (\oc8051_symbolic_cxrom1.regarray[7] [3], _13887_, clk);
  dff _27917_ (\oc8051_symbolic_cxrom1.regarray[7] [4], _13888_, clk);
  dff _27918_ (\oc8051_symbolic_cxrom1.regarray[7] [5], _13889_, clk);
  dff _27919_ (\oc8051_symbolic_cxrom1.regarray[7] [6], _13890_, clk);
  dff _27920_ (\oc8051_symbolic_cxrom1.regarray[7] [7], _13891_, clk);
  dff _27921_ (\oc8051_symbolic_cxrom1.regarray[6] [0], _09217_, clk);
  dff _27922_ (\oc8051_symbolic_cxrom1.regarray[6] [1], _09220_, clk);
  dff _27923_ (\oc8051_symbolic_cxrom1.regarray[6] [2], _09224_, clk);
  dff _27924_ (\oc8051_symbolic_cxrom1.regarray[6] [3], _09229_, clk);
  dff _27925_ (\oc8051_symbolic_cxrom1.regarray[6] [4], _09233_, clk);
  dff _27926_ (\oc8051_symbolic_cxrom1.regarray[6] [5], _09235_, clk);
  dff _27927_ (\oc8051_symbolic_cxrom1.regarray[6] [6], _09238_, clk);
  dff _27928_ (\oc8051_symbolic_cxrom1.regarray[6] [7], _09242_, clk);
  dff _27929_ (\oc8051_symbolic_cxrom1.regarray[5] [0], _09110_, clk);
  dff _27930_ (\oc8051_symbolic_cxrom1.regarray[5] [1], _09115_, clk);
  dff _27931_ (\oc8051_symbolic_cxrom1.regarray[5] [2], _09120_, clk);
  dff _27932_ (\oc8051_symbolic_cxrom1.regarray[5] [3], _09125_, clk);
  dff _27933_ (\oc8051_symbolic_cxrom1.regarray[5] [4], _09129_, clk);
  dff _27934_ (\oc8051_symbolic_cxrom1.regarray[5] [5], _09134_, clk);
  dff _27935_ (\oc8051_symbolic_cxrom1.regarray[5] [6], _09138_, clk);
  dff _27936_ (\oc8051_symbolic_cxrom1.regarray[5] [7], _09141_, clk);
  dff _27937_ (\oc8051_symbolic_cxrom1.regarray[1] [0], _08705_, clk);
  dff _27938_ (\oc8051_symbolic_cxrom1.regarray[1] [1], _08709_, clk);
  dff _27939_ (\oc8051_symbolic_cxrom1.regarray[1] [2], _08712_, clk);
  dff _27940_ (\oc8051_symbolic_cxrom1.regarray[1] [3], _08715_, clk);
  dff _27941_ (\oc8051_symbolic_cxrom1.regarray[1] [4], _08717_, clk);
  dff _27942_ (\oc8051_symbolic_cxrom1.regarray[1] [5], _08719_, clk);
  dff _27943_ (\oc8051_symbolic_cxrom1.regarray[1] [6], _08721_, clk);
  dff _27944_ (\oc8051_symbolic_cxrom1.regarray[1] [7], _08724_, clk);
  dff _27945_ (\oc8051_symbolic_cxrom1.regarray[0] [0], _08586_, clk);
  dff _27946_ (\oc8051_symbolic_cxrom1.regarray[0] [1], _08591_, clk);
  dff _27947_ (\oc8051_symbolic_cxrom1.regarray[0] [2], _08597_, clk);
  dff _27948_ (\oc8051_symbolic_cxrom1.regarray[0] [3], _08600_, clk);
  dff _27949_ (\oc8051_symbolic_cxrom1.regarray[0] [4], _08606_, clk);
  dff _27950_ (\oc8051_symbolic_cxrom1.regarray[0] [5], _08612_, clk);
  dff _27951_ (\oc8051_symbolic_cxrom1.regarray[0] [6], _08617_, clk);
  dff _27952_ (\oc8051_symbolic_cxrom1.regarray[0] [7], _08619_, clk);
  dff _27953_ (\oc8051_symbolic_cxrom1.regarray[3] [0], _13879_, clk);
  dff _27954_ (\oc8051_symbolic_cxrom1.regarray[3] [1], _08899_, clk);
  dff _27955_ (\oc8051_symbolic_cxrom1.regarray[3] [2], _08902_, clk);
  dff _27956_ (\oc8051_symbolic_cxrom1.regarray[3] [3], _08907_, clk);
  dff _27957_ (\oc8051_symbolic_cxrom1.regarray[3] [4], _08912_, clk);
  dff _27958_ (\oc8051_symbolic_cxrom1.regarray[3] [5], _08916_, clk);
  dff _27959_ (\oc8051_symbolic_cxrom1.regarray[3] [6], _08919_, clk);
  dff _27960_ (\oc8051_symbolic_cxrom1.regarray[3] [7], _08922_, clk);
  dff _27961_ (\oc8051_symbolic_cxrom1.regarray[2] [0], _08801_, clk);
  dff _27962_ (\oc8051_symbolic_cxrom1.regarray[2] [1], _08805_, clk);
  dff _27963_ (\oc8051_symbolic_cxrom1.regarray[2] [2], _08810_, clk);
  dff _27964_ (\oc8051_symbolic_cxrom1.regarray[2] [3], _08814_, clk);
  dff _27965_ (\oc8051_symbolic_cxrom1.regarray[2] [4], _08817_, clk);
  dff _27966_ (\oc8051_symbolic_cxrom1.regarray[2] [5], _13878_, clk);
  dff _27967_ (\oc8051_symbolic_cxrom1.regarray[2] [6], _08822_, clk);
  dff _27968_ (\oc8051_symbolic_cxrom1.regarray[2] [7], _08825_, clk);
  dff _27969_ (\oc8051_symbolic_cxrom1.regarray[4] [0], _09011_, clk);
  dff _27970_ (\oc8051_symbolic_cxrom1.regarray[4] [1], _09016_, clk);
  dff _27971_ (\oc8051_symbolic_cxrom1.regarray[4] [2], _13880_, clk);
  dff _27972_ (\oc8051_symbolic_cxrom1.regarray[4] [3], _13881_, clk);
  dff _27973_ (\oc8051_symbolic_cxrom1.regarray[4] [4], _13882_, clk);
  dff _27974_ (\oc8051_symbolic_cxrom1.regarray[4] [5], _13883_, clk);
  dff _27975_ (\oc8051_symbolic_cxrom1.regarray[4] [6], _09034_, clk);
  dff _27976_ (\oc8051_symbolic_cxrom1.regarray[4] [7], _09037_, clk);
  dff _27977_ (\oc8051_symbolic_cxrom1.regvalid [0], _07256_, clk);
  dff _27978_ (\oc8051_symbolic_cxrom1.regvalid [1], _07287_, clk);
  dff _27979_ (\oc8051_symbolic_cxrom1.regvalid [2], _07324_, clk);
  dff _27980_ (\oc8051_symbolic_cxrom1.regvalid [3], _07361_, clk);
  dff _27981_ (\oc8051_symbolic_cxrom1.regvalid [4], _07415_, clk);
  dff _27982_ (\oc8051_symbolic_cxrom1.regvalid [5], _07480_, clk);
  dff _27983_ (\oc8051_symbolic_cxrom1.regvalid [6], _07541_, clk);
  dff _27984_ (\oc8051_symbolic_cxrom1.regvalid [7], _07615_, clk);
  dff _27985_ (\oc8051_symbolic_cxrom1.regvalid [8], _07673_, clk);
  dff _27986_ (\oc8051_symbolic_cxrom1.regvalid [9], _07739_, clk);
  dff _27987_ (\oc8051_symbolic_cxrom1.regvalid [10], _07829_, clk);
  dff _27988_ (\oc8051_symbolic_cxrom1.regvalid [11], _07927_, clk);
  dff _27989_ (\oc8051_symbolic_cxrom1.regvalid [12], _08032_, clk);
  dff _27990_ (\oc8051_symbolic_cxrom1.regvalid [13], _08119_, clk);
  dff _27991_ (\oc8051_symbolic_cxrom1.regvalid [14], _08231_, clk);
  dff _27992_ (\oc8051_symbolic_cxrom1.regvalid [15], _07207_, clk);
  dff _27993_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _04128_, clk);
  dff _27994_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _04074_, clk);
  dff _27995_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _04054_, clk);
  dff _27996_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _04050_, clk);
  dff _27997_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4], _12807_, clk);
  dff _27998_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5], _03846_, clk);
  dff _27999_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], _03614_, clk);
  dff _28000_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1], _10695_, clk);
  dff _28001_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0], _13506_, clk);
  dff _28002_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1], _13470_, clk);
  dff _28003_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2], _00331_, clk);
  dff _28004_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3], _00235_, clk);
  dff _28005_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4], _00205_, clk);
  dff _28006_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5], _00153_, clk);
  dff _28007_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6], _00085_, clk);
  dff _28008_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7], _03883_, clk);
  dff _28009_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], _11685_, clk);
  dff _28010_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _10840_, clk);
  dff _28011_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0], _06005_, clk);
  dff _28012_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1], _06036_, clk);
  dff _28013_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2], _06017_, clk);
  dff _28014_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3], _06013_, clk);
  dff _28015_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4], _06007_, clk);
  dff _28016_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5], _11741_, clk);
  dff _28017_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6], _12386_, clk);
  dff _28018_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7], _06548_, clk);
  dff _28019_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8], _00475_, clk);
  dff _28020_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9], _00910_, clk);
  dff _28021_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10], _01737_, clk);
  dff _28022_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11], _03645_, clk);
  dff _28023_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12], _04571_, clk);
  dff _28024_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13], _03742_, clk);
  dff _28025_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [0], _06907_, clk);
  dff _28026_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [1], _06909_, clk);
  dff _28027_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [2], _06912_, clk);
  dff _28028_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [3], _06914_, clk);
  dff _28029_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [4], _06917_, clk);
  dff _28030_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [5], _06920_, clk);
  dff _28031_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [6], _06923_, clk);
  dff _28032_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [7], _06780_, clk);
  dff _28033_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [5], _12033_, clk);
  dff _28034_ (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], _01125_, clk);
  dff _28035_ (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], _12598_, clk);
  dff _28036_ (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], _04080_, clk);
  dff _28037_ (\oc8051_top_1.oc8051_decoder1.mem_act [0], _01436_, clk);
  dff _28038_ (\oc8051_top_1.oc8051_decoder1.mem_act [1], _07502_, clk);
  dff _28039_ (\oc8051_top_1.oc8051_decoder1.mem_act [2], _04142_, clk);
  dff _28040_ (\oc8051_top_1.oc8051_decoder1.state [0], _02378_, clk);
  dff _28041_ (\oc8051_top_1.oc8051_decoder1.state [1], _04144_, clk);
  dff _28042_ (\oc8051_top_1.oc8051_decoder1.op [0], _07409_, clk);
  dff _28043_ (\oc8051_top_1.oc8051_decoder1.op [1], _07268_, clk);
  dff _28044_ (\oc8051_top_1.oc8051_decoder1.op [2], _03600_, clk);
  dff _28045_ (\oc8051_top_1.oc8051_decoder1.op [3], _03347_, clk);
  dff _28046_ (\oc8051_top_1.oc8051_decoder1.op [4], _07341_, clk);
  dff _28047_ (\oc8051_top_1.oc8051_decoder1.op [5], _02850_, clk);
  dff _28048_ (\oc8051_top_1.oc8051_decoder1.op [6], _02838_, clk);
  dff _28049_ (\oc8051_top_1.oc8051_decoder1.op [7], _04168_, clk);
  dff _28050_ (\oc8051_top_1.oc8051_decoder1.src_sel3 , _04091_, clk);
  dff _28051_ (\oc8051_top_1.oc8051_decoder1.wr_sfr [0], _03548_, clk);
  dff _28052_ (\oc8051_top_1.oc8051_decoder1.wr_sfr [1], _04062_, clk);
  dff _28053_ (\oc8051_top_1.oc8051_decoder1.src_sel2 [0], _03824_, clk);
  dff _28054_ (\oc8051_top_1.oc8051_decoder1.src_sel2 [1], _04176_, clk);
  dff _28055_ (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _04490_, clk);
  dff _28056_ (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _10247_, clk);
  dff _28057_ (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], _04179_, clk);
  dff _28058_ (\oc8051_top_1.oc8051_decoder1.src_sel1 [0], _10693_, clk);
  dff _28059_ (\oc8051_top_1.oc8051_decoder1.src_sel1 [1], _10282_, clk);
  dff _28060_ (\oc8051_top_1.oc8051_decoder1.src_sel1 [2], _04181_, clk);
  dff _28061_ (\oc8051_top_1.oc8051_decoder1.cy_sel [0], _03671_, clk);
  dff _28062_ (\oc8051_top_1.oc8051_decoder1.cy_sel [1], _04184_, clk);
  dff _28063_ (\oc8051_top_1.oc8051_decoder1.alu_op [0], _11293_, clk);
  dff _28064_ (\oc8051_top_1.oc8051_decoder1.alu_op [1], _11295_, clk);
  dff _28065_ (\oc8051_top_1.oc8051_decoder1.alu_op [2], _03558_, clk);
  dff _28066_ (\oc8051_top_1.oc8051_decoder1.alu_op [3], _04186_, clk);
  dff _28067_ (\oc8051_top_1.oc8051_decoder1.psw_set [0], _11720_, clk);
  dff _28068_ (\oc8051_top_1.oc8051_decoder1.psw_set [1], _04188_, clk);
  dff _28069_ (\oc8051_top_1.oc8051_decoder1.wr , _04221_, clk);
  dff _28070_ (\oc8051_top_1.oc8051_indi_addr1.wr_bit_r , _00251_, clk);
  dff _28071_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [0], _00328_, clk);
  dff _28072_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [1], _02609_, clk);
  dff _28073_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [2], _02612_, clk);
  dff _28074_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [3], _01932_, clk);
  dff _28075_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [4], _02330_, clk);
  dff _28076_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [5], _02545_, clk);
  dff _28077_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [6], _02503_, clk);
  dff _28078_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [7], _03324_, clk);
  dff _28079_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [0], _04166_, clk);
  dff _28080_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [1], _02536_, clk);
  dff _28081_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [2], _03720_, clk);
  dff _28082_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [3], _05581_, clk);
  dff _28083_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [4], _01631_, clk);
  dff _28084_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [5], _11191_, clk);
  dff _28085_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [6], _02190_, clk);
  dff _28086_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [7], _03332_, clk);
  dff _28087_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [0], _02413_, clk);
  dff _28088_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [1], _06961_, clk);
  dff _28089_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [2], _03673_, clk);
  dff _28090_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [3], _11681_, clk);
  dff _28091_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [4], _10816_, clk);
  dff _28092_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [5], _05578_, clk);
  dff _28093_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [6], _12281_, clk);
  dff _28094_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [7], _03446_, clk);
  dff _28095_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [0], _03914_, clk);
  dff _28096_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [1], _13761_, clk);
  dff _28097_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [2], _00219_, clk);
  dff _28098_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [3], _02471_, clk);
  dff _28099_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [4], _00060_, clk);
  dff _28100_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [5], _10361_, clk);
  dff _28101_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [6], _02165_, clk);
  dff _28102_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [7], _00076_, clk);
  dff _28103_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [0], _11882_, clk);
  dff _28104_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [1], _06623_, clk);
  dff _28105_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [2], _02353_, clk);
  dff _28106_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [3], _03769_, clk);
  dff _28107_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [4], _13682_, clk);
  dff _28108_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [5], _04052_, clk);
  dff _28109_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [6], _03636_, clk);
  dff _28110_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [7], _03850_, clk);
  dff _28111_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [0], _06610_, clk);
  dff _28112_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [1], _11755_, clk);
  dff _28113_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [2], _12772_, clk);
  dff _28114_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [3], _11298_, clk);
  dff _28115_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [4], _11748_, clk);
  dff _28116_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [5], _11302_, clk);
  dff _28117_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [6], _13157_, clk);
  dff _28118_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [7], _03888_, clk);
  dff _28119_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [0], _00025_, clk);
  dff _28120_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [1], _11229_, clk);
  dff _28121_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [2], _02818_, clk);
  dff _28122_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [3], _11880_, clk);
  dff _28123_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [4], _02286_, clk);
  dff _28124_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [5], _11869_, clk);
  dff _28125_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [6], _01895_, clk);
  dff _28126_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [7], _00247_, clk);
  dff _28127_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [0], _08551_, clk);
  dff _28128_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [1], _08614_, clk);
  dff _28129_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [2], _03270_, clk);
  dff _28130_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [3], _02012_, clk);
  dff _28131_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [4], _02010_, clk);
  dff _28132_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [5], _08845_, clk);
  dff _28133_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [6], _03566_, clk);
  dff _28134_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [7], _00122_, clk);
  dff _28135_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [0], _02597_, clk);
  dff _28136_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [1], _11963_, clk);
  dff _28137_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [2], _11184_, clk);
  dff _28138_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [3], _13222_, clk);
  dff _28139_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [4], _11375_, clk);
  dff _28140_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [0], _01437_, clk);
  dff _28141_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [1], _00999_, clk);
  dff _28142_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [2], _01447_, clk);
  dff _28143_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [3], _01444_, clk);
  dff _28144_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [4], _00996_, clk);
  dff _28145_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [5], _01077_, clk);
  dff _28146_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [6], _01453_, clk);
  dff _28147_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [7], _01449_, clk);
  dff _28148_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [8], _00992_, clk);
  dff _28149_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [9], _01493_, clk);
  dff _28150_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [10], _01459_, clk);
  dff _28151_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [11], _00962_, clk);
  dff _28152_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [12], _01073_, clk);
  dff _28153_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [13], _01135_, clk);
  dff _28154_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [14], _01150_, clk);
  dff _28155_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [15], _02604_, clk);
  dff _28156_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _01569_, clk);
  dff _28157_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _01566_, clk);
  dff _28158_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _00941_, clk);
  dff _28159_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _01584_, clk);
  dff _28160_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _01571_, clk);
  dff _28161_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _00938_, clk);
  dff _28162_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _01065_, clk);
  dff _28163_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _01593_, clk);
  dff _28164_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _01587_, clk);
  dff _28165_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _00933_, clk);
  dff _28166_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _01596_, clk);
  dff _28167_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _01594_, clk);
  dff _28168_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _00925_, clk);
  dff _28169_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _01062_, clk);
  dff _28170_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _01130_, clk);
  dff _28171_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _04429_, clk);
  dff _28172_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [0], _03454_, clk);
  dff _28173_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [1], _04082_, clk);
  dff _28174_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [2], _04044_, clk);
  dff _28175_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [3], _03936_, clk);
  dff _28176_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [4], _03902_, clk);
  dff _28177_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [5], _03873_, clk);
  dff _28178_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [6], _11974_, clk);
  dff _28179_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [7], _11165_, clk);
  dff _28180_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [8], _11355_, clk);
  dff _28181_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [9], _11551_, clk);
  dff _28182_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [10], _00549_, clk);
  dff _28183_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [11], _04015_, clk);
  dff _28184_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [12], _04352_, clk);
  dff _28185_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [13], _04284_, clk);
  dff _28186_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [14], _04275_, clk);
  dff _28187_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [15], _04017_, clk);
  dff _28188_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [16], _11984_, clk);
  dff _28189_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [17], _00395_, clk);
  dff _28190_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [18], _07338_, clk);
  dff _28191_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [19], _03784_, clk);
  dff _28192_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [20], _01666_, clk);
  dff _28193_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [21], _03688_, clk);
  dff _28194_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [22], _05764_, clk);
  dff _28195_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [23], _11981_, clk);
  dff _28196_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [24], _11162_, clk);
  dff _28197_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [25], _12011_, clk);
  dff _28198_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [26], _01193_, clk);
  dff _28199_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [27], _08287_, clk);
  dff _28200_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [28], _11992_, clk);
  dff _28201_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [29], _02450_, clk);
  dff _28202_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [30], _00159_, clk);
  dff _28203_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [31], _03428_, clk);
  dff _28204_ (\oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _11259_, clk);
  dff _28205_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [0], _03750_, clk);
  dff _28206_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [1], _12003_, clk);
  dff _28207_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [2], _11156_, clk);
  dff _28208_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [3], _03441_, clk);
  dff _28209_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [4], _03439_, clk);
  dff _28210_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [5], _03436_, clk);
  dff _28211_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [6], _03433_, clk);
  dff _28212_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [7], _05672_, clk);
  dff _28213_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [7], _03424_, clk);
  dff _28214_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [7], _06468_, clk);
  dff _28215_ (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _01918_, clk);
  dff _28216_ (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _00894_, clk);
  dff _28217_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [0], _12370_, clk);
  dff _28218_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [1], _12361_, clk);
  dff _28219_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _12346_, clk);
  dff _28220_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [3], _12343_, clk);
  dff _28221_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [4], _12286_, clk);
  dff _28222_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [5], _12275_, clk);
  dff _28223_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [6], _12065_, clk);
  dff _28224_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [7], _12440_, clk);
  dff _28225_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [8], _12523_, clk);
  dff _28226_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [9], _12520_, clk);
  dff _28227_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [10], _12467_, clk);
  dff _28228_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [11], _12058_, clk);
  dff _28229_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [12], _11110_, clk);
  dff _28230_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [13], _11826_, clk);
  dff _28231_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [14], _11798_, clk);
  dff _28232_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [15], _10889_, clk);
  dff _28233_ (\oc8051_top_1.oc8051_memory_interface1.pc [0], _11168_, clk);
  dff _28234_ (\oc8051_top_1.oc8051_memory_interface1.pc [1], _11146_, clk);
  dff _28235_ (\oc8051_top_1.oc8051_memory_interface1.pc [2], _11013_, clk);
  dff _28236_ (\oc8051_top_1.oc8051_memory_interface1.pc [3], _12087_, clk);
  dff _28237_ (\oc8051_top_1.oc8051_memory_interface1.pc [4], _11588_, clk);
  dff _28238_ (\oc8051_top_1.oc8051_memory_interface1.pc [5], _11369_, clk);
  dff _28239_ (\oc8051_top_1.oc8051_memory_interface1.pc [6], _11554_, clk);
  dff _28240_ (\oc8051_top_1.oc8051_memory_interface1.pc [7], _11438_, clk);
  dff _28241_ (\oc8051_top_1.oc8051_memory_interface1.pc [8], _11435_, clk);
  dff _28242_ (\oc8051_top_1.oc8051_memory_interface1.pc [9], _11417_, clk);
  dff _28243_ (\oc8051_top_1.oc8051_memory_interface1.pc [10], _12078_, clk);
  dff _28244_ (\oc8051_top_1.oc8051_memory_interface1.pc [11], _11096_, clk);
  dff _28245_ (\oc8051_top_1.oc8051_memory_interface1.pc [12], _10302_, clk);
  dff _28246_ (\oc8051_top_1.oc8051_memory_interface1.pc [13], _10263_, clk);
  dff _28247_ (\oc8051_top_1.oc8051_memory_interface1.pc [14], _10298_, clk);
  dff _28248_ (\oc8051_top_1.oc8051_memory_interface1.pc [15], _08560_, clk);
  dff _28249_ (\oc8051_top_1.oc8051_memory_interface1.int_ack , _11498_, clk);
  dff _28250_ (\oc8051_top_1.oc8051_memory_interface1.int_ack_t , _01864_, clk);
  dff _28251_ (\oc8051_top_1.oc8051_memory_interface1.int_ack_buff , _11504_, clk);
  dff _28252_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], _00606_, clk);
  dff _28253_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], _07307_, clk);
  dff _28254_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _01713_, clk);
  dff _28255_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], _02537_, clk);
  dff _28256_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _12105_, clk);
  dff _28257_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], _07083_, clk);
  dff _28258_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _06264_, clk);
  dff _28259_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _01884_, clk);
  dff _28260_ (\oc8051_top_1.oc8051_memory_interface1.op_pos [0], _06607_, clk);
  dff _28261_ (\oc8051_top_1.oc8051_memory_interface1.op_pos [1], _12102_, clk);
  dff _28262_ (\oc8051_top_1.oc8051_memory_interface1.op_pos [2], _01887_, clk);
  dff _28263_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [0], _11143_, clk);
  dff _28264_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [1], _11350_, clk);
  dff _28265_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [2], _11047_, clk);
  dff _28266_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [3], _11319_, clk);
  dff _28267_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [4], _11517_, clk);
  dff _28268_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [5], _02376_, clk);
  dff _28269_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [6], _02382_, clk);
  dff _28270_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [0], _01899_, clk);
  dff _28271_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [1], _02089_, clk);
  dff _28272_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [2], _12110_, clk);
  dff _28273_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [3], _11044_, clk);
  dff _28274_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [4], _03705_, clk);
  dff _28275_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [6], _03467_, clk);
  dff _28276_ (\oc8051_top_1.oc8051_memory_interface1.reti , _06484_, clk);
  dff _28277_ (\oc8051_top_1.oc8051_memory_interface1.cdata [0], _11034_, clk);
  dff _28278_ (\oc8051_top_1.oc8051_memory_interface1.cdata [1], _11314_, clk);
  dff _28279_ (\oc8051_top_1.oc8051_memory_interface1.cdata [2], _03660_, clk);
  dff _28280_ (\oc8051_top_1.oc8051_memory_interface1.cdata [3], _03771_, clk);
  dff _28281_ (\oc8051_top_1.oc8051_memory_interface1.cdata [4], _03712_, clk);
  dff _28282_ (\oc8051_top_1.oc8051_memory_interface1.cdata [5], _03679_, clk);
  dff _28283_ (\oc8051_top_1.oc8051_memory_interface1.cdata [6], _12135_, clk);
  dff _28284_ (\oc8051_top_1.oc8051_memory_interface1.cdata [7], _06592_, clk);
  dff _28285_ (\oc8051_top_1.oc8051_memory_interface1.cdone , _06691_, clk);
  dff _28286_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst , _08435_, clk);
  dff _28287_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], _02706_, clk);
  dff _28288_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], _02519_, clk);
  dff _28289_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], _02238_, clk);
  dff _28290_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], _10089_, clk);
  dff _28291_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [0], _10928_, clk);
  dff _28292_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [1], _10269_, clk);
  dff _28293_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [2], _10033_, clk);
  dff _28294_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [3], _11104_, clk);
  dff _28295_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [4], _11055_, clk);
  dff _28296_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [5], _10640_, clk);
  dff _28297_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [6], _12070_, clk);
  dff _28298_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [7], _11215_, clk);
  dff _28299_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [8], _10637_, clk);
  dff _28300_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [9], _00071_, clk);
  dff _28301_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [10], _12079_, clk);
  dff _28302_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [11], _10634_, clk);
  dff _28303_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [12], _10813_, clk);
  dff _28304_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [13], _10916_, clk);
  dff _28305_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [14], _10985_, clk);
  dff _28306_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [15], _00206_, clk);
  dff _28307_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [16], _00201_, clk);
  dff _28308_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [17], _10631_, clk);
  dff _28309_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [18], _00771_, clk);
  dff _28310_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [19], _00291_, clk);
  dff _28311_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [20], _10628_, clk);
  dff _28312_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [21], _10810_, clk);
  dff _28313_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [22], _01797_, clk);
  dff _28314_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [23], _01352_, clk);
  dff _28315_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [24], _10625_, clk);
  dff _28316_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [25], _02571_, clk);
  dff _28317_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [26], _01817_, clk);
  dff _28318_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [27], _10623_, clk);
  dff _28319_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [28], _10807_, clk);
  dff _28320_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [29], _10903_, clk);
  dff _28321_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [30], _02708_, clk);
  dff _28322_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [31], _03415_, clk);
  dff _28323_ (\oc8051_top_1.oc8051_memory_interface1.dmem_wait , _02253_, clk);
  dff _28324_ (\oc8051_top_1.oc8051_memory_interface1.istb_t , _01664_, clk);
  dff _28325_ (\oc8051_top_1.oc8051_memory_interface1.imem_wait , _01761_, clk);
  dff _28326_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _03814_, clk);
  dff _28327_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _03775_, clk);
  dff _28328_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _10604_, clk);
  dff _28329_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _10731_, clk);
  dff _28330_ (\oc8051_top_1.oc8051_memory_interface1.rd_ind , _02255_, clk);
  dff _28331_ (\oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0], clk);
  dff _28332_ (\oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1], clk);
  dff _28333_ (\oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2], clk);
  dff _28334_ (\oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3], clk);
  dff _28335_ (\oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4], clk);
  dff _28336_ (\oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5], clk);
  dff _28337_ (\oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6], clk);
  dff _28338_ (\oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7], clk);
  dff _28339_ (\oc8051_top_1.oc8051_rom1.data_o [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8], clk);
  dff _28340_ (\oc8051_top_1.oc8051_rom1.data_o [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9], clk);
  dff _28341_ (\oc8051_top_1.oc8051_rom1.data_o [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10], clk);
  dff _28342_ (\oc8051_top_1.oc8051_rom1.data_o [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11], clk);
  dff _28343_ (\oc8051_top_1.oc8051_rom1.data_o [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12], clk);
  dff _28344_ (\oc8051_top_1.oc8051_rom1.data_o [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13], clk);
  dff _28345_ (\oc8051_top_1.oc8051_rom1.data_o [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14], clk);
  dff _28346_ (\oc8051_top_1.oc8051_rom1.data_o [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15], clk);
  dff _28347_ (\oc8051_top_1.oc8051_rom1.data_o [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16], clk);
  dff _28348_ (\oc8051_top_1.oc8051_rom1.data_o [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17], clk);
  dff _28349_ (\oc8051_top_1.oc8051_rom1.data_o [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18], clk);
  dff _28350_ (\oc8051_top_1.oc8051_rom1.data_o [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19], clk);
  dff _28351_ (\oc8051_top_1.oc8051_rom1.data_o [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20], clk);
  dff _28352_ (\oc8051_top_1.oc8051_rom1.data_o [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21], clk);
  dff _28353_ (\oc8051_top_1.oc8051_rom1.data_o [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22], clk);
  dff _28354_ (\oc8051_top_1.oc8051_rom1.data_o [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23], clk);
  dff _28355_ (\oc8051_top_1.oc8051_rom1.data_o [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24], clk);
  dff _28356_ (\oc8051_top_1.oc8051_rom1.data_o [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25], clk);
  dff _28357_ (\oc8051_top_1.oc8051_rom1.data_o [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26], clk);
  dff _28358_ (\oc8051_top_1.oc8051_rom1.data_o [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27], clk);
  dff _28359_ (\oc8051_top_1.oc8051_rom1.data_o [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28], clk);
  dff _28360_ (\oc8051_top_1.oc8051_rom1.data_o [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29], clk);
  dff _28361_ (\oc8051_top_1.oc8051_rom1.data_o [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30], clk);
  dff _28362_ (\oc8051_top_1.oc8051_rom1.data_o [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31], clk);
  dff _28363_ (\oc8051_top_1.oc8051_sfr1.pres_ow , _04133_, clk);
  dff _28364_ (\oc8051_top_1.oc8051_sfr1.prescaler [0], _12084_, clk);
  dff _28365_ (\oc8051_top_1.oc8051_sfr1.prescaler [1], _12115_, clk);
  dff _28366_ (\oc8051_top_1.oc8051_sfr1.prescaler [2], _12113_, clk);
  dff _28367_ (\oc8051_top_1.oc8051_sfr1.prescaler [3], _04039_, clk);
  dff _28368_ (\oc8051_top_1.oc8051_sfr1.bit_out , _04154_, clk);
  dff _28369_ (\oc8051_top_1.oc8051_sfr1.wait_data , _04147_, clk);
  dff _28370_ (\oc8051_top_1.oc8051_sfr1.dat0 [0], _11841_, clk);
  dff _28371_ (\oc8051_top_1.oc8051_sfr1.dat0 [1], _11897_, clk);
  dff _28372_ (\oc8051_top_1.oc8051_sfr1.dat0 [2], _11894_, clk);
  dff _28373_ (\oc8051_top_1.oc8051_sfr1.dat0 [3], _11888_, clk);
  dff _28374_ (\oc8051_top_1.oc8051_sfr1.dat0 [4], _11885_, clk);
  dff _28375_ (\oc8051_top_1.oc8051_sfr1.dat0 [5], _03665_, clk);
  dff _28376_ (\oc8051_top_1.oc8051_sfr1.dat0 [6], _03526_, clk);
  dff _28377_ (\oc8051_top_1.oc8051_sfr1.dat0 [7], _04036_, clk);
  dff _28378_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], _11659_, clk);
  dff _28379_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], _07973_, clk);
  dff _28380_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], _02456_, clk);
  dff _28381_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3], _11049_, clk);
  dff _28382_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4], _02458_, clk);
  dff _28383_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], _01630_, clk);
  dff _28384_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], _07968_, clk);
  dff _28385_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], _05610_, clk);
  dff _28386_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0], _03603_, clk);
  dff _28387_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1], _00815_, clk);
  dff _28388_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2], _00807_, clk);
  dff _28389_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3], _03593_, clk);
  dff _28390_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4], _00533_, clk);
  dff _28391_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5], _00530_, clk);
  dff _28392_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6], _03638_, clk);
  dff _28393_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7], _03895_, clk);
  dff _28394_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], _07113_, clk);
  dff _28395_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], _07107_, clk);
  dff _28396_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], _07109_, clk);
  dff _28397_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], _05863_, clk);
  dff _28398_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], _02168_, clk);
  dff _28399_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], _05871_, clk);
  dff _28400_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], _05866_, clk);
  dff _28401_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7], _03398_, clk);
  dff _28402_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0], _05929_, clk);
  dff _28403_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1], _07080_, clk);
  dff _28404_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2], _07085_, clk);
  dff _28405_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3], _05899_, clk);
  dff _28406_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4], _02153_, clk);
  dff _28407_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5], _04295_, clk);
  dff _28408_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6], _05932_, clk);
  dff _28409_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7], _12026_, clk);
  dff _28410_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff , _10951_, clk);
  dff _28411_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], _02677_, clk);
  dff _28412_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], _13282_, clk);
  dff _28413_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _13271_, clk);
  dff _28414_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3], _13279_, clk);
  dff _28415_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4], _13276_, clk);
  dff _28416_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], _02867_, clk);
  dff _28417_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _13296_, clk);
  dff _28418_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _02498_, clk);
  dff _28419_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], _02636_, clk);
  dff _28420_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _04077_, clk);
  dff _28421_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc , _03681_, clk);
  dff _28422_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _13262_, clk);
  dff _28423_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _13250_, clk);
  dff _28424_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], _03329_, clk);
  dff _28425_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _02668_, clk);
  dff _28426_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _13150_, clk);
  dff _28427_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], _12455_, clk);
  dff _28428_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], _13142_, clk);
  dff _28429_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _13175_, clk);
  dff _28430_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , _00274_, clk);
  dff _28431_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , _00269_, clk);
  dff _28432_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , _08444_, clk);
  dff _28433_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , _10257_, clk);
  dff _28434_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0], _13109_, clk);
  dff _28435_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1], _13106_, clk);
  dff _28436_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2], _02889_, clk);
  dff _28437_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], _10254_, clk);
  dff _28438_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0], _13569_, clk);
  dff _28439_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], _13564_, clk);
  dff _28440_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], _13558_, clk);
  dff _28441_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3], _02805_, clk);
  dff _28442_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4], _13590_, clk);
  dff _28443_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5], _13587_, clk);
  dff _28444_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6], _13580_, clk);
  dff _28445_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _00336_, clk);
  dff _28446_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0], _13543_, clk);
  dff _28447_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1], _02815_, clk);
  dff _28448_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2], _02654_, clk);
  dff _28449_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3], _13493_, clk);
  dff _28450_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4], _13490_, clk);
  dff _28451_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5], _13483_, clk);
  dff _28452_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6], _02821_, clk);
  dff _28453_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7], _04414_, clk);
  dff _28454_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0], _03138_, clk);
  dff _28455_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1], _03305_, clk);
  dff _28456_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2], _03170_, clk);
  dff _28457_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3], _03136_, clk);
  dff _28458_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4], _03309_, clk);
  dff _28459_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5], _03172_, clk);
  dff _28460_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6], _03307_, clk);
  dff _28461_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7], _03623_, clk);
  dff _28462_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0], _03283_, clk);
  dff _28463_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1], _03164_, clk);
  dff _28464_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2], _03132_, clk);
  dff _28465_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3], _03314_, clk);
  dff _28466_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4], _03167_, clk);
  dff _28467_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5], _03312_, clk);
  dff _28468_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6], _03162_, clk);
  dff _28469_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7], _05142_, clk);
  dff _28470_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0], _03134_, clk);
  dff _28471_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1], _03311_, clk);
  dff _28472_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2], _03281_, clk);
  dff _28473_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3], _03257_, clk);
  dff _28474_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4], _03256_, clk);
  dff _28475_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5], _03160_, clk);
  dff _28476_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6], _03128_, clk);
  dff _28477_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7], _02004_, clk);
  dff _28478_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0], _03126_, clk);
  dff _28479_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1], _03317_, clk);
  dff _28480_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2], _03287_, clk);
  dff _28481_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3], _03286_, clk);
  dff _28482_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4], _03322_, clk);
  dff _28483_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5], _03158_, clk);
  dff _28484_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6], _03320_, clk);
  dff _28485_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7], _03760_, clk);
  dff _28486_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1], _06900_, clk);
  dff _28487_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], _06894_, clk);
  dff _28488_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3], _10119_, clk);
  dff _28489_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4], _06964_, clk);
  dff _28490_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5], _07223_, clk);
  dff _28491_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6], _07139_, clk);
  dff _28492_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], _04069_, clk);
  dff _28493_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop , _00271_, clk);
  dff _28494_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], _13680_, clk);
  dff _28495_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], _03675_, clk);
  dff _28496_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2], _13726_, clk);
  dff _28497_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3], _13709_, clk);
  dff _28498_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4], _13720_, clk);
  dff _28499_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5], _13717_, clk);
  dff _28500_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6], _13714_, clk);
  dff _28501_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7], _03651_, clk);
  dff _28502_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , _01080_, clk);
  dff _28503_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff , _01083_, clk);
  dff _28504_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0], _13154_, clk);
  dff _28505_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1], _13163_, clk);
  dff _28506_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2], _13167_, clk);
  dff _28507_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3], _13135_, clk);
  dff _28508_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4], _13132_, clk);
  dff _28509_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], _13129_, clk);
  dff _28510_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6], _13139_, clk);
  dff _28511_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7], _01094_, clk);
  dff _28512_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0], _13197_, clk);
  dff _28513_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1], _13191_, clk);
  dff _28514_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2], _13194_, clk);
  dff _28515_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3], _13212_, clk);
  dff _28516_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4], _13203_, clk);
  dff _28517_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5], _13209_, clk);
  dff _28518_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6], _13206_, clk);
  dff _28519_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7], _01088_, clk);
  dff _28520_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , _01092_, clk);
  dff _28521_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _01090_, clk);
  dff _28522_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0], _13219_, clk);
  dff _28523_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1], _13215_, clk);
  dff _28524_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2], _13237_, clk);
  dff _28525_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3], _13245_, clk);
  dff _28526_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4], _13242_, clk);
  dff _28527_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], _13301_, clk);
  dff _28528_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6], _13293_, clk);
  dff _28529_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7], _01042_, clk);
  dff _28530_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0], _13370_, clk);
  dff _28531_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1], _13364_, clk);
  dff _28532_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2], _13338_, clk);
  dff _28533_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3], _13340_, clk);
  dff _28534_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4], _13348_, clk);
  dff _28535_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5], _13351_, clk);
  dff _28536_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6], _13330_, clk);
  dff _28537_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7], _01046_, clk);
  dff _28538_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 , _01044_, clk);
  dff _28539_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _13376_, clk);
  dff _28540_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], _13378_, clk);
  dff _28541_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2], _13396_, clk);
  dff _28542_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3], _13388_, clk);
  dff _28543_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _13393_, clk);
  dff _28544_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], _13406_, clk);
  dff _28545_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6], _13403_, clk);
  dff _28546_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7], _01057_, clk);
  dff _28547_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r , _03495_, clk);
  dff _28548_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _02435_, clk);
  dff _28549_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , _02074_, clk);
  dff _28550_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r , _01863_, clk);
  dff _28551_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0], _01549_, clk);
  dff _28552_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1], _01547_, clk);
  dff _28553_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2], _01545_, clk);
  dff _28554_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3], _01542_, clk);
  dff _28555_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4], _01539_, clk);
  dff _28556_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5], _01490_, clk);
  dff _28557_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6], _01480_, clk);
  dff _28558_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7], _09910_, clk);
  dff _28559_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0], _01421_, clk);
  dff _28560_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1], _01403_, clk);
  dff _28561_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2], _01363_, clk);
  dff _28562_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3], _01395_, clk);
  dff _28563_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4], _01391_, clk);
  dff _28564_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5], _01387_, clk);
  dff _28565_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6], _01366_, clk);
  dff _28566_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7], _01794_, clk);
  dff _28567_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 , _03966_, clk);
  dff _28568_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0], _01265_, clk);
  dff _28569_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1], _01216_, clk);
  dff _28570_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2], _01201_, clk);
  dff _28571_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3], _01211_, clk);
  dff _28572_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4], _01207_, clk);
  dff _28573_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5], _01182_, clk);
  dff _28574_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6], _01169_, clk);
  dff _28575_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7], _03493_, clk);
  dff _28576_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0], _01143_, clk);
  dff _28577_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1], _01103_, clk);
  dff _28578_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2], _01097_, clk);
  dff _28579_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3], _01086_, clk);
  dff _28580_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4], _01037_, clk);
  dff _28581_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5], _01034_, clk);
  dff _28582_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6], _01028_, clk);
  dff _28583_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7], _03078_, clk);
  dff _28584_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set , _00793_, clk);
  dff _28585_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0], _00990_, clk);
  dff _28586_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1], _00970_, clk);
  dff _28587_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2], _00966_, clk);
  dff _28588_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3], _00930_, clk);
  dff _28589_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], _00928_, clk);
  dff _28590_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], _00922_, clk);
  dff _28591_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6], _00917_, clk);
  dff _28592_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], _00514_, clk);
  dff _28593_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0], _05541_, clk);
  dff _28594_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1], _05540_, clk);
  dff _28595_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2], _05539_, clk);
  dff _28596_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _02328_, clk);
  dff _28597_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _01099_, clk);
  dff _28598_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _02117_, clk);
  dff _28599_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _01904_, clk);
  dff _28600_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _11021_, clk);
  dff _28601_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8], _03276_, clk);
  dff _28602_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9], _00342_, clk);
  dff _28603_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], _00604_, clk);
  dff _28604_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _02834_, clk);
  dff _28605_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf , _11823_, clk);
  dff _28606_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , _01686_, clk);
  dff _28607_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , _10954_, clk);
  dff _28608_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive , _02779_, clk);
  dff _28609_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _03346_, clk);
  dff _28610_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r , _01680_, clk);
  dff _28611_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], _03881_, clk);
  dff _28612_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1], _07822_, clk);
  dff _28613_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], _11357_, clk);
  dff _28614_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], _06338_, clk);
  dff _28615_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _07180_, clk);
  dff _28616_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3], _07858_, clk);
  dff _28617_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0], _02540_, clk);
  dff _28618_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1], _06460_, clk);
  dff _28619_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2], _10900_, clk);
  dff _28620_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3], _02468_, clk);
  dff _28621_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4], _02465_, clk);
  dff _28622_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5], _02474_, clk);
  dff _28623_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6], _11758_, clk);
  dff _28624_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7], _09164_, clk);
  dff _28625_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr , _02831_, clk);
  dff _28626_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr , _02739_, clk);
  dff _28627_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans , _02836_, clk);
  dff _28628_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , _02736_, clk);
  dff _28629_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0], _00684_, clk);
  dff _28630_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1], _00682_, clk);
  dff _28631_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2], _12067_, clk);
  dff _28632_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3], _02766_, clk);
  dff _28633_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0], _01355_, clk);
  dff _28634_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1], _12055_, clk);
  dff _28635_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], _03048_, clk);
  dff _28636_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3], _03014_, clk);
  dff _28637_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4], _12049_, clk);
  dff _28638_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5], _12191_, clk);
  dff _28639_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6], _12326_, clk);
  dff _28640_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7], _12358_, clk);
  dff _28641_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8], _03153_, clk);
  dff _28642_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], _03075_, clk);
  dff _28643_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10], _02853_, clk);
  dff _28644_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0], _03714_, clk);
  dff _28645_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1], _03522_, clk);
  dff _28646_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2], _12042_, clk);
  dff _28647_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3], _12158_, clk);
  dff _28648_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4], _12323_, clk);
  dff _28649_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5], _03844_, clk);
  dff _28650_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6], _03718_, clk);
  dff _28651_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], _02851_, clk);
  dff _28652_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0], _03974_, clk);
  dff _28653_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], _12023_, clk);
  dff _28654_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2], _12151_, clk);
  dff _28655_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3], _12294_, clk);
  dff _28656_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], _12356_, clk);
  dff _28657_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5], _12383_, clk);
  dff _28658_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6], _04020_, clk);
  dff _28659_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], _02726_, clk);
  buf(\oc8051_top_1.oc8051_indi_addr1.rst , rst);
  buf(\oc8051_top_1.oc8051_indi_addr1.clk , clk);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.oc8051_rom1.clk , clk);
  buf(\oc8051_top_1.oc8051_rom1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk , clk);
  buf(\oc8051_top_1.oc8051_decoder1.new_valid_pc , pc_log_change);
  buf(\oc8051_top_1.oc8051_decoder1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.oc8051_decoder1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.oc8051_decoder1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.ip [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.wr_bit_r , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_sfr1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div1 , \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div0 , \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [0], \oc8051_top_1.oc8051_memory_interface1.op2_buff [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [1], \oc8051_top_1.oc8051_memory_interface1.op2_buff [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [2], \oc8051_top_1.oc8051_memory_interface1.op2_buff [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [3], \oc8051_top_1.oc8051_memory_interface1.op2_buff [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [4], \oc8051_top_1.oc8051_memory_interface1.op2_buff [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [5], \oc8051_top_1.oc8051_memory_interface1.op2_buff [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [6], \oc8051_top_1.oc8051_memory_interface1.op2_buff [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [7], \oc8051_top_1.oc8051_memory_interface1.imm_r [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3_r [0], \oc8051_top_1.oc8051_memory_interface1.op3_buff [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3_r [1], \oc8051_top_1.oc8051_memory_interface1.op3_buff [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3_r [2], \oc8051_top_1.oc8051_memory_interface1.op3_buff [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3_r [3], \oc8051_top_1.oc8051_memory_interface1.op3_buff [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3_r [4], \oc8051_top_1.oc8051_memory_interface1.op3_buff [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3_r [6], \oc8051_top_1.oc8051_memory_interface1.op3_buff [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3_r [7], \oc8051_top_1.oc8051_memory_interface1.imm2_r [7]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_in , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_symbolic_cxrom1.clk , clk);
  buf(\oc8051_symbolic_cxrom1.rst , rst);
  buf(\oc8051_symbolic_cxrom1.word_in [0], word_in[0]);
  buf(\oc8051_symbolic_cxrom1.word_in [1], word_in[1]);
  buf(\oc8051_symbolic_cxrom1.word_in [2], word_in[2]);
  buf(\oc8051_symbolic_cxrom1.word_in [3], word_in[3]);
  buf(\oc8051_symbolic_cxrom1.word_in [4], word_in[4]);
  buf(\oc8051_symbolic_cxrom1.word_in [5], word_in[5]);
  buf(\oc8051_symbolic_cxrom1.word_in [6], word_in[6]);
  buf(\oc8051_symbolic_cxrom1.word_in [7], word_in[7]);
  buf(\oc8051_symbolic_cxrom1.word_in [8], word_in[8]);
  buf(\oc8051_symbolic_cxrom1.word_in [9], word_in[9]);
  buf(\oc8051_symbolic_cxrom1.word_in [10], word_in[10]);
  buf(\oc8051_symbolic_cxrom1.word_in [11], word_in[11]);
  buf(\oc8051_symbolic_cxrom1.word_in [12], word_in[12]);
  buf(\oc8051_symbolic_cxrom1.word_in [13], word_in[13]);
  buf(\oc8051_symbolic_cxrom1.word_in [14], word_in[14]);
  buf(\oc8051_symbolic_cxrom1.word_in [15], word_in[15]);
  buf(\oc8051_symbolic_cxrom1.word_in [16], word_in[16]);
  buf(\oc8051_symbolic_cxrom1.word_in [17], word_in[17]);
  buf(\oc8051_symbolic_cxrom1.word_in [18], word_in[18]);
  buf(\oc8051_symbolic_cxrom1.word_in [19], word_in[19]);
  buf(\oc8051_symbolic_cxrom1.word_in [20], word_in[20]);
  buf(\oc8051_symbolic_cxrom1.word_in [21], word_in[21]);
  buf(\oc8051_symbolic_cxrom1.word_in [22], word_in[22]);
  buf(\oc8051_symbolic_cxrom1.word_in [23], word_in[23]);
  buf(\oc8051_symbolic_cxrom1.word_in [24], word_in[24]);
  buf(\oc8051_symbolic_cxrom1.word_in [25], word_in[25]);
  buf(\oc8051_symbolic_cxrom1.word_in [26], word_in[26]);
  buf(\oc8051_symbolic_cxrom1.word_in [27], word_in[27]);
  buf(\oc8051_symbolic_cxrom1.word_in [28], word_in[28]);
  buf(\oc8051_symbolic_cxrom1.word_in [29], word_in[29]);
  buf(\oc8051_symbolic_cxrom1.word_in [30], word_in[30]);
  buf(\oc8051_symbolic_cxrom1.word_in [31], word_in[31]);
  buf(\oc8051_symbolic_cxrom1.pc1 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc1 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_symbolic_cxrom1.pc1 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_symbolic_cxrom1.pc1 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_symbolic_cxrom1.pc1 [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_symbolic_cxrom1.pc1 [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_symbolic_cxrom1.pc1 [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_symbolic_cxrom1.pc1 [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_symbolic_cxrom1.pc1 [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_symbolic_cxrom1.pc1 [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_symbolic_cxrom1.pc1 [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_symbolic_cxrom1.pc1 [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_symbolic_cxrom1.pc1 [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_symbolic_cxrom1.pc1 [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_symbolic_cxrom1.pc1 [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_symbolic_cxrom1.pc1 [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_symbolic_cxrom1.pc2 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_symbolic_cxrom1.pc2 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_symbolic_cxrom1.pc2 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_symbolic_cxrom1.pc2 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_symbolic_cxrom1.pc2 [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_symbolic_cxrom1.pc2 [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_symbolic_cxrom1.pc2 [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_symbolic_cxrom1.pc2 [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_symbolic_cxrom1.pc2 [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_symbolic_cxrom1.pc2 [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_symbolic_cxrom1.pc2 [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_symbolic_cxrom1.pc2 [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_symbolic_cxrom1.pc2 [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_symbolic_cxrom1.pc2 [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_symbolic_cxrom1.pc2 [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_symbolic_cxrom1.pc2 [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [0], word_in[0]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [1], word_in[1]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [2], word_in[2]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [3], word_in[3]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [4], word_in[4]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [5], word_in[5]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [6], word_in[6]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [7], word_in[7]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [0], word_in[8]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [1], word_in[9]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [2], word_in[10]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [3], word_in[11]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [4], word_in[12]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [5], word_in[13]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [6], word_in[14]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [7], word_in[15]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [0], word_in[16]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [1], word_in[17]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [2], word_in[18]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [3], word_in[19]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [4], word_in[20]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [5], word_in[21]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [6], word_in[22]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [7], word_in[23]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [0], word_in[24]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [1], word_in[25]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [2], word_in[26]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [3], word_in[27]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [4], word_in[28]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [5], word_in[29]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [6], word_in[30]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [7], word_in[31]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_symbolic_cxrom1.pc10 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc10 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_symbolic_cxrom1.pc10 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_symbolic_cxrom1.pc10 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_symbolic_cxrom1.pc12 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc12 [1], pc1_plus_2[1]);
  buf(\oc8051_symbolic_cxrom1.pc12 [2], pc1_plus_2[2]);
  buf(\oc8051_symbolic_cxrom1.pc12 [3], pc1_plus_2[3]);
  buf(\oc8051_symbolic_cxrom1.pc20 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_symbolic_cxrom1.pc20 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_symbolic_cxrom1.pc20 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_symbolic_cxrom1.pc20 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_symbolic_cxrom1.pc22 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.clk , clk);
  buf(\oc8051_top_1.oc8051_comp1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_comp1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_comp1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_comp1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_comp1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_comp1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_comp1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_comp1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_comp1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_alu1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [4], \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [5], \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.uart_int , \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.t2_int , \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.rst , rst);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_for_ajmp [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [0], \oc8051_top_1.oc8051_sfr1.psw [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.p , \oc8051_top_1.oc8051_sfr1.psw [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_out [0], \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_out [1], \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [5], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [7], \oc8051_top_1.oc8051_memory_interface1.imm2_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [7], \oc8051_top_1.oc8051_memory_interface1.imm_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [0], \oc8051_top_1.oc8051_memory_interface1.op3_buff [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [1], \oc8051_top_1.oc8051_memory_interface1.op3_buff [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [2], \oc8051_top_1.oc8051_memory_interface1.op3_buff [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [3], \oc8051_top_1.oc8051_memory_interface1.op3_buff [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [4], \oc8051_top_1.oc8051_memory_interface1.op3_buff [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [5], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [6], \oc8051_top_1.oc8051_memory_interface1.op3_buff [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [0], \oc8051_top_1.oc8051_memory_interface1.op2_buff [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [1], \oc8051_top_1.oc8051_memory_interface1.op2_buff [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [2], \oc8051_top_1.oc8051_memory_interface1.op2_buff [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [3], \oc8051_top_1.oc8051_memory_interface1.op2_buff [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [4], \oc8051_top_1.oc8051_memory_interface1.op2_buff [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [5], \oc8051_top_1.oc8051_memory_interface1.op2_buff [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [6], \oc8051_top_1.oc8051_memory_interface1.op2_buff [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.ABINPUT [0], ABINPUT[0]);
  buf(\oc8051_top_1.ABINPUT [1], ABINPUT[1]);
  buf(\oc8051_top_1.ABINPUT [2], ABINPUT[2]);
  buf(\oc8051_top_1.ABINPUT [3], ABINPUT[3]);
  buf(\oc8051_top_1.ABINPUT [4], ABINPUT[4]);
  buf(\oc8051_top_1.ABINPUT [5], ABINPUT[5]);
  buf(\oc8051_top_1.ABINPUT [6], ABINPUT[6]);
  buf(\oc8051_top_1.ABINPUT [7], ABINPUT[7]);
  buf(\oc8051_top_1.ABINPUT [8], ABINPUT[8]);
  buf(\oc8051_top_1.wb_rst_i , rst);
  buf(\oc8051_top_1.wb_clk_i , clk);
  buf(\oc8051_top_1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.bit_data , ABINPUT[0]);
  buf(\oc8051_top_1.rd_ind , \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  buf(\oc8051_top_1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.decoder_new_valid_pc , pc_log_change);
  buf(\oc8051_top_1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.sfr_out [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.sfr_out [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.sfr_out [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.sfr_out [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.sfr_out [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.sfr_out [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.sfr_out [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.sfr_out [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.ram_data [0], ABINPUT[1]);
  buf(\oc8051_top_1.ram_data [1], ABINPUT[2]);
  buf(\oc8051_top_1.ram_data [2], ABINPUT[3]);
  buf(\oc8051_top_1.ram_data [3], ABINPUT[4]);
  buf(\oc8051_top_1.ram_data [4], ABINPUT[5]);
  buf(\oc8051_top_1.ram_data [5], ABINPUT[6]);
  buf(\oc8051_top_1.ram_data [6], ABINPUT[7]);
  buf(\oc8051_top_1.ram_data [7], ABINPUT[8]);
  buf(\oc8051_top_1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.src_sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.src_sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.pc_log_change , pc_log_change);
  buf(\oc8051_top_1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_top_1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_top_1.pc_log [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_top_1.pc_log [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_top_1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_top_1.pc_log [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_top_1.pc_log [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_top_1.pc_log [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_top_1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_top_1.pc_log [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_top_1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_top_1.pc_log [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_top_1.pc_log [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_top_1.pc_log [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_top_1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_top_1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_top_1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_top_1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_top_1.pc_log_prev [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_top_1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_top_1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_top_1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_top_1.pc_log_prev [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_top_1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_top_1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_top_1.pc_log_prev [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_top_1.pc_log_prev [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_top_1.pc_log_prev [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_top_1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_top_1.pc_log_prev [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_top_1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_top_1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.t2ex_i , t2ex_i);
  buf(\oc8051_top_1.t2_i , t2_i);
  buf(\oc8051_top_1.t1_i , t1_i);
  buf(\oc8051_top_1.t0_i , t0_i);
  buf(\oc8051_top_1.rxd_i , rxd_i);
  buf(\oc8051_top_1.p3_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.p3_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.p3_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.p3_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.p3_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.p3_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.p3_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.p3_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.p3_i [0], p3_in[0]);
  buf(\oc8051_top_1.p3_i [1], p3_in[1]);
  buf(\oc8051_top_1.p3_i [2], p3_in[2]);
  buf(\oc8051_top_1.p3_i [3], p3_in[3]);
  buf(\oc8051_top_1.p3_i [4], p3_in[4]);
  buf(\oc8051_top_1.p3_i [5], p3_in[5]);
  buf(\oc8051_top_1.p3_i [6], p3_in[6]);
  buf(\oc8051_top_1.p3_i [7], p3_in[7]);
  buf(\oc8051_top_1.p2_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.p2_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.p2_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.p2_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.p2_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.p2_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.p2_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.p2_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.p2_i [0], p2_in[0]);
  buf(\oc8051_top_1.p2_i [1], p2_in[1]);
  buf(\oc8051_top_1.p2_i [2], p2_in[2]);
  buf(\oc8051_top_1.p2_i [3], p2_in[3]);
  buf(\oc8051_top_1.p2_i [4], p2_in[4]);
  buf(\oc8051_top_1.p2_i [5], p2_in[5]);
  buf(\oc8051_top_1.p2_i [6], p2_in[6]);
  buf(\oc8051_top_1.p2_i [7], p2_in[7]);
  buf(\oc8051_top_1.p1_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.p1_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.p1_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.p1_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.p1_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.p1_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.p1_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.p1_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.p1_i [0], p1_in[0]);
  buf(\oc8051_top_1.p1_i [1], p1_in[1]);
  buf(\oc8051_top_1.p1_i [2], p1_in[2]);
  buf(\oc8051_top_1.p1_i [3], p1_in[3]);
  buf(\oc8051_top_1.p1_i [4], p1_in[4]);
  buf(\oc8051_top_1.p1_i [5], p1_in[5]);
  buf(\oc8051_top_1.p1_i [6], p1_in[6]);
  buf(\oc8051_top_1.p1_i [7], p1_in[7]);
  buf(\oc8051_top_1.p0_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.p0_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.p0_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.p0_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.p0_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.p0_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.p0_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.p0_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.p0_i [0], p0_in[0]);
  buf(\oc8051_top_1.p0_i [1], p0_in[1]);
  buf(\oc8051_top_1.p0_i [2], p0_in[2]);
  buf(\oc8051_top_1.p0_i [3], p0_in[3]);
  buf(\oc8051_top_1.p0_i [4], p0_in[4]);
  buf(\oc8051_top_1.p0_i [5], p0_in[5]);
  buf(\oc8051_top_1.p0_i [6], p0_in[6]);
  buf(\oc8051_top_1.p0_i [7], p0_in[7]);
  buf(\oc8051_top_1.cxrom_data_out [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.cxrom_data_out [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.cxrom_data_out [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.cxrom_data_out [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.cxrom_data_out [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.cxrom_data_out [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.cxrom_data_out [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.cxrom_data_out [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.cxrom_data_out [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.cxrom_data_out [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.cxrom_data_out [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.cxrom_data_out [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.cxrom_data_out [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.cxrom_data_out [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.cxrom_data_out [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.cxrom_data_out [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.cxrom_data_out [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.cxrom_data_out [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.cxrom_data_out [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.cxrom_data_out [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.cxrom_data_out [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.cxrom_data_out [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.cxrom_data_out [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.cxrom_data_out [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.cxrom_data_out [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.cxrom_data_out [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.cxrom_data_out [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.cxrom_data_out [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.cxrom_data_out [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.cxrom_data_out [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.cxrom_data_out [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.cxrom_data_out [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.decoder_new_valid_pc , pc_log_change);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [0], ABINPUT[1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [1], ABINPUT[2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [2], ABINPUT[3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [3], ABINPUT[4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [4], ABINPUT[5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [5], ABINPUT[6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [6], ABINPUT[7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [7], ABINPUT[8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.oc8051_memory_interface1.bit_in , ABINPUT[0]);
  buf(cy, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(pc1[0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(pc1[1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(pc1[2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(pc1[3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(pc1[4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(pc1[5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(pc1[6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(pc1[7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(pc1[8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(pc1[9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(pc1[10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(pc1[11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(pc1[12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(pc1[13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(pc1[14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(pc1[15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(pc2[0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(pc2[1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(pc2[2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(pc2[3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(pc2[4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(pc2[5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(pc2[6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(pc2[7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(pc2[8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(pc2[9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(pc2[10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(pc2[11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(pc2[12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(pc2[13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(pc2[14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(pc2[15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(cxrom_data_out[0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(cxrom_data_out[1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(cxrom_data_out[2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(cxrom_data_out[3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(cxrom_data_out[4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(cxrom_data_out[5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(cxrom_data_out[6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(cxrom_data_out[7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(cxrom_data_out[8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(cxrom_data_out[9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(cxrom_data_out[10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(cxrom_data_out[11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(cxrom_data_out[12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(cxrom_data_out[13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(cxrom_data_out[14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(cxrom_data_out[15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(cxrom_data_out[16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(cxrom_data_out[17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(cxrom_data_out[18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(cxrom_data_out[19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(cxrom_data_out[20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(cxrom_data_out[21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(cxrom_data_out[22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(cxrom_data_out[23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(cxrom_data_out[24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(cxrom_data_out[25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(cxrom_data_out[26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(cxrom_data_out[27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(cxrom_data_out[28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(cxrom_data_out[29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(cxrom_data_out[30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(cxrom_data_out[31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk , clk);
  buf(pc1_plus_2[0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(p3_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(p3_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(p3_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(p3_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(p3_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(p3_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(p3_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(p3_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(p2_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(p2_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(p2_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(p2_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(p2_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(p2_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(p2_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(p2_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(p1_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(p1_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(p1_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(p1_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(p1_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(p1_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(p1_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(p1_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(p0_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(p0_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(p0_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(p0_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(p0_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(p0_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(p0_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(p0_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
endmodule
