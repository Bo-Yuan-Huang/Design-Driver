
module oc8051_fv_top(clk, rst, word_in, p0_in, p1_in, p2_in, p3_in, rxd_i, t0_i, t1_i, t2_i, t2ex_i, property_invalid, ABINPUT);
  wire _00000_;
  wire _00001_;
  wire _00002_;
  wire _00003_;
  wire _00004_;
  wire _00005_;
  wire _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  wire _08001_;
  wire _08002_;
  wire _08003_;
  wire _08004_;
  wire _08005_;
  wire _08006_;
  wire _08007_;
  wire _08008_;
  wire _08009_;
  wire _08010_;
  wire _08011_;
  wire _08012_;
  wire _08013_;
  wire _08014_;
  wire _08015_;
  wire _08016_;
  wire _08017_;
  wire _08018_;
  wire _08019_;
  wire _08020_;
  wire _08021_;
  wire _08022_;
  wire _08023_;
  wire _08024_;
  wire _08025_;
  wire _08026_;
  wire _08027_;
  wire _08028_;
  wire _08029_;
  wire _08030_;
  wire _08031_;
  wire _08032_;
  wire _08033_;
  wire _08034_;
  wire _08035_;
  wire _08036_;
  wire _08037_;
  wire _08038_;
  wire _08039_;
  wire _08040_;
  wire _08041_;
  wire _08042_;
  wire _08043_;
  wire _08044_;
  wire _08045_;
  wire _08046_;
  wire _08047_;
  wire _08048_;
  wire _08049_;
  wire _08050_;
  wire _08051_;
  wire _08052_;
  wire _08053_;
  wire _08054_;
  wire _08055_;
  wire _08056_;
  wire _08057_;
  wire _08058_;
  wire _08059_;
  wire _08060_;
  wire _08061_;
  wire _08062_;
  wire _08063_;
  wire _08064_;
  wire _08065_;
  wire _08066_;
  wire _08067_;
  wire _08068_;
  wire _08069_;
  wire _08070_;
  wire _08071_;
  wire _08072_;
  wire _08073_;
  wire _08074_;
  wire _08075_;
  wire _08076_;
  wire _08077_;
  wire _08078_;
  wire _08079_;
  wire _08080_;
  wire _08081_;
  wire _08082_;
  wire _08083_;
  wire _08084_;
  wire _08085_;
  wire _08086_;
  wire _08087_;
  wire _08088_;
  wire _08089_;
  wire _08090_;
  wire _08091_;
  wire _08092_;
  wire _08093_;
  wire _08094_;
  wire _08095_;
  wire _08096_;
  wire _08097_;
  wire _08098_;
  wire _08099_;
  wire _08100_;
  wire _08101_;
  wire _08102_;
  wire _08103_;
  wire _08104_;
  wire _08105_;
  wire _08106_;
  wire _08107_;
  wire _08108_;
  wire _08109_;
  wire _08110_;
  wire _08111_;
  wire _08112_;
  wire _08113_;
  wire _08114_;
  wire _08115_;
  wire _08116_;
  wire _08117_;
  wire _08118_;
  wire _08119_;
  wire _08120_;
  wire _08121_;
  wire _08122_;
  wire _08123_;
  wire _08124_;
  wire _08125_;
  wire _08126_;
  wire _08127_;
  wire _08128_;
  wire _08129_;
  wire _08130_;
  wire _08131_;
  wire _08132_;
  wire _08133_;
  wire _08134_;
  wire _08135_;
  wire _08136_;
  wire _08137_;
  wire _08138_;
  wire _08139_;
  wire _08140_;
  wire _08141_;
  wire _08142_;
  wire _08143_;
  wire _08144_;
  wire _08145_;
  wire _08146_;
  wire _08147_;
  wire _08148_;
  wire _08149_;
  wire _08150_;
  wire _08151_;
  wire _08152_;
  wire _08153_;
  wire _08154_;
  wire _08155_;
  wire _08156_;
  wire _08157_;
  wire _08158_;
  wire _08159_;
  wire _08160_;
  wire _08161_;
  wire _08162_;
  wire _08163_;
  wire _08164_;
  wire _08165_;
  wire _08166_;
  wire _08167_;
  wire _08168_;
  wire _08169_;
  wire _08170_;
  wire _08171_;
  wire _08172_;
  wire _08173_;
  wire _08174_;
  wire _08175_;
  wire _08176_;
  wire _08177_;
  wire _08178_;
  wire _08179_;
  wire _08180_;
  wire _08181_;
  wire _08182_;
  wire _08183_;
  wire _08184_;
  wire _08185_;
  wire _08186_;
  wire _08187_;
  wire _08188_;
  wire _08189_;
  wire _08190_;
  wire _08191_;
  wire _08192_;
  wire _08193_;
  wire _08194_;
  wire _08195_;
  wire _08196_;
  wire _08197_;
  wire _08198_;
  wire _08199_;
  wire _08200_;
  wire _08201_;
  wire _08202_;
  wire _08203_;
  wire _08204_;
  wire _08205_;
  wire _08206_;
  wire _08207_;
  wire _08208_;
  wire _08209_;
  wire _08210_;
  wire _08211_;
  wire _08212_;
  wire _08213_;
  wire _08214_;
  wire _08215_;
  wire _08216_;
  wire _08217_;
  wire _08218_;
  wire _08219_;
  wire _08220_;
  wire _08221_;
  wire _08222_;
  wire _08223_;
  wire _08224_;
  wire _08225_;
  wire _08226_;
  wire _08227_;
  wire _08228_;
  wire _08229_;
  wire _08230_;
  wire _08231_;
  wire _08232_;
  wire _08233_;
  wire _08234_;
  wire _08235_;
  wire _08236_;
  wire _08237_;
  wire _08238_;
  wire _08239_;
  wire _08240_;
  wire _08241_;
  wire _08242_;
  wire _08243_;
  wire _08244_;
  wire _08245_;
  wire _08246_;
  wire _08247_;
  wire _08248_;
  wire _08249_;
  wire _08250_;
  wire _08251_;
  wire _08252_;
  wire _08253_;
  wire _08254_;
  wire _08255_;
  wire _08256_;
  wire _08257_;
  wire _08258_;
  wire _08259_;
  wire _08260_;
  wire _08261_;
  wire _08262_;
  wire _08263_;
  wire _08264_;
  wire _08265_;
  wire _08266_;
  wire _08267_;
  wire _08268_;
  wire _08269_;
  wire _08270_;
  wire _08271_;
  wire _08272_;
  wire _08273_;
  wire _08274_;
  wire _08275_;
  wire _08276_;
  wire _08277_;
  wire _08278_;
  wire _08279_;
  wire _08280_;
  wire _08281_;
  wire _08282_;
  wire _08283_;
  wire _08284_;
  wire _08285_;
  wire _08286_;
  wire _08287_;
  wire _08288_;
  wire _08289_;
  wire _08290_;
  wire _08291_;
  wire _08292_;
  wire _08293_;
  wire _08294_;
  wire _08295_;
  wire _08296_;
  wire _08297_;
  wire _08298_;
  wire _08299_;
  wire _08300_;
  wire _08301_;
  wire _08302_;
  wire _08303_;
  wire _08304_;
  wire _08305_;
  wire _08306_;
  wire _08307_;
  wire _08308_;
  wire _08309_;
  wire _08310_;
  wire _08311_;
  wire _08312_;
  wire _08313_;
  wire _08314_;
  wire _08315_;
  wire _08316_;
  wire _08317_;
  wire _08318_;
  wire _08319_;
  wire _08320_;
  wire _08321_;
  wire _08322_;
  wire _08323_;
  wire _08324_;
  wire _08325_;
  wire _08326_;
  wire _08327_;
  wire _08328_;
  wire _08329_;
  wire _08330_;
  wire _08331_;
  wire _08332_;
  wire _08333_;
  wire _08334_;
  wire _08335_;
  wire _08336_;
  wire _08337_;
  wire _08338_;
  wire _08339_;
  wire _08340_;
  wire _08341_;
  wire _08342_;
  wire _08343_;
  wire _08344_;
  wire _08345_;
  wire _08346_;
  wire _08347_;
  wire _08348_;
  wire _08349_;
  wire _08350_;
  wire _08351_;
  wire _08352_;
  wire _08353_;
  wire _08354_;
  wire _08355_;
  wire _08356_;
  wire _08357_;
  wire _08358_;
  wire _08359_;
  wire _08360_;
  wire _08361_;
  wire _08362_;
  wire _08363_;
  wire _08364_;
  wire _08365_;
  wire _08366_;
  wire _08367_;
  wire _08368_;
  wire _08369_;
  wire _08370_;
  wire _08371_;
  wire _08372_;
  wire _08373_;
  wire _08374_;
  wire _08375_;
  wire _08376_;
  wire _08377_;
  wire _08378_;
  wire _08379_;
  wire _08380_;
  wire _08381_;
  wire _08382_;
  wire _08383_;
  wire _08384_;
  wire _08385_;
  wire _08386_;
  wire _08387_;
  wire _08388_;
  wire _08389_;
  wire _08390_;
  wire _08391_;
  wire _08392_;
  wire _08393_;
  wire _08394_;
  wire _08395_;
  wire _08396_;
  wire _08397_;
  wire _08398_;
  wire _08399_;
  wire _08400_;
  wire _08401_;
  wire _08402_;
  wire _08403_;
  wire _08404_;
  wire _08405_;
  wire _08406_;
  wire _08407_;
  wire _08408_;
  wire _08409_;
  wire _08410_;
  wire _08411_;
  wire _08412_;
  wire _08413_;
  wire _08414_;
  wire _08415_;
  wire _08416_;
  wire _08417_;
  wire _08418_;
  wire _08419_;
  wire _08420_;
  wire _08421_;
  wire _08422_;
  wire _08423_;
  wire _08424_;
  wire _08425_;
  wire _08426_;
  wire _08427_;
  wire _08428_;
  wire _08429_;
  wire _08430_;
  wire _08431_;
  wire _08432_;
  wire _08433_;
  wire _08434_;
  wire _08435_;
  wire _08436_;
  wire _08437_;
  wire _08438_;
  wire _08439_;
  wire _08440_;
  wire _08441_;
  wire _08442_;
  wire _08443_;
  wire _08444_;
  wire _08445_;
  wire _08446_;
  wire _08447_;
  wire _08448_;
  wire _08449_;
  wire _08450_;
  wire _08451_;
  wire _08452_;
  wire _08453_;
  wire _08454_;
  wire _08455_;
  wire _08456_;
  wire _08457_;
  wire _08458_;
  wire _08459_;
  wire _08460_;
  wire _08461_;
  wire _08462_;
  wire _08463_;
  wire _08464_;
  wire _08465_;
  wire _08466_;
  wire _08467_;
  wire _08468_;
  wire _08469_;
  wire _08470_;
  wire _08471_;
  wire _08472_;
  wire _08473_;
  wire _08474_;
  wire _08475_;
  wire _08476_;
  wire _08477_;
  wire _08478_;
  wire _08479_;
  wire _08480_;
  wire _08481_;
  wire _08482_;
  wire _08483_;
  wire _08484_;
  wire _08485_;
  wire _08486_;
  wire _08487_;
  wire _08488_;
  wire _08489_;
  wire _08490_;
  wire _08491_;
  wire _08492_;
  wire _08493_;
  wire _08494_;
  wire _08495_;
  wire _08496_;
  wire _08497_;
  wire _08498_;
  wire _08499_;
  wire _08500_;
  wire _08501_;
  wire _08502_;
  wire _08503_;
  wire _08504_;
  wire _08505_;
  wire _08506_;
  wire _08507_;
  wire _08508_;
  wire _08509_;
  wire _08510_;
  wire _08511_;
  wire _08512_;
  wire _08513_;
  wire _08514_;
  wire _08515_;
  wire _08516_;
  wire _08517_;
  wire _08518_;
  wire _08519_;
  wire _08520_;
  wire _08521_;
  wire _08522_;
  wire _08523_;
  wire _08524_;
  wire _08525_;
  wire _08526_;
  wire _08527_;
  wire _08528_;
  wire _08529_;
  wire _08530_;
  wire _08531_;
  wire _08532_;
  wire _08533_;
  wire _08534_;
  wire _08535_;
  wire _08536_;
  wire _08537_;
  wire _08538_;
  wire _08539_;
  wire _08540_;
  wire _08541_;
  wire _08542_;
  wire _08543_;
  wire _08544_;
  wire _08545_;
  wire _08546_;
  wire _08547_;
  wire _08548_;
  wire _08549_;
  wire _08550_;
  wire _08551_;
  wire _08552_;
  wire _08553_;
  wire _08554_;
  wire _08555_;
  wire _08556_;
  wire _08557_;
  wire _08558_;
  wire _08559_;
  wire _08560_;
  wire _08561_;
  wire _08562_;
  wire _08563_;
  wire _08564_;
  wire _08565_;
  wire _08566_;
  wire _08567_;
  wire _08568_;
  wire _08569_;
  wire _08570_;
  wire _08571_;
  wire _08572_;
  wire _08573_;
  wire _08574_;
  wire _08575_;
  wire _08576_;
  wire _08577_;
  wire _08578_;
  wire _08579_;
  wire _08580_;
  wire _08581_;
  wire _08582_;
  wire _08583_;
  wire _08584_;
  wire _08585_;
  wire _08586_;
  wire _08587_;
  wire _08588_;
  wire _08589_;
  wire _08590_;
  wire _08591_;
  wire _08592_;
  wire _08593_;
  wire _08594_;
  wire _08595_;
  wire _08596_;
  wire _08597_;
  wire _08598_;
  wire _08599_;
  wire _08600_;
  wire _08601_;
  wire _08602_;
  wire _08603_;
  wire _08604_;
  wire _08605_;
  wire _08606_;
  wire _08607_;
  wire _08608_;
  wire _08609_;
  wire _08610_;
  wire _08611_;
  wire _08612_;
  wire _08613_;
  wire _08614_;
  wire _08615_;
  wire _08616_;
  wire _08617_;
  wire _08618_;
  wire _08619_;
  wire _08620_;
  wire _08621_;
  wire _08622_;
  wire _08623_;
  wire _08624_;
  wire _08625_;
  wire _08626_;
  wire _08627_;
  wire _08628_;
  wire _08629_;
  wire _08630_;
  wire _08631_;
  wire _08632_;
  wire _08633_;
  wire _08634_;
  wire _08635_;
  wire _08636_;
  wire _08637_;
  wire _08638_;
  wire _08639_;
  wire _08640_;
  wire _08641_;
  wire _08642_;
  wire _08643_;
  wire _08644_;
  wire _08645_;
  wire _08646_;
  wire _08647_;
  wire _08648_;
  wire _08649_;
  wire _08650_;
  wire _08651_;
  wire _08652_;
  wire _08653_;
  wire _08654_;
  wire _08655_;
  wire _08656_;
  wire _08657_;
  wire _08658_;
  wire _08659_;
  wire _08660_;
  wire _08661_;
  wire _08662_;
  wire _08663_;
  wire _08664_;
  wire _08665_;
  wire _08666_;
  wire _08667_;
  wire _08668_;
  wire _08669_;
  wire _08670_;
  wire _08671_;
  wire _08672_;
  wire _08673_;
  wire _08674_;
  wire _08675_;
  wire _08676_;
  wire _08677_;
  wire _08678_;
  wire _08679_;
  wire _08680_;
  wire _08681_;
  wire _08682_;
  wire _08683_;
  wire _08684_;
  wire _08685_;
  wire _08686_;
  wire _08687_;
  wire _08688_;
  wire _08689_;
  wire _08690_;
  wire _08691_;
  wire _08692_;
  wire _08693_;
  wire _08694_;
  wire _08695_;
  wire _08696_;
  wire _08697_;
  wire _08698_;
  wire _08699_;
  wire _08700_;
  wire _08701_;
  wire _08702_;
  wire _08703_;
  wire _08704_;
  wire _08705_;
  wire _08706_;
  wire _08707_;
  wire _08708_;
  wire _08709_;
  wire _08710_;
  wire _08711_;
  wire _08712_;
  wire _08713_;
  wire _08714_;
  wire _08715_;
  wire _08716_;
  wire _08717_;
  wire _08718_;
  wire _08719_;
  wire _08720_;
  wire _08721_;
  wire _08722_;
  wire _08723_;
  wire _08724_;
  wire _08725_;
  wire _08726_;
  wire _08727_;
  wire _08728_;
  wire _08729_;
  wire _08730_;
  wire _08731_;
  wire _08732_;
  wire _08733_;
  wire _08734_;
  wire _08735_;
  wire _08736_;
  wire _08737_;
  wire _08738_;
  wire _08739_;
  wire _08740_;
  wire _08741_;
  wire _08742_;
  wire _08743_;
  wire _08744_;
  wire _08745_;
  wire _08746_;
  wire _08747_;
  wire _08748_;
  wire _08749_;
  wire _08750_;
  wire _08751_;
  wire _08752_;
  wire _08753_;
  wire _08754_;
  wire _08755_;
  wire _08756_;
  wire _08757_;
  wire _08758_;
  wire _08759_;
  wire _08760_;
  wire _08761_;
  wire _08762_;
  wire _08763_;
  wire _08764_;
  wire _08765_;
  wire _08766_;
  wire _08767_;
  wire _08768_;
  wire _08769_;
  wire _08770_;
  wire _08771_;
  wire _08772_;
  wire _08773_;
  wire _08774_;
  wire _08775_;
  wire _08776_;
  wire _08777_;
  wire _08778_;
  wire _08779_;
  wire _08780_;
  wire _08781_;
  wire _08782_;
  wire _08783_;
  wire _08784_;
  wire _08785_;
  wire _08786_;
  wire _08787_;
  wire _08788_;
  wire _08789_;
  wire _08790_;
  wire _08791_;
  wire _08792_;
  wire _08793_;
  wire _08794_;
  wire _08795_;
  wire _08796_;
  wire _08797_;
  wire _08798_;
  wire _08799_;
  wire _08800_;
  wire _08801_;
  wire _08802_;
  wire _08803_;
  wire _08804_;
  wire _08805_;
  wire _08806_;
  wire _08807_;
  wire _08808_;
  wire _08809_;
  wire _08810_;
  wire _08811_;
  wire _08812_;
  wire _08813_;
  wire _08814_;
  wire _08815_;
  wire _08816_;
  wire _08817_;
  wire _08818_;
  wire _08819_;
  wire _08820_;
  wire _08821_;
  wire _08822_;
  wire _08823_;
  wire _08824_;
  wire _08825_;
  wire _08826_;
  wire _08827_;
  wire _08828_;
  wire _08829_;
  wire _08830_;
  wire _08831_;
  wire _08832_;
  wire _08833_;
  wire _08834_;
  wire _08835_;
  wire _08836_;
  wire _08837_;
  wire _08838_;
  wire _08839_;
  wire _08840_;
  wire _08841_;
  wire _08842_;
  wire _08843_;
  wire _08844_;
  wire _08845_;
  wire _08846_;
  wire _08847_;
  wire _08848_;
  wire _08849_;
  wire _08850_;
  wire _08851_;
  wire _08852_;
  wire _08853_;
  wire _08854_;
  wire _08855_;
  wire _08856_;
  wire _08857_;
  wire _08858_;
  wire _08859_;
  wire _08860_;
  wire _08861_;
  wire _08862_;
  wire _08863_;
  wire _08864_;
  wire _08865_;
  wire _08866_;
  wire _08867_;
  wire _08868_;
  wire _08869_;
  wire _08870_;
  wire _08871_;
  wire _08872_;
  wire _08873_;
  wire _08874_;
  wire _08875_;
  wire _08876_;
  wire _08877_;
  wire _08878_;
  wire _08879_;
  wire _08880_;
  wire _08881_;
  wire _08882_;
  wire _08883_;
  wire _08884_;
  wire _08885_;
  wire _08886_;
  wire _08887_;
  wire _08888_;
  wire _08889_;
  wire _08890_;
  wire _08891_;
  wire _08892_;
  wire _08893_;
  wire _08894_;
  wire _08895_;
  wire _08896_;
  wire _08897_;
  wire _08898_;
  wire _08899_;
  wire _08900_;
  wire _08901_;
  wire _08902_;
  wire _08903_;
  wire _08904_;
  wire _08905_;
  wire _08906_;
  wire _08907_;
  wire _08908_;
  wire _08909_;
  wire _08910_;
  wire _08911_;
  wire _08912_;
  wire _08913_;
  wire _08914_;
  wire _08915_;
  wire _08916_;
  wire _08917_;
  wire _08918_;
  wire _08919_;
  wire _08920_;
  wire _08921_;
  wire _08922_;
  wire _08923_;
  wire _08924_;
  wire _08925_;
  wire _08926_;
  wire _08927_;
  wire _08928_;
  wire _08929_;
  wire _08930_;
  wire _08931_;
  wire _08932_;
  wire _08933_;
  wire _08934_;
  wire _08935_;
  wire _08936_;
  wire _08937_;
  wire _08938_;
  wire _08939_;
  wire _08940_;
  wire _08941_;
  wire _08942_;
  wire _08943_;
  wire _08944_;
  wire _08945_;
  wire _08946_;
  wire _08947_;
  wire _08948_;
  wire _08949_;
  wire _08950_;
  wire _08951_;
  wire _08952_;
  wire _08953_;
  wire _08954_;
  wire _08955_;
  wire _08956_;
  wire _08957_;
  wire _08958_;
  wire _08959_;
  wire _08960_;
  wire _08961_;
  wire _08962_;
  wire _08963_;
  wire _08964_;
  wire _08965_;
  wire _08966_;
  wire _08967_;
  wire _08968_;
  wire _08969_;
  wire _08970_;
  wire _08971_;
  wire _08972_;
  wire _08973_;
  wire _08974_;
  wire _08975_;
  wire _08976_;
  wire _08977_;
  wire _08978_;
  wire _08979_;
  wire _08980_;
  wire _08981_;
  wire _08982_;
  wire _08983_;
  wire _08984_;
  wire _08985_;
  wire _08986_;
  wire _08987_;
  wire _08988_;
  wire _08989_;
  wire _08990_;
  wire _08991_;
  wire _08992_;
  wire _08993_;
  wire _08994_;
  wire _08995_;
  wire _08996_;
  wire _08997_;
  wire _08998_;
  wire _08999_;
  wire _09000_;
  wire _09001_;
  wire _09002_;
  wire _09003_;
  wire _09004_;
  wire _09005_;
  wire _09006_;
  wire _09007_;
  wire _09008_;
  wire _09009_;
  wire _09010_;
  wire _09011_;
  wire _09012_;
  wire _09013_;
  wire _09014_;
  wire _09015_;
  wire _09016_;
  wire _09017_;
  wire _09018_;
  wire _09019_;
  wire _09020_;
  wire _09021_;
  wire _09022_;
  wire _09023_;
  wire _09024_;
  wire _09025_;
  wire _09026_;
  wire _09027_;
  wire _09028_;
  wire _09029_;
  wire _09030_;
  wire _09031_;
  wire _09032_;
  wire _09033_;
  wire _09034_;
  wire _09035_;
  wire _09036_;
  wire _09037_;
  wire _09038_;
  wire _09039_;
  wire _09040_;
  wire _09041_;
  wire _09042_;
  wire _09043_;
  wire _09044_;
  wire _09045_;
  wire _09046_;
  wire _09047_;
  wire _09048_;
  wire _09049_;
  wire _09050_;
  wire _09051_;
  wire _09052_;
  wire _09053_;
  wire _09054_;
  wire _09055_;
  wire _09056_;
  wire _09057_;
  wire _09058_;
  wire _09059_;
  wire _09060_;
  wire _09061_;
  wire _09062_;
  wire _09063_;
  wire _09064_;
  wire _09065_;
  wire _09066_;
  wire _09067_;
  wire _09068_;
  wire _09069_;
  wire _09070_;
  wire _09071_;
  wire _09072_;
  wire _09073_;
  wire _09074_;
  wire _09075_;
  wire _09076_;
  wire _09077_;
  wire _09078_;
  wire _09079_;
  wire _09080_;
  wire _09081_;
  wire _09082_;
  wire _09083_;
  wire _09084_;
  wire _09085_;
  wire _09086_;
  wire _09087_;
  wire _09088_;
  wire _09089_;
  wire _09090_;
  wire _09091_;
  wire _09092_;
  wire _09093_;
  wire _09094_;
  wire _09095_;
  wire _09096_;
  wire _09097_;
  wire _09098_;
  wire _09099_;
  wire _09100_;
  wire _09101_;
  wire _09102_;
  wire _09103_;
  wire _09104_;
  wire _09105_;
  wire _09106_;
  wire _09107_;
  wire _09108_;
  wire _09109_;
  wire _09110_;
  wire _09111_;
  wire _09112_;
  wire _09113_;
  wire _09114_;
  wire _09115_;
  wire _09116_;
  wire _09117_;
  wire _09118_;
  wire _09119_;
  wire _09120_;
  wire _09121_;
  wire _09122_;
  wire _09123_;
  wire _09124_;
  wire _09125_;
  wire _09126_;
  wire _09127_;
  wire _09128_;
  wire _09129_;
  wire _09130_;
  wire _09131_;
  wire _09132_;
  wire _09133_;
  wire _09134_;
  wire _09135_;
  wire _09136_;
  wire _09137_;
  wire _09138_;
  wire _09139_;
  wire _09140_;
  wire _09141_;
  wire _09142_;
  wire _09143_;
  wire _09144_;
  wire _09145_;
  wire _09146_;
  wire _09147_;
  wire _09148_;
  wire _09149_;
  wire _09150_;
  wire _09151_;
  wire _09152_;
  wire _09153_;
  wire _09154_;
  wire _09155_;
  wire _09156_;
  wire _09157_;
  wire _09158_;
  wire _09159_;
  wire _09160_;
  wire _09161_;
  wire _09162_;
  wire _09163_;
  wire _09164_;
  wire _09165_;
  wire _09166_;
  wire _09167_;
  wire _09168_;
  wire _09169_;
  wire _09170_;
  wire _09171_;
  wire _09172_;
  wire _09173_;
  wire _09174_;
  wire _09175_;
  wire _09176_;
  wire _09177_;
  wire _09178_;
  wire _09179_;
  wire _09180_;
  wire _09181_;
  wire _09182_;
  wire _09183_;
  wire _09184_;
  wire _09185_;
  wire _09186_;
  wire _09187_;
  wire _09188_;
  wire _09189_;
  wire _09190_;
  wire _09191_;
  wire _09192_;
  wire _09193_;
  wire _09194_;
  wire _09195_;
  wire _09196_;
  wire _09197_;
  wire _09198_;
  wire _09199_;
  wire _09200_;
  wire _09201_;
  wire _09202_;
  wire _09203_;
  wire _09204_;
  wire _09205_;
  wire _09206_;
  wire _09207_;
  wire _09208_;
  wire _09209_;
  wire _09210_;
  wire _09211_;
  wire _09212_;
  wire _09213_;
  wire _09214_;
  wire _09215_;
  wire _09216_;
  wire _09217_;
  wire _09218_;
  wire _09219_;
  wire _09220_;
  wire _09221_;
  wire _09222_;
  wire _09223_;
  wire _09224_;
  wire _09225_;
  wire _09226_;
  wire _09227_;
  wire _09228_;
  wire _09229_;
  wire _09230_;
  wire _09231_;
  wire _09232_;
  wire _09233_;
  wire _09234_;
  wire _09235_;
  wire _09236_;
  wire _09237_;
  wire _09238_;
  wire _09239_;
  wire _09240_;
  wire _09241_;
  wire _09242_;
  wire _09243_;
  wire _09244_;
  wire _09245_;
  wire _09246_;
  wire _09247_;
  wire _09248_;
  wire _09249_;
  wire _09250_;
  wire _09251_;
  wire _09252_;
  wire _09253_;
  wire _09254_;
  wire _09255_;
  wire _09256_;
  wire _09257_;
  wire _09258_;
  wire _09259_;
  wire _09260_;
  wire _09261_;
  wire _09262_;
  wire _09263_;
  wire _09264_;
  wire _09265_;
  wire _09266_;
  wire _09267_;
  wire _09268_;
  wire _09269_;
  wire _09270_;
  wire _09271_;
  wire _09272_;
  wire _09273_;
  wire _09274_;
  wire _09275_;
  wire _09276_;
  wire _09277_;
  wire _09278_;
  wire _09279_;
  wire _09280_;
  wire _09281_;
  wire _09282_;
  wire _09283_;
  wire _09284_;
  wire _09285_;
  wire _09286_;
  wire _09287_;
  wire _09288_;
  wire _09289_;
  wire _09290_;
  wire _09291_;
  wire _09292_;
  wire _09293_;
  wire _09294_;
  wire _09295_;
  wire _09296_;
  wire _09297_;
  wire _09298_;
  wire _09299_;
  wire _09300_;
  wire _09301_;
  wire _09302_;
  wire _09303_;
  wire _09304_;
  wire _09305_;
  wire _09306_;
  wire _09307_;
  wire _09308_;
  wire _09309_;
  wire _09310_;
  wire _09311_;
  wire _09312_;
  wire _09313_;
  wire _09314_;
  wire _09315_;
  wire _09316_;
  wire _09317_;
  wire _09318_;
  wire _09319_;
  wire _09320_;
  wire _09321_;
  wire _09322_;
  wire _09323_;
  wire _09324_;
  wire _09325_;
  wire _09326_;
  wire _09327_;
  wire _09328_;
  wire _09329_;
  wire _09330_;
  wire _09331_;
  wire _09332_;
  wire _09333_;
  wire _09334_;
  wire _09335_;
  wire _09336_;
  wire _09337_;
  wire _09338_;
  wire _09339_;
  wire _09340_;
  wire _09341_;
  wire _09342_;
  wire _09343_;
  wire _09344_;
  wire _09345_;
  wire _09346_;
  wire _09347_;
  wire _09348_;
  wire _09349_;
  wire _09350_;
  wire _09351_;
  wire _09352_;
  wire _09353_;
  wire _09354_;
  wire _09355_;
  wire _09356_;
  wire _09357_;
  wire _09358_;
  wire _09359_;
  wire _09360_;
  wire _09361_;
  wire _09362_;
  wire _09363_;
  wire _09364_;
  wire _09365_;
  wire _09366_;
  wire _09367_;
  wire _09368_;
  wire _09369_;
  wire _09370_;
  wire _09371_;
  wire _09372_;
  wire _09373_;
  wire _09374_;
  wire _09375_;
  wire _09376_;
  wire _09377_;
  wire _09378_;
  wire _09379_;
  wire _09380_;
  wire _09381_;
  wire _09382_;
  wire _09383_;
  wire _09384_;
  wire _09385_;
  wire _09386_;
  wire _09387_;
  wire _09388_;
  wire _09389_;
  wire _09390_;
  wire _09391_;
  wire _09392_;
  wire _09393_;
  wire _09394_;
  wire _09395_;
  wire _09396_;
  wire _09397_;
  wire _09398_;
  wire _09399_;
  wire _09400_;
  wire _09401_;
  wire _09402_;
  wire _09403_;
  wire _09404_;
  wire _09405_;
  wire _09406_;
  wire _09407_;
  wire _09408_;
  wire _09409_;
  wire _09410_;
  wire _09411_;
  wire _09412_;
  wire _09413_;
  wire _09414_;
  wire _09415_;
  wire _09416_;
  wire _09417_;
  wire _09418_;
  wire _09419_;
  wire _09420_;
  wire _09421_;
  wire _09422_;
  wire _09423_;
  wire _09424_;
  wire _09425_;
  wire _09426_;
  wire _09427_;
  wire _09428_;
  wire _09429_;
  wire _09430_;
  wire _09431_;
  wire _09432_;
  wire _09433_;
  wire _09434_;
  wire _09435_;
  wire _09436_;
  wire _09437_;
  wire _09438_;
  wire _09439_;
  wire _09440_;
  wire _09441_;
  wire _09442_;
  wire _09443_;
  wire _09444_;
  wire _09445_;
  wire _09446_;
  wire _09447_;
  wire _09448_;
  wire _09449_;
  wire _09450_;
  wire _09451_;
  wire _09452_;
  wire _09453_;
  wire _09454_;
  wire _09455_;
  wire _09456_;
  wire _09457_;
  wire _09458_;
  wire _09459_;
  wire _09460_;
  wire _09461_;
  wire _09462_;
  wire _09463_;
  wire _09464_;
  wire _09465_;
  wire _09466_;
  wire _09467_;
  wire _09468_;
  wire _09469_;
  wire _09470_;
  wire _09471_;
  wire _09472_;
  wire _09473_;
  wire _09474_;
  wire _09475_;
  wire _09476_;
  wire _09477_;
  wire _09478_;
  wire _09479_;
  wire _09480_;
  wire _09481_;
  wire _09482_;
  wire _09483_;
  wire _09484_;
  wire _09485_;
  wire _09486_;
  wire _09487_;
  wire _09488_;
  wire _09489_;
  wire _09490_;
  wire _09491_;
  wire _09492_;
  wire _09493_;
  wire _09494_;
  wire _09495_;
  wire _09496_;
  wire _09497_;
  wire _09498_;
  wire _09499_;
  wire _09500_;
  wire _09501_;
  wire _09502_;
  wire _09503_;
  wire _09504_;
  wire _09505_;
  wire _09506_;
  wire _09507_;
  wire _09508_;
  wire _09509_;
  wire _09510_;
  wire _09511_;
  wire _09512_;
  wire _09513_;
  wire _09514_;
  wire _09515_;
  wire _09516_;
  wire _09517_;
  wire _09518_;
  wire _09519_;
  wire _09520_;
  wire _09521_;
  wire _09522_;
  wire _09523_;
  wire _09524_;
  wire _09525_;
  wire _09526_;
  wire _09527_;
  wire _09528_;
  wire _09529_;
  wire _09530_;
  wire _09531_;
  wire _09532_;
  wire _09533_;
  wire _09534_;
  wire _09535_;
  wire _09536_;
  wire _09537_;
  wire _09538_;
  wire _09539_;
  wire _09540_;
  wire _09541_;
  wire _09542_;
  wire _09543_;
  wire _09544_;
  wire _09545_;
  wire _09546_;
  wire _09547_;
  wire _09548_;
  wire _09549_;
  wire _09550_;
  wire _09551_;
  wire _09552_;
  wire _09553_;
  wire _09554_;
  wire _09555_;
  wire _09556_;
  wire _09557_;
  wire _09558_;
  wire _09559_;
  wire _09560_;
  wire _09561_;
  wire _09562_;
  wire _09563_;
  wire _09564_;
  wire _09565_;
  wire _09566_;
  wire _09567_;
  wire _09568_;
  wire _09569_;
  wire _09570_;
  wire _09571_;
  wire _09572_;
  wire _09573_;
  wire _09574_;
  wire _09575_;
  wire _09576_;
  wire _09577_;
  wire _09578_;
  wire _09579_;
  wire _09580_;
  wire _09581_;
  wire _09582_;
  wire _09583_;
  wire _09584_;
  wire _09585_;
  wire _09586_;
  wire _09587_;
  wire _09588_;
  wire _09589_;
  wire _09590_;
  wire _09591_;
  wire _09592_;
  wire _09593_;
  wire _09594_;
  wire _09595_;
  wire _09596_;
  wire _09597_;
  wire _09598_;
  wire _09599_;
  wire _09600_;
  wire _09601_;
  wire _09602_;
  wire _09603_;
  wire _09604_;
  wire _09605_;
  wire _09606_;
  wire _09607_;
  wire _09608_;
  wire _09609_;
  wire _09610_;
  wire _09611_;
  wire _09612_;
  wire _09613_;
  wire _09614_;
  wire _09615_;
  wire _09616_;
  wire _09617_;
  wire _09618_;
  wire _09619_;
  wire _09620_;
  wire _09621_;
  wire _09622_;
  wire _09623_;
  wire _09624_;
  wire _09625_;
  wire _09626_;
  wire _09627_;
  wire _09628_;
  wire _09629_;
  wire _09630_;
  wire _09631_;
  wire _09632_;
  wire _09633_;
  wire _09634_;
  wire _09635_;
  wire _09636_;
  wire _09637_;
  wire _09638_;
  wire _09639_;
  wire _09640_;
  wire _09641_;
  wire _09642_;
  wire _09643_;
  wire _09644_;
  wire _09645_;
  wire _09646_;
  wire _09647_;
  wire _09648_;
  wire _09649_;
  wire _09650_;
  wire _09651_;
  wire _09652_;
  wire _09653_;
  wire _09654_;
  wire _09655_;
  wire _09656_;
  wire _09657_;
  wire _09658_;
  wire _09659_;
  wire _09660_;
  wire _09661_;
  wire _09662_;
  wire _09663_;
  wire _09664_;
  wire _09665_;
  wire _09666_;
  wire _09667_;
  wire _09668_;
  wire _09669_;
  wire _09670_;
  wire _09671_;
  wire _09672_;
  wire _09673_;
  wire _09674_;
  wire _09675_;
  wire _09676_;
  wire _09677_;
  wire _09678_;
  wire _09679_;
  wire _09680_;
  wire _09681_;
  wire _09682_;
  wire _09683_;
  wire _09684_;
  wire _09685_;
  wire _09686_;
  wire _09687_;
  wire _09688_;
  wire _09689_;
  wire _09690_;
  wire _09691_;
  wire _09692_;
  wire _09693_;
  wire _09694_;
  wire _09695_;
  wire _09696_;
  wire _09697_;
  wire _09698_;
  wire _09699_;
  wire _09700_;
  wire _09701_;
  wire _09702_;
  wire _09703_;
  wire _09704_;
  wire _09705_;
  wire _09706_;
  wire _09707_;
  wire _09708_;
  wire _09709_;
  wire _09710_;
  wire _09711_;
  wire _09712_;
  wire _09713_;
  wire _09714_;
  wire _09715_;
  wire _09716_;
  wire _09717_;
  wire _09718_;
  wire _09719_;
  wire _09720_;
  wire _09721_;
  wire _09722_;
  wire _09723_;
  wire _09724_;
  wire _09725_;
  wire _09726_;
  wire _09727_;
  wire _09728_;
  wire _09729_;
  wire _09730_;
  wire _09731_;
  wire _09732_;
  wire _09733_;
  wire _09734_;
  wire _09735_;
  wire _09736_;
  wire _09737_;
  wire _09738_;
  wire _09739_;
  wire _09740_;
  wire _09741_;
  wire _09742_;
  wire _09743_;
  wire _09744_;
  wire _09745_;
  wire _09746_;
  wire _09747_;
  wire _09748_;
  wire _09749_;
  wire _09750_;
  wire _09751_;
  wire _09752_;
  wire _09753_;
  wire _09754_;
  wire _09755_;
  wire _09756_;
  wire _09757_;
  wire _09758_;
  wire _09759_;
  wire _09760_;
  wire _09761_;
  wire _09762_;
  wire _09763_;
  wire _09764_;
  wire _09765_;
  wire _09766_;
  wire _09767_;
  wire _09768_;
  wire _09769_;
  wire _09770_;
  wire _09771_;
  wire _09772_;
  wire _09773_;
  wire _09774_;
  wire _09775_;
  wire _09776_;
  wire _09777_;
  wire _09778_;
  wire _09779_;
  wire _09780_;
  wire _09781_;
  wire _09782_;
  wire _09783_;
  wire _09784_;
  wire _09785_;
  wire _09786_;
  wire _09787_;
  wire _09788_;
  wire _09789_;
  wire _09790_;
  wire _09791_;
  wire _09792_;
  wire _09793_;
  wire _09794_;
  wire _09795_;
  wire _09796_;
  wire _09797_;
  wire _09798_;
  wire _09799_;
  wire _09800_;
  wire _09801_;
  wire _09802_;
  wire _09803_;
  wire _09804_;
  wire _09805_;
  wire _09806_;
  wire _09807_;
  wire _09808_;
  wire _09809_;
  wire _09810_;
  wire _09811_;
  wire _09812_;
  wire _09813_;
  wire _09814_;
  wire _09815_;
  wire _09816_;
  wire _09817_;
  wire _09818_;
  wire _09819_;
  wire _09820_;
  wire _09821_;
  wire _09822_;
  wire _09823_;
  wire _09824_;
  wire _09825_;
  wire _09826_;
  wire _09827_;
  wire _09828_;
  wire _09829_;
  wire _09830_;
  wire _09831_;
  wire _09832_;
  wire _09833_;
  wire _09834_;
  wire _09835_;
  wire _09836_;
  wire _09837_;
  wire _09838_;
  wire _09839_;
  wire _09840_;
  wire _09841_;
  wire _09842_;
  wire _09843_;
  wire _09844_;
  wire _09845_;
  wire _09846_;
  wire _09847_;
  wire _09848_;
  wire _09849_;
  wire _09850_;
  wire _09851_;
  wire _09852_;
  wire _09853_;
  wire _09854_;
  wire _09855_;
  wire _09856_;
  wire _09857_;
  wire _09858_;
  wire _09859_;
  wire _09860_;
  wire _09861_;
  wire _09862_;
  wire _09863_;
  wire _09864_;
  wire _09865_;
  wire _09866_;
  wire _09867_;
  wire _09868_;
  wire _09869_;
  wire _09870_;
  wire _09871_;
  wire _09872_;
  wire _09873_;
  wire _09874_;
  wire _09875_;
  wire _09876_;
  wire _09877_;
  wire _09878_;
  wire _09879_;
  wire _09880_;
  wire _09881_;
  wire _09882_;
  wire _09883_;
  wire _09884_;
  wire _09885_;
  wire _09886_;
  wire _09887_;
  wire _09888_;
  wire _09889_;
  wire _09890_;
  wire _09891_;
  wire _09892_;
  wire _09893_;
  wire _09894_;
  wire _09895_;
  wire _09896_;
  wire _09897_;
  wire _09898_;
  wire _09899_;
  wire _09900_;
  wire _09901_;
  wire _09902_;
  wire _09903_;
  wire _09904_;
  wire _09905_;
  wire _09906_;
  wire _09907_;
  wire _09908_;
  wire _09909_;
  wire _09910_;
  wire _09911_;
  wire _09912_;
  wire _09913_;
  wire _09914_;
  wire _09915_;
  wire _09916_;
  wire _09917_;
  wire _09918_;
  wire _09919_;
  wire _09920_;
  wire _09921_;
  wire _09922_;
  wire _09923_;
  wire _09924_;
  wire _09925_;
  wire _09926_;
  wire _09927_;
  wire _09928_;
  wire _09929_;
  wire _09930_;
  wire _09931_;
  wire _09932_;
  wire _09933_;
  wire _09934_;
  wire _09935_;
  wire _09936_;
  wire _09937_;
  wire _09938_;
  wire _09939_;
  wire _09940_;
  wire _09941_;
  wire _09942_;
  wire _09943_;
  wire _09944_;
  wire _09945_;
  wire _09946_;
  wire _09947_;
  wire _09948_;
  wire _09949_;
  wire _09950_;
  wire _09951_;
  wire _09952_;
  wire _09953_;
  wire _09954_;
  wire _09955_;
  wire _09956_;
  wire _09957_;
  wire _09958_;
  wire _09959_;
  wire _09960_;
  wire _09961_;
  wire _09962_;
  wire _09963_;
  wire _09964_;
  wire _09965_;
  wire _09966_;
  wire _09967_;
  wire _09968_;
  wire _09969_;
  wire _09970_;
  wire _09971_;
  wire _09972_;
  wire _09973_;
  wire _09974_;
  wire _09975_;
  wire _09976_;
  wire _09977_;
  wire _09978_;
  wire _09979_;
  wire _09980_;
  wire _09981_;
  wire _09982_;
  wire _09983_;
  wire _09984_;
  wire _09985_;
  wire _09986_;
  wire _09987_;
  wire _09988_;
  wire _09989_;
  wire _09990_;
  wire _09991_;
  wire _09992_;
  wire _09993_;
  wire _09994_;
  wire _09995_;
  wire _09996_;
  wire _09997_;
  wire _09998_;
  wire _09999_;
  wire _10000_;
  wire _10001_;
  wire _10002_;
  wire _10003_;
  wire _10004_;
  wire _10005_;
  wire _10006_;
  wire _10007_;
  wire _10008_;
  wire _10009_;
  wire _10010_;
  wire _10011_;
  wire _10012_;
  wire _10013_;
  wire _10014_;
  wire _10015_;
  wire _10016_;
  wire _10017_;
  wire _10018_;
  wire _10019_;
  wire _10020_;
  wire _10021_;
  wire _10022_;
  wire _10023_;
  wire _10024_;
  wire _10025_;
  wire _10026_;
  wire _10027_;
  wire _10028_;
  wire _10029_;
  wire _10030_;
  wire _10031_;
  wire _10032_;
  wire _10033_;
  wire _10034_;
  wire _10035_;
  wire _10036_;
  wire _10037_;
  wire _10038_;
  wire _10039_;
  wire _10040_;
  wire _10041_;
  wire _10042_;
  wire _10043_;
  wire _10044_;
  wire _10045_;
  wire _10046_;
  wire _10047_;
  wire _10048_;
  wire _10049_;
  wire _10050_;
  wire _10051_;
  wire _10052_;
  wire _10053_;
  wire _10054_;
  wire _10055_;
  wire _10056_;
  wire _10057_;
  wire _10058_;
  wire _10059_;
  wire _10060_;
  wire _10061_;
  wire _10062_;
  wire _10063_;
  wire _10064_;
  wire _10065_;
  wire _10066_;
  wire _10067_;
  wire _10068_;
  wire _10069_;
  wire _10070_;
  wire _10071_;
  wire _10072_;
  wire _10073_;
  wire _10074_;
  wire _10075_;
  wire _10076_;
  wire _10077_;
  wire _10078_;
  wire _10079_;
  wire _10080_;
  wire _10081_;
  wire _10082_;
  wire _10083_;
  wire _10084_;
  wire _10085_;
  wire _10086_;
  wire _10087_;
  wire _10088_;
  wire _10089_;
  wire _10090_;
  wire _10091_;
  wire _10092_;
  wire _10093_;
  wire _10094_;
  wire _10095_;
  wire _10096_;
  wire _10097_;
  wire _10098_;
  wire _10099_;
  wire _10100_;
  wire _10101_;
  wire _10102_;
  wire _10103_;
  wire _10104_;
  wire _10105_;
  wire _10106_;
  wire _10107_;
  wire _10108_;
  wire _10109_;
  wire _10110_;
  wire _10111_;
  wire _10112_;
  wire _10113_;
  wire _10114_;
  wire _10115_;
  wire _10116_;
  wire _10117_;
  wire _10118_;
  wire _10119_;
  wire _10120_;
  wire _10121_;
  wire _10122_;
  wire _10123_;
  wire _10124_;
  wire _10125_;
  wire _10126_;
  wire _10127_;
  wire _10128_;
  wire _10129_;
  wire _10130_;
  wire _10131_;
  wire _10132_;
  wire _10133_;
  wire _10134_;
  wire _10135_;
  wire _10136_;
  wire _10137_;
  wire _10138_;
  wire _10139_;
  wire _10140_;
  wire _10141_;
  wire _10142_;
  wire _10143_;
  wire _10144_;
  wire _10145_;
  wire _10146_;
  wire _10147_;
  wire _10148_;
  wire _10149_;
  wire _10150_;
  wire _10151_;
  wire _10152_;
  wire _10153_;
  wire _10154_;
  wire _10155_;
  wire _10156_;
  wire _10157_;
  wire _10158_;
  wire _10159_;
  wire _10160_;
  wire _10161_;
  wire _10162_;
  wire _10163_;
  wire _10164_;
  wire _10165_;
  wire _10166_;
  wire _10167_;
  wire _10168_;
  wire _10169_;
  wire _10170_;
  wire _10171_;
  wire _10172_;
  wire _10173_;
  wire _10174_;
  wire _10175_;
  wire _10176_;
  wire _10177_;
  wire _10178_;
  wire _10179_;
  wire _10180_;
  wire _10181_;
  wire _10182_;
  wire _10183_;
  wire _10184_;
  wire _10185_;
  wire _10186_;
  wire _10187_;
  wire _10188_;
  wire _10189_;
  wire _10190_;
  wire _10191_;
  wire _10192_;
  wire _10193_;
  wire _10194_;
  wire _10195_;
  wire _10196_;
  wire _10197_;
  wire _10198_;
  wire _10199_;
  wire _10200_;
  wire _10201_;
  wire _10202_;
  wire _10203_;
  wire _10204_;
  wire _10205_;
  wire _10206_;
  wire _10207_;
  wire _10208_;
  wire _10209_;
  wire _10210_;
  wire _10211_;
  wire _10212_;
  wire _10213_;
  wire _10214_;
  wire _10215_;
  wire _10216_;
  wire _10217_;
  wire _10218_;
  wire _10219_;
  wire _10220_;
  wire _10221_;
  wire _10222_;
  wire _10223_;
  wire _10224_;
  wire _10225_;
  wire _10226_;
  wire _10227_;
  wire _10228_;
  wire _10229_;
  wire _10230_;
  wire _10231_;
  wire _10232_;
  wire _10233_;
  wire _10234_;
  wire _10235_;
  wire _10236_;
  wire _10237_;
  wire _10238_;
  wire _10239_;
  wire _10240_;
  wire _10241_;
  wire _10242_;
  wire _10243_;
  wire _10244_;
  wire _10245_;
  wire _10246_;
  wire _10247_;
  wire _10248_;
  wire _10249_;
  wire _10250_;
  wire _10251_;
  wire _10252_;
  wire _10253_;
  wire _10254_;
  wire _10255_;
  wire _10256_;
  wire _10257_;
  wire _10258_;
  wire _10259_;
  wire _10260_;
  wire _10261_;
  wire _10262_;
  wire _10263_;
  wire _10264_;
  wire _10265_;
  wire _10266_;
  wire _10267_;
  wire _10268_;
  wire _10269_;
  wire _10270_;
  wire _10271_;
  wire _10272_;
  wire _10273_;
  wire _10274_;
  wire _10275_;
  wire _10276_;
  wire _10277_;
  wire _10278_;
  wire _10279_;
  wire _10280_;
  wire _10281_;
  wire _10282_;
  wire _10283_;
  wire _10284_;
  wire _10285_;
  wire _10286_;
  wire _10287_;
  wire _10288_;
  wire _10289_;
  wire _10290_;
  wire _10291_;
  wire _10292_;
  wire _10293_;
  wire _10294_;
  wire _10295_;
  wire _10296_;
  wire _10297_;
  wire _10298_;
  wire _10299_;
  wire _10300_;
  wire _10301_;
  wire _10302_;
  wire _10303_;
  wire _10304_;
  wire _10305_;
  wire _10306_;
  wire _10307_;
  wire _10308_;
  wire _10309_;
  wire _10310_;
  wire _10311_;
  wire _10312_;
  wire _10313_;
  wire _10314_;
  wire _10315_;
  wire _10316_;
  wire _10317_;
  wire _10318_;
  wire _10319_;
  wire _10320_;
  wire _10321_;
  wire _10322_;
  wire _10323_;
  wire _10324_;
  wire _10325_;
  wire _10326_;
  wire _10327_;
  wire _10328_;
  wire _10329_;
  wire _10330_;
  wire _10331_;
  wire _10332_;
  wire _10333_;
  wire _10334_;
  wire _10335_;
  wire _10336_;
  wire _10337_;
  wire _10338_;
  wire _10339_;
  wire _10340_;
  wire _10341_;
  wire _10342_;
  wire _10343_;
  wire _10344_;
  wire _10345_;
  wire _10346_;
  wire _10347_;
  wire _10348_;
  wire _10349_;
  wire _10350_;
  wire _10351_;
  wire _10352_;
  wire _10353_;
  wire _10354_;
  wire _10355_;
  wire _10356_;
  wire _10357_;
  wire _10358_;
  wire _10359_;
  wire _10360_;
  wire _10361_;
  wire _10362_;
  wire _10363_;
  wire _10364_;
  wire _10365_;
  wire _10366_;
  wire _10367_;
  wire _10368_;
  wire _10369_;
  wire _10370_;
  wire _10371_;
  wire _10372_;
  wire _10373_;
  wire _10374_;
  wire _10375_;
  wire _10376_;
  wire _10377_;
  wire _10378_;
  wire _10379_;
  wire _10380_;
  wire _10381_;
  wire _10382_;
  wire _10383_;
  wire _10384_;
  wire _10385_;
  wire _10386_;
  wire _10387_;
  wire _10388_;
  wire _10389_;
  wire _10390_;
  wire _10391_;
  wire _10392_;
  wire _10393_;
  wire _10394_;
  wire _10395_;
  wire _10396_;
  wire _10397_;
  wire _10398_;
  wire _10399_;
  wire _10400_;
  wire _10401_;
  wire _10402_;
  wire _10403_;
  wire _10404_;
  wire _10405_;
  wire _10406_;
  wire _10407_;
  wire _10408_;
  wire _10409_;
  wire _10410_;
  wire _10411_;
  wire _10412_;
  wire _10413_;
  wire _10414_;
  wire _10415_;
  wire _10416_;
  wire _10417_;
  wire _10418_;
  wire _10419_;
  wire _10420_;
  wire _10421_;
  wire _10422_;
  wire _10423_;
  wire _10424_;
  wire _10425_;
  wire _10426_;
  wire _10427_;
  wire _10428_;
  wire _10429_;
  wire _10430_;
  wire _10431_;
  wire _10432_;
  wire _10433_;
  wire _10434_;
  wire _10435_;
  wire _10436_;
  wire _10437_;
  wire _10438_;
  wire _10439_;
  wire _10440_;
  wire _10441_;
  wire _10442_;
  wire _10443_;
  wire _10444_;
  wire _10445_;
  wire _10446_;
  wire _10447_;
  wire _10448_;
  wire _10449_;
  wire _10450_;
  wire _10451_;
  wire _10452_;
  wire _10453_;
  wire _10454_;
  wire _10455_;
  wire _10456_;
  wire _10457_;
  wire _10458_;
  wire _10459_;
  wire _10460_;
  wire _10461_;
  wire _10462_;
  wire _10463_;
  wire _10464_;
  wire _10465_;
  wire _10466_;
  wire _10467_;
  wire _10468_;
  wire _10469_;
  wire _10470_;
  wire _10471_;
  wire _10472_;
  wire _10473_;
  wire _10474_;
  wire _10475_;
  wire _10476_;
  wire _10477_;
  wire _10478_;
  wire _10479_;
  wire _10480_;
  wire _10481_;
  wire _10482_;
  wire _10483_;
  wire _10484_;
  wire _10485_;
  wire _10486_;
  wire _10487_;
  wire _10488_;
  wire _10489_;
  wire _10490_;
  wire _10491_;
  wire _10492_;
  wire _10493_;
  wire _10494_;
  wire _10495_;
  wire _10496_;
  wire _10497_;
  wire _10498_;
  wire _10499_;
  wire _10500_;
  wire _10501_;
  wire _10502_;
  wire _10503_;
  wire _10504_;
  wire _10505_;
  wire _10506_;
  wire _10507_;
  wire _10508_;
  wire _10509_;
  wire _10510_;
  wire _10511_;
  wire _10512_;
  wire _10513_;
  wire _10514_;
  wire _10515_;
  wire _10516_;
  wire _10517_;
  wire _10518_;
  wire _10519_;
  wire _10520_;
  wire _10521_;
  wire _10522_;
  wire _10523_;
  wire _10524_;
  wire _10525_;
  wire _10526_;
  wire _10527_;
  wire _10528_;
  wire _10529_;
  wire _10530_;
  wire _10531_;
  wire _10532_;
  wire _10533_;
  wire _10534_;
  wire _10535_;
  wire _10536_;
  wire _10537_;
  wire _10538_;
  wire _10539_;
  wire _10540_;
  wire _10541_;
  wire _10542_;
  wire _10543_;
  wire _10544_;
  wire _10545_;
  wire _10546_;
  wire _10547_;
  wire _10548_;
  wire _10549_;
  wire _10550_;
  wire _10551_;
  wire _10552_;
  wire _10553_;
  wire _10554_;
  wire _10555_;
  wire _10556_;
  wire _10557_;
  wire _10558_;
  wire _10559_;
  wire _10560_;
  wire _10561_;
  wire _10562_;
  wire _10563_;
  wire _10564_;
  wire _10565_;
  wire _10566_;
  wire _10567_;
  wire _10568_;
  wire _10569_;
  wire _10570_;
  wire _10571_;
  wire _10572_;
  wire _10573_;
  wire _10574_;
  wire _10575_;
  wire _10576_;
  wire _10577_;
  wire _10578_;
  wire _10579_;
  wire _10580_;
  wire _10581_;
  wire _10582_;
  wire _10583_;
  wire _10584_;
  wire _10585_;
  wire _10586_;
  wire _10587_;
  wire _10588_;
  wire _10589_;
  wire _10590_;
  wire _10591_;
  wire _10592_;
  wire _10593_;
  wire _10594_;
  wire _10595_;
  wire _10596_;
  wire _10597_;
  wire _10598_;
  wire _10599_;
  wire _10600_;
  wire _10601_;
  wire _10602_;
  wire _10603_;
  wire _10604_;
  wire _10605_;
  wire _10606_;
  wire _10607_;
  wire _10608_;
  wire _10609_;
  wire _10610_;
  wire _10611_;
  wire _10612_;
  wire _10613_;
  wire _10614_;
  wire _10615_;
  wire _10616_;
  wire _10617_;
  wire _10618_;
  wire _10619_;
  wire _10620_;
  wire _10621_;
  wire _10622_;
  wire _10623_;
  wire _10624_;
  wire _10625_;
  wire _10626_;
  wire _10627_;
  wire _10628_;
  wire _10629_;
  wire _10630_;
  wire _10631_;
  wire _10632_;
  wire _10633_;
  wire _10634_;
  wire _10635_;
  wire _10636_;
  wire _10637_;
  wire _10638_;
  wire _10639_;
  wire _10640_;
  wire _10641_;
  wire _10642_;
  wire _10643_;
  wire _10644_;
  wire _10645_;
  wire _10646_;
  wire _10647_;
  wire _10648_;
  wire _10649_;
  wire _10650_;
  wire _10651_;
  wire _10652_;
  wire _10653_;
  wire _10654_;
  wire _10655_;
  wire _10656_;
  wire _10657_;
  wire _10658_;
  wire _10659_;
  wire _10660_;
  wire _10661_;
  wire _10662_;
  wire _10663_;
  wire _10664_;
  wire _10665_;
  wire _10666_;
  wire _10667_;
  wire _10668_;
  wire _10669_;
  wire _10670_;
  wire _10671_;
  wire _10672_;
  wire _10673_;
  wire _10674_;
  wire _10675_;
  wire _10676_;
  wire _10677_;
  wire _10678_;
  wire _10679_;
  wire _10680_;
  wire _10681_;
  wire _10682_;
  wire _10683_;
  wire _10684_;
  wire _10685_;
  wire _10686_;
  wire _10687_;
  wire _10688_;
  wire _10689_;
  wire _10690_;
  wire _10691_;
  wire _10692_;
  wire _10693_;
  wire _10694_;
  wire _10695_;
  wire _10696_;
  wire _10697_;
  wire _10698_;
  wire _10699_;
  wire _10700_;
  wire _10701_;
  wire _10702_;
  wire _10703_;
  wire _10704_;
  wire _10705_;
  wire _10706_;
  wire _10707_;
  wire _10708_;
  wire _10709_;
  wire _10710_;
  wire _10711_;
  wire _10712_;
  wire _10713_;
  wire _10714_;
  wire _10715_;
  wire _10716_;
  wire _10717_;
  wire _10718_;
  wire _10719_;
  wire _10720_;
  wire _10721_;
  wire _10722_;
  wire _10723_;
  wire _10724_;
  wire _10725_;
  wire _10726_;
  wire _10727_;
  wire _10728_;
  wire _10729_;
  wire _10730_;
  wire _10731_;
  wire _10732_;
  wire _10733_;
  wire _10734_;
  wire _10735_;
  wire _10736_;
  wire _10737_;
  wire _10738_;
  wire _10739_;
  wire _10740_;
  wire _10741_;
  wire _10742_;
  wire _10743_;
  wire _10744_;
  wire _10745_;
  wire _10746_;
  wire _10747_;
  wire _10748_;
  wire _10749_;
  wire _10750_;
  wire _10751_;
  wire _10752_;
  wire _10753_;
  wire _10754_;
  wire _10755_;
  wire _10756_;
  wire _10757_;
  wire _10758_;
  wire _10759_;
  wire _10760_;
  wire _10761_;
  wire _10762_;
  wire _10763_;
  wire _10764_;
  wire _10765_;
  wire _10766_;
  wire _10767_;
  wire _10768_;
  wire _10769_;
  wire _10770_;
  wire _10771_;
  wire _10772_;
  wire _10773_;
  wire _10774_;
  wire _10775_;
  wire _10776_;
  wire _10777_;
  wire _10778_;
  wire _10779_;
  wire _10780_;
  wire _10781_;
  wire _10782_;
  wire _10783_;
  wire _10784_;
  wire _10785_;
  wire _10786_;
  wire _10787_;
  wire _10788_;
  wire _10789_;
  wire _10790_;
  wire _10791_;
  wire _10792_;
  wire _10793_;
  wire _10794_;
  wire _10795_;
  wire _10796_;
  wire _10797_;
  wire _10798_;
  wire _10799_;
  wire _10800_;
  wire _10801_;
  wire _10802_;
  wire _10803_;
  wire _10804_;
  wire _10805_;
  wire _10806_;
  wire _10807_;
  wire _10808_;
  wire _10809_;
  wire _10810_;
  wire _10811_;
  wire _10812_;
  wire _10813_;
  wire _10814_;
  wire _10815_;
  wire _10816_;
  wire _10817_;
  wire _10818_;
  wire _10819_;
  wire _10820_;
  wire _10821_;
  wire _10822_;
  wire _10823_;
  wire _10824_;
  wire _10825_;
  wire _10826_;
  wire _10827_;
  wire _10828_;
  wire _10829_;
  wire _10830_;
  wire _10831_;
  wire _10832_;
  wire _10833_;
  wire _10834_;
  wire _10835_;
  wire _10836_;
  wire _10837_;
  wire _10838_;
  wire _10839_;
  wire _10840_;
  wire _10841_;
  wire _10842_;
  wire _10843_;
  wire _10844_;
  wire _10845_;
  wire _10846_;
  wire _10847_;
  wire _10848_;
  wire _10849_;
  wire _10850_;
  wire _10851_;
  wire _10852_;
  wire _10853_;
  wire _10854_;
  wire _10855_;
  wire _10856_;
  wire _10857_;
  wire _10858_;
  wire _10859_;
  wire _10860_;
  wire _10861_;
  wire _10862_;
  wire _10863_;
  wire _10864_;
  wire _10865_;
  wire _10866_;
  wire _10867_;
  wire _10868_;
  wire _10869_;
  wire _10870_;
  wire _10871_;
  wire _10872_;
  wire _10873_;
  wire _10874_;
  wire _10875_;
  wire _10876_;
  wire _10877_;
  wire _10878_;
  wire _10879_;
  wire _10880_;
  wire _10881_;
  wire _10882_;
  wire _10883_;
  wire _10884_;
  wire _10885_;
  wire _10886_;
  wire _10887_;
  wire _10888_;
  wire _10889_;
  wire _10890_;
  wire _10891_;
  wire _10892_;
  wire _10893_;
  wire _10894_;
  wire _10895_;
  wire _10896_;
  wire _10897_;
  wire _10898_;
  wire _10899_;
  wire _10900_;
  wire _10901_;
  wire _10902_;
  wire _10903_;
  wire _10904_;
  wire _10905_;
  wire _10906_;
  wire _10907_;
  wire _10908_;
  wire _10909_;
  wire _10910_;
  wire _10911_;
  wire _10912_;
  wire _10913_;
  wire _10914_;
  wire _10915_;
  wire _10916_;
  wire _10917_;
  wire _10918_;
  wire _10919_;
  wire _10920_;
  wire _10921_;
  wire _10922_;
  wire _10923_;
  wire _10924_;
  wire _10925_;
  wire _10926_;
  wire _10927_;
  wire _10928_;
  wire _10929_;
  wire _10930_;
  wire _10931_;
  wire _10932_;
  wire _10933_;
  wire _10934_;
  wire _10935_;
  wire _10936_;
  wire _10937_;
  wire _10938_;
  wire _10939_;
  wire _10940_;
  wire _10941_;
  wire _10942_;
  wire _10943_;
  wire _10944_;
  wire _10945_;
  wire _10946_;
  wire _10947_;
  wire _10948_;
  wire _10949_;
  wire _10950_;
  wire _10951_;
  wire _10952_;
  wire _10953_;
  wire _10954_;
  wire _10955_;
  wire _10956_;
  wire _10957_;
  wire _10958_;
  wire _10959_;
  wire _10960_;
  wire _10961_;
  wire _10962_;
  wire _10963_;
  wire _10964_;
  wire _10965_;
  wire _10966_;
  wire _10967_;
  wire _10968_;
  wire _10969_;
  wire _10970_;
  wire _10971_;
  wire _10972_;
  wire _10973_;
  wire _10974_;
  wire _10975_;
  wire _10976_;
  wire _10977_;
  wire _10978_;
  wire _10979_;
  wire _10980_;
  wire _10981_;
  wire _10982_;
  wire _10983_;
  wire _10984_;
  wire _10985_;
  wire _10986_;
  wire _10987_;
  wire _10988_;
  wire _10989_;
  wire _10990_;
  wire _10991_;
  wire _10992_;
  wire _10993_;
  wire _10994_;
  wire _10995_;
  wire _10996_;
  wire _10997_;
  wire _10998_;
  wire _10999_;
  wire _11000_;
  wire _11001_;
  wire _11002_;
  wire _11003_;
  wire _11004_;
  wire _11005_;
  wire _11006_;
  wire _11007_;
  wire _11008_;
  wire _11009_;
  wire _11010_;
  wire _11011_;
  wire _11012_;
  wire _11013_;
  wire _11014_;
  wire _11015_;
  wire _11016_;
  wire _11017_;
  wire _11018_;
  wire _11019_;
  wire _11020_;
  wire _11021_;
  wire _11022_;
  wire _11023_;
  wire _11024_;
  wire _11025_;
  wire _11026_;
  wire _11027_;
  wire _11028_;
  wire _11029_;
  wire _11030_;
  wire _11031_;
  wire _11032_;
  wire _11033_;
  wire _11034_;
  wire _11035_;
  wire _11036_;
  wire _11037_;
  wire _11038_;
  wire _11039_;
  wire _11040_;
  wire _11041_;
  wire _11042_;
  wire _11043_;
  wire _11044_;
  wire _11045_;
  wire _11046_;
  wire _11047_;
  wire _11048_;
  wire _11049_;
  wire _11050_;
  wire _11051_;
  wire _11052_;
  wire _11053_;
  wire _11054_;
  wire _11055_;
  wire _11056_;
  wire _11057_;
  wire _11058_;
  wire _11059_;
  wire _11060_;
  wire _11061_;
  wire _11062_;
  wire _11063_;
  wire _11064_;
  wire _11065_;
  wire _11066_;
  wire _11067_;
  wire _11068_;
  wire _11069_;
  wire _11070_;
  wire _11071_;
  wire _11072_;
  wire _11073_;
  wire _11074_;
  wire _11075_;
  wire _11076_;
  wire _11077_;
  wire _11078_;
  wire _11079_;
  wire _11080_;
  wire _11081_;
  wire _11082_;
  wire _11083_;
  wire _11084_;
  wire _11085_;
  wire _11086_;
  wire _11087_;
  wire _11088_;
  wire _11089_;
  wire _11090_;
  wire _11091_;
  wire _11092_;
  wire _11093_;
  wire _11094_;
  wire _11095_;
  wire _11096_;
  wire _11097_;
  wire _11098_;
  wire _11099_;
  wire _11100_;
  wire _11101_;
  wire _11102_;
  wire _11103_;
  wire _11104_;
  wire _11105_;
  wire _11106_;
  wire _11107_;
  wire _11108_;
  wire _11109_;
  wire _11110_;
  wire _11111_;
  wire _11112_;
  wire _11113_;
  wire _11114_;
  wire _11115_;
  wire _11116_;
  wire _11117_;
  wire _11118_;
  wire _11119_;
  wire _11120_;
  wire _11121_;
  wire _11122_;
  wire _11123_;
  wire _11124_;
  wire _11125_;
  wire _11126_;
  wire _11127_;
  wire _11128_;
  wire _11129_;
  wire _11130_;
  wire _11131_;
  wire _11132_;
  wire _11133_;
  wire _11134_;
  wire _11135_;
  wire _11136_;
  wire _11137_;
  wire _11138_;
  wire _11139_;
  wire _11140_;
  wire _11141_;
  wire _11142_;
  wire _11143_;
  wire _11144_;
  wire _11145_;
  wire _11146_;
  wire _11147_;
  wire _11148_;
  wire _11149_;
  wire _11150_;
  wire _11151_;
  wire _11152_;
  wire _11153_;
  wire _11154_;
  wire _11155_;
  wire _11156_;
  wire _11157_;
  wire _11158_;
  wire _11159_;
  wire _11160_;
  wire _11161_;
  wire _11162_;
  wire _11163_;
  wire _11164_;
  wire _11165_;
  wire _11166_;
  wire _11167_;
  wire _11168_;
  wire _11169_;
  wire _11170_;
  wire _11171_;
  wire _11172_;
  wire _11173_;
  wire _11174_;
  wire _11175_;
  wire _11176_;
  wire _11177_;
  wire _11178_;
  wire _11179_;
  wire _11180_;
  wire _11181_;
  wire _11182_;
  wire _11183_;
  wire _11184_;
  wire _11185_;
  wire _11186_;
  wire _11187_;
  wire _11188_;
  wire _11189_;
  wire _11190_;
  wire _11191_;
  wire _11192_;
  wire _11193_;
  wire _11194_;
  wire _11195_;
  wire _11196_;
  wire _11197_;
  wire _11198_;
  wire _11199_;
  wire _11200_;
  wire _11201_;
  wire _11202_;
  wire _11203_;
  wire _11204_;
  wire _11205_;
  wire _11206_;
  wire _11207_;
  wire _11208_;
  wire _11209_;
  wire _11210_;
  wire _11211_;
  wire _11212_;
  wire _11213_;
  wire _11214_;
  wire _11215_;
  wire _11216_;
  wire _11217_;
  wire _11218_;
  wire _11219_;
  wire _11220_;
  wire _11221_;
  wire _11222_;
  wire _11223_;
  wire _11224_;
  wire _11225_;
  wire _11226_;
  wire _11227_;
  wire _11228_;
  wire _11229_;
  wire _11230_;
  wire _11231_;
  wire _11232_;
  wire _11233_;
  wire _11234_;
  wire _11235_;
  wire _11236_;
  wire _11237_;
  wire _11238_;
  wire _11239_;
  wire _11240_;
  wire _11241_;
  wire _11242_;
  wire _11243_;
  wire _11244_;
  wire _11245_;
  wire _11246_;
  wire _11247_;
  wire _11248_;
  wire _11249_;
  wire _11250_;
  wire _11251_;
  wire _11252_;
  wire _11253_;
  wire _11254_;
  wire _11255_;
  wire _11256_;
  wire _11257_;
  wire _11258_;
  wire _11259_;
  wire _11260_;
  wire _11261_;
  wire _11262_;
  wire _11263_;
  wire _11264_;
  wire _11265_;
  wire _11266_;
  wire _11267_;
  wire _11268_;
  wire _11269_;
  wire _11270_;
  wire _11271_;
  wire _11272_;
  wire _11273_;
  wire _11274_;
  wire _11275_;
  wire _11276_;
  wire _11277_;
  wire _11278_;
  wire _11279_;
  wire _11280_;
  wire _11281_;
  wire _11282_;
  wire _11283_;
  wire _11284_;
  wire _11285_;
  wire _11286_;
  wire _11287_;
  wire _11288_;
  wire _11289_;
  wire _11290_;
  wire _11291_;
  wire _11292_;
  wire _11293_;
  wire _11294_;
  wire _11295_;
  wire _11296_;
  wire _11297_;
  wire _11298_;
  wire _11299_;
  wire _11300_;
  wire _11301_;
  wire _11302_;
  wire _11303_;
  wire _11304_;
  wire _11305_;
  wire _11306_;
  wire _11307_;
  wire _11308_;
  wire _11309_;
  wire _11310_;
  wire _11311_;
  wire _11312_;
  wire _11313_;
  wire _11314_;
  wire _11315_;
  wire _11316_;
  wire _11317_;
  wire _11318_;
  wire _11319_;
  wire _11320_;
  wire _11321_;
  wire _11322_;
  wire _11323_;
  wire _11324_;
  wire _11325_;
  wire _11326_;
  wire _11327_;
  wire _11328_;
  wire _11329_;
  wire _11330_;
  wire _11331_;
  wire _11332_;
  wire _11333_;
  wire _11334_;
  wire _11335_;
  wire _11336_;
  wire _11337_;
  wire _11338_;
  wire _11339_;
  wire _11340_;
  wire _11341_;
  wire _11342_;
  wire _11343_;
  wire _11344_;
  wire _11345_;
  wire _11346_;
  wire _11347_;
  wire _11348_;
  wire _11349_;
  wire _11350_;
  wire _11351_;
  wire _11352_;
  wire _11353_;
  wire _11354_;
  wire _11355_;
  wire _11356_;
  wire _11357_;
  wire _11358_;
  wire _11359_;
  wire _11360_;
  wire _11361_;
  wire _11362_;
  wire _11363_;
  wire _11364_;
  wire _11365_;
  wire _11366_;
  wire _11367_;
  wire _11368_;
  wire _11369_;
  wire _11370_;
  wire _11371_;
  wire _11372_;
  wire _11373_;
  wire _11374_;
  wire _11375_;
  wire _11376_;
  wire _11377_;
  wire _11378_;
  wire _11379_;
  wire _11380_;
  wire _11381_;
  wire _11382_;
  wire _11383_;
  wire _11384_;
  wire _11385_;
  wire _11386_;
  wire _11387_;
  wire _11388_;
  wire _11389_;
  wire _11390_;
  wire _11391_;
  wire _11392_;
  wire _11393_;
  wire _11394_;
  wire _11395_;
  wire _11396_;
  wire _11397_;
  wire _11398_;
  wire _11399_;
  wire _11400_;
  wire _11401_;
  wire _11402_;
  wire _11403_;
  wire _11404_;
  wire _11405_;
  wire _11406_;
  wire _11407_;
  wire _11408_;
  wire _11409_;
  wire _11410_;
  wire _11411_;
  wire _11412_;
  wire _11413_;
  wire _11414_;
  wire _11415_;
  wire _11416_;
  wire _11417_;
  wire _11418_;
  wire _11419_;
  wire _11420_;
  wire _11421_;
  wire _11422_;
  wire _11423_;
  wire _11424_;
  wire _11425_;
  wire _11426_;
  wire _11427_;
  wire _11428_;
  wire _11429_;
  wire _11430_;
  wire _11431_;
  wire _11432_;
  wire _11433_;
  wire _11434_;
  wire _11435_;
  wire _11436_;
  wire _11437_;
  wire _11438_;
  wire _11439_;
  wire _11440_;
  wire _11441_;
  wire _11442_;
  wire _11443_;
  wire _11444_;
  wire _11445_;
  wire _11446_;
  wire _11447_;
  wire _11448_;
  wire _11449_;
  wire _11450_;
  wire _11451_;
  wire _11452_;
  wire _11453_;
  wire _11454_;
  wire _11455_;
  wire _11456_;
  wire _11457_;
  wire _11458_;
  wire _11459_;
  wire _11460_;
  wire _11461_;
  wire _11462_;
  wire _11463_;
  wire _11464_;
  wire _11465_;
  wire _11466_;
  wire _11467_;
  wire _11468_;
  wire _11469_;
  wire _11470_;
  wire _11471_;
  wire _11472_;
  wire _11473_;
  wire _11474_;
  wire _11475_;
  wire _11476_;
  wire _11477_;
  wire _11478_;
  wire _11479_;
  wire _11480_;
  wire _11481_;
  wire _11482_;
  wire _11483_;
  wire _11484_;
  wire _11485_;
  wire _11486_;
  wire _11487_;
  wire _11488_;
  wire _11489_;
  wire _11490_;
  wire _11491_;
  wire _11492_;
  wire _11493_;
  wire _11494_;
  wire _11495_;
  wire _11496_;
  wire _11497_;
  wire _11498_;
  wire _11499_;
  wire _11500_;
  wire _11501_;
  wire _11502_;
  wire _11503_;
  wire _11504_;
  wire _11505_;
  wire _11506_;
  wire _11507_;
  wire _11508_;
  wire _11509_;
  wire _11510_;
  wire _11511_;
  wire _11512_;
  wire _11513_;
  wire _11514_;
  wire _11515_;
  wire _11516_;
  wire _11517_;
  wire _11518_;
  wire _11519_;
  wire _11520_;
  wire _11521_;
  wire _11522_;
  wire _11523_;
  wire _11524_;
  wire _11525_;
  wire _11526_;
  wire _11527_;
  wire _11528_;
  wire _11529_;
  wire _11530_;
  wire _11531_;
  wire _11532_;
  wire _11533_;
  wire _11534_;
  wire _11535_;
  wire _11536_;
  wire _11537_;
  wire _11538_;
  wire _11539_;
  wire _11540_;
  wire _11541_;
  wire _11542_;
  wire _11543_;
  wire _11544_;
  wire _11545_;
  wire _11546_;
  wire _11547_;
  wire _11548_;
  wire _11549_;
  wire _11550_;
  wire _11551_;
  wire _11552_;
  wire _11553_;
  wire _11554_;
  wire _11555_;
  wire _11556_;
  wire _11557_;
  wire _11558_;
  wire _11559_;
  wire _11560_;
  wire _11561_;
  wire _11562_;
  wire _11563_;
  wire _11564_;
  wire _11565_;
  wire _11566_;
  wire _11567_;
  wire _11568_;
  wire _11569_;
  wire _11570_;
  wire _11571_;
  wire _11572_;
  wire _11573_;
  wire _11574_;
  wire _11575_;
  wire _11576_;
  wire _11577_;
  wire _11578_;
  wire _11579_;
  wire _11580_;
  wire _11581_;
  wire _11582_;
  wire _11583_;
  wire _11584_;
  wire _11585_;
  wire _11586_;
  wire _11587_;
  wire _11588_;
  wire _11589_;
  wire _11590_;
  wire _11591_;
  wire _11592_;
  wire _11593_;
  wire _11594_;
  wire _11595_;
  wire _11596_;
  wire _11597_;
  wire _11598_;
  wire _11599_;
  wire _11600_;
  wire _11601_;
  wire _11602_;
  wire _11603_;
  wire _11604_;
  wire _11605_;
  wire _11606_;
  wire _11607_;
  wire _11608_;
  wire _11609_;
  wire _11610_;
  wire _11611_;
  wire _11612_;
  wire _11613_;
  wire _11614_;
  wire _11615_;
  wire _11616_;
  wire _11617_;
  wire _11618_;
  wire _11619_;
  wire _11620_;
  wire _11621_;
  wire _11622_;
  wire _11623_;
  wire _11624_;
  wire _11625_;
  wire _11626_;
  wire _11627_;
  wire _11628_;
  wire _11629_;
  wire _11630_;
  wire _11631_;
  wire _11632_;
  wire _11633_;
  wire _11634_;
  wire _11635_;
  wire _11636_;
  wire _11637_;
  wire _11638_;
  wire _11639_;
  wire _11640_;
  wire _11641_;
  wire _11642_;
  wire _11643_;
  wire _11644_;
  wire _11645_;
  wire _11646_;
  wire _11647_;
  wire _11648_;
  wire _11649_;
  wire _11650_;
  wire _11651_;
  wire _11652_;
  wire _11653_;
  wire _11654_;
  wire _11655_;
  wire _11656_;
  wire _11657_;
  wire _11658_;
  wire _11659_;
  wire _11660_;
  wire _11661_;
  wire _11662_;
  wire _11663_;
  wire _11664_;
  wire _11665_;
  wire _11666_;
  wire _11667_;
  wire _11668_;
  wire _11669_;
  wire _11670_;
  wire _11671_;
  wire _11672_;
  wire _11673_;
  wire _11674_;
  wire _11675_;
  wire _11676_;
  wire _11677_;
  wire _11678_;
  wire _11679_;
  wire _11680_;
  wire _11681_;
  wire _11682_;
  wire _11683_;
  wire _11684_;
  wire _11685_;
  wire _11686_;
  wire _11687_;
  wire _11688_;
  wire _11689_;
  wire _11690_;
  wire _11691_;
  wire _11692_;
  wire _11693_;
  wire _11694_;
  wire _11695_;
  wire _11696_;
  wire _11697_;
  wire _11698_;
  wire _11699_;
  wire _11700_;
  wire _11701_;
  wire _11702_;
  wire _11703_;
  wire _11704_;
  wire _11705_;
  wire _11706_;
  wire _11707_;
  wire _11708_;
  wire _11709_;
  wire _11710_;
  wire _11711_;
  wire _11712_;
  wire _11713_;
  wire _11714_;
  wire _11715_;
  wire _11716_;
  wire _11717_;
  wire _11718_;
  wire _11719_;
  wire _11720_;
  wire _11721_;
  wire _11722_;
  wire _11723_;
  wire _11724_;
  wire _11725_;
  wire _11726_;
  wire _11727_;
  wire _11728_;
  wire _11729_;
  wire _11730_;
  wire _11731_;
  wire _11732_;
  wire _11733_;
  wire _11734_;
  wire _11735_;
  wire _11736_;
  wire _11737_;
  wire _11738_;
  wire _11739_;
  wire _11740_;
  wire _11741_;
  wire _11742_;
  wire _11743_;
  wire _11744_;
  wire _11745_;
  wire _11746_;
  wire _11747_;
  wire _11748_;
  wire _11749_;
  wire _11750_;
  wire _11751_;
  wire _11752_;
  wire _11753_;
  wire _11754_;
  wire _11755_;
  wire _11756_;
  wire _11757_;
  wire _11758_;
  wire _11759_;
  wire _11760_;
  wire _11761_;
  wire _11762_;
  wire _11763_;
  wire _11764_;
  wire _11765_;
  wire _11766_;
  wire _11767_;
  wire _11768_;
  wire _11769_;
  wire _11770_;
  wire _11771_;
  wire _11772_;
  wire _11773_;
  wire _11774_;
  wire _11775_;
  wire _11776_;
  wire _11777_;
  wire _11778_;
  wire _11779_;
  wire _11780_;
  wire _11781_;
  wire _11782_;
  wire _11783_;
  wire _11784_;
  wire _11785_;
  wire _11786_;
  wire _11787_;
  wire _11788_;
  wire _11789_;
  wire _11790_;
  wire _11791_;
  wire _11792_;
  wire _11793_;
  wire _11794_;
  wire _11795_;
  wire _11796_;
  wire _11797_;
  wire _11798_;
  wire _11799_;
  wire _11800_;
  wire _11801_;
  wire _11802_;
  wire _11803_;
  wire _11804_;
  wire _11805_;
  wire _11806_;
  wire _11807_;
  wire _11808_;
  wire _11809_;
  wire _11810_;
  wire _11811_;
  wire _11812_;
  wire _11813_;
  wire _11814_;
  wire _11815_;
  wire _11816_;
  wire _11817_;
  wire _11818_;
  wire _11819_;
  wire _11820_;
  wire _11821_;
  wire _11822_;
  wire _11823_;
  wire _11824_;
  wire _11825_;
  wire _11826_;
  wire _11827_;
  wire _11828_;
  wire _11829_;
  wire _11830_;
  wire _11831_;
  wire _11832_;
  wire _11833_;
  wire _11834_;
  wire _11835_;
  wire _11836_;
  wire _11837_;
  wire _11838_;
  wire _11839_;
  wire _11840_;
  wire _11841_;
  wire _11842_;
  wire _11843_;
  wire _11844_;
  wire _11845_;
  wire _11846_;
  wire _11847_;
  wire _11848_;
  wire _11849_;
  wire _11850_;
  wire _11851_;
  wire _11852_;
  wire _11853_;
  wire _11854_;
  wire _11855_;
  wire _11856_;
  wire _11857_;
  wire _11858_;
  wire _11859_;
  wire _11860_;
  wire _11861_;
  wire _11862_;
  wire _11863_;
  wire _11864_;
  wire _11865_;
  wire _11866_;
  wire _11867_;
  wire _11868_;
  wire _11869_;
  wire _11870_;
  wire _11871_;
  wire _11872_;
  wire _11873_;
  wire _11874_;
  wire _11875_;
  wire _11876_;
  wire _11877_;
  wire _11878_;
  wire _11879_;
  wire _11880_;
  wire _11881_;
  wire _11882_;
  wire _11883_;
  wire _11884_;
  wire _11885_;
  wire _11886_;
  wire _11887_;
  wire _11888_;
  wire _11889_;
  wire _11890_;
  wire _11891_;
  wire _11892_;
  wire _11893_;
  wire _11894_;
  wire _11895_;
  wire _11896_;
  wire _11897_;
  wire _11898_;
  wire _11899_;
  wire _11900_;
  wire _11901_;
  wire _11902_;
  wire _11903_;
  wire _11904_;
  wire _11905_;
  wire _11906_;
  wire _11907_;
  wire _11908_;
  wire _11909_;
  wire _11910_;
  wire _11911_;
  wire _11912_;
  wire _11913_;
  wire _11914_;
  wire _11915_;
  wire _11916_;
  wire _11917_;
  wire _11918_;
  wire _11919_;
  wire _11920_;
  wire _11921_;
  wire _11922_;
  wire _11923_;
  wire _11924_;
  wire _11925_;
  wire _11926_;
  wire _11927_;
  wire _11928_;
  wire _11929_;
  wire _11930_;
  wire _11931_;
  wire _11932_;
  wire _11933_;
  wire _11934_;
  wire _11935_;
  wire _11936_;
  wire _11937_;
  wire _11938_;
  wire _11939_;
  wire _11940_;
  wire _11941_;
  wire _11942_;
  wire _11943_;
  wire _11944_;
  wire _11945_;
  wire _11946_;
  wire _11947_;
  wire _11948_;
  wire _11949_;
  wire _11950_;
  wire _11951_;
  wire _11952_;
  wire _11953_;
  wire _11954_;
  wire _11955_;
  wire _11956_;
  wire _11957_;
  wire _11958_;
  wire _11959_;
  wire _11960_;
  wire _11961_;
  wire _11962_;
  wire _11963_;
  wire _11964_;
  wire _11965_;
  wire _11966_;
  wire _11967_;
  wire _11968_;
  wire _11969_;
  wire _11970_;
  wire _11971_;
  wire _11972_;
  wire _11973_;
  wire _11974_;
  wire _11975_;
  wire _11976_;
  wire _11977_;
  wire _11978_;
  wire _11979_;
  wire _11980_;
  wire _11981_;
  wire _11982_;
  wire _11983_;
  wire _11984_;
  wire _11985_;
  wire _11986_;
  wire _11987_;
  wire _11988_;
  wire _11989_;
  wire _11990_;
  wire _11991_;
  wire _11992_;
  wire _11993_;
  wire _11994_;
  wire _11995_;
  wire _11996_;
  wire _11997_;
  wire _11998_;
  wire _11999_;
  wire _12000_;
  wire _12001_;
  wire _12002_;
  wire _12003_;
  wire _12004_;
  wire _12005_;
  wire _12006_;
  wire _12007_;
  wire _12008_;
  wire _12009_;
  wire _12010_;
  wire _12011_;
  wire _12012_;
  wire _12013_;
  wire _12014_;
  wire _12015_;
  wire _12016_;
  wire _12017_;
  wire _12018_;
  wire _12019_;
  wire _12020_;
  wire _12021_;
  wire _12022_;
  wire _12023_;
  wire _12024_;
  wire _12025_;
  wire _12026_;
  wire _12027_;
  wire _12028_;
  wire _12029_;
  wire _12030_;
  wire _12031_;
  wire _12032_;
  wire _12033_;
  wire _12034_;
  wire _12035_;
  wire _12036_;
  wire _12037_;
  wire _12038_;
  wire _12039_;
  wire _12040_;
  wire _12041_;
  wire _12042_;
  wire _12043_;
  wire _12044_;
  wire _12045_;
  wire _12046_;
  wire _12047_;
  wire _12048_;
  wire _12049_;
  wire _12050_;
  wire _12051_;
  wire _12052_;
  wire _12053_;
  wire _12054_;
  wire _12055_;
  wire _12056_;
  wire _12057_;
  wire _12058_;
  wire _12059_;
  wire _12060_;
  wire _12061_;
  wire _12062_;
  wire _12063_;
  wire _12064_;
  wire _12065_;
  wire _12066_;
  wire _12067_;
  wire _12068_;
  wire _12069_;
  wire _12070_;
  wire _12071_;
  wire _12072_;
  wire _12073_;
  wire _12074_;
  wire _12075_;
  wire _12076_;
  wire _12077_;
  wire _12078_;
  wire _12079_;
  wire _12080_;
  wire _12081_;
  wire _12082_;
  wire _12083_;
  wire _12084_;
  wire _12085_;
  wire _12086_;
  wire _12087_;
  wire _12088_;
  wire _12089_;
  wire _12090_;
  wire _12091_;
  wire _12092_;
  wire _12093_;
  wire _12094_;
  wire _12095_;
  wire _12096_;
  wire _12097_;
  wire _12098_;
  wire _12099_;
  wire _12100_;
  wire _12101_;
  wire _12102_;
  wire _12103_;
  wire _12104_;
  wire _12105_;
  wire _12106_;
  wire _12107_;
  wire _12108_;
  wire _12109_;
  wire _12110_;
  wire _12111_;
  wire _12112_;
  wire _12113_;
  wire _12114_;
  wire _12115_;
  wire _12116_;
  wire _12117_;
  wire _12118_;
  wire _12119_;
  wire _12120_;
  wire _12121_;
  wire _12122_;
  wire _12123_;
  wire _12124_;
  wire _12125_;
  wire _12126_;
  wire _12127_;
  wire _12128_;
  wire _12129_;
  wire _12130_;
  wire _12131_;
  wire _12132_;
  wire _12133_;
  wire _12134_;
  wire _12135_;
  wire _12136_;
  wire _12137_;
  wire _12138_;
  wire _12139_;
  wire _12140_;
  wire _12141_;
  wire _12142_;
  wire _12143_;
  wire _12144_;
  wire _12145_;
  wire _12146_;
  wire _12147_;
  wire _12148_;
  wire _12149_;
  wire _12150_;
  wire _12151_;
  wire _12152_;
  wire _12153_;
  wire _12154_;
  wire _12155_;
  wire _12156_;
  wire _12157_;
  wire _12158_;
  wire _12159_;
  wire _12160_;
  wire _12161_;
  wire _12162_;
  wire _12163_;
  wire _12164_;
  wire _12165_;
  wire _12166_;
  wire _12167_;
  wire _12168_;
  wire _12169_;
  wire _12170_;
  wire _12171_;
  wire _12172_;
  wire _12173_;
  wire _12174_;
  wire _12175_;
  wire _12176_;
  wire _12177_;
  wire _12178_;
  wire _12179_;
  wire _12180_;
  wire _12181_;
  wire _12182_;
  wire _12183_;
  wire _12184_;
  wire _12185_;
  wire _12186_;
  wire _12187_;
  wire _12188_;
  wire _12189_;
  wire _12190_;
  wire _12191_;
  wire _12192_;
  wire _12193_;
  wire _12194_;
  wire _12195_;
  wire _12196_;
  wire _12197_;
  wire _12198_;
  wire _12199_;
  wire _12200_;
  wire _12201_;
  wire _12202_;
  wire _12203_;
  wire _12204_;
  wire _12205_;
  wire _12206_;
  wire _12207_;
  wire _12208_;
  wire _12209_;
  wire _12210_;
  wire _12211_;
  wire _12212_;
  wire _12213_;
  wire _12214_;
  wire _12215_;
  wire _12216_;
  wire _12217_;
  wire _12218_;
  wire _12219_;
  wire _12220_;
  wire _12221_;
  wire _12222_;
  wire _12223_;
  wire _12224_;
  wire _12225_;
  wire _12226_;
  wire _12227_;
  wire _12228_;
  wire _12229_;
  wire _12230_;
  wire _12231_;
  wire _12232_;
  wire _12233_;
  wire _12234_;
  wire _12235_;
  wire _12236_;
  wire _12237_;
  wire _12238_;
  wire _12239_;
  wire _12240_;
  wire _12241_;
  wire _12242_;
  wire _12243_;
  wire _12244_;
  wire _12245_;
  wire _12246_;
  wire _12247_;
  wire _12248_;
  wire _12249_;
  wire _12250_;
  wire _12251_;
  wire _12252_;
  wire _12253_;
  wire _12254_;
  wire _12255_;
  wire _12256_;
  wire _12257_;
  wire _12258_;
  wire _12259_;
  wire _12260_;
  wire _12261_;
  wire _12262_;
  wire _12263_;
  wire _12264_;
  wire _12265_;
  wire _12266_;
  wire _12267_;
  wire _12268_;
  wire _12269_;
  wire _12270_;
  wire _12271_;
  wire _12272_;
  wire _12273_;
  wire _12274_;
  wire _12275_;
  wire _12276_;
  wire _12277_;
  wire _12278_;
  wire _12279_;
  wire _12280_;
  wire _12281_;
  wire _12282_;
  wire _12283_;
  wire _12284_;
  wire _12285_;
  wire _12286_;
  wire _12287_;
  wire _12288_;
  wire _12289_;
  wire _12290_;
  wire _12291_;
  wire _12292_;
  wire _12293_;
  wire _12294_;
  wire _12295_;
  wire _12296_;
  wire _12297_;
  wire _12298_;
  wire _12299_;
  wire _12300_;
  wire _12301_;
  wire _12302_;
  wire _12303_;
  wire _12304_;
  wire _12305_;
  wire _12306_;
  wire _12307_;
  wire _12308_;
  wire _12309_;
  wire _12310_;
  wire _12311_;
  wire _12312_;
  wire _12313_;
  wire _12314_;
  wire _12315_;
  wire _12316_;
  wire _12317_;
  wire _12318_;
  wire _12319_;
  wire _12320_;
  wire _12321_;
  wire _12322_;
  wire _12323_;
  wire _12324_;
  wire _12325_;
  wire _12326_;
  wire _12327_;
  wire _12328_;
  wire _12329_;
  wire _12330_;
  wire _12331_;
  wire _12332_;
  wire _12333_;
  wire _12334_;
  wire _12335_;
  wire _12336_;
  wire _12337_;
  wire _12338_;
  wire _12339_;
  wire _12340_;
  wire _12341_;
  wire _12342_;
  wire _12343_;
  wire _12344_;
  wire _12345_;
  wire _12346_;
  wire _12347_;
  wire _12348_;
  wire _12349_;
  wire _12350_;
  wire _12351_;
  wire _12352_;
  wire _12353_;
  wire _12354_;
  wire _12355_;
  wire _12356_;
  wire _12357_;
  wire _12358_;
  wire _12359_;
  wire _12360_;
  wire _12361_;
  wire _12362_;
  wire _12363_;
  wire _12364_;
  wire _12365_;
  wire _12366_;
  wire _12367_;
  wire _12368_;
  wire _12369_;
  wire _12370_;
  wire _12371_;
  wire _12372_;
  wire _12373_;
  wire _12374_;
  wire _12375_;
  wire _12376_;
  wire _12377_;
  wire _12378_;
  wire _12379_;
  wire _12380_;
  wire _12381_;
  wire _12382_;
  wire _12383_;
  wire _12384_;
  wire _12385_;
  wire _12386_;
  wire _12387_;
  wire _12388_;
  wire _12389_;
  wire _12390_;
  wire _12391_;
  wire _12392_;
  wire _12393_;
  wire _12394_;
  wire _12395_;
  wire _12396_;
  wire _12397_;
  wire _12398_;
  wire _12399_;
  wire _12400_;
  wire _12401_;
  wire _12402_;
  wire _12403_;
  wire _12404_;
  wire _12405_;
  wire _12406_;
  wire _12407_;
  wire _12408_;
  wire _12409_;
  wire _12410_;
  wire _12411_;
  wire _12412_;
  wire _12413_;
  wire _12414_;
  wire _12415_;
  wire _12416_;
  wire _12417_;
  wire _12418_;
  wire _12419_;
  wire _12420_;
  wire _12421_;
  wire _12422_;
  wire _12423_;
  wire _12424_;
  wire _12425_;
  wire _12426_;
  wire _12427_;
  wire _12428_;
  wire _12429_;
  wire _12430_;
  wire _12431_;
  wire _12432_;
  wire _12433_;
  wire _12434_;
  wire _12435_;
  wire _12436_;
  wire _12437_;
  wire _12438_;
  wire _12439_;
  wire _12440_;
  wire _12441_;
  wire _12442_;
  wire _12443_;
  wire _12444_;
  wire _12445_;
  wire _12446_;
  wire _12447_;
  wire _12448_;
  wire _12449_;
  wire _12450_;
  wire _12451_;
  wire _12452_;
  wire _12453_;
  wire _12454_;
  wire _12455_;
  wire _12456_;
  wire _12457_;
  wire _12458_;
  wire _12459_;
  wire _12460_;
  wire _12461_;
  wire _12462_;
  wire _12463_;
  wire _12464_;
  wire _12465_;
  wire _12466_;
  wire _12467_;
  wire _12468_;
  wire _12469_;
  wire _12470_;
  wire _12471_;
  wire _12472_;
  wire _12473_;
  wire _12474_;
  wire _12475_;
  wire _12476_;
  wire _12477_;
  wire _12478_;
  wire _12479_;
  wire _12480_;
  wire _12481_;
  wire _12482_;
  wire _12483_;
  wire _12484_;
  wire _12485_;
  wire _12486_;
  wire _12487_;
  wire _12488_;
  wire _12489_;
  wire _12490_;
  wire _12491_;
  wire _12492_;
  wire _12493_;
  wire _12494_;
  wire _12495_;
  wire _12496_;
  wire _12497_;
  wire _12498_;
  wire _12499_;
  wire _12500_;
  wire _12501_;
  wire _12502_;
  wire _12503_;
  wire _12504_;
  wire _12505_;
  wire _12506_;
  wire _12507_;
  wire _12508_;
  wire _12509_;
  wire _12510_;
  wire _12511_;
  wire _12512_;
  wire _12513_;
  wire _12514_;
  wire _12515_;
  wire _12516_;
  wire _12517_;
  wire _12518_;
  wire _12519_;
  wire _12520_;
  wire _12521_;
  wire _12522_;
  wire _12523_;
  wire _12524_;
  wire _12525_;
  wire _12526_;
  wire _12527_;
  wire _12528_;
  wire _12529_;
  wire _12530_;
  wire _12531_;
  wire _12532_;
  wire _12533_;
  wire _12534_;
  wire _12535_;
  wire _12536_;
  wire _12537_;
  wire _12538_;
  wire _12539_;
  wire _12540_;
  wire _12541_;
  wire _12542_;
  wire _12543_;
  wire _12544_;
  wire _12545_;
  wire _12546_;
  wire _12547_;
  wire _12548_;
  wire _12549_;
  wire _12550_;
  wire _12551_;
  wire _12552_;
  wire _12553_;
  wire _12554_;
  wire _12555_;
  wire _12556_;
  wire _12557_;
  wire _12558_;
  wire _12559_;
  wire _12560_;
  wire _12561_;
  wire _12562_;
  wire _12563_;
  wire _12564_;
  wire _12565_;
  wire _12566_;
  wire _12567_;
  wire _12568_;
  wire _12569_;
  wire _12570_;
  wire _12571_;
  wire _12572_;
  wire _12573_;
  wire _12574_;
  wire _12575_;
  wire _12576_;
  wire _12577_;
  wire _12578_;
  wire _12579_;
  wire _12580_;
  wire _12581_;
  wire _12582_;
  wire _12583_;
  wire _12584_;
  wire _12585_;
  wire _12586_;
  wire _12587_;
  wire _12588_;
  wire _12589_;
  wire _12590_;
  wire _12591_;
  wire _12592_;
  wire _12593_;
  wire _12594_;
  wire _12595_;
  wire _12596_;
  wire _12597_;
  wire _12598_;
  wire _12599_;
  wire _12600_;
  wire _12601_;
  wire _12602_;
  wire _12603_;
  wire _12604_;
  wire _12605_;
  wire _12606_;
  wire _12607_;
  wire _12608_;
  wire _12609_;
  wire _12610_;
  wire _12611_;
  wire _12612_;
  wire _12613_;
  wire _12614_;
  wire _12615_;
  wire _12616_;
  wire _12617_;
  wire _12618_;
  wire _12619_;
  wire _12620_;
  wire _12621_;
  wire _12622_;
  wire _12623_;
  wire _12624_;
  wire _12625_;
  wire _12626_;
  wire _12627_;
  wire _12628_;
  wire _12629_;
  wire _12630_;
  wire _12631_;
  wire _12632_;
  wire _12633_;
  wire _12634_;
  wire _12635_;
  wire _12636_;
  wire _12637_;
  wire _12638_;
  wire _12639_;
  wire _12640_;
  wire _12641_;
  wire _12642_;
  wire _12643_;
  wire _12644_;
  wire _12645_;
  wire _12646_;
  wire _12647_;
  wire _12648_;
  wire _12649_;
  wire _12650_;
  wire _12651_;
  wire _12652_;
  wire _12653_;
  wire _12654_;
  wire _12655_;
  wire _12656_;
  wire _12657_;
  wire _12658_;
  wire _12659_;
  wire _12660_;
  wire _12661_;
  wire _12662_;
  wire _12663_;
  wire _12664_;
  wire _12665_;
  wire _12666_;
  wire _12667_;
  wire _12668_;
  wire _12669_;
  wire _12670_;
  wire _12671_;
  wire _12672_;
  wire _12673_;
  wire _12674_;
  wire _12675_;
  wire _12676_;
  wire _12677_;
  wire _12678_;
  wire _12679_;
  wire _12680_;
  wire _12681_;
  wire _12682_;
  wire _12683_;
  wire _12684_;
  wire _12685_;
  wire _12686_;
  wire _12687_;
  wire _12688_;
  wire _12689_;
  wire _12690_;
  wire _12691_;
  wire _12692_;
  wire _12693_;
  wire _12694_;
  wire _12695_;
  wire _12696_;
  wire _12697_;
  wire _12698_;
  wire _12699_;
  wire _12700_;
  wire _12701_;
  wire _12702_;
  wire _12703_;
  wire _12704_;
  wire _12705_;
  wire _12706_;
  wire _12707_;
  wire _12708_;
  wire _12709_;
  wire _12710_;
  wire _12711_;
  wire _12712_;
  wire _12713_;
  wire _12714_;
  wire _12715_;
  wire _12716_;
  wire _12717_;
  wire _12718_;
  wire _12719_;
  wire _12720_;
  wire _12721_;
  wire _12722_;
  wire _12723_;
  wire _12724_;
  wire _12725_;
  wire _12726_;
  wire _12727_;
  wire _12728_;
  wire _12729_;
  wire _12730_;
  wire _12731_;
  wire _12732_;
  wire _12733_;
  wire _12734_;
  wire _12735_;
  wire _12736_;
  wire _12737_;
  wire _12738_;
  wire _12739_;
  wire _12740_;
  wire _12741_;
  wire _12742_;
  wire _12743_;
  wire _12744_;
  wire _12745_;
  wire _12746_;
  wire _12747_;
  wire _12748_;
  wire _12749_;
  wire _12750_;
  wire _12751_;
  wire _12752_;
  wire _12753_;
  wire _12754_;
  wire _12755_;
  wire _12756_;
  wire _12757_;
  wire _12758_;
  wire _12759_;
  wire _12760_;
  wire _12761_;
  wire _12762_;
  wire _12763_;
  wire _12764_;
  wire _12765_;
  wire _12766_;
  wire _12767_;
  wire _12768_;
  wire _12769_;
  wire _12770_;
  wire _12771_;
  wire _12772_;
  wire _12773_;
  wire _12774_;
  wire _12775_;
  wire _12776_;
  wire _12777_;
  wire _12778_;
  wire _12779_;
  wire _12780_;
  wire _12781_;
  wire _12782_;
  wire _12783_;
  wire _12784_;
  wire _12785_;
  wire _12786_;
  wire _12787_;
  wire _12788_;
  wire _12789_;
  wire _12790_;
  wire _12791_;
  wire _12792_;
  wire _12793_;
  wire _12794_;
  wire _12795_;
  wire _12796_;
  wire _12797_;
  wire _12798_;
  wire _12799_;
  wire _12800_;
  wire _12801_;
  wire _12802_;
  wire _12803_;
  wire _12804_;
  wire _12805_;
  wire _12806_;
  wire _12807_;
  wire _12808_;
  wire _12809_;
  wire _12810_;
  wire _12811_;
  wire _12812_;
  wire _12813_;
  wire _12814_;
  wire _12815_;
  wire _12816_;
  wire _12817_;
  wire _12818_;
  wire _12819_;
  wire _12820_;
  wire _12821_;
  wire _12822_;
  wire _12823_;
  wire _12824_;
  wire _12825_;
  wire _12826_;
  wire _12827_;
  wire _12828_;
  wire _12829_;
  wire _12830_;
  wire _12831_;
  wire _12832_;
  wire _12833_;
  wire _12834_;
  wire _12835_;
  wire _12836_;
  wire _12837_;
  wire _12838_;
  wire _12839_;
  wire _12840_;
  wire _12841_;
  wire _12842_;
  wire _12843_;
  wire _12844_;
  wire _12845_;
  wire _12846_;
  wire _12847_;
  wire _12848_;
  wire _12849_;
  wire _12850_;
  wire _12851_;
  wire _12852_;
  wire _12853_;
  wire _12854_;
  wire _12855_;
  wire _12856_;
  wire _12857_;
  wire _12858_;
  wire _12859_;
  wire _12860_;
  wire _12861_;
  wire _12862_;
  wire _12863_;
  wire _12864_;
  wire _12865_;
  wire _12866_;
  wire _12867_;
  wire _12868_;
  wire _12869_;
  wire _12870_;
  wire _12871_;
  wire _12872_;
  wire _12873_;
  wire _12874_;
  wire _12875_;
  wire _12876_;
  wire _12877_;
  wire _12878_;
  wire _12879_;
  wire _12880_;
  wire _12881_;
  wire _12882_;
  wire _12883_;
  wire _12884_;
  wire _12885_;
  wire _12886_;
  wire _12887_;
  wire _12888_;
  wire _12889_;
  wire _12890_;
  wire _12891_;
  wire _12892_;
  wire _12893_;
  wire _12894_;
  wire _12895_;
  wire _12896_;
  wire _12897_;
  wire _12898_;
  wire _12899_;
  wire _12900_;
  wire _12901_;
  wire _12902_;
  wire _12903_;
  wire _12904_;
  wire _12905_;
  wire _12906_;
  wire _12907_;
  wire _12908_;
  wire _12909_;
  wire _12910_;
  wire _12911_;
  wire _12912_;
  wire _12913_;
  wire _12914_;
  wire _12915_;
  wire _12916_;
  wire _12917_;
  wire _12918_;
  wire _12919_;
  wire _12920_;
  wire _12921_;
  wire _12922_;
  wire _12923_;
  wire _12924_;
  wire _12925_;
  wire _12926_;
  wire _12927_;
  wire _12928_;
  wire _12929_;
  wire _12930_;
  wire _12931_;
  wire _12932_;
  wire _12933_;
  wire _12934_;
  wire _12935_;
  wire _12936_;
  wire _12937_;
  wire _12938_;
  wire _12939_;
  wire _12940_;
  wire _12941_;
  wire _12942_;
  wire _12943_;
  wire _12944_;
  wire _12945_;
  wire _12946_;
  wire _12947_;
  wire _12948_;
  wire _12949_;
  wire _12950_;
  wire _12951_;
  wire _12952_;
  wire _12953_;
  wire _12954_;
  wire _12955_;
  wire _12956_;
  wire _12957_;
  wire _12958_;
  wire _12959_;
  wire _12960_;
  wire _12961_;
  wire _12962_;
  wire _12963_;
  wire _12964_;
  wire _12965_;
  wire _12966_;
  wire _12967_;
  wire _12968_;
  wire _12969_;
  wire _12970_;
  wire _12971_;
  wire _12972_;
  wire _12973_;
  wire _12974_;
  wire _12975_;
  wire _12976_;
  wire _12977_;
  wire _12978_;
  wire _12979_;
  wire _12980_;
  wire _12981_;
  wire _12982_;
  wire _12983_;
  wire _12984_;
  wire _12985_;
  wire _12986_;
  wire _12987_;
  wire _12988_;
  wire _12989_;
  wire _12990_;
  wire _12991_;
  wire _12992_;
  wire _12993_;
  wire _12994_;
  wire _12995_;
  wire _12996_;
  wire _12997_;
  wire _12998_;
  wire _12999_;
  wire _13000_;
  wire _13001_;
  wire _13002_;
  wire _13003_;
  wire _13004_;
  wire _13005_;
  wire _13006_;
  wire _13007_;
  wire _13008_;
  wire _13009_;
  wire _13010_;
  wire _13011_;
  wire _13012_;
  wire _13013_;
  wire _13014_;
  wire _13015_;
  wire _13016_;
  wire _13017_;
  wire _13018_;
  wire _13019_;
  wire _13020_;
  wire _13021_;
  wire _13022_;
  wire _13023_;
  wire _13024_;
  wire _13025_;
  wire _13026_;
  wire _13027_;
  wire _13028_;
  wire _13029_;
  wire _13030_;
  wire _13031_;
  wire _13032_;
  wire _13033_;
  wire _13034_;
  wire _13035_;
  wire _13036_;
  wire _13037_;
  wire _13038_;
  wire _13039_;
  wire _13040_;
  wire _13041_;
  wire _13042_;
  wire _13043_;
  wire _13044_;
  wire _13045_;
  wire _13046_;
  wire _13047_;
  wire _13048_;
  wire _13049_;
  wire _13050_;
  wire _13051_;
  wire _13052_;
  wire _13053_;
  wire _13054_;
  wire _13055_;
  wire _13056_;
  wire _13057_;
  wire _13058_;
  wire _13059_;
  wire _13060_;
  wire _13061_;
  wire _13062_;
  wire _13063_;
  wire _13064_;
  wire _13065_;
  wire _13066_;
  wire _13067_;
  wire _13068_;
  wire _13069_;
  wire _13070_;
  wire _13071_;
  wire _13072_;
  wire _13073_;
  wire _13074_;
  wire _13075_;
  wire _13076_;
  wire _13077_;
  wire _13078_;
  wire _13079_;
  wire _13080_;
  wire _13081_;
  wire _13082_;
  wire _13083_;
  wire _13084_;
  wire _13085_;
  wire _13086_;
  wire _13087_;
  wire _13088_;
  wire _13089_;
  wire _13090_;
  wire _13091_;
  wire _13092_;
  wire _13093_;
  wire _13094_;
  wire _13095_;
  wire _13096_;
  wire _13097_;
  wire _13098_;
  wire _13099_;
  wire _13100_;
  wire _13101_;
  wire _13102_;
  wire _13103_;
  wire _13104_;
  wire _13105_;
  wire _13106_;
  wire _13107_;
  wire _13108_;
  wire _13109_;
  wire _13110_;
  wire _13111_;
  wire _13112_;
  wire _13113_;
  wire _13114_;
  wire _13115_;
  wire _13116_;
  wire _13117_;
  wire _13118_;
  wire _13119_;
  wire _13120_;
  wire _13121_;
  wire _13122_;
  wire _13123_;
  wire _13124_;
  wire _13125_;
  wire _13126_;
  wire _13127_;
  wire _13128_;
  wire _13129_;
  wire _13130_;
  wire _13131_;
  wire _13132_;
  wire _13133_;
  wire _13134_;
  wire _13135_;
  wire _13136_;
  wire _13137_;
  wire _13138_;
  wire _13139_;
  wire _13140_;
  wire _13141_;
  wire _13142_;
  wire _13143_;
  wire _13144_;
  wire _13145_;
  wire _13146_;
  wire _13147_;
  wire _13148_;
  wire _13149_;
  wire _13150_;
  wire _13151_;
  wire _13152_;
  wire _13153_;
  wire _13154_;
  wire _13155_;
  wire _13156_;
  wire _13157_;
  wire _13158_;
  wire _13159_;
  wire _13160_;
  wire _13161_;
  wire _13162_;
  wire _13163_;
  wire _13164_;
  wire _13165_;
  wire _13166_;
  wire _13167_;
  wire _13168_;
  wire _13169_;
  wire _13170_;
  wire _13171_;
  wire _13172_;
  wire _13173_;
  wire _13174_;
  wire _13175_;
  wire _13176_;
  wire _13177_;
  wire _13178_;
  wire _13179_;
  wire _13180_;
  wire _13181_;
  wire _13182_;
  wire _13183_;
  wire _13184_;
  wire _13185_;
  wire _13186_;
  wire _13187_;
  wire _13188_;
  wire _13189_;
  wire _13190_;
  wire _13191_;
  wire _13192_;
  wire _13193_;
  wire _13194_;
  wire _13195_;
  wire _13196_;
  wire _13197_;
  wire _13198_;
  wire _13199_;
  wire _13200_;
  wire _13201_;
  wire _13202_;
  wire _13203_;
  wire _13204_;
  wire _13205_;
  wire _13206_;
  wire _13207_;
  wire _13208_;
  wire _13209_;
  wire _13210_;
  wire _13211_;
  wire _13212_;
  wire _13213_;
  wire _13214_;
  wire _13215_;
  wire _13216_;
  wire _13217_;
  wire _13218_;
  wire _13219_;
  wire _13220_;
  wire _13221_;
  wire _13222_;
  wire _13223_;
  wire _13224_;
  wire _13225_;
  wire _13226_;
  wire _13227_;
  wire _13228_;
  wire _13229_;
  wire _13230_;
  wire _13231_;
  wire _13232_;
  wire _13233_;
  wire _13234_;
  wire _13235_;
  wire _13236_;
  wire _13237_;
  wire _13238_;
  wire _13239_;
  wire _13240_;
  wire _13241_;
  wire _13242_;
  wire _13243_;
  wire _13244_;
  wire _13245_;
  wire _13246_;
  wire _13247_;
  wire _13248_;
  wire _13249_;
  wire _13250_;
  wire _13251_;
  wire _13252_;
  wire _13253_;
  wire _13254_;
  wire _13255_;
  wire _13256_;
  wire _13257_;
  wire _13258_;
  wire _13259_;
  wire _13260_;
  wire _13261_;
  wire _13262_;
  wire _13263_;
  wire _13264_;
  wire _13265_;
  wire _13266_;
  wire _13267_;
  wire _13268_;
  wire _13269_;
  wire _13270_;
  wire _13271_;
  wire _13272_;
  wire _13273_;
  wire _13274_;
  wire _13275_;
  wire _13276_;
  wire _13277_;
  wire _13278_;
  wire _13279_;
  wire _13280_;
  wire _13281_;
  wire _13282_;
  wire _13283_;
  wire _13284_;
  wire _13285_;
  wire _13286_;
  wire _13287_;
  wire _13288_;
  wire _13289_;
  wire _13290_;
  wire _13291_;
  wire _13292_;
  wire _13293_;
  wire _13294_;
  wire _13295_;
  wire _13296_;
  wire _13297_;
  wire _13298_;
  wire _13299_;
  wire _13300_;
  wire _13301_;
  wire _13302_;
  wire _13303_;
  wire _13304_;
  wire _13305_;
  wire _13306_;
  wire _13307_;
  wire _13308_;
  wire _13309_;
  wire _13310_;
  wire _13311_;
  wire _13312_;
  wire _13313_;
  wire _13314_;
  wire _13315_;
  wire _13316_;
  wire _13317_;
  wire _13318_;
  wire _13319_;
  wire _13320_;
  wire _13321_;
  wire _13322_;
  wire _13323_;
  wire _13324_;
  wire _13325_;
  wire _13326_;
  wire _13327_;
  wire _13328_;
  wire _13329_;
  wire _13330_;
  wire _13331_;
  wire _13332_;
  wire _13333_;
  wire _13334_;
  wire _13335_;
  wire _13336_;
  wire _13337_;
  wire _13338_;
  wire _13339_;
  wire _13340_;
  wire _13341_;
  wire _13342_;
  wire _13343_;
  wire _13344_;
  wire _13345_;
  wire _13346_;
  wire _13347_;
  wire _13348_;
  wire _13349_;
  wire _13350_;
  wire _13351_;
  wire _13352_;
  wire _13353_;
  wire _13354_;
  wire _13355_;
  wire _13356_;
  wire _13357_;
  wire _13358_;
  wire _13359_;
  wire _13360_;
  wire _13361_;
  wire _13362_;
  wire _13363_;
  wire _13364_;
  wire _13365_;
  wire _13366_;
  wire _13367_;
  wire _13368_;
  wire _13369_;
  wire _13370_;
  wire _13371_;
  wire _13372_;
  wire _13373_;
  wire _13374_;
  wire _13375_;
  wire _13376_;
  wire _13377_;
  wire _13378_;
  wire _13379_;
  wire _13380_;
  wire _13381_;
  wire _13382_;
  wire _13383_;
  wire _13384_;
  wire _13385_;
  wire _13386_;
  wire _13387_;
  wire _13388_;
  wire _13389_;
  wire _13390_;
  wire _13391_;
  wire _13392_;
  wire _13393_;
  wire _13394_;
  wire _13395_;
  wire _13396_;
  wire _13397_;
  wire _13398_;
  wire _13399_;
  wire _13400_;
  wire _13401_;
  wire _13402_;
  wire _13403_;
  wire _13404_;
  wire _13405_;
  wire _13406_;
  wire _13407_;
  wire _13408_;
  wire _13409_;
  wire _13410_;
  wire _13411_;
  wire _13412_;
  wire _13413_;
  wire _13414_;
  wire _13415_;
  wire _13416_;
  wire _13417_;
  wire _13418_;
  wire _13419_;
  wire _13420_;
  wire _13421_;
  wire _13422_;
  wire _13423_;
  wire _13424_;
  wire _13425_;
  wire _13426_;
  wire _13427_;
  wire _13428_;
  wire _13429_;
  wire _13430_;
  wire _13431_;
  wire _13432_;
  wire _13433_;
  wire _13434_;
  wire _13435_;
  wire _13436_;
  wire _13437_;
  wire _13438_;
  wire _13439_;
  wire _13440_;
  wire _13441_;
  wire _13442_;
  wire _13443_;
  wire _13444_;
  wire _13445_;
  wire _13446_;
  wire _13447_;
  wire _13448_;
  wire _13449_;
  wire _13450_;
  wire _13451_;
  wire _13452_;
  wire _13453_;
  wire _13454_;
  wire _13455_;
  wire _13456_;
  wire _13457_;
  wire _13458_;
  wire _13459_;
  wire _13460_;
  wire _13461_;
  wire _13462_;
  wire _13463_;
  wire _13464_;
  wire _13465_;
  wire _13466_;
  wire _13467_;
  wire _13468_;
  wire _13469_;
  wire _13470_;
  wire _13471_;
  wire _13472_;
  wire _13473_;
  wire _13474_;
  wire _13475_;
  wire _13476_;
  wire _13477_;
  wire _13478_;
  wire _13479_;
  wire _13480_;
  wire _13481_;
  wire _13482_;
  wire _13483_;
  wire _13484_;
  wire _13485_;
  wire _13486_;
  wire _13487_;
  wire _13488_;
  wire _13489_;
  wire _13490_;
  wire _13491_;
  wire _13492_;
  wire _13493_;
  wire _13494_;
  wire _13495_;
  wire _13496_;
  wire _13497_;
  wire _13498_;
  wire _13499_;
  wire _13500_;
  wire _13501_;
  wire _13502_;
  wire _13503_;
  wire _13504_;
  wire _13505_;
  wire _13506_;
  wire _13507_;
  wire _13508_;
  wire _13509_;
  wire _13510_;
  wire _13511_;
  wire _13512_;
  wire _13513_;
  wire _13514_;
  wire _13515_;
  wire _13516_;
  wire _13517_;
  wire _13518_;
  wire _13519_;
  wire _13520_;
  wire _13521_;
  wire _13522_;
  wire _13523_;
  wire _13524_;
  wire _13525_;
  wire _13526_;
  wire _13527_;
  wire _13528_;
  wire _13529_;
  wire _13530_;
  wire _13531_;
  wire _13532_;
  wire _13533_;
  wire _13534_;
  wire _13535_;
  wire _13536_;
  wire _13537_;
  wire _13538_;
  wire _13539_;
  wire _13540_;
  wire _13541_;
  wire _13542_;
  wire _13543_;
  wire _13544_;
  wire _13545_;
  wire _13546_;
  wire _13547_;
  wire _13548_;
  wire _13549_;
  wire _13550_;
  wire _13551_;
  wire _13552_;
  wire _13553_;
  wire _13554_;
  wire _13555_;
  wire _13556_;
  wire _13557_;
  wire _13558_;
  wire _13559_;
  wire _13560_;
  wire _13561_;
  wire _13562_;
  wire _13563_;
  wire _13564_;
  wire _13565_;
  wire _13566_;
  wire _13567_;
  wire _13568_;
  wire _13569_;
  wire _13570_;
  wire _13571_;
  wire _13572_;
  wire _13573_;
  wire _13574_;
  wire _13575_;
  wire _13576_;
  wire _13577_;
  wire _13578_;
  wire _13579_;
  wire _13580_;
  wire _13581_;
  wire _13582_;
  wire _13583_;
  wire _13584_;
  wire _13585_;
  wire _13586_;
  wire _13587_;
  wire _13588_;
  wire _13589_;
  wire _13590_;
  wire _13591_;
  wire _13592_;
  wire _13593_;
  wire _13594_;
  wire _13595_;
  wire _13596_;
  wire _13597_;
  wire _13598_;
  wire _13599_;
  wire _13600_;
  wire _13601_;
  wire _13602_;
  wire _13603_;
  wire _13604_;
  wire _13605_;
  wire _13606_;
  wire _13607_;
  wire _13608_;
  wire _13609_;
  wire _13610_;
  wire _13611_;
  wire _13612_;
  wire _13613_;
  wire _13614_;
  wire _13615_;
  wire _13616_;
  wire _13617_;
  wire _13618_;
  wire _13619_;
  wire _13620_;
  wire _13621_;
  wire _13622_;
  wire _13623_;
  wire _13624_;
  wire _13625_;
  wire _13626_;
  wire _13627_;
  wire _13628_;
  wire _13629_;
  wire _13630_;
  wire _13631_;
  wire _13632_;
  wire _13633_;
  wire _13634_;
  wire _13635_;
  wire _13636_;
  wire _13637_;
  wire _13638_;
  wire _13639_;
  wire _13640_;
  wire _13641_;
  wire _13642_;
  wire _13643_;
  wire _13644_;
  wire _13645_;
  wire _13646_;
  wire _13647_;
  wire _13648_;
  wire _13649_;
  wire _13650_;
  wire _13651_;
  wire _13652_;
  wire _13653_;
  wire _13654_;
  wire _13655_;
  wire _13656_;
  wire _13657_;
  wire _13658_;
  wire _13659_;
  wire _13660_;
  wire _13661_;
  wire _13662_;
  wire _13663_;
  wire _13664_;
  wire _13665_;
  wire _13666_;
  wire _13667_;
  wire _13668_;
  wire _13669_;
  wire _13670_;
  wire _13671_;
  wire _13672_;
  wire _13673_;
  wire _13674_;
  wire _13675_;
  wire _13676_;
  wire _13677_;
  wire _13678_;
  wire _13679_;
  wire _13680_;
  wire _13681_;
  wire _13682_;
  wire _13683_;
  wire _13684_;
  wire _13685_;
  wire _13686_;
  wire _13687_;
  wire _13688_;
  wire _13689_;
  wire _13690_;
  wire _13691_;
  wire _13692_;
  wire _13693_;
  wire _13694_;
  wire _13695_;
  wire _13696_;
  wire _13697_;
  wire _13698_;
  wire _13699_;
  wire _13700_;
  wire _13701_;
  wire _13702_;
  wire _13703_;
  wire _13704_;
  wire _13705_;
  wire _13706_;
  wire _13707_;
  wire _13708_;
  wire _13709_;
  wire _13710_;
  wire _13711_;
  wire _13712_;
  wire _13713_;
  wire _13714_;
  wire _13715_;
  wire _13716_;
  wire _13717_;
  wire _13718_;
  wire _13719_;
  wire _13720_;
  wire _13721_;
  wire _13722_;
  wire _13723_;
  wire _13724_;
  wire _13725_;
  wire _13726_;
  wire _13727_;
  wire _13728_;
  wire _13729_;
  wire _13730_;
  wire _13731_;
  wire _13732_;
  wire _13733_;
  wire _13734_;
  wire _13735_;
  wire _13736_;
  wire _13737_;
  wire _13738_;
  wire _13739_;
  wire _13740_;
  wire _13741_;
  wire _13742_;
  wire _13743_;
  wire _13744_;
  wire _13745_;
  wire _13746_;
  wire _13747_;
  wire _13748_;
  wire _13749_;
  wire _13750_;
  wire _13751_;
  wire _13752_;
  wire _13753_;
  wire _13754_;
  wire _13755_;
  wire _13756_;
  wire _13757_;
  wire _13758_;
  wire _13759_;
  wire _13760_;
  wire _13761_;
  wire _13762_;
  wire _13763_;
  wire _13764_;
  wire _13765_;
  wire _13766_;
  wire _13767_;
  wire _13768_;
  wire _13769_;
  wire _13770_;
  wire _13771_;
  wire _13772_;
  wire _13773_;
  wire _13774_;
  wire _13775_;
  wire _13776_;
  wire _13777_;
  wire _13778_;
  wire _13779_;
  wire _13780_;
  wire _13781_;
  wire _13782_;
  wire _13783_;
  wire _13784_;
  wire _13785_;
  wire _13786_;
  wire _13787_;
  wire _13788_;
  wire _13789_;
  wire _13790_;
  wire _13791_;
  wire _13792_;
  wire _13793_;
  wire _13794_;
  wire _13795_;
  wire _13796_;
  wire _13797_;
  wire _13798_;
  wire _13799_;
  wire _13800_;
  wire _13801_;
  wire _13802_;
  wire _13803_;
  wire _13804_;
  wire _13805_;
  wire _13806_;
  wire _13807_;
  wire _13808_;
  wire _13809_;
  wire _13810_;
  wire _13811_;
  wire _13812_;
  wire _13813_;
  wire _13814_;
  wire _13815_;
  wire _13816_;
  wire _13817_;
  wire _13818_;
  wire _13819_;
  wire _13820_;
  wire _13821_;
  wire _13822_;
  wire _13823_;
  wire _13824_;
  wire _13825_;
  wire _13826_;
  wire _13827_;
  wire _13828_;
  wire _13829_;
  wire _13830_;
  wire _13831_;
  wire _13832_;
  wire _13833_;
  wire _13834_;
  wire _13835_;
  wire _13836_;
  wire _13837_;
  wire _13838_;
  wire _13839_;
  wire _13840_;
  wire _13841_;
  wire _13842_;
  wire _13843_;
  wire _13844_;
  wire _13845_;
  wire _13846_;
  wire _13847_;
  wire _13848_;
  wire _13849_;
  wire _13850_;
  wire _13851_;
  wire _13852_;
  wire _13853_;
  wire _13854_;
  wire _13855_;
  wire _13856_;
  wire _13857_;
  wire _13858_;
  wire _13859_;
  wire _13860_;
  wire _13861_;
  wire _13862_;
  wire _13863_;
  wire _13864_;
  wire _13865_;
  wire _13866_;
  wire _13867_;
  wire _13868_;
  wire _13869_;
  wire _13870_;
  wire _13871_;
  wire _13872_;
  wire _13873_;
  wire _13874_;
  wire _13875_;
  wire _13876_;
  wire _13877_;
  wire _13878_;
  wire _13879_;
  wire _13880_;
  wire _13881_;
  wire _13882_;
  wire _13883_;
  wire _13884_;
  wire _13885_;
  wire _13886_;
  wire _13887_;
  wire _13888_;
  wire _13889_;
  wire _13890_;
  wire _13891_;
  wire _13892_;
  wire _13893_;
  wire _13894_;
  wire _13895_;
  wire _13896_;
  wire _13897_;
  wire _13898_;
  wire _13899_;
  wire _13900_;
  wire _13901_;
  wire _13902_;
  wire _13903_;
  wire _13904_;
  wire _13905_;
  wire _13906_;
  wire _13907_;
  wire _13908_;
  wire _13909_;
  wire _13910_;
  wire _13911_;
  wire _13912_;
  wire _13913_;
  wire _13914_;
  wire _13915_;
  wire _13916_;
  wire _13917_;
  wire _13918_;
  wire _13919_;
  wire _13920_;
  wire _13921_;
  wire _13922_;
  wire _13923_;
  wire _13924_;
  wire _13925_;
  wire _13926_;
  wire _13927_;
  wire _13928_;
  wire _13929_;
  wire _13930_;
  wire _13931_;
  wire _13932_;
  wire _13933_;
  wire _13934_;
  wire _13935_;
  wire _13936_;
  wire _13937_;
  wire _13938_;
  wire _13939_;
  wire _13940_;
  wire _13941_;
  wire _13942_;
  wire _13943_;
  wire _13944_;
  wire _13945_;
  wire _13946_;
  wire _13947_;
  wire _13948_;
  wire _13949_;
  wire _13950_;
  wire _13951_;
  wire _13952_;
  wire _13953_;
  wire _13954_;
  wire _13955_;
  wire _13956_;
  wire _13957_;
  wire _13958_;
  wire _13959_;
  wire _13960_;
  wire _13961_;
  wire _13962_;
  wire _13963_;
  wire _13964_;
  wire _13965_;
  wire _13966_;
  wire _13967_;
  wire _13968_;
  wire _13969_;
  wire _13970_;
  wire _13971_;
  wire _13972_;
  wire _13973_;
  wire _13974_;
  wire _13975_;
  wire _13976_;
  wire _13977_;
  wire _13978_;
  wire _13979_;
  wire _13980_;
  wire _13981_;
  wire _13982_;
  wire _13983_;
  wire _13984_;
  wire _13985_;
  wire _13986_;
  wire _13987_;
  wire _13988_;
  wire _13989_;
  wire _13990_;
  wire _13991_;
  wire _13992_;
  wire _13993_;
  wire _13994_;
  wire _13995_;
  wire _13996_;
  wire _13997_;
  wire _13998_;
  wire _13999_;
  wire _14000_;
  wire _14001_;
  wire _14002_;
  wire _14003_;
  wire _14004_;
  wire _14005_;
  wire _14006_;
  wire _14007_;
  wire _14008_;
  wire _14009_;
  wire _14010_;
  wire _14011_;
  wire _14012_;
  wire _14013_;
  wire _14014_;
  wire _14015_;
  wire _14016_;
  wire _14017_;
  wire _14018_;
  wire _14019_;
  wire _14020_;
  wire _14021_;
  wire _14022_;
  wire _14023_;
  wire _14024_;
  wire _14025_;
  wire _14026_;
  wire _14027_;
  wire _14028_;
  wire _14029_;
  wire _14030_;
  wire _14031_;
  wire _14032_;
  wire _14033_;
  wire _14034_;
  wire _14035_;
  wire _14036_;
  wire _14037_;
  wire _14038_;
  wire _14039_;
  wire _14040_;
  wire _14041_;
  wire _14042_;
  wire _14043_;
  wire _14044_;
  wire _14045_;
  wire _14046_;
  wire _14047_;
  wire _14048_;
  wire _14049_;
  wire _14050_;
  wire _14051_;
  wire _14052_;
  wire _14053_;
  wire _14054_;
  wire _14055_;
  wire _14056_;
  wire _14057_;
  wire _14058_;
  wire _14059_;
  wire _14060_;
  wire _14061_;
  wire _14062_;
  wire _14063_;
  wire _14064_;
  wire _14065_;
  wire _14066_;
  wire _14067_;
  wire _14068_;
  wire _14069_;
  wire _14070_;
  wire _14071_;
  wire _14072_;
  wire _14073_;
  wire _14074_;
  wire _14075_;
  wire _14076_;
  wire _14077_;
  wire _14078_;
  wire _14079_;
  wire _14080_;
  wire _14081_;
  wire _14082_;
  wire _14083_;
  wire _14084_;
  wire _14085_;
  wire _14086_;
  wire _14087_;
  wire _14088_;
  wire _14089_;
  wire _14090_;
  wire _14091_;
  wire _14092_;
  wire _14093_;
  wire _14094_;
  wire _14095_;
  wire _14096_;
  wire _14097_;
  wire _14098_;
  wire _14099_;
  wire _14100_;
  wire _14101_;
  wire _14102_;
  wire _14103_;
  wire _14104_;
  wire _14105_;
  wire _14106_;
  wire _14107_;
  wire _14108_;
  wire _14109_;
  wire _14110_;
  wire _14111_;
  wire _14112_;
  wire _14113_;
  wire _14114_;
  wire _14115_;
  wire _14116_;
  wire _14117_;
  wire _14118_;
  wire _14119_;
  wire _14120_;
  wire _14121_;
  wire _14122_;
  wire _14123_;
  wire _14124_;
  wire _14125_;
  wire _14126_;
  wire _14127_;
  wire _14128_;
  wire _14129_;
  wire _14130_;
  wire _14131_;
  wire _14132_;
  wire _14133_;
  wire _14134_;
  wire _14135_;
  wire _14136_;
  wire _14137_;
  wire _14138_;
  wire _14139_;
  wire _14140_;
  wire _14141_;
  wire _14142_;
  wire _14143_;
  wire _14144_;
  wire _14145_;
  wire _14146_;
  wire _14147_;
  wire _14148_;
  wire _14149_;
  wire _14150_;
  wire _14151_;
  wire _14152_;
  wire _14153_;
  wire _14154_;
  wire _14155_;
  wire _14156_;
  wire _14157_;
  wire _14158_;
  wire _14159_;
  wire _14160_;
  wire _14161_;
  wire _14162_;
  wire _14163_;
  wire _14164_;
  wire _14165_;
  wire _14166_;
  wire _14167_;
  wire _14168_;
  wire _14169_;
  wire _14170_;
  wire _14171_;
  wire _14172_;
  wire _14173_;
  wire _14174_;
  wire _14175_;
  wire _14176_;
  wire _14177_;
  wire _14178_;
  wire _14179_;
  wire _14180_;
  wire _14181_;
  wire _14182_;
  wire _14183_;
  wire _14184_;
  wire _14185_;
  wire _14186_;
  wire _14187_;
  wire _14188_;
  wire _14189_;
  wire _14190_;
  wire _14191_;
  wire _14192_;
  wire _14193_;
  wire _14194_;
  wire _14195_;
  wire _14196_;
  wire _14197_;
  wire _14198_;
  wire _14199_;
  wire _14200_;
  wire _14201_;
  wire _14202_;
  wire _14203_;
  wire _14204_;
  wire _14205_;
  wire _14206_;
  wire _14207_;
  wire _14208_;
  wire _14209_;
  wire _14210_;
  wire _14211_;
  wire _14212_;
  wire _14213_;
  wire _14214_;
  wire _14215_;
  wire _14216_;
  wire _14217_;
  wire _14218_;
  wire _14219_;
  wire _14220_;
  wire _14221_;
  wire _14222_;
  wire _14223_;
  wire _14224_;
  wire _14225_;
  wire _14226_;
  wire _14227_;
  wire _14228_;
  wire _14229_;
  wire _14230_;
  wire _14231_;
  wire _14232_;
  wire _14233_;
  wire _14234_;
  wire _14235_;
  wire _14236_;
  wire _14237_;
  wire _14238_;
  wire _14239_;
  wire _14240_;
  wire _14241_;
  wire _14242_;
  wire _14243_;
  wire _14244_;
  wire _14245_;
  wire _14246_;
  wire _14247_;
  wire _14248_;
  wire _14249_;
  wire _14250_;
  wire _14251_;
  wire _14252_;
  wire _14253_;
  wire _14254_;
  wire _14255_;
  wire _14256_;
  wire _14257_;
  wire _14258_;
  wire _14259_;
  wire _14260_;
  wire _14261_;
  wire _14262_;
  wire _14263_;
  wire _14264_;
  wire _14265_;
  wire _14266_;
  wire _14267_;
  wire _14268_;
  wire _14269_;
  wire _14270_;
  wire _14271_;
  wire _14272_;
  wire _14273_;
  wire _14274_;
  wire _14275_;
  wire _14276_;
  wire _14277_;
  wire _14278_;
  wire _14279_;
  wire _14280_;
  wire _14281_;
  wire _14282_;
  wire _14283_;
  wire _14284_;
  wire _14285_;
  wire _14286_;
  wire _14287_;
  wire _14288_;
  wire _14289_;
  wire _14290_;
  wire _14291_;
  wire _14292_;
  wire _14293_;
  wire _14294_;
  wire _14295_;
  wire _14296_;
  wire _14297_;
  wire _14298_;
  wire _14299_;
  wire _14300_;
  wire _14301_;
  wire _14302_;
  wire _14303_;
  wire _14304_;
  wire _14305_;
  wire _14306_;
  wire _14307_;
  wire _14308_;
  wire _14309_;
  wire _14310_;
  wire _14311_;
  wire _14312_;
  wire _14313_;
  wire _14314_;
  wire _14315_;
  wire _14316_;
  wire _14317_;
  wire _14318_;
  wire _14319_;
  wire _14320_;
  wire _14321_;
  wire _14322_;
  wire _14323_;
  wire _14324_;
  wire _14325_;
  wire _14326_;
  wire _14327_;
  wire _14328_;
  wire _14329_;
  wire _14330_;
  wire _14331_;
  wire _14332_;
  wire _14333_;
  wire _14334_;
  wire _14335_;
  wire _14336_;
  wire _14337_;
  wire _14338_;
  wire _14339_;
  wire _14340_;
  wire _14341_;
  wire _14342_;
  wire _14343_;
  wire _14344_;
  wire _14345_;
  wire _14346_;
  wire _14347_;
  wire _14348_;
  wire _14349_;
  wire _14350_;
  wire _14351_;
  wire _14352_;
  wire _14353_;
  wire _14354_;
  wire _14355_;
  wire _14356_;
  wire _14357_;
  wire _14358_;
  wire _14359_;
  wire _14360_;
  wire _14361_;
  wire _14362_;
  wire _14363_;
  wire _14364_;
  wire _14365_;
  wire _14366_;
  wire _14367_;
  wire _14368_;
  wire _14369_;
  wire _14370_;
  wire _14371_;
  wire _14372_;
  wire _14373_;
  wire _14374_;
  wire _14375_;
  wire _14376_;
  wire _14377_;
  wire _14378_;
  wire _14379_;
  wire _14380_;
  wire _14381_;
  wire _14382_;
  wire _14383_;
  wire _14384_;
  wire _14385_;
  wire _14386_;
  wire _14387_;
  wire _14388_;
  wire _14389_;
  wire _14390_;
  wire _14391_;
  wire _14392_;
  wire _14393_;
  wire _14394_;
  wire _14395_;
  wire _14396_;
  wire _14397_;
  wire _14398_;
  wire _14399_;
  wire _14400_;
  wire _14401_;
  wire _14402_;
  wire _14403_;
  wire _14404_;
  wire _14405_;
  wire _14406_;
  wire _14407_;
  wire _14408_;
  wire _14409_;
  wire _14410_;
  wire _14411_;
  wire _14412_;
  wire _14413_;
  wire _14414_;
  wire _14415_;
  wire _14416_;
  wire _14417_;
  wire _14418_;
  wire _14419_;
  wire _14420_;
  wire _14421_;
  wire _14422_;
  wire _14423_;
  wire _14424_;
  wire _14425_;
  wire _14426_;
  wire _14427_;
  wire _14428_;
  wire _14429_;
  wire _14430_;
  wire _14431_;
  wire _14432_;
  wire _14433_;
  wire _14434_;
  wire _14435_;
  wire _14436_;
  wire _14437_;
  wire _14438_;
  wire _14439_;
  wire _14440_;
  wire _14441_;
  wire _14442_;
  wire _14443_;
  wire _14444_;
  wire _14445_;
  wire _14446_;
  wire _14447_;
  wire _14448_;
  wire _14449_;
  wire _14450_;
  wire _14451_;
  wire _14452_;
  wire _14453_;
  wire _14454_;
  wire _14455_;
  wire _14456_;
  wire _14457_;
  wire _14458_;
  wire _14459_;
  wire _14460_;
  wire _14461_;
  wire _14462_;
  wire _14463_;
  wire _14464_;
  wire _14465_;
  wire _14466_;
  wire _14467_;
  wire _14468_;
  wire _14469_;
  wire _14470_;
  wire _14471_;
  wire _14472_;
  wire _14473_;
  wire _14474_;
  wire _14475_;
  wire _14476_;
  wire _14477_;
  wire _14478_;
  wire _14479_;
  wire _14480_;
  wire _14481_;
  wire _14482_;
  wire _14483_;
  wire _14484_;
  wire _14485_;
  wire _14486_;
  wire _14487_;
  wire _14488_;
  wire _14489_;
  wire _14490_;
  wire _14491_;
  wire _14492_;
  wire _14493_;
  wire _14494_;
  wire _14495_;
  wire _14496_;
  wire _14497_;
  wire _14498_;
  wire _14499_;
  wire _14500_;
  wire _14501_;
  wire _14502_;
  wire _14503_;
  wire _14504_;
  wire _14505_;
  wire _14506_;
  wire _14507_;
  wire _14508_;
  wire _14509_;
  wire _14510_;
  wire _14511_;
  wire _14512_;
  wire _14513_;
  wire _14514_;
  wire _14515_;
  wire _14516_;
  wire _14517_;
  wire _14518_;
  wire _14519_;
  wire _14520_;
  wire _14521_;
  wire _14522_;
  wire _14523_;
  wire _14524_;
  wire _14525_;
  wire _14526_;
  wire _14527_;
  wire _14528_;
  wire _14529_;
  wire _14530_;
  wire _14531_;
  wire _14532_;
  wire _14533_;
  wire _14534_;
  wire _14535_;
  wire _14536_;
  wire _14537_;
  wire _14538_;
  wire _14539_;
  wire _14540_;
  wire _14541_;
  wire _14542_;
  wire _14543_;
  wire _14544_;
  wire _14545_;
  wire _14546_;
  wire _14547_;
  wire _14548_;
  wire _14549_;
  wire _14550_;
  wire _14551_;
  wire _14552_;
  wire _14553_;
  wire _14554_;
  wire _14555_;
  wire _14556_;
  wire _14557_;
  wire _14558_;
  wire _14559_;
  wire _14560_;
  wire _14561_;
  wire _14562_;
  wire _14563_;
  wire _14564_;
  wire _14565_;
  wire _14566_;
  wire _14567_;
  wire _14568_;
  wire _14569_;
  wire _14570_;
  wire _14571_;
  wire _14572_;
  wire _14573_;
  wire _14574_;
  wire _14575_;
  wire _14576_;
  wire _14577_;
  wire _14578_;
  wire _14579_;
  wire _14580_;
  wire _14581_;
  wire _14582_;
  wire _14583_;
  wire _14584_;
  wire _14585_;
  wire _14586_;
  wire _14587_;
  wire _14588_;
  wire _14589_;
  wire _14590_;
  wire _14591_;
  wire _14592_;
  wire _14593_;
  wire _14594_;
  wire _14595_;
  wire _14596_;
  wire _14597_;
  wire _14598_;
  wire _14599_;
  wire _14600_;
  wire _14601_;
  wire _14602_;
  wire _14603_;
  wire _14604_;
  wire _14605_;
  wire _14606_;
  wire _14607_;
  input [8:0] ABINPUT;
  input clk;
  wire [31:0] cxrom_data_out;
  wire first_instr;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein0 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein1 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein2 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein3 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout0 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout1 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout2 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout3 ;
  wire \oc8051_symbolic_cxrom1.clk ;
  wire [31:0] \oc8051_symbolic_cxrom1.cxrom_data_out ;
  wire [15:0] \oc8051_symbolic_cxrom1.pc1 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc10 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc12 ;
  wire [15:0] \oc8051_symbolic_cxrom1.pc2 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc20 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc22 ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[0] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[10] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[11] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[12] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[13] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[14] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[15] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[1] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[2] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[3] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[4] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[5] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[6] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[7] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[8] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[9] ;
  wire [15:0] \oc8051_symbolic_cxrom1.regvalid ;
  wire \oc8051_symbolic_cxrom1.rst ;
  wire [31:0] \oc8051_symbolic_cxrom1.word_in ;
  wire [8:0] \oc8051_top_1.ABINPUT ;
  wire [7:0] \oc8051_top_1.acc ;
  wire \oc8051_top_1.bit_data ;
  wire [31:0] \oc8051_top_1.cxrom_data_out ;
  wire \oc8051_top_1.cy ;
  wire [1:0] \oc8051_top_1.cy_sel ;
  wire [7:0] \oc8051_top_1.dptr_hi ;
  wire [7:0] \oc8051_top_1.dptr_lo ;
  wire [31:0] \oc8051_top_1.idat_onchip ;
  wire \oc8051_top_1.int_ack ;
  wire [7:0] \oc8051_top_1.int_src ;
  wire \oc8051_top_1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.mem_act ;
  wire \oc8051_top_1.oc8051_alu1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.divsrc2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.des2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div0 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.div_out ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.rst ;
  wire [5:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.rst ;
  wire [15:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul ;
  wire \oc8051_top_1.oc8051_alu1.rst ;
  wire \oc8051_top_1.oc8051_alu1.srcAc ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.acc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.clk ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.dptr ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op1_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op2_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op3_r ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.pc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_alu_src_sel1.sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_alu_src_sel1.sel2 ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.sel3 ;
  wire [7:0] \oc8051_top_1.oc8051_comp1.acc ;
  wire \oc8051_top_1.oc8051_comp1.cy ;
  wire \oc8051_top_1.oc8051_cy_select1.cy_in ;
  wire [1:0] \oc8051_top_1.oc8051_cy_select1.cy_sel ;
  wire [3:0] \oc8051_top_1.oc8051_decoder1.alu_op ;
  wire \oc8051_top_1.oc8051_decoder1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.cy_sel ;
  wire \oc8051_top_1.oc8051_decoder1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_decoder1.op ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.psw_set ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_wr_sel ;
  wire \oc8051_top_1.oc8051_decoder1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.src_sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.src_sel2 ;
  wire \oc8051_top_1.oc8051_decoder1.src_sel3 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.state ;
  wire \oc8051_top_1.oc8051_decoder1.wait_data ;
  wire \oc8051_top_1.oc8051_decoder1.wr ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.wr_sfr ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[7] ;
  wire \oc8051_top_1.oc8051_indi_addr1.clk ;
  wire \oc8051_top_1.oc8051_indi_addr1.rst ;
  wire \oc8051_top_1.oc8051_indi_addr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.acc ;
  wire \oc8051_top_1.oc8051_memory_interface1.bit_in ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.cdata ;
  wire \oc8051_top_1.oc8051_memory_interface1.cdone ;
  wire \oc8051_top_1.oc8051_memory_interface1.clk ;
  wire \oc8051_top_1.oc8051_memory_interface1.dmem_wait ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dptr ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.iadr_t ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_cur ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_old ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_onchip ;
  wire \oc8051_top_1.oc8051_memory_interface1.imem_wait ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm2_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.in_ram ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_t ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_v ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_vec_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.istb_t ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op2_buff ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op3_buff ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.op_pos ;
  wire \oc8051_top_1.oc8051_memory_interface1.out_of_rst ;
  wire [3:0] \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_buf ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_for_ajmp ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log_prev ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_out ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_addr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_ind ;
  wire \oc8051_top_1.oc8051_memory_interface1.reti ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ri_r ;
  wire [4:0] \oc8051_top_1.oc8051_memory_interface1.rn_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.sfr ;
  wire \oc8051_top_1.oc8051_memory_interface1.sfr_bit ;
  wire \oc8051_top_1.oc8051_rom1.clk ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.cxrom_data_out ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.data_o ;
  wire \oc8051_top_1.oc8051_rom1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.b_reg ;
  wire \oc8051_top_1.oc8051_sfr1.bit_out ;
  wire \oc8051_top_1.oc8051_sfr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.cy ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_lo ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.int_ack ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ip ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ack ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.t2_int ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.uart_int ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.p ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.set ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd ;
  wire [11:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp ;
  wire [10:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.pres_ow ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.prescaler ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.psw_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.rxd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.srcAc ;
  wire \oc8051_top_1.oc8051_sfr1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.t2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.tc2_int ;
  wire \oc8051_top_1.oc8051_sfr1.tclk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.tf0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.uart_int ;
  wire \oc8051_top_1.oc8051_sfr1.wait_data ;
  wire \oc8051_top_1.oc8051_sfr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.p0_i ;
  wire [7:0] \oc8051_top_1.p0_o ;
  wire [7:0] \oc8051_top_1.p1_i ;
  wire [7:0] \oc8051_top_1.p1_o ;
  wire [7:0] \oc8051_top_1.p2_i ;
  wire [7:0] \oc8051_top_1.p2_o ;
  wire [7:0] \oc8051_top_1.p3_i ;
  wire [7:0] \oc8051_top_1.p3_o ;
  wire [15:0] \oc8051_top_1.pc ;
  wire [15:0] \oc8051_top_1.pc_log ;
  wire [15:0] \oc8051_top_1.pc_log_prev ;
  wire [1:0] \oc8051_top_1.psw_set ;
  wire [7:0] \oc8051_top_1.ram_data ;
  wire \oc8051_top_1.rd_ind ;
  wire \oc8051_top_1.reti ;
  wire \oc8051_top_1.rxd_i ;
  wire \oc8051_top_1.sfr_bit ;
  wire [7:0] \oc8051_top_1.sfr_out ;
  wire \oc8051_top_1.srcAc ;
  wire [2:0] \oc8051_top_1.src_sel1 ;
  wire [1:0] \oc8051_top_1.src_sel2 ;
  wire \oc8051_top_1.src_sel3 ;
  wire \oc8051_top_1.t0_i ;
  wire \oc8051_top_1.t1_i ;
  wire \oc8051_top_1.t2_i ;
  wire \oc8051_top_1.t2ex_i ;
  wire \oc8051_top_1.wait_data ;
  wire \oc8051_top_1.wb_clk_i ;
  wire \oc8051_top_1.wb_rst_i ;
  input [7:0] p0_in;
  wire [7:0] p0_out;
  input [7:0] p1_in;
  wire [7:0] p1_out;
  input [7:0] p2_in;
  wire [7:0] p2_out;
  input [7:0] p3_in;
  wire [7:0] p3_out;
  wire [15:0] pc1;
  wire [15:0] pc1_plus_2;
  wire [15:0] pc2;
  output property_invalid;
  input rst;
  input rxd_i;
  input t0_i;
  input t1_i;
  input t2_i;
  input t2ex_i;
  input [31:0] word_in;
  nor _14608_ (_06295_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  not _14609_ (_06296_, _06295_);
  and _14610_ (_06297_, _06296_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr );
  and _14611_ (_06298_, _06297_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  and _14612_ (_06299_, _06298_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  nor _14613_ (_06300_, _06298_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  nor _14614_ (_06301_, _06300_, _06299_);
  and _14615_ (_06302_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and _14616_ (_06303_, _06302_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  and _14617_ (_06304_, _06303_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  and _14618_ (_06305_, _06304_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  not _14619_ (_06306_, _06305_);
  not _14620_ (_06307_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  not _14621_ (_06308_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and _14622_ (_06309_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _06308_);
  and _14623_ (_06310_, _06309_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  and _14624_ (_06311_, _06310_, _06307_);
  not _14625_ (_06312_, _06311_);
  nor _14626_ (_06313_, _06304_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  nor _14627_ (_06314_, _06313_, _06312_);
  and _14628_ (_06315_, _06314_, _06306_);
  not _14629_ (_06316_, _06315_);
  not _14630_ (_06317_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  and _14631_ (_06318_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _06308_);
  and _14632_ (_06319_, _06318_, _06317_);
  and _14633_ (_06320_, _06319_, _06307_);
  and _14634_ (_06321_, _06320_, \oc8051_top_1.oc8051_memory_interface1.imm_r [4]);
  nor _14635_ (_06322_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and _14636_ (_06323_, _06322_, _06317_);
  or _14637_ (_06324_, _06323_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and _14638_ (_06325_, _06324_, \oc8051_top_1.oc8051_memory_interface1.rn_r [4]);
  nor _14639_ (_06326_, _06325_, _06321_);
  and _14640_ (_06327_, _06319_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and _14641_ (_06328_, _06327_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [4]);
  not _14642_ (_06329_, _06328_);
  and _14643_ (_06330_, _06310_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and _14644_ (_06331_, _06322_, _06309_);
  and _14645_ (_06332_, _06331_, \oc8051_top_1.oc8051_memory_interface1.ri_r [4]);
  nor _14646_ (_06333_, _06332_, _06330_);
  and _14647_ (_06334_, _06333_, _06329_);
  and _14648_ (_06335_, _06334_, _06326_);
  and _14649_ (_06336_, _06335_, _06316_);
  not _14650_ (_06337_, _06336_);
  and _14651_ (_06338_, _06305_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  not _14652_ (_06339_, _06338_);
  nor _14653_ (_06340_, _06305_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor _14654_ (_06341_, _06340_, _06312_);
  and _14655_ (_06342_, _06341_, _06339_);
  not _14656_ (_06343_, _06342_);
  and _14657_ (_06344_, _06331_, \oc8051_top_1.oc8051_memory_interface1.ri_r [5]);
  and _14658_ (_06345_, _06327_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [5]);
  and _14659_ (_06346_, _06320_, \oc8051_top_1.oc8051_memory_interface1.imm_r [5]);
  or _14660_ (_06347_, _06346_, _06345_);
  or _14661_ (_06348_, _06347_, _06330_);
  nor _14662_ (_06349_, _06348_, _06344_);
  and _14663_ (_06350_, _06349_, _06343_);
  and _14664_ (_06351_, _06350_, _06337_);
  and _14665_ (_06352_, _06338_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  not _14666_ (_06353_, _06352_);
  nor _14667_ (_06354_, _06338_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor _14668_ (_06355_, _06354_, _06312_);
  and _14669_ (_06356_, _06355_, _06353_);
  not _14670_ (_06357_, _06356_);
  and _14671_ (_06358_, _06331_, \oc8051_top_1.oc8051_memory_interface1.ri_r [6]);
  and _14672_ (_06359_, _06320_, \oc8051_top_1.oc8051_memory_interface1.imm_r [6]);
  and _14673_ (_06360_, _06327_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  or _14674_ (_06361_, _06360_, _06359_);
  or _14675_ (_06362_, _06361_, _06330_);
  nor _14676_ (_06363_, _06362_, _06358_);
  and _14677_ (_06364_, _06363_, _06357_);
  not _14678_ (_06365_, _06364_);
  not _14679_ (_06366_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  nor _14680_ (_06367_, _06352_, _06366_);
  and _14681_ (_06368_, _06352_, _06366_);
  nor _14682_ (_06369_, _06368_, _06367_);
  nor _14683_ (_06370_, _06369_, _06312_);
  not _14684_ (_06371_, _06370_);
  and _14685_ (_06372_, _06320_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  not _14686_ (_06373_, _06372_);
  and _14687_ (_06374_, _06327_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  not _14688_ (_06375_, _06374_);
  and _14689_ (_06376_, _06331_, \oc8051_top_1.oc8051_memory_interface1.ri_r [7]);
  nor _14690_ (_06377_, _06376_, _06330_);
  and _14691_ (_06378_, _06377_, _06375_);
  and _14692_ (_06379_, _06378_, _06373_);
  and _14693_ (_06380_, _06379_, _06371_);
  nor _14694_ (_06381_, _06380_, _06365_);
  and _14695_ (_06382_, _06381_, _06351_);
  and _14696_ (_06383_, _06327_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [3]);
  and _14697_ (_06384_, _06320_, \oc8051_top_1.oc8051_memory_interface1.imm_r [3]);
  nor _14698_ (_06385_, _06384_, _06383_);
  nor _14699_ (_06386_, _06303_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor _14700_ (_06387_, _06386_, _06304_);
  and _14701_ (_06388_, _06387_, _06311_);
  not _14702_ (_06389_, _06388_);
  and _14703_ (_06390_, _06331_, \oc8051_top_1.oc8051_memory_interface1.ri_r [3]);
  and _14704_ (_06391_, _06324_, \oc8051_top_1.oc8051_memory_interface1.rn_r [3]);
  nor _14705_ (_06392_, _06391_, _06390_);
  and _14706_ (_06393_, _06392_, _06389_);
  and _14707_ (_06394_, _06393_, _06385_);
  not _14708_ (_06395_, _06394_);
  and _14709_ (_06396_, _06320_, \oc8051_top_1.oc8051_memory_interface1.imm_r [0]);
  and _14710_ (_06397_, _06331_, \oc8051_top_1.oc8051_memory_interface1.ri_r [0]);
  nor _14711_ (_06398_, _06397_, _06396_);
  and _14712_ (_06399_, _06327_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  not _14713_ (_06400_, _06399_);
  not _14714_ (_06401_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and _14715_ (_06402_, _06311_, _06401_);
  and _14716_ (_06403_, _06324_, \oc8051_top_1.oc8051_memory_interface1.rn_r [0]);
  nor _14717_ (_06404_, _06403_, _06402_);
  and _14718_ (_06405_, _06404_, _06400_);
  and _14719_ (_06406_, _06405_, _06398_);
  not _14720_ (_06407_, _06406_);
  nor _14721_ (_06408_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  nor _14722_ (_06409_, _06408_, _06302_);
  and _14723_ (_06410_, _06409_, _06311_);
  and _14724_ (_06411_, _06331_, \oc8051_top_1.oc8051_memory_interface1.ri_r [1]);
  nor _14725_ (_06412_, _06411_, _06410_);
  and _14726_ (_06413_, _06327_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [1]);
  and _14727_ (_06414_, _06320_, \oc8051_top_1.oc8051_memory_interface1.imm_r [1]);
  and _14728_ (_06415_, _06324_, \oc8051_top_1.oc8051_memory_interface1.rn_r [1]);
  or _14729_ (_06416_, _06415_, _06414_);
  nor _14730_ (_06417_, _06416_, _06413_);
  and _14731_ (_06418_, _06417_, _06412_);
  nor _14732_ (_06419_, _06302_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor _14733_ (_06420_, _06419_, _06303_);
  and _14734_ (_06421_, _06420_, _06311_);
  and _14735_ (_06422_, _06331_, \oc8051_top_1.oc8051_memory_interface1.ri_r [2]);
  nor _14736_ (_06423_, _06422_, _06421_);
  and _14737_ (_06424_, _06327_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [2]);
  and _14738_ (_06425_, _06320_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  and _14739_ (_06426_, _06324_, \oc8051_top_1.oc8051_memory_interface1.rn_r [2]);
  or _14740_ (_06427_, _06426_, _06425_);
  nor _14741_ (_06428_, _06427_, _06424_);
  and _14742_ (_06430_, _06428_, _06423_);
  and _14743_ (_06431_, _06430_, _06418_);
  and _14744_ (_06432_, _06431_, _06407_);
  and _14745_ (_06434_, _06432_, _06395_);
  and _14746_ (_06435_, _06309_, _06307_);
  not _14747_ (_06436_, _06435_);
  not _14748_ (_06437_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and _14749_ (_06438_, \oc8051_top_1.oc8051_decoder1.wr , _06308_);
  and _14750_ (_06439_, _06438_, _06437_);
  and _14751_ (_06440_, _06439_, _06436_);
  and _14752_ (_06441_, _06440_, _06434_);
  and _14753_ (_06442_, _06441_, _06382_);
  nor _14754_ (_06443_, _06442_, rst);
  and _14755_ (_14257_, _06443_, _06301_);
  not _14756_ (_06444_, rst);
  and _14757_ (_06445_, _06380_, _06364_);
  and _14758_ (_06446_, _06445_, _06351_);
  and _14759_ (_06447_, _06446_, _06434_);
  and _14760_ (_06448_, _06447_, _06439_);
  not _14761_ (_06449_, _06448_);
  and _14762_ (_06450_, _06449_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  and _14763_ (_06451_, \oc8051_top_1.oc8051_decoder1.alu_op [1], _06308_);
  and _14764_ (_06452_, _06451_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and _14765_ (_06453_, \oc8051_top_1.oc8051_decoder1.alu_op [3], _06308_);
  and _14766_ (_06454_, _06453_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and _14767_ (_06455_, _06454_, _06452_);
  and _14768_ (_06456_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  nor _14769_ (_06457_, _06456_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  not _14770_ (_06458_, \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  and _14771_ (_06459_, _06458_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r );
  nor _14772_ (_06460_, _06459_, ABINPUT[0]);
  nand _14773_ (_06461_, _06458_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r );
  nor _14774_ (_06462_, _06461_, \oc8051_top_1.oc8051_sfr1.bit_out );
  nor _14775_ (_06463_, _06462_, _06460_);
  nor _14776_ (_06464_, _06463_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  nor _14777_ (_06465_, _06464_, _06457_);
  or _14778_ (_06466_, _06459_, ABINPUT[6]);
  or _14779_ (_06467_, _06461_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  nand _14780_ (_06468_, _06467_, _06466_);
  nor _14781_ (_06469_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  not _14782_ (_06470_, _06469_);
  or _14783_ (_06472_, _06470_, _06468_);
  not _14784_ (_06474_, \oc8051_top_1.oc8051_memory_interface1.imm_r [5]);
  nand _14785_ (_06475_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  or _14786_ (_06476_, _06475_, _06474_);
  not _14787_ (_06477_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  not _14788_ (_06478_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  nand _14789_ (_06479_, _06478_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  or _14790_ (_06480_, _06479_, _06477_);
  and _14791_ (_06481_, _06480_, _06476_);
  and _14792_ (_06482_, _06481_, _06472_);
  not _14793_ (_06483_, _06482_);
  and _14794_ (_06484_, _06483_, _06465_);
  not _14795_ (_06485_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  not _14796_ (_06486_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and _14797_ (_06487_, _06486_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  and _14798_ (_06488_, _06487_, _06485_);
  nand _14799_ (_06489_, _06488_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [5]);
  nor _14800_ (_06490_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], _06485_);
  and _14801_ (_06491_, _06490_, _06486_);
  nand _14802_ (_06492_, _06491_, \oc8051_top_1.oc8051_memory_interface1.imm_r [5]);
  and _14803_ (_06493_, _06492_, _06489_);
  nor _14804_ (_06494_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and _14805_ (_06495_, _06494_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  nand _14806_ (_06496_, _06495_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and _14807_ (_06497_, _06490_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  nand _14808_ (_06498_, _06497_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and _14809_ (_06499_, _06498_, _06496_);
  and _14810_ (_06500_, _06499_, _06493_);
  and _14811_ (_06501_, _06494_, _06486_);
  not _14812_ (_06502_, _06501_);
  or _14813_ (_06503_, _06502_, _06468_);
  and _14814_ (_06504_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and _14815_ (_06505_, _06504_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  nand _14816_ (_06506_, _06505_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [5]);
  and _14817_ (_06507_, _06504_, _06486_);
  nand _14818_ (_06508_, _06507_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and _14819_ (_06509_, _06508_, _06506_);
  and _14820_ (_06510_, _06509_, _06503_);
  and _14821_ (_06511_, _06510_, _06500_);
  nor _14822_ (_06512_, _06511_, _06465_);
  or _14823_ (_06513_, _06512_, _06484_);
  and _14824_ (_06514_, _06513_, _06455_);
  not _14825_ (_06515_, _06465_);
  nand _14826_ (_06516_, _06488_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [4]);
  nand _14827_ (_06518_, _06491_, \oc8051_top_1.oc8051_memory_interface1.imm_r [4]);
  and _14828_ (_06519_, _06518_, _06516_);
  nand _14829_ (_06520_, _06495_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nand _14830_ (_06521_, _06497_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _14831_ (_06522_, _06521_, _06520_);
  and _14832_ (_06523_, _06522_, _06519_);
  or _14833_ (_06524_, _06459_, ABINPUT[5]);
  or _14834_ (_06525_, _06461_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  nand _14835_ (_06526_, _06525_, _06524_);
  or _14836_ (_06527_, _06526_, _06502_);
  nand _14837_ (_06528_, _06505_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [4]);
  nand _14838_ (_06529_, _06507_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and _14839_ (_06530_, _06529_, _06528_);
  and _14840_ (_06531_, _06530_, _06527_);
  and _14841_ (_06532_, _06531_, _06523_);
  not _14842_ (_06534_, _06532_);
  nand _14843_ (_06535_, _06488_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [3]);
  nand _14844_ (_06537_, _06491_, \oc8051_top_1.oc8051_memory_interface1.imm_r [3]);
  and _14845_ (_06538_, _06537_, _06535_);
  and _14846_ (_06539_, _06495_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _14847_ (_06540_, _06497_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nor _14848_ (_06541_, _06540_, _06539_);
  and _14849_ (_06542_, _06541_, _06538_);
  or _14850_ (_06543_, _06459_, ABINPUT[4]);
  or _14851_ (_06544_, _06461_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  nand _14852_ (_06545_, _06544_, _06543_);
  or _14853_ (_06546_, _06545_, _06502_);
  and _14854_ (_06547_, _06505_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [3]);
  and _14855_ (_06548_, _06507_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor _14856_ (_06549_, _06548_, _06547_);
  and _14857_ (_06550_, _06549_, _06546_);
  and _14858_ (_06551_, _06550_, _06542_);
  not _14859_ (_06552_, _06551_);
  nand _14860_ (_06553_, _06488_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [1]);
  nand _14861_ (_06554_, _06491_, \oc8051_top_1.oc8051_memory_interface1.imm_r [1]);
  and _14862_ (_06555_, _06554_, _06553_);
  nand _14863_ (_06556_, _06497_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nand _14864_ (_06557_, _06495_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and _14865_ (_06558_, _06557_, _06556_);
  and _14866_ (_06559_, _06558_, _06555_);
  or _14867_ (_06560_, _06459_, ABINPUT[2]);
  or _14868_ (_06561_, _06461_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  nand _14869_ (_06562_, _06561_, _06560_);
  or _14870_ (_06563_, _06562_, _06502_);
  nand _14871_ (_06564_, _06505_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [1]);
  nand _14872_ (_06565_, _06507_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and _14873_ (_06567_, _06565_, _06564_);
  and _14874_ (_06568_, _06567_, _06563_);
  and _14875_ (_06570_, _06568_, _06559_);
  and _14876_ (_06571_, _06488_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  and _14877_ (_06572_, _06491_, \oc8051_top_1.oc8051_memory_interface1.imm_r [0]);
  nor _14878_ (_06573_, _06572_, _06571_);
  and _14879_ (_06574_, _06495_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and _14880_ (_06575_, _06497_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor _14881_ (_06576_, _06575_, _06574_);
  and _14882_ (_06577_, _06576_, _06573_);
  or _14883_ (_06578_, _06459_, ABINPUT[1]);
  or _14884_ (_06579_, _06461_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  and _14885_ (_06580_, _06579_, _06578_);
  and _14886_ (_06581_, _06580_, _06501_);
  and _14887_ (_06582_, _06505_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [0]);
  and _14888_ (_06583_, _06507_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor _14889_ (_06584_, _06583_, _06582_);
  not _14890_ (_06585_, _06584_);
  nor _14891_ (_06586_, _06585_, _06581_);
  and _14892_ (_06587_, _06586_, _06577_);
  nor _14893_ (_06588_, _06587_, _06570_);
  nand _14894_ (_06589_, _06488_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [2]);
  nand _14895_ (_06590_, _06491_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  and _14896_ (_06591_, _06590_, _06589_);
  or _14897_ (_06592_, _06459_, ABINPUT[3]);
  or _14898_ (_06593_, _06461_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  nand _14899_ (_06594_, _06593_, _06592_);
  or _14900_ (_06595_, _06594_, _06502_);
  and _14901_ (_06596_, _06595_, _06591_);
  nand _14902_ (_06597_, _06497_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nand _14903_ (_06598_, _06495_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and _14904_ (_06599_, _06598_, _06597_);
  nand _14905_ (_06600_, _06507_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nand _14906_ (_06601_, _06505_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [2]);
  and _14907_ (_06602_, _06601_, _06600_);
  and _14908_ (_06603_, _06602_, _06599_);
  and _14909_ (_06604_, _06603_, _06596_);
  not _14910_ (_06605_, _06604_);
  and _14911_ (_06606_, _06605_, _06588_);
  and _14912_ (_06607_, _06606_, _06552_);
  and _14913_ (_06608_, _06607_, _06534_);
  and _14914_ (_06609_, _06608_, _06515_);
  and _14915_ (_06610_, _06604_, _06570_);
  and _14916_ (_06611_, _06610_, _06587_);
  and _14917_ (_06612_, _06611_, _06551_);
  and _14918_ (_06613_, _06612_, _06532_);
  and _14919_ (_06614_, _06613_, _06465_);
  nor _14920_ (_06615_, _06614_, _06609_);
  nor _14921_ (_06616_, _06615_, _06511_);
  not _14922_ (_06617_, _06616_);
  not _14923_ (_06618_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and _14924_ (_06619_, _06451_, _06618_);
  and _14925_ (_06620_, _06619_, _06454_);
  not _14926_ (_06621_, _06620_);
  and _14927_ (_06622_, _06615_, _06511_);
  nor _14928_ (_06623_, _06622_, _06621_);
  and _14929_ (_06624_, _06623_, _06617_);
  nor _14930_ (_06625_, _06624_, _06514_);
  and _14931_ (_06626_, \oc8051_top_1.oc8051_decoder1.alu_op [0], _06308_);
  and _14932_ (_06627_, \oc8051_top_1.oc8051_decoder1.alu_op [2], _06308_);
  nor _14933_ (_06628_, _06627_, _06453_);
  and _14934_ (_06629_, _06628_, _06626_);
  not _14935_ (_06630_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  not _14936_ (_06631_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and _14937_ (_06632_, _06627_, _06631_);
  and _14938_ (_06633_, _06632_, _06630_);
  nor _14939_ (_06634_, _06633_, _06629_);
  not _14940_ (_06635_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and _14941_ (_06636_, _06453_, _06635_);
  and _14942_ (_06637_, _06636_, _06451_);
  not _14943_ (_06638_, _06637_);
  nor _14944_ (_06639_, _06626_, _06451_);
  and _14945_ (_06640_, _06639_, _06628_);
  and _14946_ (_06641_, _06454_, _06630_);
  nor _14947_ (_06642_, _06641_, _06640_);
  and _14948_ (_06643_, _06642_, _06638_);
  and _14949_ (_06644_, _06643_, _06634_);
  nor _14950_ (_06645_, _06644_, _06511_);
  not _14951_ (_06646_, _06645_);
  and _14952_ (_06647_, _06639_, _06636_);
  nor _14953_ (_06648_, _06511_, _06482_);
  and _14954_ (_06649_, _06511_, _06482_);
  nor _14955_ (_06650_, _06649_, _06648_);
  and _14956_ (_06651_, _06650_, _06647_);
  not _14957_ (_06652_, _06651_);
  and _14958_ (_06653_, _06626_, _06630_);
  and _14959_ (_06654_, _06653_, _06636_);
  not _14960_ (_06655_, _06654_);
  nor _14961_ (_06656_, _06655_, _06649_);
  not _14962_ (_06657_, _06656_);
  and _14963_ (_06658_, _06632_, _06452_);
  and _14964_ (_06659_, _06658_, _06648_);
  and _14965_ (_06660_, _06632_, _06619_);
  and _14966_ (_06661_, _06660_, _06511_);
  nor _14967_ (_06662_, _06661_, _06659_);
  and _14968_ (_06663_, _06662_, _06657_);
  and _14969_ (_06664_, _06663_, _06652_);
  and _14970_ (_06665_, _06664_, _06646_);
  and _14971_ (_06666_, _06665_, _06625_);
  nor _14972_ (_06667_, _06666_, _06449_);
  or _14973_ (_06668_, _06667_, _06450_);
  and _14974_ (_06471_, _06668_, _06444_);
  or _14975_ (_06669_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and _14976_ (_06670_, _06395_, _06336_);
  not _14977_ (_06671_, _06350_);
  nor _14978_ (_06672_, _06364_, _06671_);
  and _14979_ (_06673_, _06438_, _06436_);
  and _14980_ (_06674_, _06673_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  not _14981_ (_06675_, _06674_);
  nor _14982_ (_06676_, _06675_, _06380_);
  and _14983_ (_06677_, _06676_, _06672_);
  and _14984_ (_06678_, _06677_, _06670_);
  or _14985_ (_06679_, _06678_, _06669_);
  and _14986_ (_06680_, _06628_, _06619_);
  not _14987_ (_06681_, _06680_);
  nand _14988_ (_06682_, _06491_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  nand _14989_ (_06683_, _06488_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  and _14990_ (_06684_, _06683_, _06682_);
  and _14991_ (_06685_, _06497_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and _14992_ (_06686_, _06495_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor _14993_ (_06687_, _06686_, _06685_);
  and _14994_ (_06688_, _06687_, _06684_);
  or _14995_ (_06689_, _06459_, ABINPUT[8]);
  or _14996_ (_06690_, _06461_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  nand _14997_ (_06691_, _06690_, _06689_);
  or _14998_ (_06692_, _06691_, _06502_);
  and _14999_ (_06693_, _06505_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [7]);
  and _15000_ (_06694_, _06507_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor _15001_ (_06695_, _06694_, _06693_);
  and _15002_ (_06696_, _06695_, _06692_);
  and _15003_ (_06697_, _06696_, _06688_);
  or _15004_ (_06698_, _06691_, _06470_);
  not _15005_ (_06699_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  or _15006_ (_06700_, _06475_, _06699_);
  not _15007_ (_06701_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or _15008_ (_06702_, _06479_, _06701_);
  and _15009_ (_06703_, _06702_, _06700_);
  and _15010_ (_06704_, _06703_, _06698_);
  not _15011_ (_06705_, _06704_);
  and _15012_ (_06706_, _06705_, _06697_);
  nor _15013_ (_06707_, _06704_, _06697_);
  and _15014_ (_06708_, _06704_, _06697_);
  nor _15015_ (_06709_, _06708_, _06707_);
  nand _15016_ (_06710_, _06488_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  nand _15017_ (_06711_, _06491_, \oc8051_top_1.oc8051_memory_interface1.imm_r [6]);
  and _15018_ (_06712_, _06711_, _06710_);
  and _15019_ (_06714_, _06497_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and _15020_ (_06716_, _06495_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor _15021_ (_06718_, _06716_, _06714_);
  and _15022_ (_06720_, _06718_, _06712_);
  or _15023_ (_06722_, _06459_, ABINPUT[7]);
  or _15024_ (_06723_, _06461_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  nand _15025_ (_06725_, _06723_, _06722_);
  or _15026_ (_06727_, _06725_, _06502_);
  and _15027_ (_06728_, _06505_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [6]);
  and _15028_ (_06729_, _06507_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor _15029_ (_06730_, _06729_, _06728_);
  and _15030_ (_06731_, _06730_, _06727_);
  and _15031_ (_06732_, _06731_, _06720_);
  or _15032_ (_06733_, _06725_, _06470_);
  not _15033_ (_06734_, \oc8051_top_1.oc8051_memory_interface1.imm_r [6]);
  or _15034_ (_06735_, _06475_, _06734_);
  not _15035_ (_06736_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or _15036_ (_06737_, _06479_, _06736_);
  and _15037_ (_06738_, _06737_, _06735_);
  and _15038_ (_06739_, _06738_, _06733_);
  not _15039_ (_06740_, _06739_);
  nor _15040_ (_06741_, _06740_, _06732_);
  nor _15041_ (_06742_, _06739_, _06732_);
  and _15042_ (_06743_, _06739_, _06732_);
  nor _15043_ (_06744_, _06743_, _06742_);
  nor _15044_ (_06745_, _06511_, _06483_);
  or _15045_ (_06746_, _06526_, _06470_);
  not _15046_ (_06747_, \oc8051_top_1.oc8051_memory_interface1.imm_r [4]);
  or _15047_ (_06748_, _06475_, _06747_);
  not _15048_ (_06749_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or _15049_ (_06750_, _06479_, _06749_);
  and _15050_ (_06751_, _06750_, _06748_);
  and _15051_ (_06752_, _06751_, _06746_);
  not _15052_ (_06753_, _06752_);
  and _15053_ (_06754_, _06753_, _06532_);
  nor _15054_ (_06755_, _06754_, _06650_);
  nor _15055_ (_06756_, _06755_, _06745_);
  nor _15056_ (_06757_, _06756_, _06744_);
  nor _15057_ (_06758_, _06757_, _06741_);
  and _15058_ (_06759_, _06756_, _06744_);
  nor _15059_ (_06760_, _06759_, _06757_);
  not _15060_ (_06761_, _06760_);
  and _15061_ (_06762_, _06754_, _06650_);
  nor _15062_ (_06763_, _06762_, _06755_);
  not _15063_ (_06764_, _06763_);
  nor _15064_ (_06765_, _06752_, _06532_);
  and _15065_ (_06766_, _06752_, _06532_);
  nor _15066_ (_06767_, _06766_, _06765_);
  not _15067_ (_06768_, _06767_);
  or _15068_ (_06769_, _06545_, _06470_);
  not _15069_ (_06770_, \oc8051_top_1.oc8051_memory_interface1.imm_r [3]);
  or _15070_ (_06771_, _06475_, _06770_);
  not _15071_ (_06772_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or _15072_ (_06773_, _06479_, _06772_);
  and _15073_ (_06774_, _06773_, _06771_);
  and _15074_ (_06775_, _06774_, _06769_);
  and _15075_ (_06776_, _06775_, _06551_);
  nor _15076_ (_06777_, _06775_, _06551_);
  nor _15077_ (_06778_, _06777_, _06776_);
  or _15078_ (_06779_, _06594_, _06470_);
  not _15079_ (_06780_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  or _15080_ (_06781_, _06475_, _06780_);
  not _15081_ (_06782_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or _15082_ (_06783_, _06479_, _06782_);
  and _15083_ (_06784_, _06783_, _06781_);
  and _15084_ (_06785_, _06784_, _06779_);
  nor _15085_ (_06786_, _06785_, _06604_);
  and _15086_ (_06787_, _06785_, _06604_);
  nor _15087_ (_06788_, _06787_, _06786_);
  or _15088_ (_06789_, _06562_, _06470_);
  not _15089_ (_06790_, \oc8051_top_1.oc8051_memory_interface1.imm_r [1]);
  or _15090_ (_06791_, _06475_, _06790_);
  not _15091_ (_06792_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or _15092_ (_06793_, _06479_, _06792_);
  and _15093_ (_06794_, _06793_, _06791_);
  nand _15094_ (_06795_, _06794_, _06789_);
  not _15095_ (_06796_, _06795_);
  nor _15096_ (_06797_, _06796_, _06570_);
  and _15097_ (_06798_, _06796_, _06570_);
  nor _15098_ (_06799_, _06798_, _06797_);
  nand _15099_ (_06800_, _06580_, _06469_);
  not _15100_ (_06801_, \oc8051_top_1.oc8051_memory_interface1.imm_r [0]);
  or _15101_ (_06802_, _06475_, _06801_);
  not _15102_ (_06803_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or _15103_ (_06804_, _06479_, _06803_);
  and _15104_ (_06805_, _06804_, _06802_);
  nand _15105_ (_06806_, _06805_, _06800_);
  and _15106_ (_06807_, _06806_, _06587_);
  nor _15107_ (_06808_, _06807_, _06799_);
  nor _15108_ (_06809_, _06795_, _06570_);
  nor _15109_ (_06810_, _06809_, _06808_);
  nor _15110_ (_06811_, _06810_, _06788_);
  not _15111_ (_06812_, _06785_);
  nor _15112_ (_06813_, _06812_, _06604_);
  nor _15113_ (_06814_, _06813_, _06811_);
  nor _15114_ (_06815_, _06814_, _06778_);
  and _15115_ (_06816_, _06814_, _06778_);
  nor _15116_ (_06817_, _06816_, _06815_);
  and _15117_ (_06818_, _06810_, _06788_);
  nor _15118_ (_06819_, _06818_, _06811_);
  not _15119_ (_06820_, _06819_);
  and _15120_ (_06821_, _06807_, _06799_);
  nor _15121_ (_06822_, _06821_, _06808_);
  not _15122_ (_06823_, _06822_);
  not _15123_ (_06824_, _06806_);
  nor _15124_ (_06825_, _06824_, _06587_);
  and _15125_ (_06826_, _06824_, _06587_);
  nor _15126_ (_06827_, _06826_, _06825_);
  nor _15127_ (_06828_, _06827_, _06515_);
  and _15128_ (_06829_, _06828_, _06823_);
  and _15129_ (_06830_, _06829_, _06820_);
  not _15130_ (_06831_, _06830_);
  nor _15131_ (_06832_, _06831_, _06817_);
  not _15132_ (_06833_, _06775_);
  or _15133_ (_06834_, _06833_, _06551_);
  and _15134_ (_06835_, _06833_, _06551_);
  or _15135_ (_06836_, _06814_, _06835_);
  and _15136_ (_06837_, _06836_, _06834_);
  or _15137_ (_06838_, _06837_, _06832_);
  and _15138_ (_06839_, _06838_, _06768_);
  and _15139_ (_06840_, _06839_, _06764_);
  and _15140_ (_06841_, _06840_, _06761_);
  nor _15141_ (_06842_, _06841_, _06758_);
  nor _15142_ (_06843_, _06842_, _06709_);
  nor _15143_ (_06844_, _06843_, _06706_);
  nor _15144_ (_06845_, _06844_, _06681_);
  not _15145_ (_06846_, _06845_);
  and _15146_ (_06847_, _06653_, _06628_);
  not _15147_ (_06848_, _06847_);
  not _15148_ (_06849_, _06744_);
  and _15149_ (_06850_, _06765_, _06650_);
  nor _15150_ (_06851_, _06850_, _06648_);
  nor _15151_ (_06852_, _06851_, _06849_);
  not _15152_ (_06853_, _06788_);
  and _15153_ (_06854_, _06825_, _06799_);
  nor _15154_ (_06855_, _06854_, _06797_);
  nor _15155_ (_06856_, _06855_, _06853_);
  nor _15156_ (_06857_, _06856_, _06786_);
  nor _15157_ (_06858_, _06857_, _06778_);
  and _15158_ (_06859_, _06857_, _06778_);
  nor _15159_ (_06860_, _06859_, _06858_);
  and _15160_ (_06861_, _06827_, _06465_);
  and _15161_ (_06862_, _06861_, _06799_);
  and _15162_ (_06863_, _06855_, _06853_);
  nor _15163_ (_06864_, _06863_, _06856_);
  and _15164_ (_06865_, _06864_, _06862_);
  not _15165_ (_06866_, _06865_);
  nor _15166_ (_06867_, _06866_, _06860_);
  nor _15167_ (_06868_, _06857_, _06776_);
  or _15168_ (_06869_, _06868_, _06777_);
  or _15169_ (_06870_, _06869_, _06867_);
  and _15170_ (_06871_, _06870_, _06767_);
  and _15171_ (_06872_, _06871_, _06650_);
  and _15172_ (_06873_, _06851_, _06849_);
  nor _15173_ (_06874_, _06873_, _06852_);
  and _15174_ (_06875_, _06874_, _06872_);
  or _15175_ (_06876_, _06875_, _06742_);
  nor _15176_ (_06877_, _06876_, _06852_);
  nor _15177_ (_06878_, _06877_, _06708_);
  nor _15178_ (_06879_, _06878_, _06707_);
  nor _15179_ (_06880_, _06879_, _06848_);
  and _15180_ (_06881_, _06732_, _06511_);
  not _15181_ (_06882_, _06881_);
  and _15182_ (_06883_, _06653_, _06632_);
  nor _15183_ (_06884_, _06610_, _06551_);
  and _15184_ (_06885_, _06884_, _06883_);
  and _15185_ (_06886_, _06885_, _06534_);
  nor _15186_ (_06887_, _06886_, _06882_);
  nor _15187_ (_06888_, _06887_, _06697_);
  nor _15188_ (_06889_, _06888_, _06465_);
  not _15189_ (_06890_, _06889_);
  not _15190_ (_06891_, _06883_);
  nor _15191_ (_06892_, _06697_, _06515_);
  not _15192_ (_06893_, _06892_);
  nor _15193_ (_06894_, _06893_, _06887_);
  nor _15194_ (_06895_, _06894_, _06891_);
  and _15195_ (_06896_, _06895_, _06890_);
  nor _15196_ (_06897_, _06465_, _06463_);
  not _15197_ (_06898_, _06647_);
  and _15198_ (_06899_, _06465_, _06463_);
  or _15199_ (_06900_, _06899_, _06898_);
  and _15200_ (_06901_, _06900_, _06655_);
  or _15201_ (_06902_, _06901_, _06897_);
  not _15202_ (_06903_, _06587_);
  and _15203_ (_06904_, _06653_, _06454_);
  and _15204_ (_06905_, _06904_, _06903_);
  and _15205_ (_06906_, _06463_, _06457_);
  and _15206_ (_06907_, _06636_, _06619_);
  and _15207_ (_06908_, _06658_, _06463_);
  nor _15208_ (_06909_, _06908_, _06907_);
  nor _15209_ (_06910_, _06909_, _06906_);
  nor _15210_ (_06911_, _06910_, _06905_);
  and _15211_ (_06912_, _06911_, _06902_);
  and _15212_ (_06913_, _06636_, _06452_);
  not _15213_ (_06914_, _06697_);
  and _15214_ (_06915_, _06914_, _06913_);
  nor _15215_ (_06916_, _06660_, _06465_);
  not _15216_ (_06917_, _06463_);
  and _15217_ (_06918_, _06639_, _06454_);
  and _15218_ (_06919_, _06918_, _06917_);
  nor _15219_ (_06920_, _06919_, _06640_);
  and _15220_ (_06921_, _06920_, _06465_);
  nor _15221_ (_06922_, _06921_, _06916_);
  or _15222_ (_06923_, _06922_, _06885_);
  nor _15223_ (_06924_, _06923_, _06915_);
  and _15224_ (_06925_, _06924_, _06912_);
  not _15225_ (_06926_, _06925_);
  nor _15226_ (_06927_, _06926_, _06896_);
  not _15227_ (_06928_, _06927_);
  nor _15228_ (_06929_, _06928_, _06880_);
  and _15229_ (_06930_, _06929_, _06846_);
  not _15230_ (_06931_, _06430_);
  nor _15231_ (_06932_, _06418_, _06406_);
  and _15232_ (_06933_, _06932_, _06931_);
  not _15233_ (_06934_, _06933_);
  nor _15234_ (_06935_, _06934_, _06930_);
  nand _15235_ (_06936_, _06934_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  nand _15236_ (_06937_, _06936_, _06678_);
  or _15237_ (_06938_, _06937_, _06935_);
  and _15238_ (_06939_, _06938_, _06679_);
  nor _15239_ (_06940_, _06380_, _06337_);
  and _15240_ (_06941_, _06940_, _06672_);
  and _15241_ (_06942_, _06431_, _06406_);
  not _15242_ (_06943_, _06440_);
  nor _15243_ (_06944_, _06943_, _06394_);
  and _15244_ (_06945_, _06944_, _06942_);
  and _15245_ (_06946_, _06945_, _06941_);
  or _15246_ (_06947_, _06946_, _06939_);
  and _15247_ (_06948_, _06697_, _06515_);
  not _15248_ (_06949_, _06948_);
  not _15249_ (_06951_, _06455_);
  and _15250_ (_06952_, _06704_, _06465_);
  nor _15251_ (_06953_, _06952_, _06951_);
  and _15252_ (_06954_, _06953_, _06949_);
  and _15253_ (_06955_, _06881_, _06613_);
  nor _15254_ (_06956_, _06955_, _06515_);
  not _15255_ (_06957_, _06732_);
  not _15256_ (_06958_, _06511_);
  and _15257_ (_06959_, _06608_, _06958_);
  and _15258_ (_06960_, _06959_, _06957_);
  nor _15259_ (_06961_, _06960_, _06465_);
  nor _15260_ (_06962_, _06961_, _06956_);
  and _15261_ (_06963_, _06962_, _06914_);
  nor _15262_ (_06964_, _06962_, _06914_);
  nor _15263_ (_06965_, _06964_, _06963_);
  and _15264_ (_06966_, _06965_, _06620_);
  nor _15265_ (_06967_, _06966_, _06954_);
  and _15266_ (_06968_, _06709_, _06647_);
  and _15267_ (_06969_, _06707_, _06658_);
  nor _15268_ (_06970_, _06708_, _06655_);
  and _15269_ (_06971_, _06697_, _06660_);
  or _15270_ (_06972_, _06971_, _06970_);
  or _15271_ (_06973_, _06972_, _06969_);
  nor _15272_ (_06974_, _06973_, _06968_);
  nor _15273_ (_06975_, _06697_, _06644_);
  not _15274_ (_06976_, _06975_);
  and _15275_ (_06977_, _06976_, _06974_);
  and _15276_ (_06978_, _06977_, _06967_);
  nand _15277_ (_06979_, _06978_, _06946_);
  and _15278_ (_06980_, _06979_, _06444_);
  and _15279_ (_09333_, _06980_, _06947_);
  not _15280_ (_06981_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and _15281_ (_06982_, _06418_, _06406_);
  and _15282_ (_06983_, _06982_, _06931_);
  and _15283_ (_06984_, _06944_, _06983_);
  and _15284_ (_06985_, _06984_, _06941_);
  and _15285_ (_06986_, _06418_, _06407_);
  and _15286_ (_06987_, _06986_, _06931_);
  and _15287_ (_06988_, _06944_, _06987_);
  and _15288_ (_06989_, _06988_, _06941_);
  nor _15289_ (_06990_, _06989_, _06985_);
  nor _15290_ (_06991_, _06990_, _06981_);
  and _15291_ (_06992_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and _15292_ (_06993_, _06992_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and _15293_ (_06994_, _06993_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and _15294_ (_06995_, _06994_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and _15295_ (_06996_, _06995_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and _15296_ (_06997_, _06996_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and _15297_ (_06998_, _06997_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and _15298_ (_06999_, _06998_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and _15299_ (_07000_, _06999_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and _15300_ (_07001_, _07000_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and _15301_ (_07002_, _07001_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and _15302_ (_07003_, _07002_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and _15303_ (_07004_, _07003_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  and _15304_ (_07005_, _07004_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  and _15305_ (_07006_, _07005_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  or _15306_ (_07007_, \oc8051_top_1.oc8051_sfr1.pres_ow , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  not _15307_ (_07008_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or _15308_ (_07009_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _07008_);
  and _15309_ (_07010_, _07009_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and _15310_ (_07011_, _07010_, _07007_);
  nor _15311_ (_07012_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  not _15312_ (_07013_, _07012_);
  not _15313_ (_07014_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and _15314_ (_07015_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and _15315_ (_07016_, _07015_, _07012_);
  and _15316_ (_07017_, _07016_, _07014_);
  nor _15317_ (_07018_, _07017_, _07013_);
  and _15318_ (_07019_, _07018_, _07011_);
  and _15319_ (_07020_, _07019_, _06990_);
  and _15320_ (_07021_, _07020_, _07006_);
  or _15321_ (_07022_, _07021_, _06991_);
  and _15322_ (_09435_, _07022_, _06444_);
  nand _15323_ (_07023_, _06989_, _06978_);
  and _15324_ (_07024_, _07011_, _07005_);
  nor _15325_ (_07025_, _07024_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  and _15326_ (_07026_, _07011_, _07006_);
  nor _15327_ (_07027_, _07026_, _07025_);
  and _15328_ (_07028_, _07012_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  not _15329_ (_07029_, _07028_);
  and _15330_ (_07030_, _07029_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  and _15331_ (_07031_, _07030_, _07011_);
  and _15332_ (_07032_, _07031_, _07006_);
  or _15333_ (_07033_, _07032_, _07017_);
  or _15334_ (_07034_, _07033_, _07027_);
  not _15335_ (_07035_, _07017_);
  nor _15336_ (_07036_, _07035_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  nor _15337_ (_07037_, _07036_, _06985_);
  and _15338_ (_07038_, _07037_, _07034_);
  and _15339_ (_07039_, _06985_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  or _15340_ (_07040_, _07039_, _06989_);
  or _15341_ (_07041_, _07040_, _07038_);
  and _15342_ (_07042_, _07041_, _06444_);
  and _15343_ (_11388_, _07042_, _07023_);
  and _15344_ (_07043_, _06432_, _06394_);
  and _15345_ (_07044_, _07043_, _06446_);
  and _15346_ (_07045_, _07044_, _06439_);
  not _15347_ (_07046_, _07045_);
  and _15348_ (_07047_, _07046_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  and _15349_ (_07048_, _06795_, _06455_);
  and _15350_ (_07049_, _06587_, _06570_);
  nor _15351_ (_07050_, _07049_, _06588_);
  and _15352_ (_07052_, _07050_, _06465_);
  nor _15353_ (_07053_, _07050_, _06465_);
  or _15354_ (_07054_, _07053_, _06621_);
  nor _15355_ (_07055_, _07054_, _07052_);
  nor _15356_ (_07056_, _07055_, _07048_);
  nor _15357_ (_07057_, _06644_, _06570_);
  not _15358_ (_07058_, _07057_);
  and _15359_ (_07059_, _06799_, _06647_);
  not _15360_ (_07060_, _07059_);
  nor _15361_ (_07061_, _06798_, _06655_);
  not _15362_ (_07062_, _07061_);
  and _15363_ (_07063_, _06797_, _06658_);
  and _15364_ (_07064_, _06660_, _06570_);
  nor _15365_ (_07065_, _07064_, _07063_);
  and _15366_ (_07066_, _07065_, _07062_);
  and _15367_ (_07067_, _07066_, _07060_);
  and _15368_ (_07068_, _07067_, _07058_);
  and _15369_ (_07069_, _07068_, _07056_);
  not _15370_ (_07070_, _07069_);
  and _15371_ (_07071_, _07070_, _07045_);
  or _15372_ (_07072_, _07071_, _07047_);
  and _15373_ (_11722_, _07072_, _06444_);
  and _15374_ (_07073_, \oc8051_top_1.oc8051_memory_interface1.reti , \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  and _15375_ (_07074_, _06444_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  and _15376_ (_12487_, _07074_, _07073_);
  not _15377_ (_07075_, _07073_);
  not _15378_ (_07076_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  not _15379_ (_07077_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and _15380_ (_07078_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _07077_);
  and _15381_ (_07079_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _15382_ (_07080_, _07079_, _07078_);
  and _15383_ (_07081_, _07080_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  nor _15384_ (_07082_, _07081_, _07076_);
  and _15385_ (_07083_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and _15386_ (_07084_, _07083_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  not _15387_ (_07085_, _07084_);
  and _15388_ (_07086_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and _15389_ (_07087_, _07086_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and _15390_ (_07088_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and _15391_ (_07089_, _07088_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  nor _15392_ (_07090_, _07089_, _07087_);
  and _15393_ (_07091_, _07090_, _07085_);
  not _15394_ (_07092_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  nor _15395_ (_07093_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  nor _15396_ (_07094_, _07093_, _07092_);
  and _15397_ (_07095_, _07094_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  not _15398_ (_07096_, _07095_);
  not _15399_ (_07098_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  nor _15400_ (_07099_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  nor _15401_ (_07100_, _07099_, _07098_);
  nand _15402_ (_07101_, _07100_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and _15403_ (_07102_, _07101_, _07096_);
  and _15404_ (_07103_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and _15405_ (_07104_, _07103_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  not _15406_ (_07105_, _07104_);
  and _15407_ (_07106_, _07105_, _07102_);
  and _15408_ (_07107_, _07106_, _07091_);
  nor _15409_ (_07108_, _07107_, _07082_);
  and _15410_ (_07109_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _07076_);
  not _15411_ (_07110_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and _15412_ (_07111_, _07094_, _07110_);
  not _15413_ (_07112_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and _15414_ (_07113_, _07100_, _07112_);
  nor _15415_ (_07114_, _07113_, _07111_);
  not _15416_ (_07115_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and _15417_ (_07116_, _07103_, _07115_);
  not _15418_ (_07117_, _07116_);
  not _15419_ (_07118_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and _15420_ (_07119_, _07083_, _07118_);
  not _15421_ (_07120_, _07119_);
  not _15422_ (_07121_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and _15423_ (_07122_, _07086_, _07121_);
  not _15424_ (_07123_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and _15425_ (_07124_, _07088_, _07123_);
  nor _15426_ (_07125_, _07124_, _07122_);
  and _15427_ (_07126_, _07125_, _07120_);
  and _15428_ (_07127_, _07126_, _07117_);
  nand _15429_ (_07128_, _07127_, _07114_);
  nand _15430_ (_07130_, _07128_, _07109_);
  not _15431_ (_07131_, _07130_);
  nor _15432_ (_07132_, _07131_, _07108_);
  and _15433_ (_07133_, _07132_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  not _15434_ (_07134_, _07108_);
  nor _15435_ (_07135_, _07077_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  and _15436_ (_07136_, _07077_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  nor _15437_ (_07137_, _07136_, _07135_);
  nor _15438_ (_07138_, _07137_, _07134_);
  or _15439_ (_07139_, _07138_, _07133_);
  and _15440_ (_07140_, _07139_, _07075_);
  and _15441_ (_07141_, _07137_, _07073_);
  or _15442_ (_07142_, _07141_, _07140_);
  and _15443_ (_12749_, _07142_, _06444_);
  nand _15444_ (_07143_, _07130_, _07076_);
  or _15445_ (_07144_, _07143_, _07108_);
  nand _15446_ (_07145_, _07135_, _07073_);
  and _15447_ (_07146_, _07145_, _06444_);
  and _15448_ (_12769_, _07146_, _07144_);
  and _15449_ (_07147_, _06942_, _06395_);
  and _15450_ (_07148_, _07147_, _06446_);
  not _15451_ (_07149_, _07044_);
  and _15452_ (_07150_, _06942_, _06394_);
  and _15453_ (_07151_, _07150_, _06446_);
  and _15454_ (_07152_, _06350_, _06336_);
  and _15455_ (_07153_, _07152_, _06445_);
  and _15456_ (_07154_, _07153_, _06434_);
  nor _15457_ (_07155_, _07154_, _07151_);
  nand _15458_ (_07156_, _07155_, _07149_);
  nor _15459_ (_07157_, _07156_, _07148_);
  not _15460_ (_07158_, _06439_);
  and _15461_ (_07159_, _07153_, _07150_);
  or _15462_ (_07160_, _07159_, _07158_);
  or _15463_ (_07161_, _07160_, _07157_);
  and _15464_ (_07162_, _07161_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  and _15465_ (_07163_, _06439_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  and _15466_ (_07164_, _07163_, _07156_);
  nor _15467_ (_07166_, _06532_, _06465_);
  and _15468_ (_07167_, _06753_, _06465_);
  or _15469_ (_07168_, _07167_, _07166_);
  and _15470_ (_07169_, _07168_, _06455_);
  nor _15471_ (_07170_, _06607_, _06465_);
  nor _15472_ (_07171_, _06612_, _06515_);
  nor _15473_ (_07172_, _07171_, _07170_);
  nor _15474_ (_07173_, _07172_, _06534_);
  and _15475_ (_07174_, _07172_, _06534_);
  nor _15476_ (_07175_, _07174_, _07173_);
  and _15477_ (_07176_, _07175_, _06620_);
  nor _15478_ (_07177_, _07176_, _07169_);
  nor _15479_ (_07178_, _06644_, _06532_);
  not _15480_ (_07179_, _07178_);
  and _15481_ (_07180_, _06767_, _06647_);
  and _15482_ (_07181_, _06765_, _06658_);
  nor _15483_ (_07182_, _06766_, _06655_);
  and _15484_ (_07183_, _06660_, _06532_);
  or _15485_ (_07184_, _07183_, _07182_);
  or _15486_ (_07185_, _07184_, _07181_);
  nor _15487_ (_07186_, _07185_, _07180_);
  and _15488_ (_07187_, _07186_, _07179_);
  and _15489_ (_07188_, _07187_, _07177_);
  and _15490_ (_07189_, _07148_, _06439_);
  not _15491_ (_07190_, _07189_);
  nor _15492_ (_07191_, _07190_, _07188_);
  or _15493_ (_07192_, _07191_, _07164_);
  or _15494_ (_07193_, _07192_, _07162_);
  and _15495_ (_13150_, _07193_, _06444_);
  or _15496_ (_07194_, _07091_, _07082_);
  nor _15497_ (_07195_, _07130_, _07108_);
  not _15498_ (_07196_, _07195_);
  or _15499_ (_07197_, _07196_, _07126_);
  and _15500_ (_07198_, _07197_, _07194_);
  nor _15501_ (_07199_, _07073_, _07077_);
  not _15502_ (_07200_, _07199_);
  or _15503_ (_07201_, _07200_, _07198_);
  not _15504_ (_07202_, _07114_);
  and _15505_ (_07203_, _07202_, _07109_);
  and _15506_ (_07204_, _07116_, _07109_);
  or _15507_ (_07205_, _07204_, _07203_);
  or _15508_ (_07206_, _07205_, _07108_);
  not _15509_ (_07207_, _07106_);
  or _15510_ (_07208_, _07194_, _07207_);
  and _15511_ (_07209_, _07208_, _07199_);
  and _15512_ (_07210_, _07209_, _07206_);
  or _15513_ (_07211_, _07210_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  and _15514_ (_07213_, _07211_, _06444_);
  and _15515_ (_13339_, _07213_, _07201_);
  and _15516_ (_07214_, _06440_, _06394_);
  and _15517_ (_07215_, _07214_, _06942_);
  nor _15518_ (_07216_, _06380_, _06364_);
  and _15519_ (_07217_, _07216_, _06351_);
  and _15520_ (_07218_, _07217_, _07215_);
  not _15521_ (_07219_, _07218_);
  and _15522_ (_07220_, _07219_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  nor _15523_ (_07221_, _07219_, _07188_);
  nor _15524_ (_07222_, _07221_, _07220_);
  nor _15525_ (_07223_, _07222_, _06337_);
  and _15526_ (_07224_, _07222_, _06337_);
  nor _15527_ (_07225_, _07224_, _07223_);
  not _15528_ (_07226_, \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  nor _15529_ (_07227_, \oc8051_top_1.oc8051_memory_interface1.imem_wait , \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  and _15530_ (_07228_, _07227_, _07226_);
  nor _15531_ (_07229_, \oc8051_top_1.oc8051_decoder1.state [1], \oc8051_top_1.oc8051_decoder1.state [0]);
  and _15532_ (_07230_, _07229_, _06308_);
  and _15533_ (_07231_, _07230_, _07228_);
  not _15534_ (_07232_, _07231_);
  not _15535_ (_07233_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  not _15536_ (_07234_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  not _15537_ (_07235_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  not _15538_ (_07236_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  nor _15539_ (_07237_, _07236_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _15540_ (_07238_, _07237_, _07235_);
  nand _15541_ (_07239_, _07238_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  and _15542_ (_07240_, _07236_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nand _15543_ (_07241_, _07240_, _07235_);
  not _15544_ (_07242_, _07241_);
  nand _15545_ (_07243_, _07242_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  and _15546_ (_07244_, _07243_, _07239_);
  nor _15547_ (_07245_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor _15548_ (_07246_, _07245_, _07235_);
  nand _15549_ (_07247_, _07246_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and _15550_ (_07248_, _07245_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nand _15551_ (_07249_, _07248_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and _15552_ (_07250_, _07249_, _07247_);
  and _15553_ (_07251_, _07245_, _07235_);
  nand _15554_ (_07252_, _07251_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  and _15555_ (_07253_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _15556_ (_07254_, _07253_, _07235_);
  nand _15557_ (_07255_, _07254_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  and _15558_ (_07256_, _07255_, _07252_);
  and _15559_ (_07257_, _07256_, _07250_);
  nand _15560_ (_07258_, _07257_, _07244_);
  nand _15561_ (_07259_, _07258_, _07234_);
  nand _15562_ (_07260_, _07259_, _07233_);
  nor _15563_ (_07261_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], _07233_);
  not _15564_ (_07262_, _07261_);
  and _15565_ (_07263_, _07262_, _07260_);
  or _15566_ (_07264_, _07263_, _07232_);
  not _15567_ (_07265_, _07228_);
  nor _15568_ (_07266_, _07230_, \oc8051_top_1.oc8051_decoder1.op [0]);
  nor _15569_ (_07267_, _07266_, _07265_);
  and _15570_ (_07268_, _07267_, _07264_);
  and _15571_ (_07269_, _07268_, _06406_);
  not _15572_ (_07270_, _07269_);
  and _15573_ (_07271_, _06439_, _06431_);
  and _15574_ (_07272_, _07271_, _06350_);
  and _15575_ (_07273_, _07272_, _06445_);
  nor _15576_ (_07274_, _07268_, _06406_);
  not _15577_ (_07275_, _07274_);
  and _15578_ (_07276_, _07275_, _07273_);
  and _15579_ (_07277_, _07276_, _07270_);
  and _15580_ (_07278_, _07219_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  nor _15581_ (_07280_, _06775_, _06951_);
  nor _15582_ (_07281_, _06611_, _06515_);
  nor _15583_ (_07282_, _06606_, _06465_);
  nor _15584_ (_07283_, _07282_, _07281_);
  and _15585_ (_07284_, _07283_, _06552_);
  not _15586_ (_07285_, _07284_);
  nor _15587_ (_07286_, _07283_, _06552_);
  nor _15588_ (_07287_, _07286_, _06621_);
  and _15589_ (_07288_, _07287_, _07285_);
  nor _15590_ (_07289_, _07288_, _07280_);
  nor _15591_ (_07290_, _06776_, _06655_);
  and _15592_ (_07291_, _06778_, _06647_);
  nor _15593_ (_07292_, _07291_, _07290_);
  and _15594_ (_07293_, _06777_, _06658_);
  and _15595_ (_07294_, _06660_, _06551_);
  nor _15596_ (_07295_, _07294_, _07293_);
  nor _15597_ (_07296_, _06644_, _06551_);
  not _15598_ (_07297_, _07296_);
  and _15599_ (_07298_, _07297_, _07295_);
  and _15600_ (_07299_, _07298_, _07292_);
  and _15601_ (_07300_, _07299_, _07289_);
  nor _15602_ (_07301_, _07300_, _07219_);
  nor _15603_ (_07302_, _07301_, _07278_);
  and _15604_ (_07303_, _07302_, _06395_);
  nor _15605_ (_07304_, _07302_, _06395_);
  nor _15606_ (_07305_, _07304_, _07303_);
  and _15607_ (_07306_, _07305_, _07277_);
  and _15608_ (_07307_, _07306_, _07225_);
  nor _15609_ (_07308_, _07268_, _07302_);
  and _15610_ (_07309_, _07308_, _07222_);
  and _15611_ (_07310_, _07309_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  not _15612_ (_07311_, _07268_);
  and _15613_ (_07312_, _07311_, _07302_);
  and _15614_ (_07313_, _07312_, _07222_);
  and _15615_ (_07314_, _07313_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  nor _15616_ (_07315_, _07314_, _07310_);
  not _15617_ (_07316_, _07222_);
  and _15618_ (_07317_, _07268_, _07302_);
  and _15619_ (_07318_, _07317_, _07316_);
  and _15620_ (_07319_, _07318_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  nor _15621_ (_07320_, _07311_, _07302_);
  and _15622_ (_07321_, _07320_, _07316_);
  and _15623_ (_07322_, _07321_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  nor _15624_ (_07323_, _07322_, _07319_);
  and _15625_ (_07324_, _07323_, _07315_);
  and _15626_ (_07325_, _07308_, _07316_);
  and _15627_ (_07326_, _07325_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  and _15628_ (_07327_, _07312_, _07316_);
  and _15629_ (_07329_, _07327_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  nor _15630_ (_07330_, _07329_, _07326_);
  and _15631_ (_07331_, _07320_, _07222_);
  and _15632_ (_07332_, _07331_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  and _15633_ (_07333_, _07317_, _07222_);
  and _15634_ (_07334_, _07333_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  nor _15635_ (_07335_, _07334_, _07332_);
  and _15636_ (_07336_, _07335_, _07330_);
  and _15637_ (_07338_, _07336_, _07324_);
  nor _15638_ (_07339_, _07338_, _07307_);
  not _15639_ (_07340_, _07300_);
  and _15640_ (_07341_, _07307_, _07340_);
  nor _15641_ (_07342_, _07341_, _07339_);
  nor _15642_ (_14055_, _07342_, rst);
  and _15643_ (_07343_, _07309_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  and _15644_ (_07344_, _07313_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  nor _15645_ (_07345_, _07344_, _07343_);
  and _15646_ (_07346_, _07327_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  and _15647_ (_07347_, _07321_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  nor _15648_ (_07348_, _07347_, _07346_);
  and _15649_ (_07349_, _07348_, _07345_);
  and _15650_ (_07350_, _07325_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  and _15651_ (_07351_, _07318_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  nor _15652_ (_07352_, _07351_, _07350_);
  and _15653_ (_07353_, _07331_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  and _15654_ (_07354_, _07333_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  nor _15655_ (_07355_, _07354_, _07353_);
  and _15656_ (_07356_, _07355_, _07352_);
  and _15657_ (_07357_, _07356_, _07349_);
  nor _15658_ (_07358_, _07357_, _07307_);
  not _15659_ (_07359_, _07188_);
  and _15660_ (_07360_, _07307_, _07359_);
  nor _15661_ (_07361_, _07360_, _07358_);
  nor _15662_ (_14295_, _07361_, rst);
  and _15663_ (_07362_, _07321_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  and _15664_ (_07363_, _07325_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  nor _15665_ (_07364_, _07363_, _07362_);
  and _15666_ (_07365_, _07327_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  and _15667_ (_07366_, _07333_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  nor _15668_ (_07367_, _07366_, _07365_);
  and _15669_ (_07368_, _07367_, _07364_);
  and _15670_ (_07369_, _07313_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  and _15671_ (_07370_, _07331_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  nor _15672_ (_07371_, _07370_, _07369_);
  and _15673_ (_07372_, _07309_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  and _15674_ (_07373_, _07318_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  nor _15675_ (_07374_, _07373_, _07372_);
  and _15676_ (_07375_, _07374_, _07371_);
  and _15677_ (_07376_, _07375_, _07368_);
  nor _15678_ (_07377_, _07376_, _07307_);
  not _15679_ (_07378_, _06666_);
  and _15680_ (_07379_, _07307_, _07378_);
  nor _15681_ (_07380_, _07379_, _07377_);
  nor _15682_ (_01145_, _07380_, rst);
  nor _15683_ (_07381_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  nor _15684_ (_07382_, _07381_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf );
  not _15685_ (_07383_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  and _15686_ (_07384_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  and _15687_ (_07385_, _07077_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  nor _15688_ (_07386_, _07385_, _07384_);
  nor _15689_ (_07387_, _07386_, _07076_);
  or _15690_ (_07388_, _07387_, _07383_);
  and _15691_ (_07389_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], _07077_);
  and _15692_ (_07390_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  nor _15693_ (_07391_, _07390_, _07389_);
  nor _15694_ (_07392_, _07391_, _07076_);
  and _15695_ (_07393_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and _15696_ (_07394_, _07077_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  nor _15697_ (_07396_, _07394_, _07393_);
  nand _15698_ (_07397_, _07396_, _07392_);
  or _15699_ (_07398_, _07397_, _07388_);
  and _15700_ (_07399_, _07398_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or _15701_ (_07400_, _07399_, _07382_);
  and _15702_ (_07401_, _06364_, _06350_);
  and _15703_ (_07402_, _07401_, _06940_);
  nor _15704_ (_07403_, _06675_, _06394_);
  and _15705_ (_07404_, _07403_, _06933_);
  and _15706_ (_07405_, _07404_, _07402_);
  or _15707_ (_07406_, _07405_, _07400_);
  and _15708_ (_07407_, _07402_, _06945_);
  not _15709_ (_07408_, _07407_);
  and _15710_ (_07409_, _07408_, _07406_);
  nand _15711_ (_07410_, _07405_, _06930_);
  and _15712_ (_07411_, _07410_, _07409_);
  nor _15713_ (_07412_, _07408_, _06978_);
  or _15714_ (_07413_, _07412_, _07411_);
  and _15715_ (_01342_, _07413_, _06444_);
  and _15716_ (_07414_, _07153_, _07043_);
  nor _15717_ (_07415_, _07159_, _07414_);
  and _15718_ (_07416_, _07153_, _07147_);
  not _15719_ (_07417_, _07416_);
  and _15720_ (_07418_, _07155_, _07417_);
  and _15721_ (_07419_, _07418_, _07415_);
  or _15722_ (_07420_, _07419_, _07158_);
  and _15723_ (_07421_, _07420_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  and _15724_ (_07422_, _07153_, _06431_);
  and _15725_ (_07423_, _06439_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  and _15726_ (_07424_, _07423_, _07422_);
  and _15727_ (_07425_, _07151_, _06439_);
  and _15728_ (_07426_, _07425_, _07340_);
  or _15729_ (_07427_, _07426_, _07424_);
  or _15730_ (_07428_, _07427_, _07421_);
  and _15731_ (_01560_, _07428_, _06444_);
  not _15732_ (_07429_, _07230_);
  nor _15733_ (_07430_, _07253_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor _15734_ (_07431_, _07430_, _07429_);
  nor _15735_ (_07432_, _07431_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  and _15736_ (_07433_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  not _15737_ (_07434_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  nor _15738_ (_07435_, _07432_, _07434_);
  or _15739_ (_07436_, _07435_, _07433_);
  and _15740_ (_01936_, _07436_, _06444_);
  not _15741_ (_07437_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and _15742_ (_07438_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], _06308_);
  and _15743_ (_07439_, _07438_, _07437_);
  and _15744_ (_07440_, _06795_, _06640_);
  and _15745_ (_07441_, _06913_, _06958_);
  and _15746_ (_07442_, _06955_, _06697_);
  and _15747_ (_07443_, _07442_, _06824_);
  and _15748_ (_07444_, _07443_, _06465_);
  nor _15749_ (_07445_, _06824_, _06697_);
  and _15750_ (_07446_, _07445_, _06960_);
  and _15751_ (_07447_, _07446_, _06515_);
  nor _15752_ (_07448_, _07447_, _07444_);
  nor _15753_ (_07450_, _07448_, _06795_);
  and _15754_ (_07451_, _07448_, _06795_);
  nor _15755_ (_07453_, _07451_, _07450_);
  nor _15756_ (_07454_, _07453_, _06621_);
  nor _15757_ (_07456_, _06570_, _06951_);
  or _15758_ (_07457_, _07456_, _07454_);
  or _15759_ (_07458_, _07457_, _07441_);
  and _15760_ (_07459_, _06639_, _06632_);
  nor _15761_ (_07460_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nand _15762_ (_07461_, _07460_, _06697_);
  nor _15763_ (_07462_, _07460_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7]);
  not _15764_ (_07463_, _07462_);
  and _15765_ (_07464_, _07463_, _07461_);
  not _15766_ (_07465_, _07464_);
  or _15767_ (_07466_, _06806_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand _15768_ (_07467_, _06785_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  and _15769_ (_07468_, _07467_, _07466_);
  or _15770_ (_07470_, _07468_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not _15771_ (_07471_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not _15772_ (_07472_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand _15773_ (_07473_, _06752_, _07472_);
  nand _15774_ (_07474_, _06739_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  and _15775_ (_07475_, _07474_, _07473_);
  or _15776_ (_07476_, _07475_, _07471_);
  and _15777_ (_07477_, _07476_, _07470_);
  nor _15778_ (_07478_, _07477_, _07465_);
  and _15779_ (_07479_, _07477_, _07465_);
  nand _15780_ (_07480_, _07460_, _06732_);
  nor _15781_ (_07481_, _07460_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6]);
  not _15782_ (_07482_, _07481_);
  and _15783_ (_07483_, _07482_, _07480_);
  not _15784_ (_07484_, _07483_);
  and _15785_ (_07486_, _06795_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or _15786_ (_07487_, _07486_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nand _15787_ (_07488_, _06775_, _07472_);
  nand _15788_ (_07489_, _06482_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  and _15789_ (_07490_, _07489_, _07488_);
  or _15790_ (_07491_, _07490_, _07471_);
  and _15791_ (_07492_, _07491_, _07487_);
  or _15792_ (_07493_, _07492_, _07484_);
  nor _15793_ (_07495_, _07493_, _07479_);
  nor _15794_ (_07496_, _07495_, _07478_);
  nor _15795_ (_07497_, _07479_, _07478_);
  nand _15796_ (_07499_, _07492_, _07484_);
  and _15797_ (_07500_, _07499_, _07493_);
  and _15798_ (_07501_, _07500_, _07497_);
  nand _15799_ (_07502_, _07460_, _06511_);
  nor _15800_ (_07503_, _07460_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5]);
  not _15801_ (_07504_, _07503_);
  and _15802_ (_07505_, _07504_, _07502_);
  not _15803_ (_07506_, _07505_);
  and _15804_ (_07507_, _06806_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or _15805_ (_07508_, _07507_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nand _15806_ (_07509_, _06785_, _07472_);
  nand _15807_ (_07510_, _06752_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  and _15808_ (_07511_, _07510_, _07509_);
  or _15809_ (_07512_, _07511_, _07471_);
  and _15810_ (_07513_, _07512_, _07508_);
  nor _15811_ (_07515_, _07513_, _07506_);
  not _15812_ (_07516_, _07515_);
  or _15813_ (_07517_, _06795_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand _15814_ (_07518_, _06775_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  and _15815_ (_07519_, _07518_, _07517_);
  and _15816_ (_07520_, _07519_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not _15817_ (_07521_, _07520_);
  nor _15818_ (_07522_, _07460_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4]);
  not _15819_ (_07523_, _07522_);
  nand _15820_ (_07524_, _07460_, _06532_);
  and _15821_ (_07525_, _07524_, _07523_);
  and _15822_ (_07526_, _07525_, _07521_);
  and _15823_ (_07527_, _07513_, _07506_);
  nor _15824_ (_07528_, _07527_, _07515_);
  nand _15825_ (_07529_, _07528_, _07526_);
  nand _15826_ (_07530_, _07529_, _07516_);
  nand _15827_ (_07531_, _07530_, _07501_);
  and _15828_ (_07532_, _07531_, _07496_);
  and _15829_ (_07533_, _07468_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nor _15830_ (_07534_, _07460_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3]);
  not _15831_ (_07535_, _07534_);
  nand _15832_ (_07536_, _07460_, _06551_);
  and _15833_ (_07537_, _07536_, _07535_);
  not _15834_ (_07538_, _07537_);
  or _15835_ (_07539_, _07538_, _07533_);
  not _15836_ (_07540_, _07533_);
  or _15837_ (_07541_, _07537_, _07540_);
  nand _15838_ (_07542_, _07541_, _07539_);
  and _15839_ (_07543_, _07486_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not _15840_ (_07544_, _07543_);
  nand _15841_ (_07545_, _07460_, _06604_);
  nor _15842_ (_07546_, _07460_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2]);
  not _15843_ (_07547_, _07546_);
  and _15844_ (_07548_, _07547_, _07545_);
  nand _15845_ (_07549_, _07548_, _07544_);
  and _15846_ (_07550_, _07507_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not _15847_ (_07551_, _07550_);
  nand _15848_ (_07552_, _07460_, _06570_);
  nor _15849_ (_07553_, _07460_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1]);
  not _15850_ (_07554_, _07553_);
  and _15851_ (_07555_, _07554_, _07552_);
  nor _15852_ (_07556_, _07555_, _07551_);
  or _15853_ (_07557_, _07548_, _07544_);
  nand _15854_ (_07558_, _07557_, _07549_);
  or _15855_ (_07559_, _07558_, _07556_);
  and _15856_ (_07560_, _07559_, _07549_);
  or _15857_ (_07561_, _07560_, _07542_);
  nand _15858_ (_07562_, _07561_, _07539_);
  not _15859_ (_07564_, _07525_);
  and _15860_ (_07565_, _07564_, _07520_);
  nor _15861_ (_07566_, _07565_, _07526_);
  and _15862_ (_07567_, _07528_, _07566_);
  and _15863_ (_07568_, _07567_, _07501_);
  nand _15864_ (_07569_, _07568_, _07562_);
  nand _15865_ (_07570_, _07569_, _07532_);
  nor _15866_ (_07571_, _07519_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and _15867_ (_07572_, _06482_, _07472_);
  and _15868_ (_07573_, _06704_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _15869_ (_07574_, _07573_, _07572_);
  nor _15870_ (_07575_, _07574_, _07471_);
  nor _15871_ (_07576_, _07575_, _07571_);
  not _15872_ (_07577_, _07576_);
  and _15873_ (_07578_, _06739_, _06704_);
  nor _15874_ (_07579_, _07578_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _15875_ (_07580_, _07490_, _07475_);
  nor _15876_ (_07581_, _07574_, _07511_);
  and _15877_ (_07582_, _07581_, _07580_);
  nor _15878_ (_07583_, _07582_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nor _15879_ (_07584_, _07583_, _07579_);
  and _15880_ (_07585_, _07584_, _07577_);
  and _15881_ (_07586_, _07585_, _07570_);
  and _15882_ (_07587_, _07586_, _07459_);
  nor _15883_ (_07588_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  not _15884_ (_07589_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and _15885_ (_07590_, _07589_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _15886_ (_07591_, _07590_, _07588_);
  not _15887_ (_07592_, _07591_);
  nor _15888_ (_07593_, _07592_, _06879_);
  nor _15889_ (_07594_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  not _15890_ (_07595_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and _15891_ (_07596_, _07595_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _15892_ (_07597_, _07596_, _07594_);
  nor _15893_ (_07598_, _07597_, _07593_);
  and _15894_ (_07599_, _07597_, _07593_);
  nor _15895_ (_07600_, _07599_, _07598_);
  and _15896_ (_07601_, _07600_, _06847_);
  and _15897_ (_07602_, _06628_, _06452_);
  not _15898_ (_07603_, _06570_);
  nor _15899_ (_07604_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  nand _15900_ (_07605_, _07604_, _06704_);
  not _15901_ (_07606_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  or _15902_ (_07607_, _07606_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  or _15903_ (_07608_, _07607_, _06482_);
  not _15904_ (_07609_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  or _15905_ (_07610_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], _07609_);
  or _15906_ (_07611_, _07610_, _06775_);
  and _15907_ (_07612_, _07611_, _07608_);
  and _15908_ (_07613_, _07610_, _07607_);
  or _15909_ (_07614_, _06795_, _07609_);
  nand _15910_ (_07615_, _07614_, _07613_);
  nand _15911_ (_07616_, _07615_, _07612_);
  and _15912_ (_07617_, _07616_, _07605_);
  and _15913_ (_07618_, _07617_, _07603_);
  nand _15914_ (_07619_, _07604_, _06739_);
  or _15915_ (_07620_, _07607_, _06752_);
  or _15916_ (_07621_, _07610_, _06785_);
  and _15917_ (_07622_, _07621_, _07620_);
  or _15918_ (_07624_, _06806_, _07609_);
  nand _15919_ (_07625_, _07624_, _07613_);
  nand _15920_ (_07626_, _07625_, _07622_);
  and _15921_ (_07627_, _07626_, _07619_);
  and _15922_ (_07628_, _07627_, _06903_);
  and _15923_ (_07629_, _07628_, _07618_);
  nand _15924_ (_07630_, _07626_, _07619_);
  or _15925_ (_07631_, _07630_, _06570_);
  and _15926_ (_07632_, _07617_, _06903_);
  not _15927_ (_07633_, _07632_);
  and _15928_ (_07634_, _07633_, _07631_);
  nor _15929_ (_07635_, _07634_, _07629_);
  and _15930_ (_07636_, _07635_, _07602_);
  or _15931_ (_07637_, _07636_, _07601_);
  or _15932_ (_07638_, _07637_, _07587_);
  or _15933_ (_07639_, _07638_, _07458_);
  nor _15934_ (_07640_, _07639_, _07440_);
  and _15935_ (_07641_, _07640_, _07439_);
  not _15936_ (_07642_, _07641_);
  not _15937_ (_07643_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1]);
  and _15938_ (_07644_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], _06308_);
  and _15939_ (_07646_, _07644_, _07643_);
  and _15940_ (_07647_, _06671_, _06336_);
  and _15941_ (_07649_, _07647_, _07216_);
  and _15942_ (_07650_, _07649_, _07150_);
  and _15943_ (_07651_, _07650_, _06440_);
  nor _15944_ (_07652_, _07651_, _07646_);
  not _15945_ (_07653_, _07652_);
  nor _15946_ (_07654_, _07586_, _07465_);
  not _15947_ (_07655_, _07654_);
  not _15948_ (_07656_, _07500_);
  and _15949_ (_07657_, _07566_, _07562_);
  nor _15950_ (_07659_, _07657_, _07526_);
  or _15951_ (_07660_, _07659_, _07527_);
  and _15952_ (_07661_, _07660_, _07516_);
  or _15953_ (_07662_, _07661_, _07656_);
  and _15954_ (_07664_, _07662_, _07493_);
  nand _15955_ (_07665_, _07664_, _07497_);
  or _15956_ (_07666_, _07664_, _07497_);
  nand _15957_ (_07667_, _07666_, _07665_);
  nand _15958_ (_07668_, _07667_, _07586_);
  and _15959_ (_07669_, _07668_, _07655_);
  or _15960_ (_07670_, _07669_, _07576_);
  nand _15961_ (_07671_, _07669_, _07576_);
  not _15962_ (_07672_, _07477_);
  not _15963_ (_07673_, _07586_);
  and _15964_ (_07674_, _07661_, _07656_);
  not _15965_ (_07675_, _07674_);
  and _15966_ (_07676_, _07675_, _07662_);
  nor _15967_ (_07677_, _07676_, _07673_);
  nor _15968_ (_07679_, _07586_, _07483_);
  nor _15969_ (_07680_, _07679_, _07677_);
  and _15970_ (_07681_, _07680_, _07672_);
  nand _15971_ (_07682_, _07681_, _07671_);
  and _15972_ (_07683_, _07682_, _07670_);
  and _15973_ (_07684_, _07671_, _07670_);
  nor _15974_ (_07685_, _07680_, _07672_);
  nor _15975_ (_07686_, _07685_, _07681_);
  and _15976_ (_07687_, _07686_, _07684_);
  not _15977_ (_07688_, _07492_);
  nor _15978_ (_07689_, _07528_, _07659_);
  and _15979_ (_07690_, _07528_, _07659_);
  or _15980_ (_07691_, _07690_, _07689_);
  nor _15981_ (_07692_, _07691_, _07673_);
  nor _15982_ (_07693_, _07586_, _07505_);
  nor _15983_ (_07694_, _07693_, _07692_);
  and _15984_ (_07695_, _07694_, _07688_);
  not _15985_ (_07696_, _07513_);
  nor _15986_ (_07697_, _07566_, _07562_);
  or _15987_ (_07698_, _07697_, _07657_);
  and _15988_ (_07699_, _07698_, _07586_);
  nor _15989_ (_07700_, _07586_, _07525_);
  nor _15990_ (_07701_, _07700_, _07699_);
  and _15991_ (_07703_, _07701_, _07696_);
  not _15992_ (_07704_, _07703_);
  nor _15993_ (_07706_, _07694_, _07688_);
  or _15994_ (_07707_, _07695_, _07706_);
  nor _15995_ (_07708_, _07707_, _07704_);
  nor _15996_ (_07709_, _07708_, _07695_);
  not _15997_ (_07711_, _07709_);
  nor _15998_ (_07712_, _07586_, _07538_);
  and _15999_ (_07713_, _07560_, _07542_);
  not _16000_ (_07714_, _07713_);
  and _16001_ (_07715_, _07714_, _07561_);
  and _16002_ (_07716_, _07715_, _07586_);
  or _16003_ (_07717_, _07716_, _07712_);
  nor _16004_ (_07718_, _07717_, _07521_);
  not _16005_ (_07719_, _07718_);
  nand _16006_ (_07720_, _07673_, _07555_);
  nor _16007_ (_07721_, _07555_, _07550_);
  and _16008_ (_07722_, _07555_, _07550_);
  nor _16009_ (_07723_, _07722_, _07721_);
  nand _16010_ (_07724_, _07586_, _07723_);
  nand _16011_ (_07725_, _07724_, _07720_);
  nand _16012_ (_07726_, _07725_, _07544_);
  or _16013_ (_07727_, _07725_, _07544_);
  nand _16014_ (_07728_, _07727_, _07726_);
  nor _16015_ (_07729_, _07460_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0]);
  and _16016_ (_07730_, _07460_, _06587_);
  nor _16017_ (_07731_, _07730_, _07729_);
  nor _16018_ (_07732_, _07731_, _07551_);
  or _16019_ (_07733_, _07732_, _07728_);
  and _16020_ (_07734_, _07733_, _07726_);
  or _16021_ (_07735_, _07586_, _07548_);
  and _16022_ (_07736_, _07558_, _07556_);
  not _16023_ (_07737_, _07736_);
  and _16024_ (_07738_, _07737_, _07559_);
  or _16025_ (_07739_, _07738_, _07673_);
  and _16026_ (_07740_, _07739_, _07735_);
  and _16027_ (_07741_, _07740_, _07540_);
  nor _16028_ (_07742_, _07740_, _07540_);
  or _16029_ (_07743_, _07742_, _07741_);
  or _16030_ (_07744_, _07743_, _07734_);
  and _16031_ (_07745_, _07717_, _07521_);
  nor _16032_ (_07746_, _07745_, _07741_);
  nand _16033_ (_07747_, _07746_, _07744_);
  and _16034_ (_07748_, _07747_, _07719_);
  nor _16035_ (_07749_, _07701_, _07696_);
  nor _16036_ (_07750_, _07749_, _07703_);
  not _16037_ (_07751_, _07750_);
  nor _16038_ (_07752_, _07707_, _07751_);
  and _16039_ (_07753_, _07752_, _07748_);
  or _16040_ (_07754_, _07753_, _07711_);
  nand _16041_ (_07755_, _07754_, _07687_);
  nand _16042_ (_07756_, _07755_, _07683_);
  and _16043_ (_07757_, _07756_, _07584_);
  not _16044_ (_07758_, _07757_);
  and _16045_ (_07760_, _07732_, _07728_);
  not _16046_ (_07761_, _07760_);
  and _16047_ (_07762_, _07761_, _07733_);
  or _16048_ (_07763_, _07762_, _07758_);
  or _16049_ (_07764_, _07757_, _07725_);
  and _16050_ (_07765_, _07764_, _07763_);
  nand _16051_ (_07766_, _07765_, _07459_);
  not _16052_ (_07767_, _07604_);
  and _16053_ (_07768_, _07767_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6]);
  and _16054_ (_07769_, _07617_, _06534_);
  and _16055_ (_07770_, _07627_, _06552_);
  and _16056_ (_07771_, _07770_, _07769_);
  and _16057_ (_07772_, _07627_, _06534_);
  and _16058_ (_07773_, _07617_, _06958_);
  nand _16059_ (_07774_, _07773_, _07772_);
  and _16060_ (_07775_, _07627_, _06958_);
  or _16061_ (_07776_, _07775_, _07769_);
  and _16062_ (_07777_, _07776_, _07774_);
  and _16063_ (_07778_, _07777_, _07771_);
  or _16064_ (_07779_, _07774_, _06732_);
  and _16065_ (_07780_, _07627_, _06957_);
  not _16066_ (_07781_, _07780_);
  nand _16067_ (_07782_, _07781_, _07774_);
  and _16068_ (_07783_, _07782_, _07779_);
  nand _16069_ (_07784_, _07783_, _07773_);
  or _16070_ (_07785_, _07780_, _07773_);
  and _16071_ (_07786_, _07785_, _07784_);
  nand _16072_ (_07787_, _07786_, _07778_);
  not _16073_ (_07788_, _07787_);
  not _16074_ (_07789_, _07779_);
  and _16075_ (_07790_, _07783_, _07773_);
  or _16076_ (_07791_, _07630_, _06697_);
  nand _16077_ (_07792_, _07616_, _07605_);
  or _16078_ (_07793_, _07792_, _06732_);
  or _16079_ (_07794_, _07793_, _07791_);
  nand _16080_ (_07795_, _07793_, _07791_);
  and _16081_ (_07796_, _07795_, _07794_);
  nand _16082_ (_07797_, _07796_, _07790_);
  or _16083_ (_07798_, _07796_, _07790_);
  and _16084_ (_07799_, _07798_, _07797_);
  nand _16085_ (_07800_, _07799_, _07789_);
  or _16086_ (_07801_, _07799_, _07789_);
  and _16087_ (_07802_, _07801_, _07800_);
  nand _16088_ (_07803_, _07802_, _07788_);
  or _16089_ (_07804_, _07802_, _07788_);
  nand _16090_ (_07805_, _07804_, _07803_);
  not _16091_ (_07806_, _07805_);
  and _16092_ (_07807_, _07627_, _06605_);
  nand _16093_ (_07808_, _07807_, _07618_);
  and _16094_ (_07810_, _07617_, _06605_);
  and _16095_ (_07811_, _07810_, _07631_);
  nand _16096_ (_07812_, _07811_, _07770_);
  nand _16097_ (_07813_, _07812_, _07808_);
  not _16098_ (_07814_, _07771_);
  and _16099_ (_07815_, _07617_, _06552_);
  or _16100_ (_07816_, _07815_, _07772_);
  and _16101_ (_07817_, _07816_, _07814_);
  nand _16102_ (_07818_, _07817_, _07813_);
  not _16103_ (_07819_, _07818_);
  not _16104_ (_07820_, _07778_);
  or _16105_ (_07821_, _07777_, _07771_);
  and _16106_ (_07822_, _07821_, _07820_);
  and _16107_ (_07823_, _07822_, _07819_);
  or _16108_ (_07825_, _07786_, _07778_);
  and _16109_ (_07826_, _07825_, _07787_);
  nand _16110_ (_07827_, _07826_, _07823_);
  or _16111_ (_07828_, _07807_, _07618_);
  and _16112_ (_07829_, _07828_, _07808_);
  and _16113_ (_07830_, _07829_, _07629_);
  or _16114_ (_07831_, _07811_, _07770_);
  and _16115_ (_07832_, _07831_, _07812_);
  nand _16116_ (_07833_, _07832_, _07830_);
  not _16117_ (_07834_, _07833_);
  or _16118_ (_07835_, _07817_, _07813_);
  and _16119_ (_07836_, _07835_, _07818_);
  nand _16120_ (_07837_, _07836_, _07834_);
  not _16121_ (_07838_, _07837_);
  nand _16122_ (_07839_, _07822_, _07819_);
  or _16123_ (_07840_, _07822_, _07819_);
  and _16124_ (_07841_, _07840_, _07839_);
  nand _16125_ (_07842_, _07841_, _07838_);
  not _16126_ (_07843_, _07842_);
  or _16127_ (_07844_, _07826_, _07823_);
  and _16128_ (_07845_, _07844_, _07827_);
  nand _16129_ (_07846_, _07845_, _07843_);
  nand _16130_ (_07847_, _07846_, _07827_);
  nand _16131_ (_07848_, _07847_, _07806_);
  nand _16132_ (_07850_, _07848_, _07803_);
  and _16133_ (_07851_, _07617_, _06914_);
  and _16134_ (_07853_, _07851_, _07781_);
  and _16135_ (_07854_, _07800_, _07797_);
  not _16136_ (_07856_, _07854_);
  nand _16137_ (_07857_, _07856_, _07853_);
  or _16138_ (_07858_, _07856_, _07853_);
  and _16139_ (_07859_, _07858_, _07857_);
  nand _16140_ (_07861_, _07859_, _07850_);
  or _16141_ (_07862_, _07859_, _07850_);
  and _16142_ (_07864_, _07862_, _07861_);
  nand _16143_ (_07865_, _07864_, _07768_);
  and _16144_ (_07866_, _07767_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5]);
  or _16145_ (_07868_, _07847_, _07806_);
  and _16146_ (_07869_, _07868_, _07848_);
  nand _16147_ (_07870_, _07869_, _07866_);
  or _16148_ (_07871_, _07869_, _07866_);
  nand _16149_ (_07872_, _07871_, _07870_);
  and _16150_ (_07873_, _07767_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4]);
  or _16151_ (_07874_, _07845_, _07843_);
  and _16152_ (_07875_, _07874_, _07846_);
  nand _16153_ (_07877_, _07875_, _07873_);
  or _16154_ (_07879_, _07875_, _07873_);
  nand _16155_ (_07880_, _07879_, _07877_);
  and _16156_ (_07881_, _07767_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3]);
  or _16157_ (_07882_, _07841_, _07838_);
  and _16158_ (_07883_, _07882_, _07842_);
  nand _16159_ (_07884_, _07883_, _07881_);
  or _16160_ (_07885_, _07883_, _07881_);
  and _16161_ (_07886_, _07885_, _07884_);
  and _16162_ (_07887_, _07767_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2]);
  or _16163_ (_07888_, _07836_, _07834_);
  and _16164_ (_07889_, _07888_, _07837_);
  nand _16165_ (_07890_, _07889_, _07887_);
  and _16166_ (_07891_, _07767_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1]);
  or _16167_ (_07892_, _07832_, _07830_);
  and _16168_ (_07893_, _07892_, _07833_);
  nand _16169_ (_07894_, _07893_, _07891_);
  and _16170_ (_07895_, _07767_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0]);
  nand _16171_ (_07896_, _07829_, _07629_);
  or _16172_ (_07897_, _07829_, _07629_);
  and _16173_ (_07898_, _07897_, _07896_);
  and _16174_ (_07899_, _07898_, _07895_);
  or _16175_ (_07900_, _07893_, _07891_);
  and _16176_ (_07901_, _07900_, _07894_);
  nand _16177_ (_07902_, _07901_, _07899_);
  nand _16178_ (_07903_, _07902_, _07894_);
  or _16179_ (_07904_, _07889_, _07887_);
  and _16180_ (_07905_, _07904_, _07890_);
  nand _16181_ (_07906_, _07905_, _07903_);
  nand _16182_ (_07907_, _07906_, _07890_);
  nand _16183_ (_07908_, _07907_, _07886_);
  and _16184_ (_07910_, _07908_, _07884_);
  or _16185_ (_07911_, _07910_, _07880_);
  and _16186_ (_07912_, _07911_, _07877_);
  or _16187_ (_07913_, _07912_, _07872_);
  and _16188_ (_07914_, _07913_, _07870_);
  or _16189_ (_07915_, _07864_, _07768_);
  nand _16190_ (_07916_, _07915_, _07865_);
  or _16191_ (_07917_, _07916_, _07914_);
  and _16192_ (_07918_, _07917_, _07865_);
  and _16193_ (_07919_, _07767_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7]);
  and _16194_ (_07920_, _07857_, _07794_);
  nand _16195_ (_07921_, _07920_, _07861_);
  nand _16196_ (_07922_, _07921_, _07919_);
  or _16197_ (_07923_, _07921_, _07919_);
  nand _16198_ (_07924_, _07923_, _07922_);
  or _16199_ (_07925_, _07924_, _07918_);
  nand _16200_ (_07926_, _07924_, _07918_);
  and _16201_ (_07927_, _07926_, _07925_);
  nand _16202_ (_07928_, _07927_, _07602_);
  nor _16203_ (_07929_, _06828_, _06823_);
  nor _16204_ (_07930_, _07929_, _06829_);
  nor _16205_ (_07931_, _07930_, _06681_);
  not _16206_ (_07932_, _07931_);
  not _16207_ (_07933_, _06641_);
  nor _16208_ (_07935_, _07933_, _06604_);
  not _16209_ (_07936_, _07935_);
  and _16210_ (_07937_, _06640_, _07603_);
  nor _16211_ (_07938_, _06638_, _06587_);
  nor _16212_ (_07939_, _07938_, _07937_);
  and _16213_ (_07940_, _07939_, _07936_);
  and _16214_ (_07941_, _07940_, _07067_);
  and _16215_ (_07942_, _07941_, _07056_);
  nor _16216_ (_07943_, _06884_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and _16217_ (_07944_, _07943_, _07603_);
  nor _16218_ (_07945_, _07943_, _07603_);
  nor _16219_ (_07946_, _07945_, _07944_);
  nor _16220_ (_07947_, _07946_, _06891_);
  nor _16221_ (_07948_, _06825_, _06799_);
  or _16222_ (_07949_, _07948_, _06854_);
  and _16223_ (_07950_, _07949_, _06861_);
  nor _16224_ (_07951_, _07949_, _06861_);
  or _16225_ (_07952_, _07951_, _07950_);
  and _16226_ (_07953_, _07952_, _06847_);
  nor _16227_ (_07955_, _07953_, _07947_);
  and _16228_ (_07956_, _07955_, _07942_);
  and _16229_ (_07957_, _07956_, _07932_);
  and _16230_ (_07958_, _07957_, _07928_);
  nand _16231_ (_07959_, _07958_, _07766_);
  nand _16232_ (_07960_, _07959_, _07653_);
  not _16233_ (_07961_, _07439_);
  and _16234_ (_07962_, _06940_, _06394_);
  nor _16235_ (_07963_, _06364_, _06350_);
  and _16236_ (_07965_, _07963_, _06674_);
  and _16237_ (_07966_, _07965_, _07962_);
  and _16238_ (_07967_, _07966_, _06432_);
  and _16239_ (_07968_, _07967_, _06930_);
  nor _16240_ (_07969_, _07967_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or _16241_ (_07971_, _07969_, _07653_);
  or _16242_ (_07972_, _07971_, _07968_);
  and _16243_ (_07974_, _07972_, _07961_);
  nand _16244_ (_07975_, _07974_, _07960_);
  and _16245_ (_07976_, _07975_, _07642_);
  and _16246_ (_06429_, _07976_, _06444_);
  not _16247_ (_07978_, _07731_);
  and _16248_ (_07979_, _07757_, _07550_);
  nor _16249_ (_07980_, _07979_, _07978_);
  and _16250_ (_07981_, _07979_, _07978_);
  or _16251_ (_07982_, _07981_, _07980_);
  nand _16252_ (_07984_, _07982_, _07459_);
  not _16253_ (_07985_, _07917_);
  and _16254_ (_07986_, _07916_, _07914_);
  nor _16255_ (_07987_, _07986_, _07985_);
  and _16256_ (_07988_, _07987_, _07602_);
  nor _16257_ (_07989_, _06827_, _06465_);
  nor _16258_ (_07990_, _07989_, _06861_);
  not _16259_ (_07991_, _07990_);
  nor _16260_ (_07993_, _06847_, _06680_);
  nor _16261_ (_07994_, _07993_, _07991_);
  not _16262_ (_07995_, _07994_);
  nor _16263_ (_07996_, _06825_, _06898_);
  nor _16264_ (_07997_, _07996_, _06654_);
  or _16265_ (_07998_, _07997_, _06826_);
  and _16266_ (_07999_, _06825_, _06658_);
  and _16267_ (_08000_, _06806_, _06455_);
  or _16268_ (_08001_, _06660_, _06620_);
  and _16269_ (_08002_, _08001_, _06587_);
  or _16270_ (_08003_, _08002_, _08000_);
  nor _16271_ (_08004_, _08003_, _07999_);
  and _16272_ (_08005_, _06914_, _06907_);
  and _16273_ (_08006_, _06913_, _06465_);
  nor _16274_ (_08007_, _08006_, _08005_);
  or _16275_ (_08008_, _07933_, _06570_);
  nor _16276_ (_08009_, _06883_, _06640_);
  nor _16277_ (_08010_, _08009_, _06587_);
  not _16278_ (_08011_, _08010_);
  and _16279_ (_08012_, _08011_, _08008_);
  and _16280_ (_08013_, _08012_, _08007_);
  and _16281_ (_08014_, _08013_, _08004_);
  and _16282_ (_08015_, _08014_, _07998_);
  and _16283_ (_08016_, _08015_, _07995_);
  not _16284_ (_08017_, _08016_);
  nor _16285_ (_08018_, _08017_, _07988_);
  nand _16286_ (_08019_, _08018_, _07984_);
  nand _16287_ (_08020_, _08019_, _07653_);
  not _16288_ (_08021_, _06942_);
  nor _16289_ (_08022_, _06930_, _08021_);
  nor _16290_ (_08023_, _06942_, _06803_);
  nor _16291_ (_08024_, _08023_, _08022_);
  or _16292_ (_08025_, _07646_, _07439_);
  nor _16293_ (_08026_, _08025_, _07651_);
  and _16294_ (_08027_, _08026_, _07966_);
  not _16295_ (_08028_, _08027_);
  nor _16296_ (_08029_, _08028_, _08024_);
  not _16297_ (_08030_, _06380_);
  and _16298_ (_08031_, _06394_, _06336_);
  and _16299_ (_08032_, _08031_, _07963_);
  and _16300_ (_08033_, _08032_, _08030_);
  and _16301_ (_08034_, _08033_, _06674_);
  not _16302_ (_08035_, _08034_);
  and _16303_ (_08036_, _08035_, _08026_);
  and _16304_ (_08037_, _08036_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or _16305_ (_08038_, _08037_, _07439_);
  nor _16306_ (_08039_, _08038_, _08029_);
  nand _16307_ (_08040_, _08039_, _08020_);
  and _16308_ (_08041_, _06806_, _06640_);
  and _16309_ (_08042_, _06913_, _06534_);
  nor _16310_ (_08043_, _06948_, _06892_);
  and _16311_ (_08044_, _08043_, _06962_);
  nor _16312_ (_08045_, _08044_, _06806_);
  and _16313_ (_08046_, _08044_, _06806_);
  nor _16314_ (_08047_, _08046_, _08045_);
  and _16315_ (_08048_, _08047_, _06620_);
  nor _16316_ (_08049_, _06587_, _06951_);
  or _16317_ (_08050_, _08049_, _08048_);
  or _16318_ (_08051_, _08050_, _08042_);
  and _16319_ (_08052_, _07757_, _07459_);
  and _16320_ (_08053_, _07592_, _06879_);
  nor _16321_ (_08054_, _08053_, _07593_);
  and _16322_ (_08055_, _08054_, _06847_);
  and _16323_ (_08056_, _07628_, _07602_);
  or _16324_ (_08057_, _08056_, _08055_);
  or _16325_ (_08058_, _08057_, _08052_);
  or _16326_ (_08059_, _08058_, _08051_);
  nor _16327_ (_08060_, _08059_, _08041_);
  and _16328_ (_08061_, _08060_, _07439_);
  not _16329_ (_08062_, _08061_);
  and _16330_ (_08063_, _08062_, _08040_);
  and _16331_ (_06433_, _08063_, _06444_);
  and _16332_ (_08064_, _07231_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  and _16333_ (_08065_, _08064_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  not _16334_ (_08066_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  nor _16335_ (_08067_, _08064_, _08066_);
  or _16336_ (_08069_, _08067_, _08065_);
  and _16337_ (_06473_, _08069_, _06444_);
  and _16338_ (_08070_, _07758_, _07694_);
  nand _16339_ (_08071_, _07750_, _07748_);
  nand _16340_ (_08072_, _08071_, _07704_);
  nor _16341_ (_08073_, _08072_, _07707_);
  and _16342_ (_08074_, _08072_, _07707_);
  or _16343_ (_08076_, _08074_, _08073_);
  and _16344_ (_08077_, _08076_, _07757_);
  or _16345_ (_08078_, _08077_, _08070_);
  and _16346_ (_08079_, _08078_, _07459_);
  or _16347_ (_08080_, _07924_, _07865_);
  nand _16348_ (_08081_, _08080_, _07922_);
  and _16349_ (_08082_, _07767_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8]);
  and _16350_ (_08083_, _07767_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  and _16351_ (_08084_, _08083_, _08082_);
  and _16352_ (_08085_, _08084_, _08081_);
  nor _16353_ (_08086_, _07924_, _07916_);
  nand _16354_ (_08087_, _08084_, _08086_);
  nor _16355_ (_08088_, _08087_, _07914_);
  or _16356_ (_08089_, _08088_, _08085_);
  and _16357_ (_08090_, _07767_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10]);
  and _16358_ (_08091_, _07767_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  and _16359_ (_08092_, _08091_, _08090_);
  nand _16360_ (_08093_, _08092_, _08089_);
  nand _16361_ (_08094_, _08089_, _08090_);
  not _16362_ (_08095_, _08091_);
  nand _16363_ (_08096_, _08095_, _08094_);
  and _16364_ (_08097_, _08096_, _08093_);
  and _16365_ (_08098_, _08097_, _07602_);
  nor _16366_ (_08099_, _06765_, _06650_);
  nor _16367_ (_08100_, _08099_, _06850_);
  or _16368_ (_08101_, _08100_, _06871_);
  nor _16369_ (_08102_, _06872_, _06848_);
  and _16370_ (_08103_, _08102_, _08101_);
  nor _16371_ (_08104_, _06839_, _06764_);
  or _16372_ (_08105_, _08104_, _06840_);
  and _16373_ (_08106_, _08105_, _06680_);
  nor _16374_ (_08107_, _06881_, _06697_);
  or _16375_ (_08108_, _06885_, _06465_);
  nor _16376_ (_08109_, _08108_, _08107_);
  nor _16377_ (_08110_, _08109_, _06886_);
  and _16378_ (_08111_, _08110_, _06511_);
  nor _16379_ (_08112_, _08110_, _06511_);
  or _16380_ (_08113_, _08112_, _08111_);
  and _16381_ (_08114_, _08113_, _06883_);
  and _16382_ (_08115_, _06640_, _06958_);
  nor _16383_ (_08116_, _06638_, _06532_);
  nor _16384_ (_08117_, _06732_, _07933_);
  or _16385_ (_08119_, _08117_, _08116_);
  nor _16386_ (_08120_, _08119_, _08115_);
  nand _16387_ (_08121_, _08120_, _06664_);
  nor _16388_ (_08122_, _08121_, _08114_);
  nand _16389_ (_08123_, _08122_, _06625_);
  or _16390_ (_08124_, _08123_, _08106_);
  or _16391_ (_08125_, _08124_, _08103_);
  or _16392_ (_08126_, _08125_, _08098_);
  or _16393_ (_08127_, _08126_, _08079_);
  and _16394_ (_08128_, _08127_, _07653_);
  nand _16395_ (_08129_, _06987_, _06930_);
  or _16396_ (_08130_, _06987_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and _16397_ (_08131_, _08130_, _08027_);
  and _16398_ (_08132_, _08131_, _08129_);
  and _16399_ (_08133_, _08036_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or _16400_ (_08134_, _08133_, _07439_);
  or _16401_ (_08135_, _08134_, _08132_);
  or _16402_ (_08136_, _08135_, _08128_);
  nor _16403_ (_08137_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  not _16404_ (_08138_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _16405_ (_08139_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _08138_);
  nor _16406_ (_08141_, _08139_, _08137_);
  nor _16407_ (_08142_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  not _16408_ (_08143_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and _16409_ (_08144_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _08143_);
  nor _16410_ (_08145_, _08144_, _08142_);
  and _16411_ (_08146_, _08145_, _07599_);
  and _16412_ (_08147_, _08146_, _08141_);
  nor _16413_ (_08148_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  not _16414_ (_08150_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _16415_ (_08151_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _08150_);
  nor _16416_ (_08152_, _08151_, _08148_);
  and _16417_ (_08153_, _08152_, _08147_);
  nor _16418_ (_08154_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  not _16419_ (_08155_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and _16420_ (_08156_, _08155_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _16421_ (_08157_, _08156_, _08154_);
  or _16422_ (_08158_, _08157_, _08153_);
  and _16423_ (_08159_, _08157_, _08153_);
  nor _16424_ (_08160_, _08159_, _06848_);
  and _16425_ (_08161_, _08160_, _08158_);
  or _16426_ (_08162_, _07907_, _07886_);
  and _16427_ (_08163_, _08162_, _07908_);
  and _16428_ (_08164_, _08163_, _07602_);
  nor _16429_ (_08165_, _06806_, _06795_);
  and _16430_ (_08166_, _06785_, _06775_);
  and _16431_ (_08167_, _08166_, _08165_);
  and _16432_ (_08168_, _08167_, _07442_);
  and _16433_ (_08169_, _08168_, _06752_);
  nor _16434_ (_08170_, _08169_, _06515_);
  and _16435_ (_08171_, _07446_, _06795_);
  and _16436_ (_08172_, _08171_, _06812_);
  nand _16437_ (_08173_, _08172_, _06833_);
  nor _16438_ (_08174_, _08173_, _06752_);
  nor _16439_ (_08175_, _08174_, _06465_);
  nor _16440_ (_08176_, _08175_, _08170_);
  or _16441_ (_08177_, _08176_, _06483_);
  nand _16442_ (_08178_, _08176_, _06483_);
  and _16443_ (_08179_, _08178_, _06620_);
  and _16444_ (_08180_, _08179_, _08177_);
  and _16445_ (_08181_, _06913_, _07603_);
  nor _16446_ (_08182_, _06465_, _06951_);
  nor _16447_ (_08183_, _08182_, _06640_);
  nor _16448_ (_08184_, _08183_, _06482_);
  and _16449_ (_08185_, _07459_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  nand _16450_ (_08186_, _06465_, _06455_);
  nor _16451_ (_08187_, _08186_, _06511_);
  or _16452_ (_08188_, _08187_, _08185_);
  or _16453_ (_08190_, _08188_, _08184_);
  or _16454_ (_08191_, _08190_, _08181_);
  or _16455_ (_08192_, _08191_, _08180_);
  or _16456_ (_08193_, _08192_, _08164_);
  or _16457_ (_08194_, _08193_, _08161_);
  or _16458_ (_08195_, _08194_, _07961_);
  and _16459_ (_08196_, _08195_, _08136_);
  and _16460_ (_06517_, _08196_, _06444_);
  or _16461_ (_08197_, _07750_, _07748_);
  nand _16462_ (_08198_, _08197_, _08071_);
  nand _16463_ (_08199_, _08198_, _07757_);
  or _16464_ (_08200_, _07757_, _07701_);
  and _16465_ (_08201_, _08200_, _08199_);
  and _16466_ (_08202_, _08201_, _07459_);
  or _16467_ (_08203_, _08089_, _08090_);
  and _16468_ (_08205_, _08203_, _08094_);
  and _16469_ (_08206_, _08205_, _07602_);
  nor _16470_ (_08207_, _06838_, _06767_);
  and _16471_ (_08208_, _06838_, _06767_);
  nor _16472_ (_08209_, _08208_, _08207_);
  and _16473_ (_08210_, _08209_, _06680_);
  or _16474_ (_08211_, _06870_, _06767_);
  nor _16475_ (_08212_, _06871_, _06848_);
  and _16476_ (_08213_, _08212_, _08211_);
  nor _16477_ (_08214_, _06884_, _06891_);
  and _16478_ (_08215_, _08214_, _06534_);
  and _16479_ (_08216_, _06885_, _06532_);
  and _16480_ (_08217_, _06640_, _06534_);
  nor _16481_ (_08218_, _07933_, _06511_);
  nor _16482_ (_08220_, _06638_, _06551_);
  or _16483_ (_08221_, _08220_, _08218_);
  or _16484_ (_08222_, _08221_, _08217_);
  or _16485_ (_08223_, _08222_, _08216_);
  nor _16486_ (_08224_, _08223_, _08215_);
  and _16487_ (_08225_, _08224_, _07186_);
  nand _16488_ (_08226_, _08225_, _07177_);
  or _16489_ (_08227_, _08226_, _08213_);
  or _16490_ (_08228_, _08227_, _08210_);
  or _16491_ (_08229_, _08228_, _08206_);
  or _16492_ (_08230_, _08229_, _08202_);
  and _16493_ (_08231_, _08230_, _07653_);
  not _16494_ (_08232_, _06930_);
  and _16495_ (_08233_, _06983_, _08232_);
  nor _16496_ (_08234_, _06983_, _06749_);
  or _16497_ (_08235_, _08234_, _08233_);
  and _16498_ (_08236_, _08235_, _08027_);
  and _16499_ (_08237_, _08036_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or _16500_ (_08238_, _08237_, _07439_);
  or _16501_ (_08239_, _08238_, _08236_);
  or _16502_ (_08241_, _08239_, _08231_);
  or _16503_ (_08242_, _08152_, _08147_);
  nor _16504_ (_08243_, _08153_, _06848_);
  and _16505_ (_08244_, _08243_, _08242_);
  or _16506_ (_08245_, _07905_, _07903_);
  and _16507_ (_08246_, _08245_, _07906_);
  and _16508_ (_08247_, _08246_, _07602_);
  and _16509_ (_08248_, _08173_, _06515_);
  nor _16510_ (_08249_, _08168_, _06515_);
  or _16511_ (_08250_, _08249_, _08248_);
  nand _16512_ (_08251_, _08250_, _06752_);
  or _16513_ (_08252_, _08250_, _06752_);
  and _16514_ (_08253_, _08252_, _06620_);
  and _16515_ (_08254_, _08253_, _08251_);
  and _16516_ (_08255_, _06913_, _06903_);
  nand _16517_ (_08256_, _06532_, _06465_);
  or _16518_ (_08257_, _06753_, _06465_);
  and _16519_ (_08258_, _08257_, _06455_);
  and _16520_ (_08259_, _08258_, _08256_);
  and _16521_ (_08260_, _06753_, _06640_);
  and _16522_ (_08261_, _07459_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  or _16523_ (_08262_, _08261_, _08260_);
  or _16524_ (_08263_, _08262_, _08259_);
  or _16525_ (_08264_, _08263_, _08255_);
  or _16526_ (_08265_, _08264_, _08254_);
  or _16527_ (_08266_, _08265_, _08247_);
  or _16528_ (_08267_, _08266_, _08244_);
  or _16529_ (_08268_, _08267_, _07961_);
  and _16530_ (_08269_, _08268_, _08241_);
  and _16531_ (_06533_, _08269_, _06444_);
  and _16532_ (_08270_, _07758_, _07717_);
  or _16533_ (_08271_, _07745_, _07718_);
  not _16534_ (_08272_, _07741_);
  and _16535_ (_08273_, _07744_, _08272_);
  nand _16536_ (_08274_, _08273_, _08271_);
  or _16537_ (_08275_, _08273_, _08271_);
  and _16538_ (_08276_, _08275_, _08274_);
  and _16539_ (_08277_, _08276_, _07757_);
  or _16540_ (_08278_, _08277_, _08270_);
  and _16541_ (_08279_, _08278_, _07459_);
  nand _16542_ (_08280_, _07925_, _07922_);
  nand _16543_ (_08281_, _08280_, _08082_);
  not _16544_ (_08282_, _08083_);
  and _16545_ (_08283_, _08282_, _08281_);
  nor _16546_ (_08284_, _08283_, _08089_);
  and _16547_ (_08285_, _08284_, _07602_);
  and _16548_ (_08286_, _06831_, _06817_);
  nor _16549_ (_08287_, _08286_, _06832_);
  nor _16550_ (_08288_, _08287_, _06681_);
  nand _16551_ (_08289_, _06866_, _06860_);
  nor _16552_ (_08290_, _06867_, _06848_);
  and _16553_ (_08291_, _08290_, _08289_);
  or _16554_ (_08292_, _08214_, _06640_);
  and _16555_ (_08293_, _08292_, _06552_);
  not _16556_ (_08294_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor _16557_ (_08295_, _06610_, _08294_);
  and _16558_ (_08296_, _08295_, _08214_);
  nor _16559_ (_08297_, _07933_, _06532_);
  nor _16560_ (_08298_, _06638_, _06604_);
  nor _16561_ (_08299_, _08298_, _08297_);
  and _16562_ (_08300_, _08299_, _07295_);
  nand _16563_ (_08301_, _08300_, _07292_);
  or _16564_ (_08302_, _08301_, _08296_);
  nor _16565_ (_08303_, _08302_, _08293_);
  nand _16566_ (_08304_, _08303_, _07289_);
  or _16567_ (_08305_, _08304_, _08291_);
  or _16568_ (_08306_, _08305_, _08288_);
  or _16569_ (_08307_, _08306_, _08285_);
  or _16570_ (_08308_, _08307_, _08279_);
  and _16571_ (_08309_, _08308_, _07653_);
  and _16572_ (_08310_, _06932_, _06430_);
  nand _16573_ (_08311_, _08310_, _06930_);
  or _16574_ (_08312_, _08310_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and _16575_ (_08313_, _08312_, _08027_);
  and _16576_ (_08314_, _08313_, _08311_);
  and _16577_ (_08315_, _08036_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or _16578_ (_08316_, _08315_, _07439_);
  or _16579_ (_08317_, _08316_, _08314_);
  or _16580_ (_08318_, _08317_, _08309_);
  or _16581_ (_08319_, _08146_, _08141_);
  nor _16582_ (_08320_, _08147_, _06848_);
  and _16583_ (_08321_, _08320_, _08319_);
  and _16584_ (_08322_, _08165_, _07442_);
  and _16585_ (_08323_, _08322_, _06785_);
  nor _16586_ (_08324_, _08323_, _06515_);
  nor _16587_ (_08325_, _08172_, _06465_);
  nor _16588_ (_08326_, _08325_, _08324_);
  nand _16589_ (_08327_, _08326_, _06833_);
  or _16590_ (_08328_, _08326_, _06833_);
  and _16591_ (_08329_, _08328_, _06620_);
  and _16592_ (_08330_, _08329_, _08327_);
  or _16593_ (_08331_, _07901_, _07899_);
  and _16594_ (_08332_, _08331_, _07902_);
  and _16595_ (_08333_, _08332_, _07602_);
  nor _16596_ (_08334_, _06551_, _06951_);
  and _16597_ (_08335_, _06833_, _06640_);
  and _16598_ (_08336_, _07459_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  or _16599_ (_08337_, _08336_, _08335_);
  or _16600_ (_08338_, _08337_, _06915_);
  or _16601_ (_08339_, _08338_, _08334_);
  or _16602_ (_08340_, _08339_, _08333_);
  or _16603_ (_08341_, _08340_, _08330_);
  or _16604_ (_08342_, _08341_, _08321_);
  or _16605_ (_08343_, _08342_, _07961_);
  and _16606_ (_08344_, _08343_, _08318_);
  and _16607_ (_06536_, _08344_, _06444_);
  nand _16608_ (_08345_, _07251_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  nand _16609_ (_08346_, _07238_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  and _16610_ (_08347_, _08346_, _08345_);
  nand _16611_ (_08348_, _07246_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nand _16612_ (_08349_, _07248_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and _16613_ (_08350_, _08349_, _08348_);
  nand _16614_ (_08351_, _07254_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nand _16615_ (_08352_, _07242_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  and _16616_ (_08353_, _08352_, _08351_);
  and _16617_ (_08354_, _08353_, _08350_);
  nand _16618_ (_08355_, _08354_, _08347_);
  nand _16619_ (_08356_, _08355_, _07234_);
  nand _16620_ (_08357_, _08356_, _07233_);
  nor _16621_ (_08358_, \oc8051_top_1.oc8051_memory_interface1.cdata [7], _07233_);
  not _16622_ (_08359_, _08358_);
  and _16623_ (_08360_, _08359_, _08357_);
  and _16624_ (_06566_, _08360_, _06444_);
  nor _16625_ (_08361_, _07230_, _06699_);
  and _16626_ (_08362_, _07254_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and _16627_ (_08363_, _07238_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor _16628_ (_08364_, _08363_, _08362_);
  and _16629_ (_08365_, _07246_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and _16630_ (_08366_, _07242_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor _16631_ (_08367_, _08366_, _08365_);
  and _16632_ (_08368_, _07251_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  and _16633_ (_08369_, _07248_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nor _16634_ (_08370_, _08369_, _08368_);
  and _16635_ (_08371_, _08370_, _08367_);
  and _16636_ (_08372_, _08371_, _08364_);
  and _16637_ (_08373_, _07230_, _07234_);
  not _16638_ (_08374_, _08373_);
  nor _16639_ (_08375_, _08374_, _08372_);
  nor _16640_ (_08376_, _08375_, _08361_);
  nor _16641_ (_06569_, _08376_, rst);
  and _16642_ (_06713_, _07263_, _06444_);
  nand _16643_ (_08377_, _07248_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nand _16644_ (_08378_, _07254_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  and _16645_ (_08379_, _08378_, _08377_);
  nand _16646_ (_08380_, _07238_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  and _16647_ (_08381_, _08380_, _08379_);
  nand _16648_ (_08382_, _07242_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  and _16649_ (_08383_, _08382_, _07234_);
  nand _16650_ (_08384_, _07246_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nand _16651_ (_08385_, _07251_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  and _16652_ (_08386_, _08385_, _08384_);
  and _16653_ (_08387_, _08386_, _08383_);
  nand _16654_ (_08388_, _08387_, _08381_);
  or _16655_ (_08389_, _08388_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor _16656_ (_08390_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], _07233_);
  not _16657_ (_08391_, _08390_);
  and _16658_ (_08392_, _08391_, _08389_);
  and _16659_ (_06715_, _08392_, _06444_);
  and _16660_ (_08393_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], \oc8051_top_1.oc8051_memory_interface1.cdone );
  not _16661_ (_08394_, _08393_);
  nand _16662_ (_08395_, _07248_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nand _16663_ (_08396_, _07242_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  and _16664_ (_08397_, _08396_, _08395_);
  nand _16665_ (_08398_, _07254_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nand _16666_ (_08399_, _07238_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  and _16667_ (_08400_, _08399_, _08398_);
  and _16668_ (_08401_, _08400_, _08397_);
  nand _16669_ (_08402_, _07246_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nand _16670_ (_08403_, _07251_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  and _16671_ (_08404_, _08403_, _08402_);
  and _16672_ (_08405_, _08404_, _08401_);
  or _16673_ (_08406_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  or _16674_ (_08407_, _08406_, _08405_);
  and _16675_ (_08408_, _08407_, _08394_);
  nor _16676_ (_06717_, _08408_, rst);
  nand _16677_ (_08410_, _07251_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  nand _16678_ (_08411_, _07238_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  and _16679_ (_08412_, _08411_, _08410_);
  nand _16680_ (_08413_, _07246_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nand _16681_ (_08414_, _07248_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and _16682_ (_08415_, _08414_, _08413_);
  nand _16683_ (_08416_, _07254_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nand _16684_ (_08417_, _07242_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  and _16685_ (_08418_, _08417_, _08416_);
  and _16686_ (_08419_, _08418_, _08415_);
  nand _16687_ (_08420_, _08419_, _08412_);
  nand _16688_ (_08421_, _08420_, _07234_);
  nand _16689_ (_08422_, _08421_, _07233_);
  nor _16690_ (_08423_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], _07233_);
  not _16691_ (_08424_, _08423_);
  and _16692_ (_08425_, _08424_, _08422_);
  and _16693_ (_06719_, _08425_, _06444_);
  and _16694_ (_08426_, _07246_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and _16695_ (_08427_, _07251_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  and _16696_ (_08428_, _07248_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and _16697_ (_08429_, _07254_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor _16698_ (_08430_, _08429_, _08428_);
  and _16699_ (_08431_, _07238_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  and _16700_ (_08432_, _07242_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  nor _16701_ (_08433_, _08432_, _08431_);
  nand _16702_ (_08434_, _08433_, _08430_);
  or _16703_ (_08435_, _08434_, _08427_);
  or _16704_ (_08436_, _08435_, _08426_);
  or _16705_ (_08437_, _08436_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  or _16706_ (_08438_, _08437_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor _16707_ (_08439_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], _07233_);
  not _16708_ (_08440_, _08439_);
  and _16709_ (_08441_, _08440_, _08438_);
  and _16710_ (_06721_, _08441_, _06444_);
  nand _16711_ (_08442_, _07251_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  nand _16712_ (_08443_, _07238_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  and _16713_ (_08444_, _08443_, _08442_);
  nand _16714_ (_08445_, _07246_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  nand _16715_ (_08446_, _07248_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and _16716_ (_08447_, _08446_, _08445_);
  nand _16717_ (_08448_, _07254_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nand _16718_ (_08449_, _07242_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  and _16719_ (_08450_, _08449_, _08448_);
  and _16720_ (_08451_, _08450_, _08447_);
  nand _16721_ (_08452_, _08451_, _08444_);
  and _16722_ (_08453_, _08452_, _07234_);
  or _16723_ (_08454_, _08453_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor _16724_ (_08455_, _07233_, \oc8051_top_1.oc8051_memory_interface1.cdata [5]);
  not _16725_ (_08456_, _08455_);
  and _16726_ (_08457_, _08456_, _08454_);
  and _16727_ (_06724_, _08457_, _06444_);
  nand _16728_ (_08458_, _07242_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nand _16729_ (_08459_, _07238_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  and _16730_ (_08460_, _08459_, _08458_);
  nand _16731_ (_08461_, _07246_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nand _16732_ (_08462_, _07248_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and _16733_ (_08463_, _08462_, _08461_);
  nand _16734_ (_08464_, _07251_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  nand _16735_ (_08465_, _07254_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  and _16736_ (_08466_, _08465_, _08464_);
  and _16737_ (_08467_, _08466_, _08463_);
  and _16738_ (_08468_, _08467_, _08460_);
  or _16739_ (_08469_, _08468_, _08406_);
  and _16740_ (_08470_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], \oc8051_top_1.oc8051_memory_interface1.cdone );
  not _16741_ (_08471_, _08470_);
  and _16742_ (_08472_, _08471_, _08469_);
  nor _16743_ (_06726_, _08472_, rst);
  and _16744_ (_08473_, _06299_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  and _16745_ (_08474_, _08473_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  nor _16746_ (_08475_, _08473_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  nor _16747_ (_08476_, _08475_, _08474_);
  and _16748_ (_06950_, _08476_, _06443_);
  nor _16749_ (_08477_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  not _16750_ (_08478_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor _16751_ (_08479_, _08478_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  nor _16752_ (_08480_, _08479_, _08477_);
  not _16753_ (_08481_, \oc8051_symbolic_cxrom1.regvalid [13]);
  not _16754_ (_08482_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor _16755_ (_08483_, _07432_, _08482_);
  and _16756_ (_08484_, _08483_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor _16757_ (_08485_, _08483_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor _16758_ (_08486_, _08485_, _08484_);
  nor _16759_ (_08487_, _08486_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor _16760_ (_08488_, _08478_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3]);
  nor _16761_ (_08489_, _08488_, _08487_);
  and _16762_ (_08490_, _08489_, _08481_);
  nor _16763_ (_08491_, _08489_, \oc8051_symbolic_cxrom1.regvalid [5]);
  or _16764_ (_08492_, _08491_, _08490_);
  not _16765_ (_08493_, _08492_);
  nor _16766_ (_08494_, \oc8051_top_1.oc8051_memory_interface1.istb_t , \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  nor _16767_ (_08495_, _08478_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1]);
  nor _16768_ (_08496_, _08495_, _08494_);
  not _16769_ (_08497_, _08496_);
  and _16770_ (_08498_, _07432_, _08482_);
  nor _16771_ (_08499_, _08498_, _08483_);
  nor _16772_ (_08500_, _08499_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor _16773_ (_08501_, _08478_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2]);
  nor _16774_ (_08502_, _08501_, _08500_);
  and _16775_ (_08503_, _08502_, _08497_);
  nand _16776_ (_08504_, _08503_, _08493_);
  and _16777_ (_08505_, _08504_, _08480_);
  nor _16778_ (_08506_, _08502_, _08497_);
  not _16779_ (_08507_, _08506_);
  not _16780_ (_08508_, \oc8051_symbolic_cxrom1.regvalid [3]);
  nor _16781_ (_08509_, _08489_, _08508_);
  and _16782_ (_08510_, _08489_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor _16783_ (_08511_, _08510_, _08509_);
  nor _16784_ (_08512_, _08511_, _08507_);
  and _16785_ (_08513_, _08502_, _08496_);
  not _16786_ (_08514_, _08513_);
  not _16787_ (_08515_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and _16788_ (_08516_, _08489_, _08515_);
  nor _16789_ (_08517_, _08489_, \oc8051_symbolic_cxrom1.regvalid [7]);
  or _16790_ (_08518_, _08517_, _08516_);
  nor _16791_ (_08519_, _08518_, _08514_);
  nor _16792_ (_08520_, _08519_, _08512_);
  not _16793_ (_08521_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and _16794_ (_08522_, _08489_, _08521_);
  nor _16795_ (_08523_, _08502_, _08496_);
  not _16796_ (_08524_, _08523_);
  nor _16797_ (_08525_, _08489_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or _16798_ (_08526_, _08525_, _08524_);
  or _16799_ (_08527_, _08526_, _08522_);
  and _16800_ (_08528_, _08527_, _08520_);
  and _16801_ (_08529_, _08528_, _08505_);
  not _16802_ (_08530_, _08502_);
  and _16803_ (_08531_, _08489_, \oc8051_symbolic_cxrom1.regvalid [12]);
  not _16804_ (_08532_, _08489_);
  and _16805_ (_08533_, _08532_, \oc8051_symbolic_cxrom1.regvalid [4]);
  nor _16806_ (_08534_, _08533_, _08531_);
  nor _16807_ (_08535_, _08534_, _08530_);
  nor _16808_ (_08536_, _08502_, _08489_);
  and _16809_ (_08537_, _08536_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and _16810_ (_08538_, _08530_, _08489_);
  and _16811_ (_08539_, _08538_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor _16812_ (_08540_, _08539_, _08537_);
  not _16813_ (_08541_, _08540_);
  nor _16814_ (_08542_, _08541_, _08535_);
  nor _16815_ (_08543_, _08542_, _08496_);
  and _16816_ (_08544_, _08536_, _08496_);
  and _16817_ (_08545_, _08544_, \oc8051_symbolic_cxrom1.regvalid [2]);
  not _16818_ (_08546_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and _16819_ (_08547_, _08489_, _08546_);
  nor _16820_ (_08548_, _08489_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or _16821_ (_08549_, _08548_, _08547_);
  nor _16822_ (_08550_, _08549_, _08514_);
  and _16823_ (_08551_, _08489_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and _16824_ (_08552_, _08551_, _08506_);
  or _16825_ (_08553_, _08552_, _08480_);
  or _16826_ (_08554_, _08553_, _08550_);
  or _16827_ (_08555_, _08554_, _08545_);
  nor _16828_ (_08556_, _08555_, _08543_);
  nor _16829_ (_08557_, _08556_, _08529_);
  not _16830_ (_08558_, _08557_);
  and _16831_ (_08559_, _08558_, word_in[7]);
  not _16832_ (_08560_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  nand _16833_ (_08561_, _08480_, _08560_);
  or _16834_ (_08562_, _08480_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  and _16835_ (_08563_, _08562_, _08561_);
  and _16836_ (_08564_, _08563_, _08513_);
  not _16837_ (_08565_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  nand _16838_ (_08566_, _08480_, _08565_);
  or _16839_ (_08567_, _08480_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  and _16840_ (_08568_, _08567_, _08566_);
  and _16841_ (_08569_, _08568_, _08506_);
  or _16842_ (_08570_, _08569_, _08564_);
  not _16843_ (_08571_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  nand _16844_ (_08572_, _08480_, _08571_);
  or _16845_ (_08573_, _08480_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  and _16846_ (_08574_, _08573_, _08572_);
  and _16847_ (_08575_, _08574_, _08503_);
  not _16848_ (_08576_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  nand _16849_ (_08577_, _08480_, _08576_);
  or _16850_ (_08578_, _08480_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  and _16851_ (_08579_, _08578_, _08577_);
  and _16852_ (_08580_, _08579_, _08523_);
  or _16853_ (_08581_, _08580_, _08575_);
  or _16854_ (_08582_, _08581_, _08570_);
  and _16855_ (_08583_, _08582_, _08489_);
  not _16856_ (_08584_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  nand _16857_ (_08585_, _08480_, _08584_);
  or _16858_ (_08586_, _08480_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  and _16859_ (_08587_, _08586_, _08585_);
  and _16860_ (_08588_, _08587_, _08544_);
  and _16861_ (_08589_, _08513_, _08532_);
  not _16862_ (_08590_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  nand _16863_ (_08591_, _08480_, _08590_);
  or _16864_ (_08592_, _08480_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  and _16865_ (_08593_, _08592_, _08591_);
  and _16866_ (_08594_, _08593_, _08589_);
  not _16867_ (_08595_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  nand _16868_ (_08596_, _08480_, _08595_);
  or _16869_ (_08597_, _08480_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  and _16870_ (_08598_, _08597_, _08596_);
  and _16871_ (_08599_, _08598_, _08503_);
  not _16872_ (_08600_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  nand _16873_ (_08601_, _08480_, _08600_);
  or _16874_ (_08602_, _08480_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  and _16875_ (_08603_, _08602_, _08601_);
  and _16876_ (_08604_, _08603_, _08523_);
  or _16877_ (_08605_, _08604_, _08599_);
  and _16878_ (_08606_, _08605_, _08532_);
  or _16879_ (_08607_, _08606_, _08594_);
  or _16880_ (_08608_, _08607_, _08588_);
  or _16881_ (_08609_, _08608_, _08583_);
  and _16882_ (_08610_, _08609_, _08557_);
  or _16883_ (\oc8051_symbolic_cxrom1.cxrom_data_out [7], _08610_, _08559_);
  nor _16884_ (_08611_, _08496_, _08480_);
  not _16885_ (_08612_, _08611_);
  and _16886_ (_08613_, _08496_, _08480_);
  nor _16887_ (_08614_, _08613_, _08502_);
  and _16888_ (_08615_, _08613_, _08502_);
  nor _16889_ (_08616_, _08615_, _08614_);
  not _16890_ (_08617_, _08616_);
  nor _16891_ (_08618_, _08617_, _08492_);
  nor _16892_ (_08619_, _08615_, _08532_);
  and _16893_ (_08620_, _08615_, _08532_);
  nor _16894_ (_08622_, _08620_, _08619_);
  nor _16895_ (_08623_, _08622_, _08616_);
  and _16896_ (_08624_, _08623_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and _16897_ (_08626_, _08622_, _08617_);
  and _16898_ (_08627_, _08626_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or _16899_ (_08628_, _08627_, _08624_);
  nor _16900_ (_08630_, _08628_, _08618_);
  nor _16901_ (_08631_, _08630_, _08612_);
  not _16902_ (_08632_, _08631_);
  not _16903_ (_08634_, _08613_);
  nor _16904_ (_08635_, _08617_, _08534_);
  and _16905_ (_08636_, _08626_, \oc8051_symbolic_cxrom1.regvalid [0]);
  nor _16906_ (_08638_, _08636_, _08635_);
  or _16907_ (_08639_, _08638_, _08634_);
  nand _16908_ (_08640_, _08620_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and _16909_ (_08642_, _08640_, _08639_);
  and _16910_ (_08643_, _08642_, _08632_);
  and _16911_ (_08644_, _08497_, _08480_);
  not _16912_ (_08645_, _08644_);
  nor _16913_ (_08646_, _08617_, _08549_);
  and _16914_ (_08648_, _08623_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and _16915_ (_08649_, _08626_, \oc8051_symbolic_cxrom1.regvalid [2]);
  or _16916_ (_08651_, _08649_, _08648_);
  nor _16917_ (_08652_, _08651_, _08646_);
  nor _16918_ (_08653_, _08652_, _08645_);
  not _16919_ (_08654_, _08480_);
  and _16920_ (_08655_, _08496_, _08654_);
  not _16921_ (_08656_, _08655_);
  nor _16922_ (_08657_, _08617_, _08518_);
  and _16923_ (_08658_, _08623_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and _16924_ (_08659_, _08626_, \oc8051_symbolic_cxrom1.regvalid [3]);
  or _16925_ (_08660_, _08659_, _08658_);
  nor _16926_ (_08661_, _08660_, _08657_);
  nor _16927_ (_08662_, _08661_, _08656_);
  nor _16928_ (_08663_, _08662_, _08653_);
  and _16929_ (_08664_, _08663_, _08643_);
  or _16930_ (_08665_, _08613_, _08611_);
  not _16931_ (_08666_, _08665_);
  not _16932_ (_08667_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  nand _16933_ (_08668_, _08480_, _08667_);
  or _16934_ (_08669_, _08480_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  and _16935_ (_08670_, _08669_, _08668_);
  and _16936_ (_08671_, _08670_, _08666_);
  not _16937_ (_08672_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  nand _16938_ (_08673_, _08480_, _08672_);
  or _16939_ (_08674_, _08480_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  and _16940_ (_08675_, _08674_, _08673_);
  and _16941_ (_08676_, _08675_, _08665_);
  or _16942_ (_08677_, _08676_, _08671_);
  and _16943_ (_08678_, _08677_, _08623_);
  and _16944_ (_08679_, _08616_, _08489_);
  not _16945_ (_08680_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  nand _16946_ (_08681_, _08480_, _08680_);
  or _16947_ (_08682_, _08480_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  and _16948_ (_08683_, _08682_, _08681_);
  and _16949_ (_08684_, _08683_, _08666_);
  not _16950_ (_08685_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  nand _16951_ (_08686_, _08480_, _08685_);
  or _16952_ (_08687_, _08480_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  and _16953_ (_08688_, _08687_, _08686_);
  and _16954_ (_08689_, _08688_, _08665_);
  or _16955_ (_08691_, _08689_, _08684_);
  and _16956_ (_08692_, _08691_, _08679_);
  or _16957_ (_08693_, _08692_, _08678_);
  not _16958_ (_08695_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  nand _16959_ (_08696_, _08480_, _08695_);
  or _16960_ (_08697_, _08480_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  and _16961_ (_08698_, _08697_, _08696_);
  and _16962_ (_08699_, _08698_, _08665_);
  not _16963_ (_08700_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  nand _16964_ (_08702_, _08480_, _08700_);
  or _16965_ (_08703_, _08480_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  and _16966_ (_08704_, _08703_, _08702_);
  and _16967_ (_08705_, _08704_, _08666_);
  or _16968_ (_08706_, _08705_, _08699_);
  and _16969_ (_08707_, _08706_, _08626_);
  and _16970_ (_08708_, _08616_, _08532_);
  not _16971_ (_08709_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  nand _16972_ (_08710_, _08480_, _08709_);
  or _16973_ (_08711_, _08480_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  and _16974_ (_08712_, _08711_, _08710_);
  and _16975_ (_08713_, _08712_, _08665_);
  not _16976_ (_08714_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  nand _16977_ (_08715_, _08480_, _08714_);
  or _16978_ (_08716_, _08480_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  and _16979_ (_08717_, _08716_, _08715_);
  and _16980_ (_08718_, _08717_, _08666_);
  or _16981_ (_08720_, _08718_, _08713_);
  and _16982_ (_08721_, _08720_, _08708_);
  or _16983_ (_08722_, _08721_, _08707_);
  nor _16984_ (_08723_, _08722_, _08693_);
  nor _16985_ (_08724_, _08723_, _08664_);
  and _16986_ (_08725_, _08664_, word_in[15]);
  or _16987_ (\oc8051_symbolic_cxrom1.cxrom_data_out [15], _08725_, _08724_);
  nor _16988_ (_08726_, _08513_, _08523_);
  not _16989_ (_08727_, _08726_);
  nor _16990_ (_08728_, _08727_, _08492_);
  and _16991_ (_08729_, _08513_, _08489_);
  nor _16992_ (_08730_, _08513_, _08489_);
  nor _16993_ (_08731_, _08730_, _08729_);
  nor _16994_ (_08732_, _08726_, _08731_);
  and _16995_ (_08733_, _08732_, \oc8051_symbolic_cxrom1.regvalid [1]);
  and _16996_ (_08734_, _08727_, _08731_);
  and _16997_ (_08735_, _08734_, \oc8051_symbolic_cxrom1.regvalid [9]);
  or _16998_ (_08736_, _08735_, _08733_);
  nor _16999_ (_08737_, _08736_, _08728_);
  nor _17000_ (_08738_, _08737_, _08634_);
  and _17001_ (_08739_, _08732_, \oc8051_symbolic_cxrom1.regvalid [3]);
  not _17002_ (_08740_, _08739_);
  nor _17003_ (_08742_, _08727_, _08518_);
  and _17004_ (_08744_, _08734_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor _17005_ (_08746_, _08744_, _08742_);
  and _17006_ (_08747_, _08746_, _08740_);
  nor _17007_ (_08748_, _08747_, _08645_);
  nor _17008_ (_08749_, _08748_, _08738_);
  nor _17009_ (_08751_, _08727_, _08549_);
  and _17010_ (_08752_, _08734_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and _17011_ (_08753_, _08732_, \oc8051_symbolic_cxrom1.regvalid [2]);
  or _17012_ (_08754_, _08753_, _08752_);
  nor _17013_ (_08756_, _08754_, _08751_);
  nor _17014_ (_08758_, _08756_, _08612_);
  and _17015_ (_08759_, _08732_, \oc8051_symbolic_cxrom1.regvalid [0]);
  not _17016_ (_08760_, _08759_);
  nor _17017_ (_08761_, _08727_, _08534_);
  and _17018_ (_08763_, _08734_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor _17019_ (_08764_, _08763_, _08761_);
  and _17020_ (_08765_, _08764_, _08760_);
  nor _17021_ (_08766_, _08765_, _08656_);
  nor _17022_ (_08768_, _08766_, _08758_);
  and _17023_ (_08769_, _08768_, _08749_);
  not _17024_ (_08770_, _08731_);
  and _17025_ (_08771_, _08593_, _08503_);
  and _17026_ (_08772_, _08603_, _08489_);
  or _17027_ (_08773_, _08772_, _08771_);
  and _17028_ (_08774_, _08598_, _08506_);
  and _17029_ (_08775_, _08587_, _08523_);
  or _17030_ (_08776_, _08775_, _08774_);
  or _17031_ (_08777_, _08776_, _08773_);
  and _17032_ (_08778_, _08777_, _08770_);
  and _17033_ (_08779_, _08574_, _08506_);
  and _17034_ (_08780_, _08568_, _08523_);
  or _17035_ (_08781_, _08780_, _08779_);
  and _17036_ (_08782_, _08563_, _08503_);
  and _17037_ (_08783_, _08579_, _08513_);
  or _17038_ (_08784_, _08783_, _08782_);
  or _17039_ (_08785_, _08784_, _08781_);
  and _17040_ (_08786_, _08785_, _08731_);
  nor _17041_ (_08787_, _08786_, _08778_);
  nor _17042_ (_08788_, _08787_, _08769_);
  and _17043_ (_08789_, _08769_, word_in[23]);
  or _17044_ (\oc8051_symbolic_cxrom1.cxrom_data_out [23], _08789_, _08788_);
  and _17045_ (_08790_, _08729_, _08654_);
  and _17046_ (_08791_, _08790_, \oc8051_symbolic_cxrom1.regvalid [1]);
  and _17047_ (_08792_, _08612_, _08502_);
  nor _17048_ (_08793_, _08612_, _08502_);
  nor _17049_ (_08794_, _08793_, _08792_);
  not _17050_ (_08795_, _08794_);
  nor _17051_ (_08796_, _08795_, _08518_);
  and _17052_ (_08797_, _08792_, _08489_);
  nor _17053_ (_08798_, _08792_, _08489_);
  nor _17054_ (_08799_, _08798_, _08797_);
  and _17055_ (_08800_, _08799_, _08795_);
  and _17056_ (_08801_, _08800_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor _17057_ (_08802_, _08801_, _08796_);
  nor _17058_ (_08803_, _08802_, _08612_);
  nor _17059_ (_08804_, _08803_, _08791_);
  nor _17060_ (_08805_, _08795_, _08492_);
  and _17061_ (_08806_, _08800_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor _17062_ (_08807_, _08806_, _08805_);
  nor _17063_ (_08808_, _08807_, _08656_);
  and _17064_ (_08809_, _08793_, _08509_);
  nor _17065_ (_08810_, _08809_, _08808_);
  and _17066_ (_08811_, _08810_, _08804_);
  nor _17067_ (_08812_, _08549_, _08795_);
  and _17068_ (_08813_, _08800_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor _17069_ (_08814_, _08799_, _08794_);
  and _17070_ (_08815_, _08814_, \oc8051_symbolic_cxrom1.regvalid [2]);
  or _17071_ (_08816_, _08815_, _08813_);
  nor _17072_ (_08817_, _08816_, _08812_);
  nor _17073_ (_08818_, _08817_, _08634_);
  and _17074_ (_08819_, _08502_, _08489_);
  and _17075_ (_08820_, _08644_, _08819_);
  and _17076_ (_08821_, _08820_, \oc8051_symbolic_cxrom1.regvalid [0]);
  nor _17077_ (_08822_, _08795_, _08534_);
  and _17078_ (_08823_, _08800_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor _17079_ (_08824_, _08823_, _08822_);
  nor _17080_ (_08825_, _08824_, _08645_);
  or _17081_ (_08826_, _08825_, _08821_);
  nor _17082_ (_08827_, _08826_, _08818_);
  and _17083_ (_08828_, _08827_, _08811_);
  and _17084_ (_08829_, _08675_, _08666_);
  and _17085_ (_08830_, _08670_, _08665_);
  or _17086_ (_08831_, _08830_, _08829_);
  and _17087_ (_08832_, _08831_, _08800_);
  and _17088_ (_08833_, _08698_, _08666_);
  and _17089_ (_08834_, _08704_, _08665_);
  or _17090_ (_08835_, _08834_, _08833_);
  and _17091_ (_08836_, _08835_, _08814_);
  and _17092_ (_08837_, _08794_, _08532_);
  and _17093_ (_08838_, _08712_, _08666_);
  and _17094_ (_08839_, _08717_, _08665_);
  or _17095_ (_08840_, _08839_, _08838_);
  and _17096_ (_08841_, _08840_, _08837_);
  and _17097_ (_08842_, _08794_, _08489_);
  and _17098_ (_08843_, _08688_, _08666_);
  and _17099_ (_08844_, _08683_, _08665_);
  or _17100_ (_08845_, _08844_, _08843_);
  and _17101_ (_08846_, _08845_, _08842_);
  or _17102_ (_08847_, _08846_, _08841_);
  or _17103_ (_08848_, _08847_, _08836_);
  nor _17104_ (_08849_, _08848_, _08832_);
  nor _17105_ (_08850_, _08849_, _08828_);
  and _17106_ (_08852_, _08828_, word_in[31]);
  or _17107_ (\oc8051_symbolic_cxrom1.cxrom_data_out [31], _08852_, _08850_);
  or _17108_ (_08853_, _08819_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and _17109_ (_07051_, _08853_, _06444_);
  and _17110_ (_08855_, _08828_, _06444_);
  and _17111_ (_08856_, _08855_, word_in[31]);
  and _17112_ (_08857_, _08819_, _08611_);
  and _17113_ (_08859_, _08855_, _08857_);
  and _17114_ (_08860_, _08859_, _08856_);
  not _17115_ (_08862_, _08859_);
  and _17116_ (_08863_, _08769_, _06444_);
  and _17117_ (_08865_, _08863_, _08726_);
  and _17118_ (_08866_, _08865_, _08731_);
  and _17119_ (_08867_, _08866_, _08644_);
  not _17120_ (_08868_, _08867_);
  and _17121_ (_08869_, _08664_, _06444_);
  and _17122_ (_08870_, _08869_, _08655_);
  and _17123_ (_08871_, _08870_, _08679_);
  and _17124_ (_08872_, _08529_, _06444_);
  and _17125_ (_08874_, _08872_, _08496_);
  nor _17126_ (_08875_, _08557_, rst);
  and _17127_ (_08877_, _08875_, _08819_);
  and _17128_ (_08878_, _08877_, _08874_);
  and _17129_ (_08879_, _08878_, word_in[7]);
  nor _17130_ (_08880_, _08878_, _08560_);
  nor _17131_ (_08881_, _08880_, _08879_);
  nor _17132_ (_08882_, _08881_, _08871_);
  and _17133_ (_08883_, _08871_, word_in[15]);
  or _17134_ (_08884_, _08883_, _08882_);
  and _17135_ (_08885_, _08884_, _08868_);
  and _17136_ (_08886_, _08863_, word_in[23]);
  and _17137_ (_08887_, _08886_, _08867_);
  or _17138_ (_08888_, _08887_, _08885_);
  and _17139_ (_08889_, _08888_, _08862_);
  or _17140_ (_14579_, _08889_, _08860_);
  or _17141_ (_08890_, _08814_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and _17142_ (_07097_, _08890_, _06444_);
  and _17143_ (_08891_, _08523_, _08532_);
  or _17144_ (_08892_, _08891_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or _17145_ (_08893_, _08892_, _08729_);
  and _17146_ (_07129_, _08893_, _06444_);
  and _17147_ (_08894_, _08615_, _08489_);
  or _17148_ (_08895_, _08894_, _08891_);
  or _17149_ (_08896_, _08645_, _08502_);
  nor _17150_ (_08897_, _08896_, _08489_);
  and _17151_ (_08898_, _08837_, _08655_);
  nor _17152_ (_08899_, _08898_, \oc8051_symbolic_cxrom1.regvalid [2]);
  nor _17153_ (_08900_, _08899_, _08897_);
  or _17154_ (_08901_, _08900_, _08895_);
  and _17155_ (_07165_, _08901_, _06444_);
  or _17156_ (_08902_, _08536_, \oc8051_symbolic_cxrom1.regvalid [3]);
  and _17157_ (_07212_, _08902_, _06444_);
  not _17158_ (_08903_, _08536_);
  nor _17159_ (_08904_, _08530_, _08489_);
  and _17160_ (_08905_, _08904_, _08611_);
  or _17161_ (_08906_, _08905_, \oc8051_symbolic_cxrom1.regvalid [4]);
  and _17162_ (_08907_, _08906_, _08903_);
  and _17163_ (_08908_, _08793_, _08533_);
  or _17164_ (_08909_, _08897_, _08544_);
  or _17165_ (_08910_, _08909_, _08908_);
  or _17166_ (_08911_, _08910_, _08907_);
  and _17167_ (_07279_, _08911_, _06444_);
  and _17168_ (_08912_, _06364_, _06671_);
  and _17169_ (_08913_, _08912_, _07962_);
  and _17170_ (_08914_, _08913_, _06933_);
  nand _17171_ (_08915_, _08914_, _06930_);
  or _17172_ (_08916_, _08914_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and _17173_ (_08917_, _08916_, _06674_);
  and _17174_ (_08918_, _08917_, _08915_);
  and _17175_ (_08919_, _08913_, _06942_);
  not _17176_ (_08920_, _08919_);
  nor _17177_ (_08921_, _08920_, _06978_);
  and _17178_ (_08922_, _08920_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or _17179_ (_08923_, _08922_, _08921_);
  and _17180_ (_08924_, _08923_, _06440_);
  not _17181_ (_08925_, _06673_);
  and _17182_ (_08926_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or _17183_ (_08927_, _08926_, rst);
  or _17184_ (_08928_, _08927_, _08924_);
  or _17185_ (_07328_, _08928_, _08918_);
  not _17186_ (_08929_, _08730_);
  and _17187_ (_08930_, _08613_, _08536_);
  or _17188_ (_08931_, _08905_, _08930_);
  or _17189_ (_08932_, _08931_, _08929_);
  and _17190_ (_08933_, _08932_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and _17191_ (_08934_, _08904_, _08644_);
  and _17192_ (_08935_, _08898_, \oc8051_symbolic_cxrom1.regvalid [5]);
  or _17193_ (_08936_, _08935_, _08934_);
  nor _17194_ (_08937_, _08936_, _08933_);
  nor _17195_ (_08938_, _08937_, _08798_);
  and _17196_ (_08939_, _08891_, \oc8051_symbolic_cxrom1.regvalid [5]);
  or _17197_ (_08940_, _08939_, _08898_);
  or _17198_ (_08941_, _08940_, _08905_);
  or _17199_ (_08942_, _08941_, _08930_);
  or _17200_ (_08944_, _08942_, _08938_);
  and _17201_ (_07337_, _08944_, _06444_);
  and _17202_ (_08946_, _08792_, _08532_);
  or _17203_ (_08947_, _08619_, _08946_);
  or _17204_ (_08949_, _08790_, _08731_);
  or _17205_ (_08950_, _08489_, _08480_);
  nor _17206_ (_08952_, _08950_, _08514_);
  and _17207_ (_08953_, _08931_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or _17208_ (_08955_, _08953_, _08952_);
  and _17209_ (_08956_, _08903_, \oc8051_symbolic_cxrom1.regvalid [6]);
  and _17210_ (_08958_, _08956_, _08950_);
  and _17211_ (_08959_, _08898_, \oc8051_symbolic_cxrom1.regvalid [6]);
  and _17212_ (_08961_, _08891_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or _17213_ (_08962_, _08961_, _08959_);
  or _17214_ (_08963_, _08962_, _08958_);
  or _17215_ (_08964_, _08963_, _08955_);
  and _17216_ (_08965_, _08964_, _08949_);
  or _17217_ (_08966_, _08953_, _08934_);
  or _17218_ (_08967_, _08966_, _08965_);
  and _17219_ (_08968_, _08967_, _08947_);
  and _17220_ (_08969_, _08964_, _08894_);
  or _17221_ (_08970_, _08961_, _08930_);
  or _17222_ (_08971_, _08970_, _08959_);
  or _17223_ (_08972_, _08971_, _08905_);
  or _17224_ (_08973_, _08972_, _08969_);
  or _17225_ (_08974_, _08973_, _08968_);
  and _17226_ (_07395_, _08974_, _06444_);
  and _17227_ (_08975_, _07644_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1]);
  nor _17228_ (_08976_, _06418_, _06407_);
  and _17229_ (_08977_, _08976_, _06430_);
  and _17230_ (_08978_, _07402_, _07214_);
  and _17231_ (_08979_, _08978_, _08977_);
  nor _17232_ (_08980_, _08979_, _08975_);
  or _17233_ (_08981_, _08980_, _08019_);
  not _17234_ (_08982_, _08980_);
  or _17235_ (_08983_, _08982_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and _17236_ (_08984_, _08983_, _06444_);
  and _17237_ (_07449_, _08984_, _08981_);
  nand _17238_ (_08985_, _07754_, _07686_);
  or _17239_ (_08986_, _07754_, _07686_);
  nand _17240_ (_08987_, _08986_, _08985_);
  nand _17241_ (_08988_, _08987_, _07757_);
  or _17242_ (_08989_, _07757_, _07680_);
  and _17243_ (_08990_, _08989_, _08988_);
  nand _17244_ (_08991_, _08990_, _07459_);
  and _17245_ (_08992_, _08092_, _08089_);
  and _17246_ (_08993_, _07767_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12]);
  nand _17247_ (_08994_, _08993_, _08992_);
  or _17248_ (_08995_, _08993_, _08992_);
  and _17249_ (_08996_, _08995_, _08994_);
  nand _17250_ (_08997_, _08996_, _07602_);
  nor _17251_ (_08998_, _06840_, _06761_);
  nor _17252_ (_08999_, _08998_, _06841_);
  nor _17253_ (_09000_, _08999_, _06681_);
  not _17254_ (_09001_, _09000_);
  nor _17255_ (_09002_, _06874_, _06872_);
  not _17256_ (_09003_, _09002_);
  nor _17257_ (_09004_, _06875_, _06848_);
  and _17258_ (_09005_, _09004_, _09003_);
  and _17259_ (_09006_, _06740_, _06465_);
  nor _17260_ (_09007_, _06732_, _06465_);
  or _17261_ (_09008_, _09007_, _09006_);
  and _17262_ (_09009_, _09008_, _06455_);
  nor _17263_ (_09010_, _06959_, _06957_);
  not _17264_ (_09011_, _09010_);
  and _17265_ (_09012_, _09011_, _06961_);
  and _17266_ (_09013_, _06613_, _06511_);
  nor _17267_ (_09014_, _06732_, _09013_);
  nor _17268_ (_09015_, _09014_, _06955_);
  nor _17269_ (_09016_, _09015_, _06515_);
  nor _17270_ (_09017_, _09016_, _09012_);
  nor _17271_ (_09018_, _09017_, _06621_);
  nor _17272_ (_09019_, _09018_, _09009_);
  nor _17273_ (_09020_, _08111_, _06732_);
  and _17274_ (_09021_, _08111_, _06732_);
  nor _17275_ (_09022_, _09021_, _09020_);
  nor _17276_ (_09023_, _09022_, _06891_);
  and _17277_ (_09024_, _06744_, _06647_);
  and _17278_ (_09025_, _06742_, _06658_);
  nor _17279_ (_09026_, _06743_, _06655_);
  and _17280_ (_09027_, _06732_, _06660_);
  or _17281_ (_09028_, _09027_, _09026_);
  or _17282_ (_09029_, _09028_, _09025_);
  nor _17283_ (_09030_, _09029_, _09024_);
  or _17284_ (_09031_, _06697_, _07933_);
  nor _17285_ (_09032_, _06638_, _06511_);
  and _17286_ (_09033_, _06957_, _06640_);
  nor _17287_ (_09034_, _09033_, _09032_);
  and _17288_ (_09035_, _09034_, _09031_);
  and _17289_ (_09036_, _09035_, _09030_);
  not _17290_ (_09037_, _09036_);
  nor _17291_ (_09038_, _09037_, _09023_);
  and _17292_ (_09039_, _09038_, _09019_);
  not _17293_ (_09040_, _09039_);
  nor _17294_ (_09041_, _09040_, _09005_);
  and _17295_ (_09042_, _09041_, _09001_);
  and _17296_ (_09043_, _09042_, _08997_);
  and _17297_ (_09045_, _09043_, _08991_);
  nand _17298_ (_09046_, _09045_, _08982_);
  or _17299_ (_09048_, _08982_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and _17300_ (_09049_, _09048_, _06444_);
  and _17301_ (_07452_, _09049_, _09046_);
  or _17302_ (_09051_, _08980_, _08127_);
  or _17303_ (_09052_, _08982_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and _17304_ (_09053_, _09052_, _06444_);
  and _17305_ (_07455_, _09053_, _09051_);
  or _17306_ (_09054_, _08980_, _08230_);
  or _17307_ (_09055_, _08982_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and _17308_ (_09056_, _09055_, _06444_);
  and _17309_ (_07469_, _09056_, _09054_);
  not _17310_ (_09057_, _08622_);
  and _17311_ (_09059_, _08536_, \oc8051_symbolic_cxrom1.regvalid [7]);
  or _17312_ (_09060_, _08952_, _08489_);
  and _17313_ (_09062_, _09060_, \oc8051_symbolic_cxrom1.regvalid [7]);
  not _17314_ (_09063_, \oc8051_symbolic_cxrom1.regvalid [7]);
  nor _17315_ (_09064_, _08496_, _09063_);
  and _17316_ (_09065_, _09064_, _08904_);
  or _17317_ (_09066_, _09065_, _08620_);
  or _17318_ (_09067_, _09066_, _09062_);
  or _17319_ (_09068_, _09067_, _09059_);
  and _17320_ (_09069_, _09068_, _09057_);
  and _17321_ (_09070_, _08837_, \oc8051_symbolic_cxrom1.regvalid [7]);
  and _17322_ (_09071_, _09070_, _08480_);
  and _17323_ (_09072_, _08898_, \oc8051_symbolic_cxrom1.regvalid [7]);
  or _17324_ (_09073_, _09065_, _08952_);
  or _17325_ (_09074_, _09073_, _09072_);
  or _17326_ (_09075_, _09074_, _09071_);
  or _17327_ (_09076_, _09075_, _09069_);
  and _17328_ (_09077_, _09076_, _08949_);
  and _17329_ (_09078_, _09068_, _08894_);
  or _17330_ (_09079_, _09059_, _08905_);
  or _17331_ (_09080_, _09079_, _08934_);
  or _17332_ (_09081_, _09080_, _09078_);
  or _17333_ (_09082_, _09081_, _09077_);
  and _17334_ (_07485_, _09082_, _06444_);
  or _17335_ (_09083_, _08980_, _08308_);
  or _17336_ (_09084_, _08982_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and _17337_ (_09085_, _09084_, _06444_);
  and _17338_ (_07494_, _09085_, _09083_);
  not _17339_ (_09086_, _07459_);
  and _17340_ (_09087_, _07743_, _07734_);
  not _17341_ (_09088_, _09087_);
  and _17342_ (_09089_, _09088_, _07744_);
  nor _17343_ (_09090_, _09089_, _07758_);
  nor _17344_ (_09091_, _07757_, _07740_);
  or _17345_ (_09092_, _09091_, _09090_);
  or _17346_ (_09093_, _09092_, _09086_);
  or _17347_ (_09094_, _08280_, _08082_);
  and _17348_ (_09095_, _09094_, _08281_);
  nand _17349_ (_09096_, _09095_, _07602_);
  nor _17350_ (_09097_, _06829_, _06820_);
  nor _17351_ (_09098_, _09097_, _06830_);
  nor _17352_ (_09099_, _09098_, _06681_);
  not _17353_ (_09100_, _09099_);
  nor _17354_ (_09101_, _06864_, _06862_);
  not _17355_ (_09102_, _09101_);
  nor _17356_ (_09103_, _06865_, _06848_);
  and _17357_ (_09104_, _09103_, _09102_);
  not _17358_ (_09105_, _09104_);
  nor _17359_ (_09106_, _06785_, _06951_);
  and _17360_ (_09107_, _07049_, _06465_);
  and _17361_ (_09108_, _06588_, _06515_);
  nor _17362_ (_09109_, _09108_, _09107_);
  nor _17363_ (_09110_, _09109_, _06605_);
  and _17364_ (_09111_, _09109_, _06605_);
  or _17365_ (_09112_, _09111_, _09110_);
  and _17366_ (_09113_, _09112_, _06620_);
  nor _17367_ (_09114_, _09113_, _09106_);
  and _17368_ (_09115_, _06610_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor _17369_ (_09116_, _07945_, _06604_);
  nor _17370_ (_09117_, _09116_, _09115_);
  nor _17371_ (_09118_, _09117_, _06891_);
  nor _17372_ (_09119_, _06787_, _06655_);
  and _17373_ (_09120_, _06788_, _06647_);
  nor _17374_ (_09121_, _09120_, _09119_);
  and _17375_ (_09122_, _06786_, _06658_);
  and _17376_ (_09123_, _06660_, _06604_);
  nor _17377_ (_09124_, _09123_, _09122_);
  or _17378_ (_09125_, _07933_, _06551_);
  nor _17379_ (_09126_, _06638_, _06570_);
  and _17380_ (_09127_, _06640_, _06605_);
  nor _17381_ (_09128_, _09127_, _09126_);
  and _17382_ (_09129_, _09128_, _09125_);
  and _17383_ (_09130_, _09129_, _09124_);
  and _17384_ (_09131_, _09130_, _09121_);
  not _17385_ (_09132_, _09131_);
  nor _17386_ (_09133_, _09132_, _09118_);
  and _17387_ (_09134_, _09133_, _09114_);
  and _17388_ (_09135_, _09134_, _09105_);
  and _17389_ (_09136_, _09135_, _09100_);
  and _17390_ (_09137_, _09136_, _09096_);
  and _17391_ (_09138_, _09137_, _09093_);
  nand _17392_ (_09139_, _09138_, _08982_);
  or _17393_ (_09140_, _08982_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and _17394_ (_09141_, _09140_, _06444_);
  and _17395_ (_07498_, _09141_, _09139_);
  or _17396_ (_09142_, _08980_, _07959_);
  or _17397_ (_09143_, _08982_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and _17398_ (_09144_, _09143_, _06444_);
  and _17399_ (_07514_, _09144_, _09142_);
  or _17400_ (_09145_, _08800_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and _17401_ (_07563_, _09145_, _06444_);
  not _17402_ (_09146_, _07414_);
  nor _17403_ (_09147_, _09146_, _06666_);
  and _17404_ (_09149_, _09146_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  or _17405_ (_09151_, _09149_, _07158_);
  or _17406_ (_09152_, _09151_, _09147_);
  or _17407_ (_09154_, _06439_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  and _17408_ (_09155_, _09154_, _06444_);
  and _17409_ (_07623_, _09155_, _09152_);
  and _17410_ (_09157_, _08978_, _08310_);
  not _17411_ (_09158_, _09157_);
  nor _17412_ (_09160_, _09158_, _09045_);
  and _17413_ (_09161_, _09158_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or _17414_ (_09163_, _09161_, _08975_);
  or _17415_ (_09164_, _09163_, _09160_);
  and _17416_ (_09165_, _06740_, _06640_);
  and _17417_ (_09167_, _06913_, _06605_);
  or _17418_ (_09168_, _06752_, _06482_);
  and _17419_ (_09169_, _09168_, _06515_);
  or _17420_ (_09171_, _09169_, _06484_);
  or _17421_ (_09172_, _09171_, _08170_);
  nor _17422_ (_09173_, _09172_, _08248_);
  and _17423_ (_09174_, _09173_, _06739_);
  nor _17424_ (_09175_, _09173_, _06739_);
  or _17425_ (_09176_, _09175_, _09174_);
  and _17426_ (_09177_, _09176_, _06620_);
  nor _17427_ (_09178_, _06739_, _06465_);
  nor _17428_ (_09179_, _06732_, _06515_);
  or _17429_ (_09180_, _09179_, _09178_);
  and _17430_ (_09181_, _09180_, _06455_);
  or _17431_ (_09182_, _09181_, _09177_);
  or _17432_ (_09183_, _09182_, _09167_);
  and _17433_ (_09184_, _07459_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  nor _17434_ (_09185_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  not _17435_ (_09186_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and _17436_ (_09187_, _09186_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _17437_ (_09188_, _09187_, _09185_);
  nor _17438_ (_09189_, _09188_, _08159_);
  not _17439_ (_09190_, _09189_);
  and _17440_ (_09191_, _09188_, _08159_);
  nor _17441_ (_09192_, _09191_, _06848_);
  and _17442_ (_09193_, _09192_, _09190_);
  and _17443_ (_09194_, _07910_, _07880_);
  not _17444_ (_09195_, _09194_);
  and _17445_ (_09196_, _09195_, _07911_);
  and _17446_ (_09197_, _09196_, _07602_);
  or _17447_ (_09198_, _09197_, _09193_);
  or _17448_ (_09199_, _09198_, _09184_);
  or _17449_ (_09200_, _09199_, _09183_);
  nor _17450_ (_09201_, _09200_, _09165_);
  nand _17451_ (_09202_, _09201_, _08975_);
  and _17452_ (_09203_, _09202_, _06444_);
  and _17453_ (_07645_, _09203_, _09164_);
  and _17454_ (_09204_, _09157_, _08127_);
  and _17455_ (_09205_, _09158_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or _17456_ (_09206_, _09205_, _08975_);
  or _17457_ (_09207_, _09206_, _09204_);
  not _17458_ (_09208_, _08975_);
  or _17459_ (_09209_, _09208_, _08194_);
  and _17460_ (_09210_, _09209_, _06444_);
  and _17461_ (_07648_, _09210_, _09207_);
  and _17462_ (_09211_, _09157_, _08230_);
  and _17463_ (_09212_, _09158_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or _17464_ (_09213_, _09212_, _08975_);
  or _17465_ (_09214_, _09213_, _09211_);
  or _17466_ (_09215_, _09208_, _08267_);
  and _17467_ (_09216_, _09215_, _06444_);
  and _17468_ (_07658_, _09216_, _09214_);
  not _17469_ (_09217_, _08793_);
  and _17470_ (_09218_, _08619_, _09217_);
  nor _17471_ (_09219_, _08896_, _08532_);
  nor _17472_ (_09220_, _08730_, _08521_);
  or _17473_ (_09221_, _09220_, _09219_);
  and _17474_ (_09222_, _09221_, _09218_);
  and _17475_ (_09223_, _08793_, _08489_);
  nor _17476_ (_09224_, _08489_, _08521_);
  and _17477_ (_09225_, _09224_, _08513_);
  or _17478_ (_09226_, _09225_, _09223_);
  or _17479_ (_09227_, _09226_, _09222_);
  and _17480_ (_09228_, _09227_, _08619_);
  or _17481_ (_09229_, _08934_, _08837_);
  and _17482_ (_09230_, _09229_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and _17483_ (_09231_, _09221_, _08894_);
  and _17484_ (_09232_, _09224_, _08793_);
  or _17485_ (_09233_, _09232_, _08952_);
  or _17486_ (_09235_, _09233_, _09231_);
  or _17487_ (_09236_, _09235_, _09230_);
  or _17488_ (_09237_, _09236_, _08620_);
  or _17489_ (_09238_, _09237_, _09228_);
  and _17490_ (_07663_, _09238_, _06444_);
  and _17491_ (_09239_, _09157_, _08308_);
  and _17492_ (_09241_, _09158_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or _17493_ (_09242_, _09241_, _08975_);
  or _17494_ (_09243_, _09242_, _09239_);
  or _17495_ (_09244_, _09208_, _08342_);
  and _17496_ (_09246_, _09244_, _06444_);
  and _17497_ (_07678_, _09246_, _09243_);
  nor _17498_ (_09247_, _09158_, _09138_);
  and _17499_ (_09249_, _09158_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or _17500_ (_09250_, _09249_, _08975_);
  or _17501_ (_09251_, _09250_, _09247_);
  and _17502_ (_09252_, _06812_, _06640_);
  and _17503_ (_09254_, _06957_, _06913_);
  nor _17504_ (_09255_, _06604_, _06951_);
  nor _17505_ (_09256_, _08171_, _06465_);
  nor _17506_ (_09257_, _08322_, _06515_);
  or _17507_ (_09259_, _09257_, _09256_);
  and _17508_ (_09260_, _09259_, _06785_);
  nor _17509_ (_09262_, _09259_, _06785_);
  nor _17510_ (_09263_, _09262_, _09260_);
  and _17511_ (_09264_, _09263_, _06620_);
  or _17512_ (_09266_, _09264_, _09255_);
  or _17513_ (_09267_, _09266_, _09254_);
  and _17514_ (_09268_, _07459_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  nor _17515_ (_09269_, _08145_, _07599_);
  not _17516_ (_09271_, _09269_);
  nor _17517_ (_09272_, _08146_, _06848_);
  and _17518_ (_09273_, _09272_, _09271_);
  nor _17519_ (_09274_, _07898_, _07895_);
  nor _17520_ (_09275_, _09274_, _07899_);
  and _17521_ (_09276_, _09275_, _07602_);
  or _17522_ (_09277_, _09276_, _09273_);
  or _17523_ (_09278_, _09277_, _09268_);
  or _17524_ (_09279_, _09278_, _09267_);
  nor _17525_ (_09280_, _09279_, _09252_);
  nand _17526_ (_09281_, _09280_, _08975_);
  and _17527_ (_09282_, _09281_, _06444_);
  and _17528_ (_07702_, _09282_, _09251_);
  and _17529_ (_09283_, _09157_, _07959_);
  and _17530_ (_09284_, _09158_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or _17531_ (_09285_, _09284_, _08975_);
  or _17532_ (_09286_, _09285_, _09283_);
  nand _17533_ (_09287_, _08975_, _07640_);
  and _17534_ (_09288_, _09287_, _06444_);
  and _17535_ (_07705_, _09288_, _09286_);
  and _17536_ (_09289_, _09157_, _08019_);
  and _17537_ (_09290_, _09158_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or _17538_ (_09291_, _09290_, _08975_);
  or _17539_ (_09292_, _09291_, _09289_);
  nand _17540_ (_09293_, _08975_, _08060_);
  and _17541_ (_09294_, _09293_, _06444_);
  and _17542_ (_07710_, _09294_, _09292_);
  and _17543_ (_09295_, _08619_, _08524_);
  or _17544_ (_09296_, _09295_, _08894_);
  and _17545_ (_09297_, _08655_, _08842_);
  nand _17546_ (_09298_, _08614_, _08896_);
  and _17547_ (_09299_, _09298_, _08551_);
  or _17548_ (_09300_, _09299_, _09297_);
  and _17549_ (_09301_, _08708_, \oc8051_symbolic_cxrom1.regvalid [10]);
  not _17550_ (_09302_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor _17551_ (_09303_, _08665_, _09302_);
  and _17552_ (_09304_, _09303_, _08837_);
  or _17553_ (_09305_, _09304_, _09301_);
  or _17554_ (_09306_, _09305_, _09300_);
  or _17555_ (_09307_, _08620_, _09223_);
  and _17556_ (_09308_, _09307_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor _17557_ (_09309_, _08950_, _08524_);
  and _17558_ (_09310_, _09309_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or _17559_ (_09311_, _09310_, _09308_);
  or _17560_ (_09312_, _09311_, _09306_);
  and _17561_ (_09313_, _09312_, _09296_);
  and _17562_ (_09314_, _08523_, _08489_);
  and _17563_ (_09315_, _08730_, _08524_);
  and _17564_ (_09316_, _09315_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and _17565_ (_09317_, _08952_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and _17566_ (_09318_, _08891_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or _17567_ (_09319_, _09318_, _08620_);
  or _17568_ (_09320_, _09319_, _09317_);
  or _17569_ (_09321_, _09320_, _09316_);
  or _17570_ (_09322_, _09321_, _09314_);
  or _17571_ (_09323_, _09322_, _09313_);
  and _17572_ (_07759_, _09323_, _06444_);
  nand _17573_ (_09324_, _08408_, _07231_);
  nor _17574_ (_09325_, _07230_, \oc8051_top_1.oc8051_decoder1.op [2]);
  nor _17575_ (_09326_, _09325_, _07265_);
  and _17576_ (_09327_, _09326_, _09324_);
  and _17577_ (_07809_, _09327_, _06444_);
  or _17578_ (_09328_, _07420_, _07159_);
  and _17579_ (_09329_, _09328_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  not _17580_ (_09330_, _07154_);
  nor _17581_ (_09331_, _07414_, _07416_);
  nand _17582_ (_09332_, _09331_, _09330_);
  and _17583_ (_09334_, _06439_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  and _17584_ (_09335_, _09334_, _09332_);
  and _17585_ (_09336_, _07425_, _07070_);
  or _17586_ (_09337_, _09336_, _09335_);
  or _17587_ (_09338_, _09337_, _09329_);
  and _17588_ (_07824_, _09338_, _06444_);
  not _17589_ (_09339_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and _17590_ (_09340_, _06295_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  and _17591_ (_09341_, _09340_, \oc8051_top_1.oc8051_sfr1.pres_ow );
  not _17592_ (_09342_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  nor _17593_ (_09343_, _06295_, _09342_);
  and _17594_ (_09344_, _09343_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re );
  not _17595_ (_09345_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  nor _17596_ (_09346_, _09345_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  not _17597_ (_09347_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  nor _17598_ (_09348_, _09347_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  and _17599_ (_09349_, _09348_, _09346_);
  and _17600_ (_09350_, _09349_, _09344_);
  nor _17601_ (_09351_, _09350_, _09341_);
  not _17602_ (_09352_, _09351_);
  and _17603_ (_09353_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and _17604_ (_09354_, _09353_, _06296_);
  not _17605_ (_09355_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  nor _17606_ (_09356_, _09355_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  and _17607_ (_09357_, _09356_, _09342_);
  and _17608_ (_09358_, _09357_, _06295_);
  nor _17609_ (_09359_, _09358_, _09354_);
  nor _17610_ (_09360_, _09359_, _09344_);
  nor _17611_ (_09361_, _09360_, _09352_);
  nor _17612_ (_09362_, _09361_, _09339_);
  or _17613_ (_09363_, _09362_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2]);
  or _17614_ (_09364_, _09339_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  or _17615_ (_09365_, _09364_, _09351_);
  and _17616_ (_09366_, _09365_, _06444_);
  and _17617_ (_07849_, _09366_, _09363_);
  and _17618_ (_09367_, _09339_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  and _17619_ (_09368_, _09367_, _06444_);
  or _17620_ (_09369_, _09360_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  and _17621_ (_09370_, _09369_, _09351_);
  and _17622_ (_09371_, _09352_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  or _17623_ (_09372_, _09371_, _09370_);
  and _17624_ (_09373_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _06444_);
  and _17625_ (_09374_, _09373_, _09372_);
  or _17626_ (_07852_, _09374_, _09368_);
  and _17627_ (_09375_, _09339_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  and _17628_ (_09376_, _09375_, _06444_);
  or _17629_ (_09377_, _09360_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  and _17630_ (_09378_, _09377_, _09351_);
  and _17631_ (_09379_, _09352_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  or _17632_ (_09380_, _09379_, _09378_);
  and _17633_ (_09381_, _09380_, _09373_);
  or _17634_ (_07855_, _09381_, _09376_);
  and _17635_ (_09382_, _09339_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  and _17636_ (_09383_, _09382_, _06444_);
  or _17637_ (_09384_, _09352_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  or _17638_ (_09385_, _09384_, _09360_);
  or _17639_ (_09386_, _09351_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  and _17640_ (_09387_, _09386_, _09373_);
  and _17641_ (_09388_, _09387_, _09385_);
  or _17642_ (_07860_, _09388_, _09383_);
  and _17643_ (_09389_, _09339_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  and _17644_ (_09390_, _09389_, _06444_);
  or _17645_ (_09391_, _09360_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  and _17646_ (_09392_, _09391_, _09351_);
  and _17647_ (_09393_, _09352_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  or _17648_ (_09394_, _09393_, _09392_);
  and _17649_ (_09395_, _09394_, _09373_);
  or _17650_ (_07863_, _09395_, _09390_);
  or _17651_ (_09396_, _08620_, _09309_);
  and _17652_ (_09397_, _08666_, _08536_);
  or _17653_ (_09398_, _09397_, _09396_);
  and _17654_ (_09399_, _09398_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and _17655_ (_09400_, _08613_, _08842_);
  and _17656_ (_09401_, _08819_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or _17657_ (_09402_, _09401_, _09400_);
  and _17658_ (_09403_, _08708_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or _17659_ (_09404_, _09403_, _09223_);
  or _17660_ (_09405_, _09404_, _09297_);
  or _17661_ (_09406_, _09405_, _09402_);
  or _17662_ (_09407_, _09406_, _09219_);
  or _17663_ (_09408_, _09407_, _09399_);
  and _17664_ (_07867_, _09408_, _06444_);
  or _17665_ (_09409_, _09362_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1]);
  or _17666_ (_09411_, _09339_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2]);
  or _17667_ (_09412_, _09411_, _09351_);
  and _17668_ (_09413_, _09412_, _06444_);
  and _17669_ (_07876_, _09413_, _09409_);
  and _17670_ (_09414_, _07912_, _07872_);
  not _17671_ (_09415_, _09414_);
  and _17672_ (_09416_, _09415_, _07913_);
  and _17673_ (_07878_, _09416_, _06444_);
  and _17674_ (_09417_, _09339_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  and _17675_ (_09418_, _09417_, _06444_);
  or _17676_ (_09419_, _09360_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  and _17677_ (_09420_, _09419_, _09351_);
  and _17678_ (_09421_, _09352_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  or _17679_ (_09422_, _09421_, _09420_);
  and _17680_ (_09423_, _09422_, _09373_);
  or _17681_ (_07909_, _09423_, _09418_);
  and _17682_ (_09424_, _09339_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  and _17683_ (_09425_, _09424_, _06444_);
  and _17684_ (_09426_, _09352_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  nor _17685_ (_09427_, _09358_, _09344_);
  and _17686_ (_09428_, _09427_, _09354_);
  or _17687_ (_09429_, _09428_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  not _17688_ (_09430_, _09341_);
  not _17689_ (_09431_, _09349_);
  and _17690_ (_09432_, _09431_, _09344_);
  or _17691_ (_09433_, _09427_, _09432_);
  and _17692_ (_09434_, _09433_, _09430_);
  and _17693_ (_09436_, _09434_, _09429_);
  or _17694_ (_09437_, _09436_, _09426_);
  and _17695_ (_09438_, _09437_, _09373_);
  or _17696_ (_07934_, _09438_, _09425_);
  nor _17697_ (_09439_, _07188_, _06449_);
  and _17698_ (_09440_, _06449_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  or _17699_ (_09441_, _09440_, _09439_);
  and _17700_ (_07954_, _09441_, _06444_);
  nor _17701_ (_07964_, _07302_, rst);
  or _17702_ (_09442_, _09362_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  or _17703_ (_09443_, _09339_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1]);
  or _17704_ (_09444_, _09443_, _09351_);
  and _17705_ (_09445_, _09444_, _06444_);
  and _17706_ (_07970_, _09445_, _09442_);
  and _17707_ (_09447_, _09349_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  and _17708_ (_09448_, _09447_, _09359_);
  or _17709_ (_09450_, _09448_, _09361_);
  and _17710_ (_09451_, _09450_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  and _17711_ (_09452_, _09339_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  nand _17712_ (_09453_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor _17713_ (_09454_, _09453_, _09351_);
  or _17714_ (_09455_, _09454_, _09452_);
  or _17715_ (_09456_, _09455_, _09451_);
  and _17716_ (_07973_, _09456_, _06444_);
  and _17717_ (_09457_, _08797_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and _17718_ (_09458_, _08544_, \oc8051_symbolic_cxrom1.regvalid [12]);
  or _17719_ (_09459_, _08897_, _08793_);
  and _17720_ (_09460_, _09459_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and _17721_ (_09461_, _08904_, \oc8051_symbolic_cxrom1.regvalid [12]);
  or _17722_ (_09462_, _09461_, _08842_);
  or _17723_ (_09463_, _09462_, _09460_);
  or _17724_ (_09464_, _09463_, _09458_);
  or _17725_ (_09465_, _09464_, _09457_);
  and _17726_ (_07977_, _09465_, _06444_);
  not _17727_ (_09466_, _09362_);
  and _17728_ (_09467_, _06444_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  and _17729_ (_09468_, _09467_, _09466_);
  and _17730_ (_09469_, _09349_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  and _17731_ (_09470_, _09469_, _09359_);
  or _17732_ (_09471_, _09470_, _09352_);
  and _17733_ (_09472_, _09373_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  and _17734_ (_09473_, _09472_, _09471_);
  or _17735_ (_07983_, _09473_, _09468_);
  or _17736_ (_09474_, _08392_, _07232_);
  nor _17737_ (_09475_, _07230_, \oc8051_top_1.oc8051_decoder1.op [1]);
  nor _17738_ (_09476_, _09475_, _07265_);
  and _17739_ (_09477_, _09476_, _09474_);
  and _17740_ (_07992_, _09477_, _06444_);
  and _17741_ (_09478_, _06944_, _08310_);
  and _17742_ (_09479_, _09478_, _06941_);
  nand _17743_ (_09480_, _09479_, _06978_);
  and _17744_ (_09481_, _07028_, _07015_);
  not _17745_ (_09482_, _09481_);
  and _17746_ (_09483_, _06944_, _08977_);
  and _17747_ (_09484_, _09483_, _06941_);
  nor _17748_ (_09485_, _09484_, _09482_);
  not _17749_ (_09486_, _09485_);
  and _17750_ (_09487_, _09486_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  and _17751_ (_09488_, _09485_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  or _17752_ (_09489_, _09488_, _09487_);
  or _17753_ (_09490_, _09489_, _09479_);
  and _17754_ (_09491_, _09490_, _06444_);
  and _17755_ (_08068_, _09491_, _09480_);
  and _17756_ (_08075_, _07268_, _06444_);
  and _17757_ (_09492_, _08726_, _08731_);
  or _17758_ (_09493_, _09492_, \oc8051_symbolic_cxrom1.regvalid [13]);
  and _17759_ (_08118_, _09493_, _06444_);
  nor _17760_ (_09494_, t2_i, rst);
  and _17761_ (_08140_, _09494_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r );
  not _17762_ (_09495_, _07006_);
  and _17763_ (_09496_, _07013_, _07011_);
  and _17764_ (_09497_, _09496_, _06990_);
  nand _17765_ (_09498_, _09497_, _09495_);
  or _17766_ (_09499_, _09497_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  and _17767_ (_09500_, _09499_, _06444_);
  and _17768_ (_08149_, _09500_, _09498_);
  nand _17769_ (_09501_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r , _06444_);
  nor _17770_ (_08189_, _09501_, t2ex_i);
  and _17771_ (_08204_, t2ex_i, _06444_);
  nand _17772_ (_09502_, _06985_, _06978_);
  not _17773_ (_09503_, _06989_);
  and _17774_ (_09504_, _07017_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and _17775_ (_09505_, _07029_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and _17776_ (_09506_, _09505_, _07026_);
  and _17777_ (_09507_, _07011_, _06997_);
  or _17778_ (_09508_, _09507_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  nand _17779_ (_09509_, _09507_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and _17780_ (_09510_, _09509_, _09508_);
  or _17781_ (_09511_, _09510_, _09506_);
  and _17782_ (_09512_, _09511_, _07035_);
  or _17783_ (_09513_, _09512_, _09504_);
  or _17784_ (_09514_, _09513_, _06985_);
  and _17785_ (_09515_, _09514_, _09503_);
  and _17786_ (_09516_, _09515_, _09502_);
  and _17787_ (_09517_, _06989_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or _17788_ (_09518_, _09517_, _09516_);
  and _17789_ (_08219_, _09518_, _06444_);
  or _17790_ (_09519_, _08679_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and _17791_ (_08240_, _09519_, _06444_);
  and _17792_ (_09520_, _09328_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  and _17793_ (_09521_, _06439_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  and _17794_ (_09522_, _09521_, _09332_);
  nor _17795_ (_09523_, _06644_, _06587_);
  not _17796_ (_09524_, _09523_);
  and _17797_ (_09525_, _09524_, _08004_);
  and _17798_ (_09526_, _09525_, _07998_);
  not _17799_ (_09527_, _09526_);
  and _17800_ (_09528_, _09527_, _07425_);
  or _17801_ (_09529_, _09528_, _09522_);
  or _17802_ (_09530_, _09529_, _09520_);
  and _17803_ (_08409_, _09530_, _06444_);
  and _17804_ (_09531_, _08875_, _08496_);
  not _17805_ (_09532_, _09531_);
  not _17806_ (_09533_, _08872_);
  and _17807_ (_09534_, _08875_, _09533_);
  and _17808_ (_09535_, _09534_, _09532_);
  and _17809_ (_09536_, _09535_, _08536_);
  not _17810_ (_09537_, _09536_);
  or _17811_ (_09538_, _09537_, word_in[0]);
  and _17812_ (_09539_, _08869_, _08894_);
  not _17813_ (_09540_, _09539_);
  or _17814_ (_09541_, _09536_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  and _17815_ (_09542_, _09541_, _09540_);
  and _17816_ (_09543_, _09542_, _09538_);
  and _17817_ (_09544_, _08863_, _08790_);
  and _17818_ (_09545_, _09539_, word_in[8]);
  or _17819_ (_09546_, _09545_, _09544_);
  or _17820_ (_09547_, _09546_, _09543_);
  and _17821_ (_09548_, _08855_, _08820_);
  not _17822_ (_09549_, _09548_);
  not _17823_ (_09550_, _09544_);
  or _17824_ (_09551_, _09550_, word_in[16]);
  and _17825_ (_09552_, _09551_, _09549_);
  and _17826_ (_09553_, _09552_, _09547_);
  and _17827_ (_09554_, _08855_, word_in[24]);
  and _17828_ (_09555_, _09554_, _09548_);
  or _17829_ (_08621_, _09555_, _09553_);
  not _17830_ (_09556_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  nor _17831_ (_09557_, _09536_, _09556_);
  and _17832_ (_09558_, _09536_, word_in[1]);
  or _17833_ (_09559_, _09558_, _09557_);
  and _17834_ (_09560_, _09559_, _09540_);
  and _17835_ (_09562_, _09539_, word_in[9]);
  or _17836_ (_09563_, _09562_, _09560_);
  and _17837_ (_09564_, _09563_, _09550_);
  and _17838_ (_09565_, _08863_, word_in[17]);
  and _17839_ (_09567_, _09565_, _09544_);
  or _17840_ (_09568_, _09567_, _09564_);
  and _17841_ (_09569_, _09568_, _09549_);
  and _17842_ (_09570_, _09548_, word_in[25]);
  or _17843_ (_08625_, _09570_, _09569_);
  or _17844_ (_09572_, _09537_, word_in[2]);
  or _17845_ (_09573_, _09536_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  and _17846_ (_09574_, _09573_, _09540_);
  and _17847_ (_09575_, _09574_, _09572_);
  and _17848_ (_09576_, _09539_, word_in[10]);
  or _17849_ (_09577_, _09576_, _09544_);
  or _17850_ (_09578_, _09577_, _09575_);
  or _17851_ (_09579_, _09550_, word_in[18]);
  and _17852_ (_09580_, _09579_, _09549_);
  and _17853_ (_09581_, _09580_, _09578_);
  and _17854_ (_09582_, _08855_, word_in[26]);
  and _17855_ (_09583_, _09582_, _09548_);
  or _17856_ (_08629_, _09583_, _09581_);
  or _17857_ (_09584_, _09537_, word_in[3]);
  or _17858_ (_09585_, _09536_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  and _17859_ (_09586_, _09585_, _09540_);
  and _17860_ (_09587_, _09586_, _09584_);
  and _17861_ (_09588_, _09539_, word_in[11]);
  or _17862_ (_09589_, _09588_, _09544_);
  or _17863_ (_09591_, _09589_, _09587_);
  or _17864_ (_09592_, _09550_, word_in[19]);
  and _17865_ (_09593_, _09592_, _09549_);
  and _17866_ (_09595_, _09593_, _09591_);
  and _17867_ (_09596_, _08855_, word_in[27]);
  and _17868_ (_09597_, _09596_, _09548_);
  or _17869_ (_08633_, _09597_, _09595_);
  or _17870_ (_09599_, _09537_, word_in[4]);
  or _17871_ (_09600_, _09536_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  and _17872_ (_09601_, _09600_, _09540_);
  and _17873_ (_09602_, _09601_, _09599_);
  and _17874_ (_09603_, _09539_, word_in[12]);
  or _17875_ (_09604_, _09603_, _09544_);
  or _17876_ (_09605_, _09604_, _09602_);
  or _17877_ (_09606_, _09550_, word_in[20]);
  and _17878_ (_09607_, _09606_, _09549_);
  and _17879_ (_09608_, _09607_, _09605_);
  and _17880_ (_09609_, _08855_, word_in[28]);
  and _17881_ (_09611_, _09609_, _09548_);
  or _17882_ (_08637_, _09611_, _09608_);
  or _17883_ (_09612_, _09537_, word_in[5]);
  or _17884_ (_09613_, _09536_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  and _17885_ (_09614_, _09613_, _09540_);
  and _17886_ (_09615_, _09614_, _09612_);
  and _17887_ (_09616_, _09539_, word_in[13]);
  or _17888_ (_09617_, _09616_, _09544_);
  or _17889_ (_09618_, _09617_, _09615_);
  or _17890_ (_09620_, _09550_, word_in[21]);
  and _17891_ (_09621_, _09620_, _09549_);
  and _17892_ (_09622_, _09621_, _09618_);
  and _17893_ (_09623_, _08855_, word_in[29]);
  and _17894_ (_09625_, _09623_, _09548_);
  or _17895_ (_08641_, _09625_, _09622_);
  and _17896_ (_09626_, _08855_, word_in[30]);
  and _17897_ (_09627_, _09626_, _09548_);
  or _17898_ (_09628_, _09537_, word_in[6]);
  or _17899_ (_09629_, _09536_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  and _17900_ (_09631_, _09629_, _09540_);
  and _17901_ (_09632_, _09631_, _09628_);
  and _17902_ (_09633_, _09539_, word_in[14]);
  or _17903_ (_09634_, _09633_, _09544_);
  or _17904_ (_09635_, _09634_, _09632_);
  or _17905_ (_09636_, _09550_, word_in[22]);
  and _17906_ (_09637_, _09636_, _09549_);
  and _17907_ (_09638_, _09637_, _09635_);
  or _17908_ (_08647_, _09638_, _09627_);
  nor _17909_ (_09639_, _09536_, _08695_);
  and _17910_ (_09640_, _08875_, word_in[7]);
  and _17911_ (_09641_, _09536_, _09640_);
  or _17912_ (_09642_, _09641_, _09639_);
  and _17913_ (_09643_, _09642_, _09540_);
  and _17914_ (_09644_, _09539_, word_in[15]);
  or _17915_ (_09645_, _09644_, _09544_);
  or _17916_ (_09646_, _09645_, _09643_);
  or _17917_ (_09647_, _09550_, word_in[23]);
  and _17918_ (_09648_, _09647_, _09549_);
  and _17919_ (_09649_, _09648_, _09646_);
  and _17920_ (_09650_, _09548_, word_in[31]);
  or _17921_ (_08650_, _09650_, _09649_);
  nor _17922_ (_09651_, _07300_, _07190_);
  and _17923_ (_09652_, _07190_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  or _17924_ (_09653_, _09652_, _09651_);
  and _17925_ (_08690_, _09653_, _06444_);
  and _17926_ (_09654_, _07429_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  and _17927_ (_09655_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and _17928_ (_09656_, _07248_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and _17929_ (_09657_, _07251_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor _17930_ (_09658_, _09657_, _09656_);
  and _17931_ (_09659_, _07246_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and _17932_ (_09660_, _07238_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor _17933_ (_09661_, _09660_, _09659_);
  not _17934_ (_09662_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor _17935_ (_09663_, _07241_, _09662_);
  and _17936_ (_09664_, _07254_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nor _17937_ (_09665_, _09664_, _09663_);
  and _17938_ (_09666_, _09665_, _09661_);
  and _17939_ (_09667_, _09666_, _09658_);
  nor _17940_ (_09669_, _09667_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _17941_ (_09670_, _09669_, _09655_);
  nor _17942_ (_09671_, _09670_, _07429_);
  nor _17943_ (_09672_, _09671_, _09654_);
  nor _17944_ (_08694_, _09672_, rst);
  nor _17945_ (_09674_, _09354_, _09344_);
  or _17946_ (_09675_, _09674_, _09339_);
  and _17947_ (_09676_, _09675_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  and _17948_ (_09677_, _09344_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and _17949_ (_09678_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  nor _17950_ (_09679_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  nor _17951_ (_09680_, _09679_, _09678_);
  and _17952_ (_09681_, _09680_, _09677_);
  or _17953_ (_09682_, _09681_, _09676_);
  and _17954_ (_08701_, _09682_, _06444_);
  nand _17955_ (_09683_, _09484_, _06978_);
  not _17956_ (_09684_, _09479_);
  and _17957_ (_09685_, _09482_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and _17958_ (_09686_, _09481_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or _17959_ (_09687_, _09686_, _09685_);
  or _17960_ (_09688_, _09687_, _09484_);
  and _17961_ (_09689_, _09688_, _09684_);
  and _17962_ (_09690_, _09689_, _09683_);
  and _17963_ (_09691_, _09479_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  or _17964_ (_09692_, _09691_, _09690_);
  and _17965_ (_08719_, _09692_, _06444_);
  and _17966_ (_09693_, _08863_, _08613_);
  and _17967_ (_09694_, _09693_, _08732_);
  and _17968_ (_09695_, _08869_, _08611_);
  and _17969_ (_09696_, _09695_, _08626_);
  not _17970_ (_09697_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  and _17971_ (_09698_, _08875_, _08903_);
  and _17972_ (_09699_, _08872_, _08497_);
  not _17973_ (_09700_, _09699_);
  nor _17974_ (_09701_, _09700_, _09698_);
  nor _17975_ (_09702_, _09701_, _09697_);
  and _17976_ (_09703_, _08875_, word_in[0]);
  and _17977_ (_09704_, _09701_, _09703_);
  or _17978_ (_09705_, _09704_, _09702_);
  or _17979_ (_09706_, _09705_, _09696_);
  not _17980_ (_09707_, _09696_);
  or _17981_ (_09709_, _09707_, word_in[8]);
  and _17982_ (_09710_, _09709_, _09706_);
  or _17983_ (_09711_, _09710_, _09694_);
  and _17984_ (_09712_, _08855_, _08790_);
  not _17985_ (_09713_, _09712_);
  not _17986_ (_09714_, _09694_);
  or _17987_ (_09715_, _09714_, word_in[16]);
  and _17988_ (_09716_, _09715_, _09713_);
  and _17989_ (_09717_, _09716_, _09711_);
  and _17990_ (_09718_, _09712_, word_in[24]);
  or _17991_ (_08741_, _09718_, _09717_);
  and _17992_ (_09719_, _09712_, word_in[25]);
  not _17993_ (_09720_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  nor _17994_ (_09721_, _09701_, _09720_);
  and _17995_ (_09722_, _08875_, word_in[1]);
  and _17996_ (_09723_, _09701_, _09722_);
  or _17997_ (_09724_, _09723_, _09721_);
  or _17998_ (_09726_, _09724_, _09696_);
  or _17999_ (_09727_, _09707_, word_in[9]);
  and _18000_ (_09728_, _09727_, _09726_);
  or _18001_ (_09729_, _09728_, _09694_);
  or _18002_ (_09731_, _09714_, word_in[17]);
  and _18003_ (_09732_, _09731_, _09713_);
  and _18004_ (_09733_, _09732_, _09729_);
  or _18005_ (_08743_, _09733_, _09719_);
  not _18006_ (_09734_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  nor _18007_ (_09735_, _09701_, _09734_);
  and _18008_ (_09736_, _08875_, word_in[2]);
  and _18009_ (_09737_, _09701_, _09736_);
  or _18010_ (_09738_, _09737_, _09735_);
  or _18011_ (_09739_, _09738_, _09696_);
  or _18012_ (_09740_, _09707_, word_in[10]);
  and _18013_ (_09741_, _09740_, _09739_);
  or _18014_ (_09743_, _09741_, _09694_);
  or _18015_ (_09744_, _09714_, word_in[18]);
  and _18016_ (_09745_, _09744_, _09713_);
  and _18017_ (_09746_, _09745_, _09743_);
  and _18018_ (_09747_, _09712_, word_in[26]);
  or _18019_ (_08745_, _09747_, _09746_);
  and _18020_ (_09748_, _09712_, word_in[27]);
  not _18021_ (_09749_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  nor _18022_ (_09750_, _09701_, _09749_);
  and _18023_ (_09751_, _08875_, word_in[3]);
  and _18024_ (_09752_, _09701_, _09751_);
  or _18025_ (_09753_, _09752_, _09750_);
  or _18026_ (_09754_, _09753_, _09696_);
  or _18027_ (_09755_, _09707_, word_in[11]);
  and _18028_ (_09756_, _09755_, _09754_);
  or _18029_ (_09757_, _09756_, _09694_);
  or _18030_ (_09758_, _09714_, word_in[19]);
  and _18031_ (_09759_, _09758_, _09713_);
  and _18032_ (_09760_, _09759_, _09757_);
  or _18033_ (_08750_, _09760_, _09748_);
  not _18034_ (_09761_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  nor _18035_ (_09762_, _09701_, _09761_);
  and _18036_ (_09763_, _08875_, word_in[4]);
  and _18037_ (_09764_, _09701_, _09763_);
  or _18038_ (_09765_, _09764_, _09762_);
  or _18039_ (_09766_, _09765_, _09696_);
  or _18040_ (_09767_, _09707_, word_in[12]);
  and _18041_ (_09768_, _09767_, _09766_);
  or _18042_ (_09769_, _09768_, _09694_);
  or _18043_ (_09770_, _09714_, word_in[20]);
  and _18044_ (_09771_, _09770_, _09713_);
  and _18045_ (_09772_, _09771_, _09769_);
  and _18046_ (_09773_, _09712_, word_in[28]);
  or _18047_ (_08755_, _09773_, _09772_);
  and _18048_ (_09774_, _09712_, word_in[29]);
  not _18049_ (_09775_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  nor _18050_ (_09776_, _09701_, _09775_);
  and _18051_ (_09777_, _08875_, word_in[5]);
  and _18052_ (_09778_, _09701_, _09777_);
  or _18053_ (_09779_, _09778_, _09776_);
  or _18054_ (_09780_, _09779_, _09696_);
  or _18055_ (_09781_, _09707_, word_in[13]);
  and _18056_ (_09782_, _09781_, _09780_);
  or _18057_ (_09783_, _09782_, _09694_);
  or _18058_ (_09785_, _09714_, word_in[21]);
  and _18059_ (_09787_, _09785_, _09713_);
  and _18060_ (_09788_, _09787_, _09783_);
  or _18061_ (_08757_, _09788_, _09774_);
  and _18062_ (_09790_, _09712_, word_in[30]);
  not _18063_ (_09792_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  nor _18064_ (_09794_, _09701_, _09792_);
  and _18065_ (_09795_, _08875_, word_in[6]);
  and _18066_ (_09797_, _09701_, _09795_);
  or _18067_ (_09798_, _09797_, _09794_);
  or _18068_ (_09800_, _09798_, _09696_);
  or _18069_ (_09802_, _09707_, word_in[14]);
  and _18070_ (_09803_, _09802_, _09800_);
  or _18071_ (_09804_, _09803_, _09694_);
  or _18072_ (_09805_, _09714_, word_in[22]);
  and _18073_ (_09806_, _09805_, _09713_);
  and _18074_ (_09807_, _09806_, _09804_);
  or _18075_ (_08762_, _09807_, _09790_);
  nor _18076_ (_09808_, _09701_, _08600_);
  and _18077_ (_09809_, _09701_, _09640_);
  or _18078_ (_09810_, _09809_, _09808_);
  or _18079_ (_09811_, _09810_, _09696_);
  or _18080_ (_09812_, _09707_, word_in[15]);
  and _18081_ (_09813_, _09812_, _09811_);
  or _18082_ (_09814_, _09813_, _09694_);
  or _18083_ (_09815_, _09714_, word_in[23]);
  and _18084_ (_09816_, _09815_, _09713_);
  and _18085_ (_09817_, _09816_, _09814_);
  and _18086_ (_09818_, _09712_, word_in[31]);
  or _18087_ (_08767_, _09818_, _09817_);
  and _18088_ (_09819_, _08869_, _08644_);
  and _18089_ (_09820_, _09819_, _08626_);
  not _18090_ (_09821_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  and _18091_ (_09822_, _09531_, _09533_);
  and _18092_ (_09823_, _09822_, _08536_);
  nor _18093_ (_09824_, _09823_, _09821_);
  and _18094_ (_09825_, _09823_, _09703_);
  or _18095_ (_09826_, _09825_, _09824_);
  or _18096_ (_09827_, _09826_, _09820_);
  and _18097_ (_09828_, _08863_, _08611_);
  and _18098_ (_09829_, _09828_, _08732_);
  not _18099_ (_09830_, _09829_);
  not _18100_ (_09831_, _09820_);
  or _18101_ (_09832_, _09831_, word_in[8]);
  and _18102_ (_09833_, _09832_, _09830_);
  and _18103_ (_09834_, _09833_, _09827_);
  and _18104_ (_09835_, _08855_, _08613_);
  and _18105_ (_09836_, _09835_, _08814_);
  and _18106_ (_09837_, _08863_, word_in[16]);
  and _18107_ (_09838_, _09829_, _09837_);
  or _18108_ (_09839_, _09838_, _09836_);
  or _18109_ (_09840_, _09839_, _09834_);
  not _18110_ (_09841_, _09836_);
  or _18111_ (_09842_, _09841_, word_in[24]);
  and _18112_ (_08851_, _09842_, _09840_);
  not _18113_ (_09843_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  nor _18114_ (_09844_, _09823_, _09843_);
  and _18115_ (_09845_, _09823_, _09722_);
  or _18116_ (_09846_, _09845_, _09844_);
  or _18117_ (_09847_, _09846_, _09820_);
  or _18118_ (_09848_, _09831_, word_in[9]);
  and _18119_ (_09850_, _09848_, _09830_);
  and _18120_ (_09851_, _09850_, _09847_);
  and _18121_ (_09853_, _09829_, word_in[17]);
  or _18122_ (_09854_, _09853_, _09836_);
  or _18123_ (_09855_, _09854_, _09851_);
  or _18124_ (_09856_, _09841_, word_in[25]);
  and _18125_ (_08854_, _09856_, _09855_);
  not _18126_ (_09857_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  nor _18127_ (_09858_, _09823_, _09857_);
  and _18128_ (_09860_, _09823_, _09736_);
  or _18129_ (_09861_, _09860_, _09858_);
  or _18130_ (_09862_, _09861_, _09820_);
  or _18131_ (_09864_, _09831_, word_in[10]);
  and _18132_ (_09865_, _09864_, _09830_);
  and _18133_ (_09866_, _09865_, _09862_);
  and _18134_ (_09867_, _09829_, word_in[18]);
  or _18135_ (_09868_, _09867_, _09866_);
  and _18136_ (_09869_, _09868_, _09841_);
  and _18137_ (_09870_, _09836_, word_in[26]);
  or _18138_ (_08858_, _09870_, _09869_);
  not _18139_ (_09871_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  nor _18140_ (_09873_, _09823_, _09871_);
  and _18141_ (_09874_, _09823_, _09751_);
  or _18142_ (_09875_, _09874_, _09873_);
  or _18143_ (_09876_, _09875_, _09820_);
  or _18144_ (_09878_, _09831_, word_in[11]);
  and _18145_ (_09879_, _09878_, _09830_);
  and _18146_ (_09881_, _09879_, _09876_);
  and _18147_ (_09882_, _09829_, word_in[19]);
  or _18148_ (_09883_, _09882_, _09836_);
  or _18149_ (_09885_, _09883_, _09881_);
  or _18150_ (_09886_, _09841_, word_in[27]);
  and _18151_ (_08861_, _09886_, _09885_);
  and _18152_ (_09888_, _09829_, word_in[20]);
  not _18153_ (_09889_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  nor _18154_ (_09891_, _09823_, _09889_);
  and _18155_ (_09892_, _09823_, _09763_);
  or _18156_ (_09893_, _09892_, _09891_);
  or _18157_ (_09895_, _09893_, _09820_);
  or _18158_ (_09896_, _09831_, word_in[12]);
  and _18159_ (_09897_, _09896_, _09830_);
  and _18160_ (_09898_, _09897_, _09895_);
  or _18161_ (_09899_, _09898_, _09888_);
  and _18162_ (_09900_, _09899_, _09841_);
  and _18163_ (_09901_, _09836_, word_in[28]);
  or _18164_ (_08864_, _09901_, _09900_);
  or _18165_ (_09902_, _09823_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  not _18166_ (_09903_, _09823_);
  or _18167_ (_09904_, _09903_, _09777_);
  and _18168_ (_09905_, _09904_, _09902_);
  or _18169_ (_09906_, _09905_, _09820_);
  or _18170_ (_09907_, _09831_, word_in[13]);
  and _18171_ (_09908_, _09907_, _09906_);
  or _18172_ (_09909_, _09908_, _09829_);
  or _18173_ (_09910_, _09830_, word_in[21]);
  and _18174_ (_09911_, _09910_, _09841_);
  and _18175_ (_09912_, _09911_, _09909_);
  and _18176_ (_09913_, _09836_, word_in[29]);
  or _18177_ (_14580_, _09913_, _09912_);
  and _18178_ (_09914_, _09829_, word_in[22]);
  not _18179_ (_09915_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  nor _18180_ (_09916_, _09823_, _09915_);
  and _18181_ (_09917_, _09823_, _09795_);
  or _18182_ (_09918_, _09917_, _09916_);
  or _18183_ (_09919_, _09918_, _09820_);
  or _18184_ (_09920_, _09831_, word_in[14]);
  and _18185_ (_09921_, _09920_, _09830_);
  and _18186_ (_09922_, _09921_, _09919_);
  or _18187_ (_09923_, _09922_, _09914_);
  and _18188_ (_09924_, _09923_, _09841_);
  and _18189_ (_09925_, _09836_, word_in[30]);
  or _18190_ (_08873_, _09925_, _09924_);
  nor _18191_ (_09926_, _09823_, _08700_);
  and _18192_ (_09927_, _09823_, _09640_);
  or _18193_ (_09928_, _09927_, _09926_);
  or _18194_ (_09929_, _09928_, _09820_);
  or _18195_ (_09930_, _09831_, word_in[15]);
  and _18196_ (_09931_, _09930_, _09830_);
  and _18197_ (_09932_, _09931_, _09929_);
  and _18198_ (_09933_, _09829_, word_in[23]);
  or _18199_ (_09934_, _09933_, _09836_);
  or _18200_ (_09935_, _09934_, _09932_);
  or _18201_ (_09936_, _09841_, word_in[31]);
  and _18202_ (_08876_, _09936_, _09935_);
  and _18203_ (_09937_, _08855_, _09309_);
  and _18204_ (_09938_, _09937_, word_in[24]);
  and _18205_ (_09939_, _08863_, _08644_);
  and _18206_ (_09940_, _09939_, _08732_);
  not _18207_ (_09941_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  not _18208_ (_09942_, _08874_);
  nor _18209_ (_09943_, _09698_, _09942_);
  nor _18210_ (_09944_, _09943_, _09941_);
  and _18211_ (_09945_, _09943_, _09703_);
  or _18212_ (_09946_, _09945_, _09944_);
  and _18213_ (_09947_, _08870_, _08626_);
  or _18214_ (_09948_, _09947_, _09946_);
  not _18215_ (_09950_, _09947_);
  or _18216_ (_09951_, _09950_, word_in[8]);
  and _18217_ (_09952_, _09951_, _09948_);
  or _18218_ (_09953_, _09952_, _09940_);
  not _18219_ (_09954_, _09937_);
  not _18220_ (_09956_, _09940_);
  or _18221_ (_09957_, _09956_, word_in[16]);
  and _18222_ (_09959_, _09957_, _09954_);
  and _18223_ (_09961_, _09959_, _09953_);
  or _18224_ (_14581_, _09961_, _09938_);
  not _18225_ (_09963_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  nor _18226_ (_09965_, _09943_, _09963_);
  and _18227_ (_09966_, _09943_, _09722_);
  or _18228_ (_09968_, _09966_, _09965_);
  or _18229_ (_09970_, _09968_, _09947_);
  or _18230_ (_09971_, _09950_, word_in[9]);
  and _18231_ (_09973_, _09971_, _09970_);
  or _18232_ (_09975_, _09973_, _09940_);
  or _18233_ (_09977_, _09956_, word_in[17]);
  and _18234_ (_09978_, _09977_, _09954_);
  and _18235_ (_09980_, _09978_, _09975_);
  and _18236_ (_09982_, _09937_, word_in[25]);
  or _18237_ (_08943_, _09982_, _09980_);
  and _18238_ (_09984_, _09937_, word_in[26]);
  not _18239_ (_09985_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  nor _18240_ (_09986_, _09943_, _09985_);
  and _18241_ (_09987_, _09943_, _09736_);
  or _18242_ (_09988_, _09987_, _09986_);
  or _18243_ (_09989_, _09988_, _09947_);
  or _18244_ (_09990_, _09950_, word_in[10]);
  and _18245_ (_09991_, _09990_, _09989_);
  or _18246_ (_09992_, _09991_, _09940_);
  or _18247_ (_09993_, _09956_, word_in[18]);
  and _18248_ (_09994_, _09993_, _09954_);
  and _18249_ (_09995_, _09994_, _09992_);
  or _18250_ (_08945_, _09995_, _09984_);
  and _18251_ (_09997_, _09937_, word_in[27]);
  not _18252_ (_09998_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  nor _18253_ (_09999_, _09943_, _09998_);
  and _18254_ (_10000_, _09943_, _09751_);
  or _18255_ (_10001_, _10000_, _09999_);
  or _18256_ (_10002_, _10001_, _09947_);
  or _18257_ (_10003_, _09950_, word_in[11]);
  and _18258_ (_10004_, _10003_, _10002_);
  or _18259_ (_10005_, _10004_, _09940_);
  or _18260_ (_10006_, _09956_, word_in[19]);
  and _18261_ (_10007_, _10006_, _09954_);
  and _18262_ (_10008_, _10007_, _10005_);
  or _18263_ (_08948_, _10008_, _09997_);
  and _18264_ (_10010_, _09943_, _09763_);
  not _18265_ (_10011_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  nor _18266_ (_10013_, _09943_, _10011_);
  nor _18267_ (_10014_, _10013_, _10010_);
  nor _18268_ (_10015_, _10014_, _09947_);
  and _18269_ (_10016_, _09947_, word_in[12]);
  or _18270_ (_10018_, _10016_, _10015_);
  and _18271_ (_10019_, _10018_, _09956_);
  and _18272_ (_10020_, _08863_, word_in[20]);
  and _18273_ (_10021_, _09940_, _10020_);
  or _18274_ (_10022_, _10021_, _09937_);
  or _18275_ (_10023_, _10022_, _10019_);
  or _18276_ (_10024_, _09954_, word_in[28]);
  and _18277_ (_08951_, _10024_, _10023_);
  and _18278_ (_10026_, _09937_, word_in[29]);
  not _18279_ (_10027_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  nor _18280_ (_10028_, _09943_, _10027_);
  and _18281_ (_10030_, _09943_, _09777_);
  or _18282_ (_10031_, _10030_, _10028_);
  or _18283_ (_10032_, _10031_, _09947_);
  or _18284_ (_10033_, _09950_, word_in[13]);
  and _18285_ (_10034_, _10033_, _10032_);
  or _18286_ (_10035_, _10034_, _09940_);
  or _18287_ (_10036_, _09956_, word_in[21]);
  and _18288_ (_10038_, _10036_, _09954_);
  and _18289_ (_10039_, _10038_, _10035_);
  or _18290_ (_08954_, _10039_, _10026_);
  and _18291_ (_10041_, _09937_, word_in[30]);
  not _18292_ (_10042_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  nor _18293_ (_10043_, _09943_, _10042_);
  and _18294_ (_10044_, _09943_, _09795_);
  or _18295_ (_10045_, _10044_, _10043_);
  or _18296_ (_10046_, _10045_, _09947_);
  or _18297_ (_10047_, _09950_, word_in[14]);
  and _18298_ (_10048_, _10047_, _10046_);
  or _18299_ (_10049_, _10048_, _09940_);
  or _18300_ (_10050_, _09956_, word_in[22]);
  and _18301_ (_10051_, _10050_, _09954_);
  and _18302_ (_10052_, _10051_, _10049_);
  or _18303_ (_08957_, _10052_, _10041_);
  nor _18304_ (_10054_, _09943_, _08584_);
  and _18305_ (_10055_, _09943_, _09640_);
  or _18306_ (_10056_, _10055_, _10054_);
  or _18307_ (_10057_, _10056_, _09947_);
  or _18308_ (_10058_, _09950_, word_in[15]);
  and _18309_ (_10059_, _10058_, _10057_);
  or _18310_ (_10060_, _10059_, _09940_);
  or _18311_ (_10061_, _09956_, word_in[23]);
  and _18312_ (_10062_, _10061_, _09954_);
  and _18313_ (_10063_, _10062_, _10060_);
  and _18314_ (_10064_, _09937_, word_in[31]);
  or _18315_ (_08960_, _10064_, _10063_);
  and _18316_ (_10065_, _08865_, _08770_);
  and _18317_ (_10066_, _10065_, _08655_);
  and _18318_ (_10067_, _08869_, _08930_);
  not _18319_ (_10068_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  nor _18320_ (_10069_, _09531_, _08872_);
  and _18321_ (_10070_, _08875_, _08904_);
  and _18322_ (_10071_, _10070_, _10069_);
  nor _18323_ (_10072_, _10071_, _10068_);
  and _18324_ (_10073_, _10071_, word_in[0]);
  or _18325_ (_10074_, _10073_, _10072_);
  or _18326_ (_10075_, _10074_, _10067_);
  not _18327_ (_10076_, _10067_);
  or _18328_ (_10077_, _10076_, word_in[8]);
  and _18329_ (_10078_, _10077_, _10075_);
  or _18330_ (_10079_, _10078_, _10066_);
  and _18331_ (_10080_, _08855_, _08897_);
  not _18332_ (_10081_, _10080_);
  not _18333_ (_10082_, _10066_);
  or _18334_ (_10083_, _10082_, _09837_);
  and _18335_ (_10084_, _10083_, _10081_);
  and _18336_ (_10085_, _10084_, _10079_);
  and _18337_ (_10086_, _10080_, word_in[24]);
  or _18338_ (_09044_, _10086_, _10085_);
  not _18339_ (_10087_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  nor _18340_ (_10088_, _10071_, _10087_);
  and _18341_ (_10089_, _10071_, word_in[1]);
  or _18342_ (_10090_, _10089_, _10088_);
  or _18343_ (_10091_, _10090_, _10067_);
  or _18344_ (_10092_, _10076_, word_in[9]);
  and _18345_ (_10093_, _10092_, _10091_);
  or _18346_ (_10094_, _10093_, _10066_);
  or _18347_ (_10095_, _10082_, _09565_);
  and _18348_ (_10096_, _10095_, _10081_);
  and _18349_ (_10097_, _10096_, _10094_);
  and _18350_ (_10098_, _10080_, word_in[25]);
  or _18351_ (_09047_, _10098_, _10097_);
  and _18352_ (_10099_, _08863_, word_in[18]);
  and _18353_ (_10100_, _10066_, _10099_);
  not _18354_ (_10101_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  nor _18355_ (_10102_, _10071_, _10101_);
  and _18356_ (_10103_, _10071_, word_in[2]);
  or _18357_ (_10104_, _10103_, _10102_);
  and _18358_ (_10105_, _10104_, _10076_);
  and _18359_ (_10106_, _10067_, word_in[10]);
  or _18360_ (_10107_, _10106_, _10105_);
  and _18361_ (_10108_, _10107_, _10082_);
  or _18362_ (_10109_, _10108_, _10100_);
  and _18363_ (_10110_, _10109_, _10081_);
  and _18364_ (_10111_, _10080_, word_in[26]);
  or _18365_ (_14582_, _10111_, _10110_);
  and _18366_ (_10112_, _07159_, _06439_);
  nand _18367_ (_10113_, _10112_, _06666_);
  or _18368_ (_10114_, _10112_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  and _18369_ (_10115_, _10114_, _06444_);
  and _18370_ (_09050_, _10115_, _10113_);
  and _18371_ (_10116_, _08863_, word_in[19]);
  and _18372_ (_10117_, _10066_, _10116_);
  not _18373_ (_10118_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  nor _18374_ (_10119_, _10071_, _10118_);
  and _18375_ (_10120_, _10071_, word_in[3]);
  or _18376_ (_10121_, _10120_, _10119_);
  and _18377_ (_10122_, _10121_, _10076_);
  and _18378_ (_10123_, _10067_, word_in[11]);
  or _18379_ (_10124_, _10123_, _10122_);
  and _18380_ (_10125_, _10124_, _10082_);
  or _18381_ (_10126_, _10125_, _10117_);
  and _18382_ (_10127_, _10126_, _10081_);
  and _18383_ (_10128_, _10080_, word_in[27]);
  or _18384_ (_14583_, _10128_, _10127_);
  not _18385_ (_10129_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  nor _18386_ (_10130_, _10071_, _10129_);
  and _18387_ (_10131_, _10071_, word_in[4]);
  or _18388_ (_10132_, _10131_, _10130_);
  or _18389_ (_10133_, _10132_, _10067_);
  or _18390_ (_10134_, _10076_, word_in[12]);
  and _18391_ (_10135_, _10134_, _10133_);
  or _18392_ (_10136_, _10135_, _10066_);
  or _18393_ (_10137_, _10082_, _10020_);
  and _18394_ (_10138_, _10137_, _10081_);
  and _18395_ (_10139_, _10138_, _10136_);
  and _18396_ (_10140_, _10080_, word_in[28]);
  or _18397_ (_14584_, _10140_, _10139_);
  not _18398_ (_10141_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  nor _18399_ (_10142_, _10071_, _10141_);
  and _18400_ (_10143_, _10071_, word_in[5]);
  or _18401_ (_10144_, _10143_, _10142_);
  or _18402_ (_10145_, _10144_, _10067_);
  or _18403_ (_10146_, _10076_, word_in[13]);
  and _18404_ (_10147_, _10146_, _10145_);
  or _18405_ (_10148_, _10147_, _10066_);
  and _18406_ (_10149_, _08863_, word_in[21]);
  or _18407_ (_10150_, _10082_, _10149_);
  and _18408_ (_10151_, _10150_, _10081_);
  and _18409_ (_10152_, _10151_, _10148_);
  and _18410_ (_10153_, _10080_, word_in[29]);
  or _18411_ (_14585_, _10153_, _10152_);
  and _18412_ (_10154_, _08863_, word_in[22]);
  and _18413_ (_10155_, _10066_, _10154_);
  not _18414_ (_10156_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  nor _18415_ (_10157_, _10071_, _10156_);
  and _18416_ (_10158_, _10071_, word_in[6]);
  or _18417_ (_10159_, _10158_, _10157_);
  and _18418_ (_10160_, _10159_, _10076_);
  and _18419_ (_10161_, _10067_, word_in[14]);
  or _18420_ (_10162_, _10161_, _10160_);
  and _18421_ (_10163_, _10162_, _10082_);
  or _18422_ (_10164_, _10163_, _10155_);
  and _18423_ (_10165_, _10164_, _10081_);
  and _18424_ (_10166_, _10080_, word_in[30]);
  or _18425_ (_09058_, _10166_, _10165_);
  nor _18426_ (_10167_, _10071_, _08709_);
  and _18427_ (_10168_, _10071_, word_in[7]);
  or _18428_ (_10169_, _10168_, _10167_);
  or _18429_ (_10170_, _10169_, _10067_);
  or _18430_ (_10171_, _10076_, word_in[15]);
  and _18431_ (_10172_, _10171_, _10170_);
  or _18432_ (_10173_, _10172_, _10066_);
  or _18433_ (_10174_, _10082_, _08886_);
  and _18434_ (_10175_, _10174_, _10081_);
  and _18435_ (_10176_, _10175_, _10173_);
  and _18436_ (_10177_, _10080_, word_in[31]);
  or _18437_ (_09061_, _10177_, _10176_);
  and _18438_ (_10178_, _10065_, _08613_);
  not _18439_ (_10179_, _10178_);
  and _18440_ (_10180_, _09695_, _08708_);
  and _18441_ (_10181_, _10070_, _09699_);
  and _18442_ (_10182_, _10181_, word_in[0]);
  not _18443_ (_10183_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  nor _18444_ (_10184_, _10181_, _10183_);
  nor _18445_ (_10185_, _10184_, _10182_);
  nor _18446_ (_10186_, _10185_, _10180_);
  and _18447_ (_10187_, _10180_, word_in[8]);
  or _18448_ (_10188_, _10187_, _10186_);
  and _18449_ (_10189_, _10188_, _10179_);
  and _18450_ (_10190_, _10178_, _09837_);
  or _18451_ (_10191_, _10190_, _10189_);
  and _18452_ (_10192_, _08855_, _08898_);
  not _18453_ (_10193_, _10192_);
  and _18454_ (_10194_, _10193_, _10191_);
  and _18455_ (_10195_, _10192_, word_in[24]);
  or _18456_ (_09148_, _10195_, _10194_);
  and _18457_ (_10196_, _10181_, word_in[1]);
  not _18458_ (_10197_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  nor _18459_ (_10198_, _10181_, _10197_);
  nor _18460_ (_10199_, _10198_, _10196_);
  nor _18461_ (_10200_, _10199_, _10180_);
  and _18462_ (_10201_, _10180_, word_in[9]);
  or _18463_ (_10202_, _10201_, _10200_);
  and _18464_ (_10203_, _10202_, _10179_);
  and _18465_ (_10204_, _10178_, _09565_);
  or _18466_ (_10205_, _10204_, _10203_);
  and _18467_ (_10206_, _10205_, _10193_);
  and _18468_ (_10207_, _10192_, word_in[25]);
  or _18469_ (_09150_, _10207_, _10206_);
  and _18470_ (_10208_, _10181_, word_in[2]);
  not _18471_ (_10209_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  nor _18472_ (_10210_, _10181_, _10209_);
  nor _18473_ (_10211_, _10210_, _10208_);
  nor _18474_ (_10212_, _10211_, _10180_);
  and _18475_ (_10213_, _10180_, word_in[10]);
  or _18476_ (_10214_, _10213_, _10212_);
  and _18477_ (_10215_, _10214_, _10179_);
  and _18478_ (_10216_, _10178_, _10099_);
  or _18479_ (_10217_, _10216_, _10215_);
  and _18480_ (_10218_, _10217_, _10193_);
  and _18481_ (_10219_, _10192_, word_in[26]);
  or _18482_ (_09153_, _10219_, _10218_);
  and _18483_ (_10220_, _10181_, word_in[3]);
  not _18484_ (_10221_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  nor _18485_ (_10222_, _10181_, _10221_);
  nor _18486_ (_10223_, _10222_, _10220_);
  nor _18487_ (_10224_, _10223_, _10180_);
  and _18488_ (_10225_, _10180_, word_in[11]);
  or _18489_ (_10226_, _10225_, _10224_);
  and _18490_ (_10227_, _10226_, _10179_);
  and _18491_ (_10228_, _10178_, _10116_);
  or _18492_ (_10229_, _10228_, _10227_);
  and _18493_ (_10230_, _10229_, _10193_);
  and _18494_ (_10231_, _10192_, word_in[27]);
  or _18495_ (_09156_, _10231_, _10230_);
  and _18496_ (_10232_, _10181_, word_in[4]);
  not _18497_ (_10233_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  nor _18498_ (_10234_, _10181_, _10233_);
  nor _18499_ (_10235_, _10234_, _10232_);
  nor _18500_ (_10236_, _10235_, _10180_);
  and _18501_ (_10237_, _10180_, word_in[12]);
  or _18502_ (_10238_, _10237_, _10236_);
  and _18503_ (_10239_, _10238_, _10179_);
  and _18504_ (_10240_, _10178_, _10020_);
  or _18505_ (_10241_, _10240_, _10239_);
  and _18506_ (_10242_, _10241_, _10193_);
  and _18507_ (_10243_, _10192_, word_in[28]);
  or _18508_ (_09159_, _10243_, _10242_);
  and _18509_ (_10244_, _10181_, word_in[5]);
  not _18510_ (_10245_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  nor _18511_ (_10246_, _10181_, _10245_);
  nor _18512_ (_10247_, _10246_, _10244_);
  nor _18513_ (_10248_, _10247_, _10180_);
  and _18514_ (_10249_, _10180_, word_in[13]);
  or _18515_ (_10250_, _10249_, _10248_);
  and _18516_ (_10251_, _10250_, _10179_);
  and _18517_ (_10252_, _10178_, _10149_);
  or _18518_ (_10253_, _10252_, _10251_);
  and _18519_ (_10254_, _10253_, _10193_);
  and _18520_ (_10255_, _10192_, word_in[29]);
  or _18521_ (_09162_, _10255_, _10254_);
  and _18522_ (_10256_, _10178_, _10154_);
  and _18523_ (_10257_, _10181_, word_in[6]);
  not _18524_ (_10258_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  nor _18525_ (_10259_, _10181_, _10258_);
  nor _18526_ (_10260_, _10259_, _10257_);
  nor _18527_ (_10261_, _10260_, _10180_);
  and _18528_ (_10262_, _10180_, word_in[14]);
  or _18529_ (_10263_, _10262_, _10261_);
  and _18530_ (_10264_, _10263_, _10179_);
  or _18531_ (_10265_, _10264_, _10256_);
  and _18532_ (_10266_, _10265_, _10193_);
  and _18533_ (_10267_, _10192_, word_in[30]);
  or _18534_ (_09166_, _10267_, _10266_);
  and _18535_ (_10268_, _10181_, word_in[7]);
  nor _18536_ (_10269_, _10181_, _08595_);
  nor _18537_ (_10270_, _10269_, _10268_);
  nor _18538_ (_10271_, _10270_, _10180_);
  and _18539_ (_10272_, _10180_, word_in[15]);
  or _18540_ (_10273_, _10272_, _10271_);
  and _18541_ (_10274_, _10273_, _10179_);
  and _18542_ (_10275_, _10178_, _08886_);
  or _18543_ (_10276_, _10275_, _10274_);
  and _18544_ (_10277_, _10276_, _10193_);
  and _18545_ (_10278_, _10192_, word_in[31]);
  or _18546_ (_09170_, _10278_, _10277_);
  nand _18547_ (_10279_, _10112_, _07300_);
  or _18548_ (_10280_, _10112_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  and _18549_ (_10281_, _10280_, _06444_);
  and _18550_ (_09234_, _10281_, _10279_);
  and _18551_ (_10282_, _08855_, _08930_);
  not _18552_ (_10283_, _10282_);
  and _18553_ (_10284_, _10065_, _08611_);
  and _18554_ (_10285_, _10284_, _09837_);
  not _18555_ (_10286_, _10284_);
  and _18556_ (_10287_, _09819_, _08708_);
  and _18557_ (_10288_, _09822_, _08904_);
  and _18558_ (_10289_, _10288_, word_in[0]);
  not _18559_ (_10290_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  nor _18560_ (_10291_, _10288_, _10290_);
  nor _18561_ (_10292_, _10291_, _10289_);
  nor _18562_ (_10293_, _10292_, _10287_);
  and _18563_ (_10294_, _10287_, word_in[8]);
  or _18564_ (_10295_, _10294_, _10293_);
  and _18565_ (_10296_, _10295_, _10286_);
  or _18566_ (_10297_, _10296_, _10285_);
  and _18567_ (_10298_, _10297_, _10283_);
  and _18568_ (_10299_, _10282_, word_in[24]);
  or _18569_ (_09240_, _10299_, _10298_);
  and _18570_ (_10300_, _10284_, _09565_);
  not _18571_ (_10301_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  nor _18572_ (_10302_, _10288_, _10301_);
  and _18573_ (_10303_, _10288_, word_in[1]);
  nor _18574_ (_10304_, _10303_, _10302_);
  nor _18575_ (_10305_, _10304_, _10287_);
  and _18576_ (_10306_, _10287_, word_in[9]);
  or _18577_ (_10307_, _10306_, _10305_);
  and _18578_ (_10308_, _10307_, _10286_);
  or _18579_ (_10309_, _10308_, _10300_);
  and _18580_ (_10310_, _10309_, _10283_);
  and _18581_ (_10311_, _10282_, word_in[25]);
  or _18582_ (_09245_, _10311_, _10310_);
  and _18583_ (_10312_, _10284_, _10099_);
  not _18584_ (_10313_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  nor _18585_ (_10314_, _10288_, _10313_);
  and _18586_ (_10315_, _10288_, word_in[2]);
  nor _18587_ (_10316_, _10315_, _10314_);
  nor _18588_ (_10317_, _10316_, _10287_);
  and _18589_ (_10318_, _10287_, word_in[10]);
  or _18590_ (_10319_, _10318_, _10317_);
  and _18591_ (_10320_, _10319_, _10286_);
  or _18592_ (_10321_, _10320_, _10312_);
  and _18593_ (_10322_, _10321_, _10283_);
  and _18594_ (_10323_, _10282_, word_in[26]);
  or _18595_ (_09248_, _10323_, _10322_);
  and _18596_ (_10324_, _10284_, _10116_);
  not _18597_ (_10325_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  nor _18598_ (_10326_, _10288_, _10325_);
  and _18599_ (_10327_, _10288_, word_in[3]);
  nor _18600_ (_10328_, _10327_, _10326_);
  nor _18601_ (_10329_, _10328_, _10287_);
  and _18602_ (_10330_, _10287_, word_in[11]);
  or _18603_ (_10331_, _10330_, _10329_);
  and _18604_ (_10332_, _10331_, _10286_);
  or _18605_ (_10333_, _10332_, _10324_);
  and _18606_ (_10334_, _10333_, _10283_);
  and _18607_ (_10335_, _10282_, word_in[27]);
  or _18608_ (_09253_, _10335_, _10334_);
  and _18609_ (_10336_, _10284_, _10020_);
  not _18610_ (_10337_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  nor _18611_ (_10338_, _10288_, _10337_);
  and _18612_ (_10339_, _10288_, word_in[4]);
  nor _18613_ (_10340_, _10339_, _10338_);
  nor _18614_ (_10341_, _10340_, _10287_);
  and _18615_ (_10342_, _10287_, word_in[12]);
  or _18616_ (_10343_, _10342_, _10341_);
  and _18617_ (_10344_, _10343_, _10286_);
  or _18618_ (_10346_, _10344_, _10336_);
  and _18619_ (_10347_, _10346_, _10283_);
  and _18620_ (_10348_, _10282_, word_in[28]);
  or _18621_ (_09258_, _10348_, _10347_);
  and _18622_ (_10349_, _10284_, _10149_);
  not _18623_ (_10350_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  nor _18624_ (_10351_, _10288_, _10350_);
  and _18625_ (_10352_, _10288_, word_in[5]);
  nor _18626_ (_10353_, _10352_, _10351_);
  nor _18627_ (_10355_, _10353_, _10287_);
  and _18628_ (_10356_, _10287_, word_in[13]);
  or _18629_ (_10358_, _10356_, _10355_);
  and _18630_ (_10359_, _10358_, _10286_);
  or _18631_ (_10360_, _10359_, _10349_);
  and _18632_ (_10361_, _10360_, _10283_);
  and _18633_ (_10363_, _10282_, word_in[29]);
  or _18634_ (_09261_, _10363_, _10361_);
  and _18635_ (_10365_, _10284_, _10154_);
  not _18636_ (_10366_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  nor _18637_ (_10367_, _10288_, _10366_);
  and _18638_ (_10368_, _10288_, word_in[6]);
  nor _18639_ (_10369_, _10368_, _10367_);
  nor _18640_ (_10370_, _10369_, _10287_);
  and _18641_ (_10371_, _10287_, word_in[14]);
  or _18642_ (_10372_, _10371_, _10370_);
  and _18643_ (_10373_, _10372_, _10286_);
  or _18644_ (_10374_, _10373_, _10365_);
  and _18645_ (_10375_, _10374_, _10283_);
  and _18646_ (_10376_, _10282_, word_in[30]);
  or _18647_ (_09265_, _10376_, _10375_);
  and _18648_ (_10377_, _10284_, _08886_);
  nor _18649_ (_10378_, _10288_, _08714_);
  and _18650_ (_10379_, _10288_, word_in[7]);
  nor _18651_ (_10380_, _10379_, _10378_);
  nor _18652_ (_10381_, _10380_, _10287_);
  and _18653_ (_10382_, _10287_, word_in[15]);
  or _18654_ (_10383_, _10382_, _10381_);
  and _18655_ (_10384_, _10383_, _10286_);
  or _18656_ (_10385_, _10384_, _10377_);
  and _18657_ (_10386_, _10385_, _10283_);
  and _18658_ (_10387_, _10282_, word_in[31]);
  or _18659_ (_09270_, _10387_, _10386_);
  and _18660_ (_10388_, _08855_, _08905_);
  not _18661_ (_10389_, _10388_);
  and _18662_ (_10390_, _10065_, _08644_);
  and _18663_ (_10391_, _10390_, _09837_);
  not _18664_ (_10392_, _10390_);
  and _18665_ (_10393_, _08870_, _08708_);
  and _18666_ (_10394_, _10070_, _08874_);
  and _18667_ (_10395_, _10394_, word_in[0]);
  not _18668_ (_10396_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  nor _18669_ (_10397_, _10394_, _10396_);
  nor _18670_ (_10398_, _10397_, _10395_);
  nor _18671_ (_10399_, _10398_, _10393_);
  and _18672_ (_10400_, _10393_, word_in[8]);
  or _18673_ (_10401_, _10400_, _10399_);
  and _18674_ (_10402_, _10401_, _10392_);
  or _18675_ (_10403_, _10402_, _10391_);
  and _18676_ (_10404_, _10403_, _10389_);
  and _18677_ (_10405_, _10388_, word_in[24]);
  or _18678_ (_14586_, _10405_, _10404_);
  not _18679_ (_10406_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  nor _18680_ (_10407_, _10394_, _10406_);
  and _18681_ (_10408_, _10394_, word_in[1]);
  nor _18682_ (_10409_, _10408_, _10407_);
  nor _18683_ (_10410_, _10409_, _10393_);
  and _18684_ (_10411_, _10393_, word_in[9]);
  or _18685_ (_10412_, _10411_, _10410_);
  and _18686_ (_10413_, _10412_, _10392_);
  and _18687_ (_10414_, _10390_, _09565_);
  or _18688_ (_10415_, _10414_, _10413_);
  and _18689_ (_10416_, _10415_, _10389_);
  and _18690_ (_10417_, _10388_, word_in[25]);
  or _18691_ (_14587_, _10417_, _10416_);
  and _18692_ (_10418_, _10390_, _10099_);
  and _18693_ (_10419_, _10394_, word_in[2]);
  not _18694_ (_10420_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  nor _18695_ (_10421_, _10394_, _10420_);
  nor _18696_ (_10422_, _10421_, _10419_);
  nor _18697_ (_10423_, _10422_, _10393_);
  and _18698_ (_10424_, _10393_, word_in[10]);
  or _18699_ (_10425_, _10424_, _10423_);
  and _18700_ (_10426_, _10425_, _10392_);
  or _18701_ (_10427_, _10426_, _10418_);
  and _18702_ (_10428_, _10427_, _10389_);
  and _18703_ (_10429_, _10388_, word_in[26]);
  or _18704_ (_14588_, _10429_, _10428_);
  and _18705_ (_10430_, _10394_, word_in[3]);
  not _18706_ (_10431_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  nor _18707_ (_10432_, _10394_, _10431_);
  nor _18708_ (_10433_, _10432_, _10430_);
  nor _18709_ (_10434_, _10433_, _10393_);
  and _18710_ (_10435_, _10393_, word_in[11]);
  or _18711_ (_10436_, _10435_, _10434_);
  and _18712_ (_10437_, _10436_, _10392_);
  and _18713_ (_10438_, _10390_, _10116_);
  or _18714_ (_10439_, _10438_, _10437_);
  and _18715_ (_10440_, _10439_, _10389_);
  and _18716_ (_10441_, _10388_, word_in[27]);
  or _18717_ (_14589_, _10441_, _10440_);
  and _18718_ (_10442_, _10394_, word_in[4]);
  not _18719_ (_10443_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  nor _18720_ (_10444_, _10394_, _10443_);
  nor _18721_ (_10445_, _10444_, _10442_);
  nor _18722_ (_10446_, _10445_, _10393_);
  and _18723_ (_10447_, _10393_, word_in[12]);
  or _18724_ (_10448_, _10447_, _10446_);
  and _18725_ (_10449_, _10448_, _10392_);
  and _18726_ (_10450_, _10390_, _10020_);
  or _18727_ (_10451_, _10450_, _10449_);
  and _18728_ (_10452_, _10451_, _10389_);
  and _18729_ (_10453_, _10388_, word_in[28]);
  or _18730_ (_14590_, _10453_, _10452_);
  not _18731_ (_10454_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  nor _18732_ (_10455_, _10394_, _10454_);
  and _18733_ (_10456_, _10394_, word_in[5]);
  or _18734_ (_10457_, _10456_, _10455_);
  or _18735_ (_10458_, _10457_, _10393_);
  not _18736_ (_10459_, _10393_);
  or _18737_ (_10460_, _10459_, word_in[13]);
  and _18738_ (_10461_, _10460_, _10458_);
  or _18739_ (_10462_, _10461_, _10390_);
  or _18740_ (_10463_, _10392_, _10149_);
  and _18741_ (_10464_, _10463_, _10462_);
  and _18742_ (_10465_, _10464_, _10389_);
  and _18743_ (_10466_, _10388_, word_in[29]);
  or _18744_ (_14591_, _10466_, _10465_);
  and _18745_ (_10467_, _10394_, word_in[6]);
  not _18746_ (_10469_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  nor _18747_ (_10470_, _10394_, _10469_);
  nor _18748_ (_10471_, _10470_, _10467_);
  nor _18749_ (_10472_, _10471_, _10393_);
  and _18750_ (_10473_, _10393_, word_in[14]);
  or _18751_ (_10474_, _10473_, _10472_);
  and _18752_ (_10475_, _10474_, _10392_);
  and _18753_ (_10476_, _10390_, _10154_);
  or _18754_ (_10477_, _10476_, _10475_);
  and _18755_ (_10478_, _10477_, _10389_);
  and _18756_ (_10479_, _10388_, word_in[30]);
  or _18757_ (_14592_, _10479_, _10478_);
  or _18758_ (_10480_, _10392_, _08886_);
  nor _18759_ (_10481_, _10394_, _08590_);
  and _18760_ (_10482_, _10394_, word_in[7]);
  or _18761_ (_10483_, _10482_, _10481_);
  or _18762_ (_10484_, _10483_, _10393_);
  or _18763_ (_10485_, _10459_, word_in[15]);
  and _18764_ (_10486_, _10485_, _10484_);
  or _18765_ (_10487_, _10486_, _10390_);
  and _18766_ (_10488_, _10487_, _10480_);
  or _18767_ (_10489_, _10488_, _10388_);
  or _18768_ (_10490_, _10389_, word_in[31]);
  and _18769_ (_14593_, _10490_, _10489_);
  nor _18770_ (_10491_, _06732_, _06644_);
  not _18771_ (_10492_, _10491_);
  and _18772_ (_10493_, _10492_, _09030_);
  and _18773_ (_10494_, _10493_, _09019_);
  nor _18774_ (_10495_, _10494_, _07190_);
  and _18775_ (_10496_, _07156_, _06439_);
  or _18776_ (_10497_, _10496_, _07161_);
  and _18777_ (_10498_, _10497_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  or _18778_ (_10499_, _10498_, _10495_);
  and _18779_ (_09410_, _10499_, _06444_);
  and _18780_ (_10500_, _08855_, _08800_);
  and _18781_ (_10501_, _10500_, _08644_);
  and _18782_ (_10502_, _08863_, _08952_);
  and _18783_ (_10503_, _08869_, _08620_);
  not _18784_ (_10504_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  and _18785_ (_10505_, _08875_, _08538_);
  and _18786_ (_10506_, _10505_, _10069_);
  nor _18787_ (_10507_, _10506_, _10504_);
  and _18788_ (_10508_, _10506_, word_in[0]);
  or _18789_ (_10509_, _10508_, _10507_);
  or _18790_ (_10510_, _10509_, _10503_);
  not _18791_ (_10511_, _10503_);
  or _18792_ (_10512_, _10511_, word_in[8]);
  and _18793_ (_10513_, _10512_, _10510_);
  or _18794_ (_10514_, _10513_, _10502_);
  not _18795_ (_10515_, _10502_);
  or _18796_ (_10516_, _10515_, word_in[16]);
  and _18797_ (_10517_, _10516_, _10514_);
  or _18798_ (_10518_, _10517_, _10501_);
  not _18799_ (_10519_, _10501_);
  or _18800_ (_10520_, _10519_, word_in[24]);
  and _18801_ (_09446_, _10520_, _10518_);
  and _18802_ (_10521_, _10502_, word_in[17]);
  not _18803_ (_10522_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  nor _18804_ (_10523_, _10506_, _10522_);
  and _18805_ (_10524_, _10506_, word_in[1]);
  or _18806_ (_10525_, _10524_, _10523_);
  and _18807_ (_10526_, _10525_, _10511_);
  and _18808_ (_10527_, _10503_, word_in[9]);
  or _18809_ (_10528_, _10527_, _10526_);
  and _18810_ (_10529_, _10528_, _10515_);
  or _18811_ (_10530_, _10529_, _10521_);
  and _18812_ (_10531_, _10530_, _10519_);
  and _18813_ (_10532_, _10501_, word_in[25]);
  or _18814_ (_09449_, _10532_, _10531_);
  and _18815_ (_10533_, _10502_, word_in[18]);
  not _18816_ (_10534_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  nor _18817_ (_10535_, _10506_, _10534_);
  and _18818_ (_10536_, _10506_, word_in[2]);
  or _18819_ (_10537_, _10536_, _10535_);
  and _18820_ (_10538_, _10537_, _10511_);
  and _18821_ (_10539_, _10503_, word_in[10]);
  or _18822_ (_10540_, _10539_, _10538_);
  and _18823_ (_10541_, _10540_, _10515_);
  or _18824_ (_10542_, _10541_, _10533_);
  and _18825_ (_10543_, _10542_, _10519_);
  and _18826_ (_10544_, _10501_, word_in[26]);
  or _18827_ (_14594_, _10544_, _10543_);
  and _18828_ (_10545_, _10502_, word_in[19]);
  not _18829_ (_10546_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  nor _18830_ (_10547_, _10506_, _10546_);
  and _18831_ (_10548_, _10506_, word_in[3]);
  or _18832_ (_10549_, _10548_, _10547_);
  and _18833_ (_10550_, _10549_, _10511_);
  and _18834_ (_10551_, _10503_, word_in[11]);
  or _18835_ (_10552_, _10551_, _10550_);
  and _18836_ (_10553_, _10552_, _10515_);
  or _18837_ (_10554_, _10553_, _10545_);
  and _18838_ (_10555_, _10554_, _10519_);
  and _18839_ (_10556_, _10501_, word_in[27]);
  or _18840_ (_14595_, _10556_, _10555_);
  and _18841_ (_10557_, _10502_, word_in[20]);
  not _18842_ (_10558_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  nor _18843_ (_10559_, _10506_, _10558_);
  and _18844_ (_10561_, _10506_, word_in[4]);
  or _18845_ (_10562_, _10561_, _10559_);
  and _18846_ (_10563_, _10562_, _10511_);
  and _18847_ (_10564_, _10503_, word_in[12]);
  or _18848_ (_10565_, _10564_, _10563_);
  and _18849_ (_10566_, _10565_, _10515_);
  or _18850_ (_10567_, _10566_, _10557_);
  and _18851_ (_10568_, _10567_, _10519_);
  and _18852_ (_10569_, _10501_, word_in[28]);
  or _18853_ (_14596_, _10569_, _10568_);
  and _18854_ (_10570_, _10502_, word_in[21]);
  not _18855_ (_10571_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  nor _18856_ (_10572_, _10506_, _10571_);
  and _18857_ (_10573_, _10506_, word_in[5]);
  or _18858_ (_10574_, _10573_, _10572_);
  and _18859_ (_10575_, _10574_, _10511_);
  and _18860_ (_10576_, _10503_, word_in[13]);
  or _18861_ (_10577_, _10576_, _10575_);
  and _18862_ (_10578_, _10577_, _10515_);
  or _18863_ (_10579_, _10578_, _10570_);
  and _18864_ (_10580_, _10579_, _10519_);
  and _18865_ (_10581_, _10501_, word_in[29]);
  or _18866_ (_14597_, _10581_, _10580_);
  and _18867_ (_10582_, _10502_, word_in[22]);
  not _18868_ (_10583_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  nor _18869_ (_10584_, _10506_, _10583_);
  and _18870_ (_10585_, _10506_, word_in[6]);
  or _18871_ (_10586_, _10585_, _10584_);
  and _18872_ (_10587_, _10586_, _10511_);
  and _18873_ (_10588_, _10503_, word_in[14]);
  or _18874_ (_10589_, _10588_, _10587_);
  and _18875_ (_10590_, _10589_, _10515_);
  or _18876_ (_10591_, _10590_, _10582_);
  and _18877_ (_10592_, _10591_, _10519_);
  and _18878_ (_10593_, _10501_, word_in[30]);
  or _18879_ (_14598_, _10593_, _10592_);
  and _18880_ (_10594_, _10502_, word_in[23]);
  nor _18881_ (_10595_, _10506_, _08672_);
  and _18882_ (_10596_, _10506_, word_in[7]);
  or _18883_ (_10597_, _10596_, _10595_);
  and _18884_ (_10598_, _10597_, _10511_);
  and _18885_ (_10599_, _10503_, word_in[15]);
  or _18886_ (_10600_, _10599_, _10598_);
  and _18887_ (_10601_, _10600_, _10515_);
  or _18888_ (_10602_, _10601_, _10594_);
  and _18889_ (_10603_, _10602_, _10519_);
  and _18890_ (_10604_, _10501_, word_in[31]);
  or _18891_ (_14599_, _10604_, _10603_);
  and _18892_ (_10605_, _10500_, _08655_);
  and _18893_ (_10606_, _09693_, _08734_);
  and _18894_ (_10607_, _09695_, _08623_);
  not _18895_ (_10608_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  and _18896_ (_10609_, _10505_, _09699_);
  nor _18897_ (_10610_, _10609_, _10608_);
  and _18898_ (_10611_, _10609_, word_in[0]);
  or _18899_ (_10612_, _10611_, _10610_);
  or _18900_ (_10613_, _10612_, _10607_);
  not _18901_ (_10614_, _10607_);
  or _18902_ (_10615_, _10614_, word_in[8]);
  and _18903_ (_10616_, _10615_, _10613_);
  or _18904_ (_10617_, _10616_, _10606_);
  not _18905_ (_10618_, _10606_);
  or _18906_ (_10619_, _10618_, _09837_);
  and _18907_ (_10620_, _10619_, _10617_);
  or _18908_ (_10621_, _10620_, _10605_);
  not _18909_ (_10622_, _10605_);
  or _18910_ (_10623_, _10622_, word_in[24]);
  and _18911_ (_14600_, _10623_, _10621_);
  not _18912_ (_10624_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  nor _18913_ (_10625_, _10609_, _10624_);
  and _18914_ (_10626_, _10609_, _09722_);
  or _18915_ (_10627_, _10626_, _10625_);
  or _18916_ (_10628_, _10627_, _10607_);
  or _18917_ (_10629_, _10614_, word_in[9]);
  and _18918_ (_10630_, _10629_, _10628_);
  or _18919_ (_10631_, _10630_, _10606_);
  or _18920_ (_10632_, _10618_, _09565_);
  and _18921_ (_10633_, _10632_, _10622_);
  and _18922_ (_10634_, _10633_, _10631_);
  and _18923_ (_10635_, _10605_, word_in[25]);
  or _18924_ (_14601_, _10635_, _10634_);
  not _18925_ (_10636_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  nor _18926_ (_10637_, _10609_, _10636_);
  and _18927_ (_10638_, _10609_, word_in[2]);
  or _18928_ (_10639_, _10638_, _10637_);
  or _18929_ (_10640_, _10639_, _10607_);
  or _18930_ (_10641_, _10614_, word_in[10]);
  and _18931_ (_10642_, _10641_, _10640_);
  or _18932_ (_10643_, _10642_, _10606_);
  or _18933_ (_10644_, _10618_, _10099_);
  and _18934_ (_10645_, _10644_, _10643_);
  or _18935_ (_10646_, _10645_, _10605_);
  or _18936_ (_10647_, _10622_, word_in[26]);
  and _18937_ (_14602_, _10647_, _10646_);
  or _18938_ (_10648_, _10618_, _10116_);
  not _18939_ (_10649_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  nor _18940_ (_10650_, _10609_, _10649_);
  and _18941_ (_10651_, _10609_, word_in[3]);
  or _18942_ (_10652_, _10651_, _10650_);
  or _18943_ (_10653_, _10652_, _10607_);
  or _18944_ (_10654_, _10614_, word_in[11]);
  and _18945_ (_10655_, _10654_, _10653_);
  or _18946_ (_10656_, _10655_, _10606_);
  and _18947_ (_10657_, _10656_, _10648_);
  or _18948_ (_10658_, _10657_, _10605_);
  or _18949_ (_10659_, _10622_, word_in[27]);
  and _18950_ (_14603_, _10659_, _10658_);
  not _18951_ (_10660_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  nor _18952_ (_10661_, _10609_, _10660_);
  and _18953_ (_10662_, _10609_, word_in[4]);
  or _18954_ (_10663_, _10662_, _10661_);
  or _18955_ (_10664_, _10663_, _10607_);
  or _18956_ (_10665_, _10614_, word_in[12]);
  and _18957_ (_10666_, _10665_, _10664_);
  or _18958_ (_10667_, _10666_, _10606_);
  or _18959_ (_10668_, _10618_, _10020_);
  and _18960_ (_10669_, _10668_, _10622_);
  and _18961_ (_10670_, _10669_, _10667_);
  and _18962_ (_10671_, _10605_, word_in[28]);
  or _18963_ (_14604_, _10671_, _10670_);
  not _18964_ (_10672_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  nor _18965_ (_10673_, _10609_, _10672_);
  and _18966_ (_10674_, _10609_, _09777_);
  or _18967_ (_10675_, _10674_, _10673_);
  or _18968_ (_10676_, _10675_, _10607_);
  or _18969_ (_10677_, _10614_, word_in[13]);
  and _18970_ (_10678_, _10677_, _10676_);
  or _18971_ (_10679_, _10678_, _10606_);
  or _18972_ (_10680_, _10618_, _10149_);
  and _18973_ (_10681_, _10680_, _10679_);
  or _18974_ (_10682_, _10681_, _10605_);
  or _18975_ (_10683_, _10622_, word_in[29]);
  and _18976_ (_14605_, _10683_, _10682_);
  or _18977_ (_10684_, _10618_, _10154_);
  not _18978_ (_10685_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  nor _18979_ (_10686_, _10609_, _10685_);
  and _18980_ (_10687_, _10609_, word_in[6]);
  or _18981_ (_10688_, _10687_, _10686_);
  or _18982_ (_10689_, _10688_, _10607_);
  or _18983_ (_10690_, _10614_, word_in[14]);
  and _18984_ (_10691_, _10690_, _10689_);
  or _18985_ (_10692_, _10691_, _10606_);
  and _18986_ (_10693_, _10692_, _10684_);
  or _18987_ (_10694_, _10693_, _10605_);
  or _18988_ (_10695_, _10622_, word_in[30]);
  and _18989_ (_14606_, _10695_, _10694_);
  nor _18990_ (_10696_, _10609_, _08576_);
  and _18991_ (_10697_, _10609_, word_in[7]);
  or _18992_ (_10698_, _10697_, _10696_);
  or _18993_ (_10699_, _10698_, _10607_);
  or _18994_ (_10700_, _10614_, word_in[15]);
  and _18995_ (_10701_, _10700_, _10699_);
  or _18996_ (_10702_, _10701_, _10606_);
  or _18997_ (_10703_, _10618_, _08886_);
  and _18998_ (_10704_, _10703_, _10702_);
  or _18999_ (_10705_, _10704_, _10605_);
  or _19000_ (_10706_, _10622_, word_in[31]);
  and _19001_ (_14607_, _10706_, _10705_);
  and _19002_ (_10707_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  not _19003_ (_10708_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  nor _19004_ (_10709_, _07432_, _10708_);
  or _19005_ (_10710_, _10709_, _10707_);
  and _19006_ (_09561_, _10710_, _06444_);
  and _19007_ (_10711_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  not _19008_ (_10712_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  nor _19009_ (_10713_, _07432_, _10712_);
  or _19010_ (_10714_, _10713_, _10711_);
  and _19011_ (_09566_, _10714_, _06444_);
  and _19012_ (_10715_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  not _19013_ (_10716_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor _19014_ (_10717_, _07432_, _10716_);
  or _19015_ (_10718_, _10717_, _10715_);
  and _19016_ (_09571_, _10718_, _06444_);
  nor _19017_ (_10719_, _07230_, _06734_);
  and _19018_ (_10720_, _07254_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and _19019_ (_10721_, _07238_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor _19020_ (_10722_, _10721_, _10720_);
  and _19021_ (_10723_, _07246_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and _19022_ (_10724_, _07251_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor _19023_ (_10725_, _10724_, _10723_);
  and _19024_ (_10726_, _07248_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  not _19025_ (_10728_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor _19026_ (_10729_, _07241_, _10728_);
  nor _19027_ (_10730_, _10729_, _10726_);
  and _19028_ (_10731_, _10730_, _10725_);
  and _19029_ (_10732_, _10731_, _10722_);
  nor _19030_ (_10733_, _10732_, _08374_);
  nor _19031_ (_10734_, _10733_, _10719_);
  nor _19032_ (_09590_, _10734_, rst);
  not _19033_ (_10735_, _08425_);
  and _19034_ (_10736_, _08472_, _08360_);
  and _19035_ (_10737_, _10736_, _08457_);
  not _19036_ (_10738_, _10737_);
  not _19037_ (_10739_, _08472_);
  and _19038_ (_10740_, _10739_, _08360_);
  not _19039_ (_10741_, _08457_);
  and _19040_ (_10742_, _10741_, _08441_);
  and _19041_ (_10743_, _10742_, _10740_);
  nor _19042_ (_10744_, _08472_, _08360_);
  and _19043_ (_10745_, _08457_, _08441_);
  and _19044_ (_10746_, _10745_, _10744_);
  nor _19045_ (_10747_, _10746_, _10743_);
  and _19046_ (_10748_, _10747_, _10738_);
  nor _19047_ (_10749_, _10748_, _10735_);
  not _19048_ (_10750_, _10749_);
  and _19049_ (_10751_, _08408_, _08392_);
  nor _19050_ (_10752_, _08425_, _07263_);
  and _19051_ (_10753_, _10752_, _10751_);
  not _19052_ (_10754_, _08392_);
  nor _19053_ (_10755_, _08425_, _08408_);
  and _19054_ (_10756_, _10755_, _10754_);
  nor _19055_ (_10757_, _10756_, _10753_);
  nor _19056_ (_10758_, _08457_, _08441_);
  and _19057_ (_10759_, _10758_, _10744_);
  and _19058_ (_10760_, _10754_, _07263_);
  and _19059_ (_10761_, _10760_, _10755_);
  and _19060_ (_10762_, _10745_, _10740_);
  and _19061_ (_10763_, _10762_, _10761_);
  nor _19062_ (_10764_, _10763_, _10759_);
  nor _19063_ (_10765_, _10764_, _10757_);
  not _19064_ (_10766_, _10765_);
  not _19065_ (_10767_, _08408_);
  nor _19066_ (_10768_, _08425_, _10767_);
  nor _19067_ (_10769_, _08392_, _07263_);
  and _19068_ (_10770_, _10769_, _10768_);
  nor _19069_ (_10771_, _10739_, _08360_);
  nor _19070_ (_10772_, _10758_, _10745_);
  and _19071_ (_10773_, _10772_, _10771_);
  and _19072_ (_10774_, _10773_, _10770_);
  and _19073_ (_10775_, _10761_, _10743_);
  nor _19074_ (_10776_, _10775_, _10774_);
  not _19075_ (_10777_, _10761_);
  and _19076_ (_10778_, _10758_, _10736_);
  nor _19077_ (_10779_, _10778_, _10746_);
  nor _19078_ (_10780_, _10779_, _10777_);
  and _19079_ (_10781_, _10745_, _10736_);
  and _19080_ (_10782_, _10769_, _10755_);
  and _19081_ (_10783_, _10782_, _10781_);
  and _19082_ (_10784_, _10771_, _10741_);
  and _19083_ (_10785_, _10784_, _10753_);
  nor _19084_ (_10786_, _10785_, _10783_);
  not _19085_ (_10787_, _10786_);
  nor _19086_ (_10788_, _10787_, _10780_);
  and _19087_ (_10789_, _10788_, _10776_);
  and _19088_ (_10790_, _10789_, _10766_);
  and _19089_ (_10791_, _10790_, _10750_);
  and _19090_ (_10792_, _10782_, _10746_);
  and _19091_ (_10793_, _10771_, _10761_);
  nor _19092_ (_10794_, _10793_, _10792_);
  and _19093_ (_10795_, _10767_, _08392_);
  nor _19094_ (_10796_, _08441_, _08425_);
  and _19095_ (_10797_, _10796_, _10795_);
  and _19096_ (_10798_, _10797_, _10736_);
  and _19097_ (_10799_, _10771_, _08457_);
  and _19098_ (_10800_, _10799_, _10782_);
  nor _19099_ (_10801_, _10800_, _10798_);
  and _19100_ (_10803_, _10801_, _10794_);
  and _19101_ (_10804_, _10770_, _10781_);
  not _19102_ (_10805_, _10778_);
  nor _19103_ (_10806_, _10753_, _08425_);
  nor _19104_ (_10807_, _10806_, _10805_);
  nor _19105_ (_10808_, _10807_, _10804_);
  and _19106_ (_10810_, _10808_, _10803_);
  not _19107_ (_10811_, _10756_);
  not _19108_ (_10812_, _08441_);
  and _19109_ (_10813_, _10744_, _08457_);
  and _19110_ (_10814_, _10813_, _10812_);
  and _19111_ (_10815_, _10742_, _10736_);
  nor _19112_ (_10816_, _10815_, _10814_);
  nor _19113_ (_10817_, _10816_, _10811_);
  and _19114_ (_10818_, _10744_, _10742_);
  and _19115_ (_10819_, _10818_, _10770_);
  and _19116_ (_10820_, _10771_, _10745_);
  and _19117_ (_10821_, _10820_, _10770_);
  nor _19118_ (_10822_, _10821_, _10819_);
  not _19119_ (_10823_, _10822_);
  nor _19120_ (_10824_, _10823_, _10817_);
  and _19121_ (_10825_, _10824_, _10810_);
  and _19122_ (_10826_, _10770_, _10759_);
  not _19123_ (_10827_, _10826_);
  and _19124_ (_10828_, _10768_, _10754_);
  not _19125_ (_10829_, _10828_);
  nor _19126_ (_10830_, _10778_, _07263_);
  nor _19127_ (_10831_, _10830_, _10829_);
  not _19128_ (_10832_, _10818_);
  nor _19129_ (_10833_, _10832_, _10757_);
  nor _19130_ (_10834_, _10833_, _10831_);
  and _19131_ (_10835_, _10834_, _10827_);
  and _19132_ (_10836_, _10740_, _08457_);
  and _19133_ (_10837_, _10836_, _10812_);
  and _19134_ (_10838_, _10837_, _10761_);
  and _19135_ (_10839_, _08441_, _10735_);
  and _19136_ (_10840_, _10839_, _10795_);
  nor _19137_ (_10841_, _10813_, _10737_);
  not _19138_ (_10842_, _10841_);
  and _19139_ (_10843_, _10842_, _10840_);
  nor _19140_ (_10844_, _10843_, _10838_);
  and _19141_ (_10845_, _10758_, _10740_);
  and _19142_ (_10846_, _10845_, _10761_);
  not _19143_ (_10847_, _10846_);
  and _19144_ (_10848_, _10761_, _10781_);
  and _19145_ (_10849_, _08392_, _07263_);
  and _19146_ (_10850_, _10849_, _10768_);
  and _19147_ (_10851_, _10850_, _10818_);
  nor _19148_ (_10852_, _10851_, _10848_);
  and _19149_ (_10853_, _10852_, _10847_);
  and _19150_ (_10854_, _10853_, _10844_);
  and _19151_ (_10855_, _10854_, _10835_);
  and _19152_ (_10856_, _10855_, _10825_);
  not _19153_ (_10857_, _10753_);
  and _19154_ (_10858_, _10737_, _10812_);
  not _19155_ (_10859_, _10858_);
  not _19156_ (_10860_, _10845_);
  nor _19157_ (_10861_, _10815_, _10781_);
  and _19158_ (_10862_, _10861_, _10860_);
  and _19159_ (_10863_, _10862_, _10859_);
  and _19160_ (_10864_, _10863_, _10747_);
  nor _19161_ (_10865_, _10864_, _10857_);
  and _19162_ (_10866_, _10850_, _10759_);
  and _19163_ (_10867_, _10815_, _10770_);
  nor _19164_ (_10868_, _10867_, _10866_);
  not _19165_ (_10869_, _10770_);
  and _19166_ (_10870_, _10740_, _10741_);
  nor _19167_ (_10871_, _10858_, _10870_);
  nor _19168_ (_10872_, _10871_, _10869_);
  not _19169_ (_10873_, _10813_);
  and _19170_ (_10874_, _10796_, _10751_);
  nor _19171_ (_10875_, _10874_, _10770_);
  nor _19172_ (_10876_, _10875_, _10873_);
  nor _19173_ (_10877_, _10876_, _10872_);
  and _19174_ (_10878_, _10877_, _10868_);
  not _19175_ (_10879_, _10878_);
  nor _19176_ (_10880_, _10879_, _10865_);
  and _19177_ (_10881_, _10880_, _10856_);
  and _19178_ (_10882_, _10881_, _10791_);
  or _19179_ (_10883_, _10795_, _08425_);
  and _19180_ (_10884_, _10883_, _10781_);
  or _19181_ (_10885_, _10884_, _10821_);
  nand _19182_ (_10886_, _10850_, _10814_);
  nand _19183_ (_10887_, _10886_, _10852_);
  nor _19184_ (_10888_, _10887_, _10885_);
  and _19185_ (_10889_, _10888_, _10868_);
  nand _19186_ (_10890_, _10889_, _10789_);
  or _19187_ (_10891_, _10890_, _10882_);
  and _19188_ (_10892_, _10891_, _07230_);
  nand _19189_ (_10893_, _10892_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor _19190_ (_10894_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , rst);
  or _19191_ (_10895_, _10892_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _19192_ (_10896_, _10895_, _10894_);
  and _19193_ (_09594_, _10896_, _10893_);
  not _19194_ (_10897_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and _19195_ (_10898_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and _19196_ (_10899_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  and _19197_ (_10900_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor _19198_ (_10901_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  nor _19199_ (_10902_, _10901_, _10899_);
  and _19200_ (_10903_, _10902_, _10900_);
  nor _19201_ (_10904_, _10903_, _10899_);
  not _19202_ (_10906_, _10904_);
  nor _19203_ (_10907_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor _19204_ (_10908_, _10907_, _10898_);
  and _19205_ (_10909_, _10908_, _10906_);
  nor _19206_ (_10910_, _10909_, _10898_);
  not _19207_ (_10911_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  not _19208_ (_10912_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor _19209_ (_10913_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3], \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and _19210_ (_10914_, _10913_, _10912_);
  and _19211_ (_10915_, _10914_, _10911_);
  and _19212_ (_10916_, _10915_, _10910_);
  nor _19213_ (_10917_, _10916_, _10897_);
  and _19214_ (_10918_, _10916_, _10897_);
  nor _19215_ (_10919_, _10918_, _10917_);
  not _19216_ (_10920_, _10919_);
  and _19217_ (_10921_, _10914_, _10910_);
  nor _19218_ (_10923_, _10921_, _10911_);
  nor _19219_ (_10924_, _10923_, _10916_);
  not _19220_ (_10925_, _10924_);
  and _19221_ (_10926_, _10913_, _10910_);
  nor _19222_ (_10927_, _10926_, _10912_);
  nor _19223_ (_10928_, _10927_, _10921_);
  not _19224_ (_10929_, _10928_);
  nor _19225_ (_10930_, _10910_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and _19226_ (_10931_, _10910_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  or _19227_ (_10932_, _10931_, _10930_);
  not _19228_ (_10933_, _10932_);
  not _19229_ (_10934_, _10882_);
  nor _19230_ (_10935_, _10902_, _10900_);
  nor _19231_ (_10936_, _10935_, _10903_);
  nand _19232_ (_10937_, _10936_, _10934_);
  nor _19233_ (_10938_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor _19234_ (_10939_, _10938_, _10900_);
  and _19235_ (_10940_, _10939_, _10891_);
  or _19236_ (_10941_, _10936_, _10934_);
  and _19237_ (_10942_, _10941_, _10937_);
  nand _19238_ (_10943_, _10942_, _10940_);
  nand _19239_ (_10944_, _10943_, _10937_);
  nor _19240_ (_10945_, _10908_, _10906_);
  nor _19241_ (_10946_, _10945_, _10909_);
  and _19242_ (_10947_, _10946_, _10944_);
  and _19243_ (_10948_, _10947_, _10933_);
  and _19244_ (_10949_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3], \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or _19245_ (_10950_, _10949_, _10913_);
  nand _19246_ (_10951_, _10950_, _10930_);
  or _19247_ (_10952_, _10950_, _10930_);
  and _19248_ (_10953_, _10952_, _10951_);
  and _19249_ (_10954_, _10953_, _10948_);
  and _19250_ (_10955_, _10954_, _10929_);
  and _19251_ (_10956_, _10955_, _10925_);
  and _19252_ (_10957_, _10956_, _10920_);
  not _19253_ (_10958_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor _19254_ (_10959_, _10918_, _10958_);
  and _19255_ (_10960_, _10915_, _10897_);
  and _19256_ (_10961_, _10960_, _10958_);
  and _19257_ (_10962_, _10961_, _10910_);
  or _19258_ (_10963_, _10962_, _10959_);
  nand _19259_ (_10964_, _10963_, _10957_);
  not _19260_ (_10965_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  nor _19261_ (_10966_, _10962_, _10965_);
  and _19262_ (_10967_, _10962_, _10965_);
  nor _19263_ (_10968_, _10967_, _10966_);
  and _19264_ (_10969_, _10968_, _10964_);
  nor _19265_ (_10970_, _10968_, _10964_);
  nor _19266_ (_10971_, _10970_, _10969_);
  or _19267_ (_10972_, _10971_, _08374_);
  or _19268_ (_10973_, _08373_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and _19269_ (_10974_, _10973_, _10894_);
  and _19270_ (_10975_, _10974_, _10972_);
  and _19271_ (_10976_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _06444_);
  and _19272_ (_10977_, _10976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  or _19273_ (_09598_, _10977_, _10975_);
  and _19274_ (_10978_, _07321_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  and _19275_ (_10979_, _07325_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  nor _19276_ (_10980_, _10979_, _10978_);
  and _19277_ (_10981_, _07333_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  and _19278_ (_10982_, _07327_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  nor _19279_ (_10983_, _10982_, _10981_);
  and _19280_ (_10984_, _10983_, _10980_);
  and _19281_ (_10985_, _07313_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  and _19282_ (_10986_, _07331_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  nor _19283_ (_10987_, _10986_, _10985_);
  and _19284_ (_10988_, _07309_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  and _19285_ (_10989_, _07318_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  nor _19286_ (_10990_, _10989_, _10988_);
  and _19287_ (_10991_, _10990_, _10987_);
  and _19288_ (_10992_, _10991_, _10984_);
  nor _19289_ (_10993_, _10992_, _07307_);
  and _19290_ (_10994_, _07307_, _07070_);
  nor _19291_ (_10995_, _10994_, _10993_);
  nor _19292_ (_09610_, _10995_, rst);
  and _19293_ (_10996_, _09828_, _08734_);
  and _19294_ (_10997_, _09819_, _08623_);
  not _19295_ (_10998_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and _19296_ (_10999_, _09822_, _08538_);
  nor _19297_ (_11000_, _10999_, _10998_);
  and _19298_ (_11001_, _10999_, word_in[0]);
  or _19299_ (_11002_, _11001_, _11000_);
  or _19300_ (_11003_, _11002_, _10997_);
  not _19301_ (_11004_, _10997_);
  or _19302_ (_11005_, _11004_, word_in[8]);
  and _19303_ (_11006_, _11005_, _11003_);
  or _19304_ (_11007_, _11006_, _10996_);
  and _19305_ (_11008_, _10500_, _08613_);
  not _19306_ (_11009_, _11008_);
  not _19307_ (_11010_, _10996_);
  or _19308_ (_11011_, _11010_, _09837_);
  and _19309_ (_11012_, _11011_, _11009_);
  and _19310_ (_11013_, _11012_, _11007_);
  and _19311_ (_11014_, _11008_, word_in[24]);
  or _19312_ (_14555_, _11014_, _11013_);
  or _19313_ (_11015_, _07432_, \oc8051_top_1.oc8051_rom1.data_o [23]);
  not _19314_ (_11016_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  nand _19315_ (_11017_, _07432_, _11016_);
  and _19316_ (_11018_, _11017_, _06444_);
  and _19317_ (_09619_, _11018_, _11015_);
  not _19318_ (_11019_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  nor _19319_ (_11020_, _10999_, _11019_);
  and _19320_ (_11021_, _10999_, word_in[1]);
  or _19321_ (_11022_, _11021_, _11020_);
  or _19322_ (_11023_, _11022_, _10997_);
  or _19323_ (_11024_, _11004_, word_in[9]);
  and _19324_ (_11025_, _11024_, _11023_);
  or _19325_ (_11026_, _11025_, _10996_);
  or _19326_ (_11027_, _11010_, _09565_);
  and _19327_ (_11028_, _11027_, _11009_);
  and _19328_ (_11029_, _11028_, _11026_);
  and _19329_ (_11030_, _11008_, word_in[25]);
  or _19330_ (_14556_, _11030_, _11029_);
  or _19331_ (_11031_, _11010_, _10099_);
  not _19332_ (_11032_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  nor _19333_ (_11033_, _10999_, _11032_);
  and _19334_ (_11034_, _10999_, word_in[2]);
  or _19335_ (_11035_, _11034_, _11033_);
  or _19336_ (_11036_, _11035_, _10997_);
  or _19337_ (_11037_, _11004_, word_in[10]);
  and _19338_ (_11038_, _11037_, _11036_);
  or _19339_ (_11039_, _11038_, _10996_);
  and _19340_ (_11040_, _11039_, _11031_);
  or _19341_ (_11041_, _11040_, _11008_);
  or _19342_ (_11042_, _11009_, word_in[26]);
  and _19343_ (_14557_, _11042_, _11041_);
  or _19344_ (_11043_, _07432_, \oc8051_top_1.oc8051_rom1.data_o [4]);
  not _19345_ (_11044_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nand _19346_ (_11045_, _07432_, _11044_);
  and _19347_ (_11046_, _11045_, _06444_);
  and _19348_ (_09624_, _11046_, _11043_);
  not _19349_ (_11047_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  nor _19350_ (_11048_, _10999_, _11047_);
  and _19351_ (_11049_, _10999_, word_in[3]);
  or _19352_ (_11050_, _11049_, _11048_);
  or _19353_ (_11051_, _11050_, _10997_);
  or _19354_ (_11052_, _11004_, word_in[11]);
  and _19355_ (_11053_, _11052_, _11051_);
  or _19356_ (_11054_, _11053_, _10996_);
  or _19357_ (_11055_, _11010_, _10116_);
  and _19358_ (_11056_, _11055_, _11009_);
  and _19359_ (_11057_, _11056_, _11054_);
  and _19360_ (_11058_, _11008_, word_in[27]);
  or _19361_ (_14558_, _11058_, _11057_);
  not _19362_ (_11059_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  nor _19363_ (_11060_, _10999_, _11059_);
  and _19364_ (_11061_, _10999_, word_in[4]);
  or _19365_ (_11062_, _11061_, _11060_);
  or _19366_ (_11063_, _11062_, _10997_);
  or _19367_ (_11064_, _11004_, word_in[12]);
  and _19368_ (_11065_, _11064_, _11063_);
  or _19369_ (_11066_, _11065_, _10996_);
  or _19370_ (_11067_, _11010_, _10020_);
  and _19371_ (_11068_, _11067_, _11066_);
  or _19372_ (_11069_, _11068_, _11008_);
  or _19373_ (_11070_, _11009_, word_in[28]);
  and _19374_ (_14559_, _11070_, _11069_);
  not _19375_ (_11071_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  nor _19376_ (_11072_, _10999_, _11071_);
  and _19377_ (_11073_, _10999_, word_in[5]);
  or _19378_ (_11074_, _11073_, _11072_);
  or _19379_ (_11075_, _11074_, _10997_);
  or _19380_ (_11076_, _11004_, word_in[13]);
  and _19381_ (_11077_, _11076_, _11075_);
  or _19382_ (_11078_, _11077_, _10996_);
  or _19383_ (_11079_, _11010_, _10149_);
  and _19384_ (_11080_, _11079_, _11078_);
  or _19385_ (_11081_, _11080_, _11008_);
  or _19386_ (_11082_, _11009_, word_in[29]);
  and _19387_ (_14560_, _11082_, _11081_);
  or _19388_ (_11083_, _11010_, _10154_);
  not _19389_ (_11084_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  nor _19390_ (_11085_, _10999_, _11084_);
  and _19391_ (_11086_, _10999_, word_in[6]);
  or _19392_ (_11087_, _11086_, _11085_);
  or _19393_ (_11088_, _11087_, _10997_);
  or _19394_ (_11089_, _11004_, word_in[14]);
  and _19395_ (_11090_, _11089_, _11088_);
  or _19396_ (_11091_, _11090_, _10996_);
  and _19397_ (_11092_, _11091_, _11083_);
  or _19398_ (_11093_, _11092_, _11008_);
  or _19399_ (_11094_, _11009_, word_in[30]);
  and _19400_ (_14561_, _11094_, _11093_);
  or _19401_ (_11095_, _07757_, _07669_);
  not _19402_ (_11096_, _07681_);
  and _19403_ (_11097_, _08985_, _11096_);
  nand _19404_ (_11098_, _11097_, _07684_);
  or _19405_ (_11099_, _11097_, _07684_);
  nand _19406_ (_11100_, _11099_, _11098_);
  nand _19407_ (_11101_, _11100_, _07757_);
  nand _19408_ (_11102_, _11101_, _11095_);
  nand _19409_ (_11103_, _11102_, _07459_);
  and _19410_ (_11104_, _07767_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  nand _19411_ (_11105_, _11104_, _08994_);
  or _19412_ (_11106_, _08994_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  nand _19413_ (_11107_, _11106_, _11105_);
  nand _19414_ (_11108_, _11107_, _07602_);
  nor _19415_ (_11109_, _08109_, _06887_);
  nor _19416_ (_11110_, _11109_, _06697_);
  and _19417_ (_11111_, _11109_, _06697_);
  nor _19418_ (_11112_, _11111_, _11110_);
  nor _19419_ (_11113_, _11112_, _06891_);
  nor _19420_ (_11114_, _06732_, _06638_);
  and _19421_ (_11115_, _06904_, _06465_);
  nor _19422_ (_11116_, _11115_, _11114_);
  and _19423_ (_11117_, _06914_, _06640_);
  and _19424_ (_11118_, _06918_, _06903_);
  nor _19425_ (_11119_, _11118_, _11117_);
  and _19426_ (_11120_, _11119_, _11116_);
  and _19427_ (_11121_, _11120_, _06974_);
  not _19428_ (_11122_, _11121_);
  nor _19429_ (_11123_, _11122_, _11113_);
  and _19430_ (_11124_, _11123_, _06967_);
  not _19431_ (_11125_, _06709_);
  and _19432_ (_11126_, _06842_, _11125_);
  nor _19433_ (_11127_, _06842_, _11125_);
  nor _19434_ (_11128_, _11127_, _11126_);
  and _19435_ (_11129_, _11128_, _06680_);
  nor _19436_ (_11130_, _06877_, _06709_);
  and _19437_ (_11131_, _06877_, _06709_);
  or _19438_ (_11132_, _11131_, _11130_);
  and _19439_ (_11133_, _11132_, _06847_);
  nor _19440_ (_11134_, _11133_, _11129_);
  and _19441_ (_11135_, _11134_, _11124_);
  and _19442_ (_11136_, _11135_, _11108_);
  nand _19443_ (_11137_, _11136_, _11103_);
  nand _19444_ (_11138_, _11137_, _07653_);
  nor _19445_ (_11139_, _06933_, _06701_);
  nor _19446_ (_11140_, _11139_, _06935_);
  nor _19447_ (_11142_, _11140_, _08028_);
  and _19448_ (_11143_, _08036_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or _19449_ (_11144_, _11143_, _07439_);
  nor _19450_ (_11145_, _11144_, _11142_);
  nand _19451_ (_11146_, _11145_, _11138_);
  and _19452_ (_11147_, _06705_, _06640_);
  and _19453_ (_11148_, _06913_, _06552_);
  nor _19454_ (_11149_, _06740_, _06465_);
  nor _19455_ (_11150_, _11149_, _09006_);
  and _19456_ (_11151_, _11150_, _09173_);
  and _19457_ (_11152_, _11151_, _06704_);
  nor _19458_ (_11153_, _11151_, _06704_);
  nor _19459_ (_11155_, _11153_, _11152_);
  nor _19460_ (_11156_, _11155_, _06621_);
  nor _19461_ (_11157_, _06704_, _06465_);
  or _19462_ (_11158_, _11157_, _06892_);
  and _19463_ (_11160_, _11158_, _06455_);
  or _19464_ (_11161_, _11160_, _11156_);
  or _19465_ (_11162_, _11161_, _11148_);
  and _19466_ (_11163_, _07459_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  nor _19467_ (_11164_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  not _19468_ (_11165_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and _19469_ (_11166_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _11165_);
  nor _19470_ (_11167_, _11166_, _11164_);
  nand _19471_ (_11168_, _11167_, _09191_);
  or _19472_ (_11169_, _11167_, _09191_);
  and _19473_ (_11170_, _11169_, _06847_);
  and _19474_ (_11171_, _11170_, _11168_);
  and _19475_ (_11172_, _09416_, _07602_);
  or _19476_ (_11173_, _11172_, _11171_);
  or _19477_ (_11174_, _11173_, _11163_);
  or _19478_ (_11175_, _11174_, _11162_);
  or _19479_ (_11177_, _11175_, _11147_);
  or _19480_ (_11178_, _11177_, _07961_);
  and _19481_ (_11179_, _11178_, _11146_);
  and _19482_ (_09630_, _11179_, _06444_);
  nor _19483_ (_11180_, _10999_, _08667_);
  and _19484_ (_11181_, _10999_, word_in[7]);
  or _19485_ (_11182_, _11181_, _11180_);
  or _19486_ (_11183_, _11182_, _10997_);
  or _19487_ (_11184_, _11004_, word_in[15]);
  and _19488_ (_11185_, _11184_, _11183_);
  or _19489_ (_11186_, _11185_, _10996_);
  or _19490_ (_11187_, _11010_, _08886_);
  and _19491_ (_11188_, _11187_, _11009_);
  and _19492_ (_11189_, _11188_, _11186_);
  and _19493_ (_11190_, _11008_, word_in[31]);
  or _19494_ (_14562_, _11190_, _11189_);
  and _19495_ (_11191_, _07429_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [2]);
  and _19496_ (_11192_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and _19497_ (_11193_, _07248_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  not _19498_ (_11194_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor _19499_ (_11195_, _07241_, _11194_);
  nor _19500_ (_11196_, _11195_, _11193_);
  and _19501_ (_11197_, _07246_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and _19502_ (_11199_, _07238_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor _19503_ (_11200_, _11199_, _11197_);
  and _19504_ (_11201_, _07251_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  and _19505_ (_11202_, _07254_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nor _19506_ (_11203_, _11202_, _11201_);
  and _19507_ (_11204_, _11203_, _11200_);
  and _19508_ (_11205_, _11204_, _11196_);
  nor _19509_ (_11206_, _11205_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _19510_ (_11207_, _11206_, _11192_);
  nor _19511_ (_11208_, _11207_, _07429_);
  nor _19512_ (_11209_, _11208_, _11191_);
  nor _19513_ (_09668_, _11209_, rst);
  nor _19514_ (_11210_, _07230_, _06790_);
  and _19515_ (_11211_, _07254_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and _19516_ (_11212_, _07238_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor _19517_ (_11213_, _11212_, _11211_);
  and _19518_ (_11215_, _07246_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and _19519_ (_11216_, _07251_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor _19520_ (_11217_, _11216_, _11215_);
  and _19521_ (_11218_, _07248_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  not _19522_ (_11220_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor _19523_ (_11221_, _07241_, _11220_);
  nor _19524_ (_11223_, _11221_, _11218_);
  and _19525_ (_11224_, _11223_, _11217_);
  and _19526_ (_11225_, _11224_, _11213_);
  nor _19527_ (_11226_, _11225_, _08374_);
  nor _19528_ (_11227_, _11226_, _11210_);
  nor _19529_ (_09673_, _11227_, rst);
  and _19530_ (_11228_, _09939_, _08734_);
  and _19531_ (_11229_, _08870_, _08623_);
  not _19532_ (_11230_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and _19533_ (_11231_, _10505_, _08874_);
  nor _19534_ (_11232_, _11231_, _11230_);
  and _19535_ (_11233_, _11231_, word_in[0]);
  or _19536_ (_11234_, _11233_, _11232_);
  or _19537_ (_11235_, _11234_, _11229_);
  not _19538_ (_11236_, _11229_);
  or _19539_ (_11237_, _11236_, word_in[8]);
  and _19540_ (_11238_, _11237_, _11235_);
  or _19541_ (_11240_, _11238_, _11228_);
  and _19542_ (_11241_, _10500_, _08611_);
  not _19543_ (_11242_, _11241_);
  not _19544_ (_11243_, _11228_);
  or _19545_ (_11244_, _11243_, _09837_);
  and _19546_ (_11245_, _11244_, _11242_);
  and _19547_ (_11246_, _11245_, _11240_);
  and _19548_ (_11247_, _11241_, _09554_);
  or _19549_ (_14563_, _11247_, _11246_);
  not _19550_ (_11249_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  nor _19551_ (_11250_, _11231_, _11249_);
  and _19552_ (_11251_, _11231_, _09722_);
  or _19553_ (_11253_, _11251_, _11250_);
  or _19554_ (_11254_, _11253_, _11229_);
  or _19555_ (_11255_, _11236_, word_in[9]);
  and _19556_ (_11256_, _11255_, _11254_);
  or _19557_ (_11257_, _11256_, _11228_);
  or _19558_ (_11258_, _11243_, _09565_);
  and _19559_ (_11259_, _11258_, _11242_);
  and _19560_ (_11260_, _11259_, _11257_);
  and _19561_ (_11261_, _08855_, word_in[25]);
  and _19562_ (_11262_, _11241_, _11261_);
  or _19563_ (_14564_, _11262_, _11260_);
  and _19564_ (_11263_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  not _19565_ (_11264_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  nor _19566_ (_11265_, _07432_, _11264_);
  or _19567_ (_11266_, _11265_, _11263_);
  and _19568_ (_09708_, _11266_, _06444_);
  not _19569_ (_11267_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  nor _19570_ (_11268_, _11231_, _11267_);
  and _19571_ (_11269_, _11231_, word_in[2]);
  or _19572_ (_11270_, _11269_, _11268_);
  or _19573_ (_11271_, _11270_, _11229_);
  or _19574_ (_11272_, _11236_, word_in[10]);
  and _19575_ (_11273_, _11272_, _11271_);
  or _19576_ (_11274_, _11273_, _11228_);
  or _19577_ (_11275_, _11243_, _10099_);
  and _19578_ (_11276_, _11275_, _11242_);
  and _19579_ (_11277_, _11276_, _11274_);
  and _19580_ (_11278_, _11241_, _09582_);
  or _19581_ (_14565_, _11278_, _11277_);
  not _19582_ (_11279_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  nor _19583_ (_11280_, _11231_, _11279_);
  and _19584_ (_11281_, _11231_, word_in[3]);
  or _19585_ (_11282_, _11281_, _11280_);
  or _19586_ (_11283_, _11282_, _11229_);
  or _19587_ (_11284_, _11236_, word_in[11]);
  and _19588_ (_11285_, _11284_, _11283_);
  or _19589_ (_11286_, _11285_, _11228_);
  or _19590_ (_11287_, _11243_, _10116_);
  and _19591_ (_11288_, _11287_, _11286_);
  or _19592_ (_11289_, _11288_, _11241_);
  or _19593_ (_11290_, _11242_, word_in[27]);
  and _19594_ (_14566_, _11290_, _11289_);
  and _19595_ (_11291_, _11228_, _10020_);
  not _19596_ (_11292_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  nor _19597_ (_11293_, _11231_, _11292_);
  and _19598_ (_11294_, _11231_, word_in[4]);
  nor _19599_ (_11295_, _11294_, _11293_);
  nor _19600_ (_11296_, _11295_, _11229_);
  and _19601_ (_11297_, _11229_, word_in[12]);
  or _19602_ (_11299_, _11297_, _11296_);
  and _19603_ (_11300_, _11299_, _11243_);
  or _19604_ (_11301_, _11300_, _11291_);
  and _19605_ (_11302_, _11301_, _11242_);
  and _19606_ (_11303_, _11241_, word_in[28]);
  or _19607_ (_14567_, _11303_, _11302_);
  not _19608_ (_11305_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  nor _19609_ (_11306_, _11231_, _11305_);
  and _19610_ (_11307_, _11231_, _09777_);
  or _19611_ (_11309_, _11307_, _11306_);
  or _19612_ (_11310_, _11309_, _11229_);
  or _19613_ (_11311_, _11236_, word_in[13]);
  and _19614_ (_11312_, _11311_, _11310_);
  or _19615_ (_11313_, _11312_, _11228_);
  or _19616_ (_11314_, _11243_, _10149_);
  and _19617_ (_11315_, _11314_, _11242_);
  and _19618_ (_11316_, _11315_, _11313_);
  and _19619_ (_11317_, _11241_, _09623_);
  or _19620_ (_14568_, _11317_, _11316_);
  not _19621_ (_11318_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  nor _19622_ (_11319_, _11231_, _11318_);
  and _19623_ (_11320_, _11231_, word_in[6]);
  or _19624_ (_11321_, _11320_, _11319_);
  or _19625_ (_11322_, _11321_, _11229_);
  or _19626_ (_11323_, _11236_, word_in[14]);
  and _19627_ (_11324_, _11323_, _11322_);
  or _19628_ (_11325_, _11324_, _11228_);
  or _19629_ (_11326_, _11243_, _10154_);
  and _19630_ (_11327_, _11326_, _11242_);
  and _19631_ (_11328_, _11327_, _11325_);
  and _19632_ (_11329_, _11241_, _09626_);
  or _19633_ (_14569_, _11329_, _11328_);
  nor _19634_ (_11330_, _11231_, _08565_);
  and _19635_ (_11331_, _11231_, word_in[7]);
  or _19636_ (_11332_, _11331_, _11330_);
  or _19637_ (_11333_, _11332_, _11229_);
  or _19638_ (_11334_, _11236_, word_in[15]);
  and _19639_ (_11335_, _11334_, _11333_);
  or _19640_ (_11336_, _11335_, _11228_);
  or _19641_ (_11337_, _11243_, _08886_);
  and _19642_ (_11338_, _11337_, _11336_);
  or _19643_ (_11339_, _11338_, _11241_);
  or _19644_ (_11340_, _11242_, word_in[31]);
  and _19645_ (_14570_, _11340_, _11339_);
  and _19646_ (_11341_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _19647_ (_11342_, _07229_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not _19648_ (_11343_, _11342_);
  or _19649_ (_11344_, _08441_, _07232_);
  nor _19650_ (_11345_, _07230_, \oc8051_top_1.oc8051_decoder1.op [4]);
  nor _19651_ (_11346_, _11345_, _07265_);
  and _19652_ (_11347_, _11346_, _11344_);
  not _19653_ (_11348_, _09327_);
  or _19654_ (_11349_, _08425_, _07232_);
  nor _19655_ (_11350_, _07230_, \oc8051_top_1.oc8051_decoder1.op [3]);
  nor _19656_ (_11351_, _11350_, _07265_);
  nand _19657_ (_11352_, _11351_, _11349_);
  and _19658_ (_11353_, _11352_, _11348_);
  and _19659_ (_11354_, _11353_, _09477_);
  and _19660_ (_11355_, _11354_, _07268_);
  and _19661_ (_11356_, _11355_, _11347_);
  or _19662_ (_11357_, _08457_, _07232_);
  nor _19663_ (_11358_, _07230_, \oc8051_top_1.oc8051_decoder1.op [5]);
  nor _19664_ (_11359_, _11358_, _07265_);
  nand _19665_ (_11360_, _11359_, _11357_);
  or _19666_ (_11361_, _08360_, _07232_);
  nor _19667_ (_11362_, _07230_, \oc8051_top_1.oc8051_decoder1.op [7]);
  nor _19668_ (_11363_, _11362_, _07265_);
  nand _19669_ (_11364_, _11363_, _11361_);
  nand _19670_ (_11365_, _08472_, _07231_);
  nor _19671_ (_11366_, _07230_, \oc8051_top_1.oc8051_decoder1.op [6]);
  nor _19672_ (_11367_, _11366_, _07265_);
  and _19673_ (_11368_, _11367_, _11365_);
  nor _19674_ (_11369_, _11368_, _11364_);
  and _19675_ (_11370_, _11369_, _11360_);
  and _19676_ (_11371_, _11370_, _11356_);
  and _19677_ (_11372_, _11359_, _11357_);
  and _19678_ (_11373_, _11368_, _11364_);
  and _19679_ (_11374_, _11373_, _11372_);
  and _19680_ (_11375_, _11356_, _11374_);
  not _19681_ (_11376_, _11347_);
  and _19682_ (_11377_, _11369_, _11372_);
  and _19683_ (_11378_, _11377_, _11376_);
  and _19684_ (_11379_, _11378_, _11355_);
  nor _19685_ (_11380_, _11379_, _11375_);
  not _19686_ (_11381_, _11380_);
  nor _19687_ (_11382_, _11381_, _11371_);
  nor _19688_ (_11383_, _11382_, _11343_);
  nor _19689_ (_11384_, _09477_, _07268_);
  and _19690_ (_11385_, _11384_, _11353_);
  not _19691_ (_11386_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and _19692_ (_11387_, \oc8051_top_1.oc8051_decoder1.state [1], _06308_);
  and _19693_ (_11389_, _11387_, _11386_);
  and _19694_ (_11390_, _11373_, _11389_);
  and _19695_ (_11391_, _11390_, _11385_);
  not _19696_ (_11392_, _11391_);
  and _19697_ (_11393_, _11352_, _09327_);
  and _19698_ (_11394_, _11384_, _11393_);
  and _19699_ (_11395_, _11370_, _11376_);
  and _19700_ (_11396_, _11395_, _11394_);
  and _19701_ (_11398_, _11378_, _11394_);
  nor _19702_ (_11399_, _11398_, _11396_);
  and _19703_ (_11400_, _11399_, _11392_);
  not _19704_ (_11401_, _11400_);
  nor _19705_ (_11402_, _11401_, _11383_);
  nor _19706_ (_11403_, _11402_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _19707_ (_11404_, _11403_, _11341_);
  and _19708_ (_11405_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  and _19709_ (_11406_, _11393_, _09477_);
  and _19710_ (_11407_, _11373_, _11360_);
  and _19711_ (_11408_, _11407_, _11376_);
  and _19712_ (_11409_, _11408_, _11406_);
  not _19713_ (_11410_, _11364_);
  and _19714_ (_11411_, _11360_, _11368_);
  and _19715_ (_11412_, _11411_, _11410_);
  and _19716_ (_11413_, _11385_, _11412_);
  and _19717_ (_11414_, _11413_, _11347_);
  nor _19718_ (_11415_, _11414_, _11409_);
  nand _19719_ (_11416_, _11395_, _11406_);
  and _19720_ (_11417_, _11372_, _11368_);
  and _19721_ (_11418_, _11417_, _11410_);
  and _19722_ (_11419_, _11418_, _11376_);
  nand _19723_ (_11420_, _11419_, _11406_);
  and _19724_ (_11421_, _11420_, _11416_);
  and _19725_ (_11422_, _11421_, _11415_);
  and _19726_ (_11423_, _11406_, _11347_);
  and _19727_ (_11424_, _11423_, _11377_);
  not _19728_ (_11425_, _11368_);
  and _19729_ (_11426_, _11425_, _11364_);
  and _19730_ (_11427_, _11426_, _11360_);
  and _19731_ (_11428_, _11406_, _11427_);
  nor _19732_ (_11429_, _11428_, _11424_);
  and _19733_ (_11430_, _11354_, _07311_);
  and _19734_ (_11431_, _11426_, _11372_);
  and _19735_ (_11432_, _11431_, _11430_);
  and _19736_ (_11433_, _11376_, _11374_);
  and _19737_ (_11434_, _11433_, _11406_);
  nor _19738_ (_11435_, _11434_, _11432_);
  and _19739_ (_11436_, _11435_, _11429_);
  and _19740_ (_11437_, _11407_, _11347_);
  and _19741_ (_11438_, _11437_, _11406_);
  and _19742_ (_11439_, _11406_, _11431_);
  or _19743_ (_11440_, _11439_, _11438_);
  not _19744_ (_11441_, _11440_);
  and _19745_ (_11442_, _11406_, _11412_);
  and _19746_ (_11443_, _11370_, _11347_);
  and _19747_ (_11444_, _11443_, _11406_);
  nor _19748_ (_11445_, _11444_, _11442_);
  and _19749_ (_11446_, _11445_, _11441_);
  and _19750_ (_11447_, _11446_, _11436_);
  and _19751_ (_11448_, _11447_, _11422_);
  and _19752_ (_11449_, _11448_, _11382_);
  nor _19753_ (_11450_, _11449_, _11343_);
  and _19754_ (_11451_, _11387_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and _19755_ (_11452_, _11432_, _11451_);
  and _19756_ (_11453_, _06308_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and _19757_ (_11454_, _11385_, _11431_);
  and _19758_ (_11455_, _11454_, _11376_);
  and _19759_ (_11456_, _11431_, _11347_);
  and _19760_ (_11457_, _11456_, _11385_);
  and _19761_ (_11458_, _11427_, _11347_);
  and _19762_ (_11459_, _11385_, _11458_);
  or _19763_ (_11460_, _11459_, _11457_);
  nor _19764_ (_11461_, _11460_, _11455_);
  and _19765_ (_11463_, _11391_, _11360_);
  not _19766_ (_11464_, _11463_);
  and _19767_ (_11465_, _11464_, _11461_);
  nor _19768_ (_11466_, _11465_, _11453_);
  nor _19769_ (_11467_, _11466_, _11392_);
  nor _19770_ (_11468_, _11467_, _11452_);
  not _19771_ (_11469_, _11468_);
  nor _19772_ (_11470_, _11469_, _11450_);
  nor _19773_ (_11471_, _11470_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _19774_ (_11472_, _11471_, _11405_);
  not _19775_ (_11473_, _11472_);
  and _19776_ (_11474_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and _19777_ (_11475_, _11347_, _11374_);
  and _19778_ (_11476_, _11475_, _11430_);
  and _19779_ (_11477_, _11408_, _11354_);
  nor _19780_ (_11478_, _11477_, _11476_);
  and _19781_ (_11479_, _11378_, _11385_);
  not _19782_ (_11480_, _09477_);
  and _19783_ (_11481_, _11480_, _07268_);
  and _19784_ (_11482_, _11393_, _11481_);
  and _19785_ (_11483_, _11408_, _11482_);
  nor _19786_ (_11484_, _11483_, _11479_);
  and _19787_ (_11485_, _11484_, _11478_);
  and _19788_ (_11486_, _11377_, _11347_);
  and _19789_ (_11487_, _11385_, _11486_);
  not _19790_ (_11488_, _11487_);
  and _19791_ (_11489_, _11486_, _11430_);
  and _19792_ (_11490_, _11412_, _11376_);
  and _19793_ (_11491_, _11490_, _11430_);
  nor _19794_ (_11492_, _11491_, _11489_);
  and _19795_ (_11493_, _11412_, _11347_);
  and _19796_ (_11494_, _11482_, _11493_);
  and _19797_ (_11495_, _11482_, _11458_);
  nor _19798_ (_11496_, _11495_, _11494_);
  and _19799_ (_11497_, _11496_, _11492_);
  and _19800_ (_11498_, _11497_, _11488_);
  and _19801_ (_11499_, _11498_, _11485_);
  not _19802_ (_11500_, _11482_);
  nor _19803_ (_11501_, _11443_, _11486_);
  or _19804_ (_11502_, _11501_, _11500_);
  and _19805_ (_11503_, _11433_, _11482_);
  and _19806_ (_11504_, _11490_, _11482_);
  nor _19807_ (_11505_, _11504_, _11503_);
  not _19808_ (_11507_, _11505_);
  or _19809_ (_11508_, _11443_, _11493_);
  and _19810_ (_11509_, _11508_, _11430_);
  nor _19811_ (_11510_, _11509_, _11507_);
  and _19812_ (_11511_, _11510_, _11502_);
  and _19813_ (_11512_, _11395_, _11430_);
  and _19814_ (_11513_, _11437_, _11354_);
  nor _19815_ (_11514_, _11513_, _11512_);
  not _19816_ (_11515_, _11514_);
  nor _19817_ (_11516_, _11437_, _11431_);
  nor _19818_ (_11517_, _11516_, _11500_);
  nor _19819_ (_11518_, _11517_, _11515_);
  nor _19820_ (_11519_, _11352_, _11347_);
  and _19821_ (_11520_, _11519_, _11377_);
  or _19822_ (_11521_, _11520_, _11413_);
  nor _19823_ (_11522_, _11521_, _11432_);
  and _19824_ (_11523_, _11427_, _11376_);
  and _19825_ (_11524_, _11482_, _11523_);
  and _19826_ (_11525_, _09477_, _09327_);
  not _19827_ (_11526_, _11352_);
  nor _19828_ (_11527_, _11526_, _11347_);
  and _19829_ (_11528_, _11527_, _11525_);
  and _19830_ (_11529_, _11528_, _11377_);
  nor _19831_ (_11530_, _11529_, _11524_);
  and _19832_ (_11531_, _11530_, _11522_);
  and _19833_ (_11532_, _11531_, _11518_);
  and _19834_ (_11533_, _11378_, _11430_);
  and _19835_ (_11534_, _11395_, _11482_);
  nor _19836_ (_11535_, _11534_, _11533_);
  and _19837_ (_11536_, _11433_, _11354_);
  and _19838_ (_11537_, _11419_, _11482_);
  nor _19839_ (_11538_, _11537_, _11536_);
  and _19840_ (_11539_, _11538_, _11535_);
  and _19841_ (_11540_, _11539_, _11461_);
  and _19842_ (_11541_, _11540_, _11532_);
  and _19843_ (_11542_, _11541_, _11511_);
  and _19844_ (_11543_, _11542_, _11499_);
  nor _19845_ (_11544_, _11543_, _11343_);
  nor _19846_ (_11545_, _11391_, _11452_);
  not _19847_ (_11546_, _11545_);
  nor _19848_ (_11547_, _11546_, _11544_);
  nor _19849_ (_11548_, _11547_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _19850_ (_11549_, _11548_, _11474_);
  and _19851_ (_11550_, _11549_, _11473_);
  and _19852_ (_11551_, _11550_, _11404_);
  and _19853_ (_11552_, _07309_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  and _19854_ (_11553_, _07331_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  nor _19855_ (_11554_, _11553_, _11552_);
  and _19856_ (_11555_, _07313_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  and _19857_ (_11556_, _07327_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  nor _19858_ (_11557_, _11556_, _11555_);
  and _19859_ (_11558_, _11557_, _11554_);
  and _19860_ (_11559_, _07325_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  and _19861_ (_11560_, _07318_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  nor _19862_ (_11561_, _11560_, _11559_);
  and _19863_ (_11562_, _07321_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  and _19864_ (_11563_, _07333_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  nor _19865_ (_11564_, _11563_, _11562_);
  and _19866_ (_11565_, _11564_, _11561_);
  and _19867_ (_11566_, _11565_, _11558_);
  nor _19868_ (_11567_, _11566_, _07307_);
  not _19869_ (_11568_, _06978_);
  and _19870_ (_11569_, _07307_, _11568_);
  nor _19871_ (_11570_, _11569_, _11567_);
  not _19872_ (_11571_, _11570_);
  and _19873_ (_11572_, _11571_, _11551_);
  not _19874_ (_11573_, _11572_);
  not _19875_ (_11574_, _11549_);
  not _19876_ (_11575_, _11404_);
  nor _19877_ (_11576_, _11472_, _11575_);
  and _19878_ (_11577_, _11576_, _11574_);
  and _19879_ (_11578_, _08978_, _06432_);
  and _19880_ (_11579_, _11578_, _06978_);
  not _19881_ (_11580_, _11578_);
  and _19882_ (_11581_, _11580_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor _19883_ (_11582_, _11580_, _07300_);
  nor _19884_ (_11583_, _11582_, _11581_);
  and _19885_ (_11584_, _11580_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor _19886_ (_11585_, _06644_, _06604_);
  not _19887_ (_11586_, _11585_);
  and _19888_ (_11587_, _11586_, _09124_);
  and _19889_ (_11588_, _11587_, _09121_);
  and _19890_ (_11589_, _11588_, _09114_);
  nor _19891_ (_11590_, _11589_, _11580_);
  nor _19892_ (_11591_, _11590_, _11584_);
  and _19893_ (_11592_, _11578_, _07070_);
  and _19894_ (_11593_, _11580_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  nor _19895_ (_11594_, _11593_, _11592_);
  nor _19896_ (_11595_, _11578_, _06401_);
  and _19897_ (_11596_, _11578_, _09527_);
  nor _19898_ (_11597_, _11596_, _11595_);
  and _19899_ (_11598_, _11597_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and _19900_ (_11599_, _11598_, _11594_);
  and _19901_ (_11600_, _11599_, _11591_);
  and _19902_ (_11601_, _11600_, _11583_);
  nor _19903_ (_11602_, _11580_, _07188_);
  and _19904_ (_11603_, _11580_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  nor _19905_ (_11604_, _11603_, _11602_);
  and _19906_ (_11605_, _11604_, _11601_);
  nor _19907_ (_11606_, _11580_, _06666_);
  and _19908_ (_11607_, _11580_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor _19909_ (_11608_, _11607_, _11606_);
  and _19910_ (_11609_, _11608_, _11605_);
  nor _19911_ (_11610_, _11580_, _10494_);
  and _19912_ (_11611_, _11580_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor _19913_ (_11612_, _11611_, _11610_);
  and _19914_ (_11613_, _11612_, _11609_);
  nor _19915_ (_11614_, _11578_, _06366_);
  nor _19916_ (_11615_, _11614_, _11613_);
  and _19917_ (_11616_, _11614_, _11613_);
  or _19918_ (_11617_, _11616_, _11615_);
  nor _19919_ (_11618_, _11617_, _06311_);
  nor _19920_ (_11619_, _11578_, _06370_);
  not _19921_ (_11620_, _11619_);
  nor _19922_ (_11621_, _11620_, _11618_);
  nor _19923_ (_11622_, _11621_, _11579_);
  and _19924_ (_11623_, _11622_, _11577_);
  not _19925_ (_11624_, _11623_);
  not _19926_ (_11625_, _08376_);
  nor _19927_ (_11626_, _11549_, _11473_);
  and _19928_ (_11627_, _11626_, _11625_);
  nor _19929_ (_11628_, _11627_, _11575_);
  and _19930_ (_11629_, _11628_, _11624_);
  and _19931_ (_11630_, _11629_, _11573_);
  nor _19932_ (_11631_, _11630_, _08030_);
  and _19933_ (_11632_, _11630_, _08030_);
  nor _19934_ (_11633_, _11632_, _11631_);
  and _19935_ (_11634_, _11472_, _11404_);
  and _19936_ (_11635_, _11634_, _11574_);
  nor _19937_ (_11636_, _07230_, _06747_);
  and _19938_ (_11637_, _07254_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and _19939_ (_11638_, _07238_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor _19940_ (_11639_, _11638_, _11637_);
  and _19941_ (_11640_, _07246_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and _19942_ (_11641_, _07251_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  nor _19943_ (_11642_, _11641_, _11640_);
  and _19944_ (_11643_, _07248_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and _19945_ (_11644_, _07242_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor _19946_ (_11645_, _11644_, _11643_);
  and _19947_ (_11646_, _11645_, _11642_);
  and _19948_ (_11647_, _11646_, _11639_);
  nor _19949_ (_11648_, _11647_, _08374_);
  nor _19950_ (_11649_, _11648_, _11636_);
  not _19951_ (_11650_, _11649_);
  and _19952_ (_11651_, _11650_, _11635_);
  and _19953_ (_11652_, _11634_, _11549_);
  and _19954_ (_11653_, _11652_, _07316_);
  nor _19955_ (_11654_, _11653_, _11651_);
  not _19956_ (_11655_, _07361_);
  and _19957_ (_11656_, _11551_, _11655_);
  not _19958_ (_11657_, _11656_);
  nor _19959_ (_11658_, _11604_, _11601_);
  nor _19960_ (_11659_, _11658_, _11605_);
  nor _19961_ (_11660_, _11659_, _06311_);
  nor _19962_ (_11661_, _11660_, _06315_);
  nor _19963_ (_11662_, _11661_, _11578_);
  nor _19964_ (_11663_, _11662_, _11602_);
  not _19965_ (_11664_, _11663_);
  and _19966_ (_11665_, _11664_, _11577_);
  and _19967_ (_11666_, _11472_, _11575_);
  nor _19968_ (_11667_, _11666_, _11665_);
  and _19969_ (_11668_, _11667_, _11657_);
  and _19970_ (_11669_, _11668_, _11654_);
  nor _19971_ (_11670_, _11669_, _06337_);
  and _19972_ (_11671_, _11669_, _06337_);
  nor _19973_ (_11672_, _11671_, _11670_);
  not _19974_ (_11673_, _07342_);
  and _19975_ (_11674_, _11551_, _11673_);
  nor _19976_ (_11675_, _07230_, _06770_);
  and _19977_ (_11676_, _07254_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and _19978_ (_11677_, _07238_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor _19979_ (_11678_, _11677_, _11676_);
  and _19980_ (_11679_, _07246_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and _19981_ (_11680_, _07242_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor _19982_ (_11681_, _11680_, _11679_);
  and _19983_ (_11682_, _07251_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  and _19984_ (_11683_, _07248_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nor _19985_ (_11684_, _11683_, _11682_);
  and _19986_ (_11685_, _11684_, _11681_);
  and _19987_ (_11686_, _11685_, _11678_);
  nor _19988_ (_11687_, _11686_, _08374_);
  nor _19989_ (_11688_, _11687_, _11675_);
  not _19990_ (_11689_, _11688_);
  and _19991_ (_11690_, _11689_, _11635_);
  nor _19992_ (_11691_, _11690_, _11674_);
  not _19993_ (_11692_, _07302_);
  and _19994_ (_11693_, _11652_, _11692_);
  nor _19995_ (_11694_, _11600_, _11583_);
  nor _19996_ (_11695_, _11694_, _11601_);
  nor _19997_ (_11696_, _11695_, _06311_);
  nor _19998_ (_11697_, _11696_, _06388_);
  nor _19999_ (_11698_, _11697_, _11578_);
  nor _20000_ (_11699_, _11698_, _11582_);
  not _20001_ (_11700_, _11699_);
  and _20002_ (_11701_, _11700_, _11577_);
  nor _20003_ (_11702_, _11701_, _11693_);
  and _20004_ (_11703_, _11702_, _11691_);
  nor _20005_ (_11704_, _11703_, _06395_);
  and _20006_ (_11705_, _11703_, _06395_);
  nor _20007_ (_11706_, _11705_, _11704_);
  and _20008_ (_11707_, _11706_, _11672_);
  not _20009_ (_11708_, _07380_);
  and _20010_ (_11709_, _11551_, _11708_);
  nor _20011_ (_11710_, _07230_, _06474_);
  and _20012_ (_11711_, _07254_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and _20013_ (_11712_, _07238_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor _20014_ (_11713_, _11712_, _11711_);
  and _20015_ (_11714_, _07246_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and _20016_ (_11715_, _07251_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor _20017_ (_11716_, _11715_, _11714_);
  and _20018_ (_11717_, _07248_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  not _20019_ (_11718_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor _20020_ (_11719_, _07241_, _11718_);
  nor _20021_ (_11720_, _11719_, _11717_);
  and _20022_ (_11721_, _11720_, _11716_);
  and _20023_ (_11723_, _11721_, _11713_);
  nor _20024_ (_11724_, _11723_, _08374_);
  nor _20025_ (_11725_, _11724_, _11710_);
  not _20026_ (_11726_, _11725_);
  and _20027_ (_11727_, _11726_, _11635_);
  nor _20028_ (_11728_, _11727_, _11709_);
  nor _20029_ (_11729_, _11608_, _11605_);
  nor _20030_ (_11730_, _11729_, _11609_);
  nor _20031_ (_11731_, _11730_, _06311_);
  nor _20032_ (_11732_, _11731_, _06342_);
  nor _20033_ (_11733_, _11732_, _11578_);
  nor _20034_ (_11734_, _11733_, _11606_);
  nor _20035_ (_11735_, _11734_, _11472_);
  nor _20036_ (_11736_, _11735_, _11575_);
  not _20037_ (_11737_, _11736_);
  nor _20038_ (_11738_, _11626_, _11550_);
  and _20039_ (_11739_, _11738_, _11737_);
  not _20040_ (_11740_, _11739_);
  and _20041_ (_11741_, _11740_, _11728_);
  and _20042_ (_11742_, _11741_, _06671_);
  nor _20043_ (_11743_, _11741_, _06671_);
  nor _20044_ (_11744_, _11743_, _11742_);
  and _20045_ (_11745_, _07321_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  and _20046_ (_11746_, _07318_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  nor _20047_ (_11747_, _11746_, _11745_);
  and _20048_ (_11749_, _07309_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  and _20049_ (_11750_, _07313_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  nor _20050_ (_11751_, _11750_, _11749_);
  and _20051_ (_11753_, _11751_, _11747_);
  and _20052_ (_11754_, _07327_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  and _20053_ (_11755_, _07333_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  nor _20054_ (_11756_, _11755_, _11754_);
  and _20055_ (_11757_, _07325_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  and _20056_ (_11758_, _07331_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  nor _20057_ (_11759_, _11758_, _11757_);
  and _20058_ (_11760_, _11759_, _11756_);
  and _20059_ (_11761_, _11760_, _11753_);
  nor _20060_ (_11762_, _11761_, _07307_);
  not _20061_ (_11763_, _10494_);
  and _20062_ (_11764_, _11763_, _07307_);
  nor _20063_ (_11765_, _11764_, _11762_);
  not _20064_ (_11766_, _11765_);
  and _20065_ (_11767_, _11766_, _11551_);
  nor _20066_ (_11769_, _11612_, _11609_);
  nor _20067_ (_11770_, _11769_, _11613_);
  nor _20068_ (_11771_, _11770_, _06311_);
  nor _20069_ (_11772_, _11771_, _06356_);
  nor _20070_ (_11773_, _11772_, _11578_);
  nor _20071_ (_11774_, _11773_, _11610_);
  not _20072_ (_11775_, _11774_);
  and _20073_ (_11776_, _11775_, _11577_);
  nor _20074_ (_11777_, _11776_, _11767_);
  not _20075_ (_11778_, _10734_);
  and _20076_ (_11779_, _11635_, _11778_);
  nor _20077_ (_11780_, _11550_, _11404_);
  nor _20078_ (_11781_, _11780_, _11779_);
  and _20079_ (_11782_, _11781_, _11777_);
  and _20080_ (_11784_, _11782_, _06365_);
  nor _20081_ (_11785_, _11782_, _06365_);
  nor _20082_ (_11786_, _11785_, _11784_);
  and _20083_ (_11787_, _11786_, _11744_);
  and _20084_ (_11788_, _11787_, _11707_);
  and _20085_ (_11789_, _11788_, _11633_);
  not _20086_ (_11790_, _10995_);
  and _20087_ (_11791_, _11551_, _11790_);
  not _20088_ (_11792_, _11791_);
  and _20089_ (_11793_, _11550_, _11575_);
  not _20090_ (_11794_, _11227_);
  and _20091_ (_11795_, _11635_, _11794_);
  nor _20092_ (_11796_, _11795_, _11793_);
  nor _20093_ (_11797_, _11598_, _11594_);
  nor _20094_ (_11798_, _11797_, _11599_);
  nor _20095_ (_11799_, _11798_, _06311_);
  nor _20096_ (_11800_, _11799_, _06410_);
  nor _20097_ (_11801_, _11800_, _11578_);
  nor _20098_ (_11802_, _11801_, _11592_);
  not _20099_ (_11803_, _11802_);
  and _20100_ (_11804_, _11803_, _11577_);
  and _20101_ (_11805_, _11652_, _09477_);
  nor _20102_ (_11807_, _11805_, _11804_);
  and _20103_ (_11808_, _11807_, _11796_);
  and _20104_ (_11809_, _11808_, _11792_);
  nor _20105_ (_11810_, _11809_, _06418_);
  and _20106_ (_11811_, _11809_, _06418_);
  nor _20107_ (_11812_, _11811_, _11810_);
  and _20108_ (_11813_, _07309_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  and _20109_ (_11814_, _07333_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  nor _20110_ (_11815_, _11814_, _11813_);
  and _20111_ (_11816_, _07313_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  and _20112_ (_11817_, _07327_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  nor _20113_ (_11818_, _11817_, _11816_);
  and _20114_ (_11819_, _11818_, _11815_);
  and _20115_ (_11820_, _07318_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  and _20116_ (_11821_, _07321_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  nor _20117_ (_11822_, _11821_, _11820_);
  and _20118_ (_11823_, _07325_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  and _20119_ (_11824_, _07331_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  nor _20120_ (_11825_, _11824_, _11823_);
  and _20121_ (_11826_, _11825_, _11822_);
  and _20122_ (_11827_, _11826_, _11819_);
  nor _20123_ (_11828_, _11827_, _07307_);
  and _20124_ (_11829_, _09527_, _07307_);
  nor _20125_ (_11830_, _11829_, _11828_);
  not _20126_ (_11831_, _11830_);
  and _20127_ (_11832_, _11831_, _11551_);
  nor _20128_ (_11833_, _07230_, _06801_);
  and _20129_ (_11834_, _07254_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and _20130_ (_11835_, _07238_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor _20131_ (_11836_, _11835_, _11834_);
  and _20132_ (_11837_, _07246_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  not _20133_ (_11838_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor _20134_ (_11839_, _07241_, _11838_);
  nor _20135_ (_11840_, _11839_, _11837_);
  and _20136_ (_11841_, _07251_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  and _20137_ (_11842_, _07248_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nor _20138_ (_11843_, _11842_, _11841_);
  and _20139_ (_11844_, _11843_, _11840_);
  and _20140_ (_11845_, _11844_, _11836_);
  nor _20141_ (_11846_, _11845_, _08374_);
  nor _20142_ (_11847_, _11846_, _11833_);
  not _20143_ (_11848_, _11847_);
  and _20144_ (_11849_, _11848_, _11635_);
  nor _20145_ (_11850_, _11849_, _11832_);
  and _20146_ (_11851_, _11652_, _07268_);
  nor _20147_ (_11852_, _11597_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  nor _20148_ (_11853_, _11852_, _11598_);
  nor _20149_ (_11854_, _11853_, _06311_);
  nor _20150_ (_11855_, _11854_, _06402_);
  nor _20151_ (_11856_, _11855_, _11578_);
  nor _20152_ (_11857_, _11856_, _11596_);
  not _20153_ (_11858_, _11857_);
  and _20154_ (_11859_, _11858_, _11577_);
  nor _20155_ (_11860_, _11859_, _11851_);
  and _20156_ (_11861_, _11860_, _11850_);
  and _20157_ (_11862_, _11861_, _06407_);
  nor _20158_ (_11863_, _11861_, _06407_);
  or _20159_ (_11864_, _11863_, _11862_);
  nor _20160_ (_11865_, _11864_, _11812_);
  and _20161_ (_11866_, _07321_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  and _20162_ (_11867_, _07327_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  nor _20163_ (_11868_, _11867_, _11866_);
  and _20164_ (_11869_, _07313_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  and _20165_ (_11870_, _07331_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  nor _20166_ (_11871_, _11870_, _11869_);
  and _20167_ (_11872_, _11871_, _11868_);
  and _20168_ (_11873_, _07318_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  and _20169_ (_11874_, _07333_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  nor _20170_ (_11875_, _11874_, _11873_);
  and _20171_ (_11876_, _07309_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  and _20172_ (_11877_, _07325_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  nor _20173_ (_11878_, _11877_, _11876_);
  and _20174_ (_11879_, _11878_, _11875_);
  and _20175_ (_11880_, _11879_, _11872_);
  nor _20176_ (_11881_, _11880_, _07307_);
  not _20177_ (_11882_, _11589_);
  and _20178_ (_11883_, _11882_, _07307_);
  nor _20179_ (_11884_, _11883_, _11881_);
  not _20180_ (_11885_, _11884_);
  and _20181_ (_11886_, _11885_, _11551_);
  not _20182_ (_11887_, _11886_);
  and _20183_ (_11888_, _11652_, _09327_);
  nor _20184_ (_11889_, _07230_, _06780_);
  and _20185_ (_11890_, _07254_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and _20186_ (_11891_, _07238_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor _20187_ (_11892_, _11891_, _11890_);
  and _20188_ (_11893_, _07246_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and _20189_ (_11895_, _07251_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  nor _20190_ (_11896_, _11895_, _11893_);
  and _20191_ (_11897_, _07248_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and _20192_ (_11899_, _07242_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor _20193_ (_11900_, _11899_, _11897_);
  and _20194_ (_11901_, _11900_, _11896_);
  and _20195_ (_11902_, _11901_, _11892_);
  nor _20196_ (_11903_, _11902_, _08374_);
  nor _20197_ (_11904_, _11903_, _11889_);
  not _20198_ (_11905_, _11904_);
  and _20199_ (_11906_, _11905_, _11635_);
  nor _20200_ (_11907_, _11599_, _11591_);
  nor _20201_ (_11908_, _11907_, _11600_);
  nor _20202_ (_11909_, _11908_, _06311_);
  nor _20203_ (_11910_, _11909_, _06421_);
  nor _20204_ (_11911_, _11910_, _11578_);
  nor _20205_ (_11912_, _11911_, _11590_);
  not _20206_ (_11914_, _11912_);
  and _20207_ (_11915_, _11914_, _11577_);
  or _20208_ (_11917_, _11915_, _11906_);
  nor _20209_ (_11918_, _11917_, _11888_);
  and _20210_ (_11919_, _11918_, _11887_);
  nor _20211_ (_11920_, _11919_, _06430_);
  and _20212_ (_11921_, _11919_, _06430_);
  nor _20213_ (_11922_, _11921_, _11920_);
  nor _20214_ (_11923_, _11922_, _08925_);
  and _20215_ (_11924_, _11923_, _11865_);
  and _20216_ (_11925_, _11924_, _11789_);
  nor _20217_ (_11926_, _06380_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and _20218_ (_11927_, _11926_, _11925_);
  not _20219_ (_11928_, _11927_);
  and _20220_ (_11929_, _11466_, _11392_);
  nor _20221_ (_11930_, _06933_, _06943_);
  and _20222_ (_11931_, _11930_, _11789_);
  and _20223_ (_11932_, _11931_, _11929_);
  and _20224_ (_11933_, _11481_, _11353_);
  and _20225_ (_11934_, _11427_, _11430_);
  nor _20226_ (_11935_, _11934_, _11933_);
  nor _20227_ (_11936_, _11935_, _11343_);
  not _20228_ (_11937_, _11128_);
  not _20229_ (_11938_, _11466_);
  nor _20230_ (_11939_, _06822_, _06763_);
  and _20231_ (_11940_, _11939_, _07991_);
  and _20232_ (_11941_, _11940_, _09098_);
  and _20233_ (_11942_, _11941_, _11392_);
  and _20234_ (_11943_, _11942_, _08287_);
  not _20235_ (_11944_, _11943_);
  nor _20236_ (_11945_, _11944_, _08209_);
  and _20237_ (_11946_, _11945_, _11938_);
  and _20238_ (_11947_, _11946_, _08999_);
  and _20239_ (_11948_, _11947_, _11937_);
  nor _20240_ (_11949_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor _20241_ (_11950_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and _20242_ (_11951_, _11950_, _11949_);
  nor _20243_ (_11952_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor _20244_ (_11953_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and _20245_ (_11954_, _11953_, _11952_);
  and _20246_ (_11955_, _11954_, _11951_);
  and _20247_ (_11957_, _11955_, _11467_);
  not _20248_ (_11958_, _11957_);
  and _20249_ (_11959_, _11929_, _06463_);
  and _20250_ (_11960_, _11463_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor _20251_ (_11961_, _11960_, _11959_);
  and _20252_ (_11962_, _11961_, _11958_);
  not _20253_ (_11963_, _11962_);
  nor _20254_ (_11964_, _11963_, _11948_);
  and _20255_ (_11965_, _11393_, _11480_);
  and _20256_ (_11966_, _11965_, _11486_);
  nor _20257_ (_11967_, _11966_, _11494_);
  and _20258_ (_11968_, _11493_, _11526_);
  not _20259_ (_11969_, _11968_);
  and _20260_ (_11970_, _11969_, _11967_);
  not _20261_ (_11971_, _11385_);
  nor _20262_ (_11972_, _11437_, _11475_);
  nor _20263_ (_11973_, _11972_, _11971_);
  not _20264_ (_11974_, _11973_);
  not _20265_ (_11975_, _11457_);
  and _20266_ (_11976_, _11526_, _11347_);
  and _20267_ (_11977_, _11976_, _11377_);
  nor _20268_ (_11978_, _11977_, _11424_);
  and _20269_ (_11979_, _11978_, _11975_);
  and _20270_ (_11980_, _11979_, _11974_);
  and _20271_ (_11981_, _11980_, _11970_);
  not _20272_ (_11982_, _11981_);
  and _20273_ (_11983_, _11982_, _11964_);
  not _20274_ (_11984_, _11432_);
  and _20275_ (_11986_, _11395_, _11385_);
  nor _20276_ (_11987_, _11986_, _11375_);
  nand _20277_ (_11989_, _11987_, _11984_);
  nor _20278_ (_11990_, _11989_, _11983_);
  and _20279_ (_11991_, _11431_, _11376_);
  and _20280_ (_11993_, _11991_, _11385_);
  nor _20281_ (_11994_, _11993_, _11459_);
  nand _20282_ (_11995_, _11376_, _11373_);
  nor _20283_ (_11996_, _11995_, _11971_);
  not _20284_ (_11997_, _11996_);
  and _20285_ (_11998_, _11997_, _11994_);
  nor _20286_ (_11999_, _11998_, _11964_);
  not _20287_ (_12001_, _11999_);
  and _20288_ (_12002_, _12001_, _11990_);
  nor _20289_ (_12003_, _11452_, _11389_);
  nor _20290_ (_12004_, _12003_, _12002_);
  nor _20291_ (_12005_, _12004_, _11936_);
  nor _20292_ (_12006_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  not _20293_ (_12008_, _12006_);
  nor _20294_ (_12009_, _12008_, _07218_);
  nor _20295_ (_12011_, _06395_, _06336_);
  and _20296_ (_12012_, _12011_, _06677_);
  not _20297_ (_12013_, _12012_);
  and _20298_ (_12014_, _12013_, _12009_);
  nor _20299_ (_12015_, _12014_, _11464_);
  not _20300_ (_12016_, _08036_);
  and _20301_ (_12017_, _11467_, _12016_);
  nor _20302_ (_12018_, _12017_, _12015_);
  not _20303_ (_12019_, _12018_);
  nor _20304_ (_12020_, _12019_, _12005_);
  not _20305_ (_12021_, _12020_);
  nor _20306_ (_12022_, _12021_, _11932_);
  and _20307_ (_12023_, _12022_, _11928_);
  not _20308_ (_12024_, _09045_);
  and _20309_ (_12025_, _11475_, _11355_);
  and _20310_ (_12026_, _12025_, _11389_);
  nor _20311_ (_12028_, _12026_, _11936_);
  and _20312_ (_12029_, _11978_, _11461_);
  nand _20313_ (_12030_, _12029_, _11967_);
  nand _20314_ (_12031_, _12030_, _11389_);
  and _20315_ (_12032_, _11934_, _11342_);
  not _20316_ (_12033_, _12032_);
  and _20317_ (_12034_, _11454_, _11342_);
  nor _20318_ (_12035_, _12034_, _11452_);
  and _20319_ (_12037_, _12035_, _12033_);
  nand _20320_ (_12038_, _12037_, _12031_);
  not _20321_ (_12039_, _11389_);
  and _20322_ (_12040_, _11385_, _11373_);
  not _20323_ (_12041_, _12040_);
  and _20324_ (_12042_, _11970_, _12041_);
  and _20325_ (_12043_, _12042_, _11987_);
  and _20326_ (_12044_, _12043_, _12029_);
  nor _20327_ (_12045_, _12044_, _12039_);
  nor _20328_ (_12046_, _12045_, _12038_);
  and _20329_ (_12047_, _12046_, _12028_);
  or _20330_ (_12048_, _12047_, _12026_);
  and _20331_ (_12050_, _12048_, _12024_);
  and _20332_ (_12051_, _11452_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or _20333_ (_12052_, _12038_, _12028_);
  nor _20334_ (_12054_, _12052_, _12045_);
  and _20335_ (_12055_, _12054_, _11778_);
  and _20336_ (_12056_, _07429_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  or _20337_ (_12058_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _07234_);
  and _20338_ (_12059_, _07248_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and _20339_ (_12060_, _07246_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  or _20340_ (_12061_, _12060_, _12059_);
  and _20341_ (_12062_, _07251_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  and _20342_ (_12063_, _07254_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and _20343_ (_12064_, _07238_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  or _20344_ (_12065_, _12064_, _12063_);
  or _20345_ (_12066_, _12065_, _12062_);
  or _20346_ (_12067_, _12066_, _12061_);
  and _20347_ (_12068_, _07242_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  or _20348_ (_12069_, _12068_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  or _20349_ (_12070_, _12069_, _12067_);
  and _20350_ (_12071_, _12070_, _07230_);
  and _20351_ (_12072_, _12071_, _12058_);
  nor _20352_ (_12073_, _12072_, _12056_);
  not _20353_ (_12074_, _12073_);
  and _20354_ (_12075_, _12074_, _12032_);
  or _20355_ (_12076_, _12075_, _12055_);
  or _20356_ (_12077_, _12076_, _12051_);
  not _20357_ (_12078_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and _20358_ (_12079_, _12037_, _12031_);
  and _20359_ (_12080_, _12079_, _11778_);
  and _20360_ (_12081_, _12074_, _12038_);
  nor _20361_ (_12082_, _12081_, _12080_);
  nor _20362_ (_12084_, _12082_, _12078_);
  and _20363_ (_12085_, _12082_, _12078_);
  nor _20364_ (_12086_, _12085_, _12084_);
  and _20365_ (_12087_, _11725_, _12079_);
  and _20366_ (_12088_, _07429_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [5]);
  and _20367_ (_12090_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and _20368_ (_12091_, _07254_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  not _20369_ (_12092_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor _20370_ (_12093_, _07241_, _12092_);
  nor _20371_ (_12094_, _12093_, _12091_);
  and _20372_ (_12095_, _07248_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and _20373_ (_12096_, _07238_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor _20374_ (_12097_, _12096_, _12095_);
  and _20375_ (_12098_, _12097_, _12094_);
  and _20376_ (_12099_, _07246_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and _20377_ (_12100_, _07251_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor _20378_ (_12101_, _12100_, _12099_);
  and _20379_ (_12102_, _12101_, _12098_);
  nor _20380_ (_12103_, _12102_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _20381_ (_12104_, _12103_, _12090_);
  nor _20382_ (_12105_, _12104_, _07429_);
  nor _20383_ (_12106_, _12105_, _12088_);
  and _20384_ (_12107_, _12106_, _12038_);
  nor _20385_ (_12108_, _12107_, _12087_);
  nor _20386_ (_12109_, _12108_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and _20387_ (_12110_, _12108_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and _20388_ (_12111_, _11649_, _12079_);
  and _20389_ (_12112_, _07429_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [4]);
  or _20390_ (_12113_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _07234_);
  and _20391_ (_12114_, _07248_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and _20392_ (_12115_, _07246_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  or _20393_ (_12116_, _12115_, _12114_);
  and _20394_ (_12117_, _07251_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  and _20395_ (_12118_, _07254_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and _20396_ (_12119_, _07238_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  or _20397_ (_12120_, _12119_, _12118_);
  or _20398_ (_12121_, _12120_, _12117_);
  or _20399_ (_12122_, _12121_, _12116_);
  and _20400_ (_12123_, _07242_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  or _20401_ (_12124_, _12123_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  or _20402_ (_12125_, _12124_, _12122_);
  and _20403_ (_12126_, _12125_, _07230_);
  and _20404_ (_12127_, _12126_, _12113_);
  nor _20405_ (_12128_, _12127_, _12112_);
  and _20406_ (_12129_, _12128_, _12038_);
  nor _20407_ (_12130_, _12129_, _12111_);
  nand _20408_ (_12131_, _12130_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _20409_ (_12132_, _11688_, _12079_);
  and _20410_ (_12134_, _07429_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [3]);
  and _20411_ (_12135_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and _20412_ (_12136_, _07254_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  not _20413_ (_12137_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor _20414_ (_12138_, _07241_, _12137_);
  nor _20415_ (_12139_, _12138_, _12136_);
  and _20416_ (_12141_, _07248_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and _20417_ (_12142_, _07238_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor _20418_ (_12144_, _12142_, _12141_);
  and _20419_ (_12145_, _12144_, _12139_);
  and _20420_ (_12146_, _07246_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and _20421_ (_12147_, _07251_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor _20422_ (_12148_, _12147_, _12146_);
  and _20423_ (_12149_, _12148_, _12145_);
  nor _20424_ (_12150_, _12149_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _20425_ (_12151_, _12150_, _12135_);
  nor _20426_ (_12152_, _12151_, _07429_);
  nor _20427_ (_12154_, _12152_, _12134_);
  and _20428_ (_12155_, _12154_, _12038_);
  nor _20429_ (_12156_, _12155_, _12132_);
  nor _20430_ (_12157_, _12156_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and _20431_ (_12158_, _12156_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  not _20432_ (_12160_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  or _20433_ (_12161_, _11905_, _12038_);
  not _20434_ (_12162_, _11209_);
  or _20435_ (_12163_, _12079_, _12162_);
  nand _20436_ (_12164_, _12163_, _12161_);
  or _20437_ (_12165_, _12164_, _12160_);
  not _20438_ (_12166_, _12165_);
  or _20439_ (_12167_, _12038_, _11794_);
  and _20440_ (_12168_, _07429_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [1]);
  and _20441_ (_12169_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and _20442_ (_12170_, _07248_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  not _20443_ (_12171_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor _20444_ (_12172_, _07241_, _12171_);
  nor _20445_ (_12173_, _12172_, _12170_);
  and _20446_ (_12174_, _07246_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and _20447_ (_12175_, _07238_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nor _20448_ (_12176_, _12175_, _12174_);
  and _20449_ (_12177_, _07251_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  and _20450_ (_12178_, _07254_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor _20451_ (_12179_, _12178_, _12177_);
  and _20452_ (_12180_, _12179_, _12176_);
  and _20453_ (_12181_, _12180_, _12173_);
  nor _20454_ (_12182_, _12181_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _20455_ (_12183_, _12182_, _12169_);
  nor _20456_ (_12184_, _12183_, _07429_);
  nor _20457_ (_12185_, _12184_, _12168_);
  not _20458_ (_12186_, _12185_);
  or _20459_ (_12187_, _12186_, _12079_);
  and _20460_ (_12188_, _12187_, _12167_);
  nand _20461_ (_12189_, _12188_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  or _20462_ (_12190_, _11848_, _12038_);
  not _20463_ (_12191_, _09672_);
  or _20464_ (_12192_, _12079_, _12191_);
  and _20465_ (_12193_, _12192_, _12190_);
  and _20466_ (_12194_, _12193_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  or _20467_ (_12195_, _12188_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and _20468_ (_12196_, _12195_, _12189_);
  and _20469_ (_12197_, _12196_, _12194_);
  not _20470_ (_12198_, _12197_);
  nand _20471_ (_12199_, _12198_, _12189_);
  nand _20472_ (_12200_, _12164_, _12160_);
  and _20473_ (_12201_, _12200_, _12165_);
  and _20474_ (_12202_, _12201_, _12199_);
  or _20475_ (_12203_, _12202_, _12166_);
  nor _20476_ (_12204_, _12203_, _12158_);
  nor _20477_ (_12205_, _12204_, _12157_);
  or _20478_ (_12206_, _12130_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _20479_ (_12207_, _12206_, _12131_);
  nand _20480_ (_12208_, _12207_, _12205_);
  nand _20481_ (_12209_, _12208_, _12131_);
  nor _20482_ (_12210_, _12209_, _12110_);
  nor _20483_ (_12211_, _12210_, _12109_);
  and _20484_ (_12212_, _12211_, _12086_);
  nor _20485_ (_12213_, _12211_, _12086_);
  nor _20486_ (_12214_, _12213_, _12212_);
  and _20487_ (_12215_, _11385_, _11342_);
  and _20488_ (_12216_, _12215_, _11431_);
  or _20489_ (_12217_, _12216_, _12045_);
  and _20490_ (_12218_, _12217_, _12052_);
  and _20491_ (_12219_, _12218_, _12214_);
  or _20492_ (_12220_, _12219_, _12077_);
  nor _20493_ (_12221_, _12220_, _12050_);
  nand _20494_ (_12222_, _12221_, _12023_);
  not _20495_ (_12223_, _07432_);
  and _20496_ (_12224_, _10949_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and _20497_ (_12225_, _12224_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and _20498_ (_12226_, _12225_, _12223_);
  and _20499_ (_12227_, _12226_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor _20500_ (_12228_, _12226_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor _20501_ (_12229_, _12228_, _12227_);
  or _20502_ (_12230_, _12229_, _12023_);
  and _20503_ (_12231_, _12230_, _06444_);
  and _20504_ (_09725_, _12231_, _12222_);
  nor _20505_ (_09730_, _11884_, rst);
  or _20506_ (_12232_, _07432_, \oc8051_top_1.oc8051_rom1.data_o [5]);
  nand _20507_ (_12233_, _07432_, _10716_);
  and _20508_ (_12234_, _12233_, _06444_);
  and _20509_ (_09742_, _12234_, _12232_);
  and _20510_ (_12235_, _08866_, _08655_);
  not _20511_ (_12236_, _12235_);
  and _20512_ (_12237_, _08869_, _09400_);
  not _20513_ (_12238_, _12237_);
  or _20514_ (_12239_, _12238_, word_in[8]);
  not _20515_ (_12240_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  and _20516_ (_12241_, _10069_, _08877_);
  nor _20517_ (_12242_, _12241_, _12240_);
  and _20518_ (_12243_, _12241_, word_in[0]);
  or _20519_ (_12244_, _12243_, _12242_);
  or _20520_ (_12245_, _12244_, _12237_);
  and _20521_ (_12246_, _12245_, _12239_);
  and _20522_ (_12247_, _12246_, _12236_);
  and _20523_ (_12248_, _08855_, _09219_);
  and _20524_ (_12249_, _12235_, _09837_);
  or _20525_ (_12250_, _12249_, _12248_);
  or _20526_ (_12251_, _12250_, _12247_);
  not _20527_ (_12252_, _12248_);
  or _20528_ (_12253_, _12252_, _09554_);
  and _20529_ (_09784_, _12253_, _12251_);
  not _20530_ (_12254_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  nor _20531_ (_12255_, _12241_, _12254_);
  and _20532_ (_12256_, _12241_, word_in[1]);
  or _20533_ (_12257_, _12256_, _12255_);
  and _20534_ (_12258_, _12257_, _12238_);
  and _20535_ (_12260_, _12237_, word_in[9]);
  or _20536_ (_12261_, _12260_, _12258_);
  and _20537_ (_12262_, _12261_, _12236_);
  and _20538_ (_12263_, _12235_, _09565_);
  or _20539_ (_12264_, _12263_, _12248_);
  or _20540_ (_12265_, _12264_, _12262_);
  or _20541_ (_12266_, _12252_, _11261_);
  and _20542_ (_09786_, _12266_, _12265_);
  not _20543_ (_12267_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  nor _20544_ (_12268_, _12241_, _12267_);
  and _20545_ (_12269_, _12241_, word_in[2]);
  or _20546_ (_12270_, _12269_, _12268_);
  and _20547_ (_12271_, _12270_, _12238_);
  and _20548_ (_12272_, _12237_, word_in[10]);
  or _20549_ (_12273_, _12272_, _12271_);
  and _20550_ (_12274_, _12273_, _12236_);
  and _20551_ (_12275_, _12235_, _10099_);
  or _20552_ (_12276_, _12275_, _12248_);
  or _20553_ (_12277_, _12276_, _12274_);
  or _20554_ (_12278_, _12252_, _09582_);
  and _20555_ (_09789_, _12278_, _12277_);
  or _20556_ (_12279_, _12238_, word_in[11]);
  not _20557_ (_12280_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  nor _20558_ (_12281_, _12241_, _12280_);
  and _20559_ (_12282_, _12241_, word_in[3]);
  or _20560_ (_12283_, _12282_, _12281_);
  or _20561_ (_12284_, _12283_, _12237_);
  and _20562_ (_12285_, _12284_, _12279_);
  and _20563_ (_12286_, _12285_, _12236_);
  and _20564_ (_12287_, _12235_, _10116_);
  or _20565_ (_12288_, _12287_, _12248_);
  or _20566_ (_12289_, _12288_, _12286_);
  or _20567_ (_12290_, _12252_, _09596_);
  and _20568_ (_09791_, _12290_, _12289_);
  or _20569_ (_12291_, _12238_, word_in[12]);
  not _20570_ (_12292_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  nor _20571_ (_12293_, _12241_, _12292_);
  and _20572_ (_12294_, _12241_, word_in[4]);
  or _20573_ (_12295_, _12294_, _12293_);
  or _20574_ (_12296_, _12295_, _12237_);
  and _20575_ (_12297_, _12296_, _12291_);
  and _20576_ (_12298_, _12297_, _12236_);
  and _20577_ (_12299_, _12235_, _10020_);
  or _20578_ (_12300_, _12299_, _12248_);
  or _20579_ (_12301_, _12300_, _12298_);
  or _20580_ (_12302_, _12252_, _09609_);
  and _20581_ (_09793_, _12302_, _12301_);
  not _20582_ (_12303_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  nor _20583_ (_12305_, _12241_, _12303_);
  and _20584_ (_12306_, _12241_, word_in[5]);
  or _20585_ (_12307_, _12306_, _12305_);
  and _20586_ (_12308_, _12307_, _12238_);
  and _20587_ (_12309_, _12237_, word_in[13]);
  or _20588_ (_12310_, _12309_, _12308_);
  and _20589_ (_12311_, _12310_, _12236_);
  and _20590_ (_12312_, _12235_, _10149_);
  or _20591_ (_12313_, _12312_, _12248_);
  or _20592_ (_12314_, _12313_, _12311_);
  or _20593_ (_12315_, _12252_, _09623_);
  and _20594_ (_09796_, _12315_, _12314_);
  or _20595_ (_12316_, _12238_, word_in[14]);
  not _20596_ (_12318_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  nor _20597_ (_12319_, _12241_, _12318_);
  and _20598_ (_12320_, _12241_, word_in[6]);
  or _20599_ (_12321_, _12320_, _12319_);
  or _20600_ (_12322_, _12321_, _12237_);
  and _20601_ (_12323_, _12322_, _12316_);
  and _20602_ (_12324_, _12323_, _12236_);
  and _20603_ (_12325_, _12235_, _10154_);
  or _20604_ (_12326_, _12325_, _12248_);
  or _20605_ (_12327_, _12326_, _12324_);
  or _20606_ (_12328_, _12252_, _09626_);
  and _20607_ (_09799_, _12328_, _12327_);
  nor _20608_ (_12329_, _12241_, _08685_);
  and _20609_ (_12330_, _12241_, word_in[7]);
  or _20610_ (_12331_, _12330_, _12329_);
  and _20611_ (_12332_, _12331_, _12238_);
  and _20612_ (_12333_, _12237_, word_in[15]);
  or _20613_ (_12335_, _12333_, _12332_);
  and _20614_ (_12336_, _12335_, _12236_);
  and _20615_ (_12337_, _12235_, _08886_);
  or _20616_ (_12338_, _12337_, _12248_);
  or _20617_ (_12339_, _12338_, _12336_);
  or _20618_ (_12340_, _12252_, _08856_);
  and _20619_ (_09801_, _12340_, _12339_);
  nor _20620_ (_09849_, _11765_, rst);
  nor _20621_ (_09852_, _11847_, rst);
  nor _20622_ (_09859_, _11649_, rst);
  nor _20623_ (_09863_, _12185_, rst);
  and _20624_ (_12342_, _08855_, _08655_);
  and _20625_ (_12343_, _12342_, _08842_);
  not _20626_ (_12344_, _12343_);
  and _20627_ (_12345_, _08866_, _08613_);
  and _20628_ (_12346_, _09695_, _08679_);
  not _20629_ (_12347_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  and _20630_ (_12348_, _09699_, _08877_);
  nor _20631_ (_12349_, _12348_, _12347_);
  and _20632_ (_12350_, _12348_, word_in[0]);
  or _20633_ (_12352_, _12350_, _12349_);
  or _20634_ (_12353_, _12352_, _12346_);
  not _20635_ (_12354_, _12346_);
  or _20636_ (_12355_, _12354_, word_in[8]);
  and _20637_ (_12357_, _12355_, _12353_);
  or _20638_ (_12358_, _12357_, _12345_);
  not _20639_ (_12359_, _12345_);
  or _20640_ (_12360_, _12359_, _09837_);
  and _20641_ (_12361_, _12360_, _12358_);
  and _20642_ (_12362_, _12361_, _12344_);
  and _20643_ (_12363_, _12343_, word_in[24]);
  or _20644_ (_14571_, _12363_, _12362_);
  and _20645_ (_12364_, _12348_, word_in[1]);
  not _20646_ (_12365_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  nor _20647_ (_12366_, _12348_, _12365_);
  nor _20648_ (_12367_, _12366_, _12364_);
  nor _20649_ (_12368_, _12367_, _12346_);
  and _20650_ (_12369_, _12346_, word_in[9]);
  or _20651_ (_12370_, _12369_, _12368_);
  and _20652_ (_12371_, _12370_, _12359_);
  and _20653_ (_12372_, _12345_, _09565_);
  or _20654_ (_12373_, _12372_, _12371_);
  and _20655_ (_12374_, _12373_, _12344_);
  and _20656_ (_12376_, _12343_, word_in[25]);
  or _20657_ (_09872_, _12376_, _12374_);
  and _20658_ (_12377_, _12348_, word_in[2]);
  not _20659_ (_12378_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  nor _20660_ (_12379_, _12348_, _12378_);
  nor _20661_ (_12381_, _12379_, _12377_);
  nor _20662_ (_12382_, _12381_, _12346_);
  and _20663_ (_12383_, _12346_, word_in[10]);
  or _20664_ (_12384_, _12383_, _12382_);
  and _20665_ (_12385_, _12384_, _12359_);
  and _20666_ (_12386_, _12345_, _10099_);
  or _20667_ (_12387_, _12386_, _12385_);
  and _20668_ (_12388_, _12387_, _12344_);
  and _20669_ (_12389_, _12343_, word_in[26]);
  or _20670_ (_09877_, _12389_, _12388_);
  and _20671_ (_12390_, _12348_, word_in[3]);
  not _20672_ (_12391_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  nor _20673_ (_12392_, _12348_, _12391_);
  nor _20674_ (_12393_, _12392_, _12390_);
  nor _20675_ (_12394_, _12393_, _12346_);
  and _20676_ (_12395_, _12346_, word_in[11]);
  or _20677_ (_12396_, _12395_, _12394_);
  and _20678_ (_12397_, _12396_, _12359_);
  and _20679_ (_12398_, _12345_, _10116_);
  or _20680_ (_12399_, _12398_, _12397_);
  and _20681_ (_12400_, _12399_, _12344_);
  and _20682_ (_12401_, _12343_, word_in[27]);
  or _20683_ (_09880_, _12401_, _12400_);
  and _20684_ (_12402_, _12348_, word_in[4]);
  not _20685_ (_12403_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  nor _20686_ (_12404_, _12348_, _12403_);
  nor _20687_ (_12405_, _12404_, _12402_);
  nor _20688_ (_12406_, _12405_, _12346_);
  and _20689_ (_12408_, _12346_, word_in[12]);
  or _20690_ (_12410_, _12408_, _12406_);
  and _20691_ (_12411_, _12410_, _12359_);
  and _20692_ (_12412_, _12345_, _10020_);
  or _20693_ (_12413_, _12412_, _12411_);
  and _20694_ (_12414_, _12413_, _12344_);
  and _20695_ (_12415_, _12343_, word_in[28]);
  or _20696_ (_09884_, _12415_, _12414_);
  not _20697_ (_12416_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  nor _20698_ (_12417_, _12348_, _12416_);
  and _20699_ (_12418_, _12348_, word_in[5]);
  nor _20700_ (_12419_, _12418_, _12417_);
  nor _20701_ (_12420_, _12419_, _12346_);
  and _20702_ (_12421_, _12346_, word_in[13]);
  or _20703_ (_12422_, _12421_, _12420_);
  and _20704_ (_12423_, _12422_, _12359_);
  and _20705_ (_12424_, _12345_, _10149_);
  or _20706_ (_12425_, _12424_, _12423_);
  and _20707_ (_12426_, _12425_, _12344_);
  and _20708_ (_12427_, _12343_, word_in[29]);
  or _20709_ (_09887_, _12427_, _12426_);
  and _20710_ (_12428_, _12348_, word_in[6]);
  not _20711_ (_12429_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  nor _20712_ (_12430_, _12348_, _12429_);
  nor _20713_ (_12431_, _12430_, _12428_);
  nor _20714_ (_12432_, _12431_, _12346_);
  and _20715_ (_12433_, _12346_, word_in[14]);
  or _20716_ (_12434_, _12433_, _12432_);
  and _20717_ (_12435_, _12434_, _12359_);
  and _20718_ (_12436_, _12345_, _10154_);
  or _20719_ (_12437_, _12436_, _12435_);
  and _20720_ (_12438_, _12437_, _12344_);
  and _20721_ (_12439_, _12343_, word_in[30]);
  or _20722_ (_09890_, _12439_, _12438_);
  nor _20723_ (_12440_, _12348_, _08571_);
  and _20724_ (_12441_, _12348_, word_in[7]);
  nor _20725_ (_12442_, _12441_, _12440_);
  nor _20726_ (_12443_, _12442_, _12346_);
  and _20727_ (_12444_, _12346_, word_in[15]);
  or _20728_ (_12445_, _12444_, _12443_);
  and _20729_ (_12446_, _12445_, _12359_);
  and _20730_ (_12447_, _12345_, _08886_);
  or _20731_ (_12448_, _12447_, _12446_);
  and _20732_ (_12449_, _12448_, _12344_);
  and _20733_ (_12450_, _12343_, word_in[31]);
  or _20734_ (_09894_, _12450_, _12449_);
  or _20735_ (_12451_, _07432_, \oc8051_top_1.oc8051_rom1.data_o [3]);
  not _20736_ (_12452_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nand _20737_ (_12453_, _07432_, _12452_);
  and _20738_ (_12454_, _12453_, _06444_);
  and _20739_ (_09949_, _12454_, _12451_);
  and _20740_ (_12455_, _09819_, _08679_);
  not _20741_ (_12456_, _12455_);
  or _20742_ (_12457_, _12456_, word_in[8]);
  and _20743_ (_12458_, _08866_, _08611_);
  not _20744_ (_12459_, _12458_);
  not _20745_ (_12460_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and _20746_ (_12461_, _09822_, _08819_);
  nor _20747_ (_12462_, _12461_, _12460_);
  and _20748_ (_12463_, _12461_, word_in[0]);
  or _20749_ (_12464_, _12463_, _12462_);
  or _20750_ (_12466_, _12464_, _12455_);
  and _20751_ (_12467_, _12466_, _12459_);
  and _20752_ (_12468_, _12467_, _12457_);
  and _20753_ (_12469_, _09835_, _08842_);
  and _20754_ (_12470_, _12458_, _09837_);
  or _20755_ (_12471_, _12470_, _12469_);
  or _20756_ (_12472_, _12471_, _12468_);
  not _20757_ (_12473_, _12469_);
  or _20758_ (_12474_, _12473_, word_in[24]);
  and _20759_ (_09955_, _12474_, _12472_);
  and _20760_ (_12475_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and _20761_ (_12476_, _12223_, \oc8051_top_1.oc8051_rom1.data_o [12]);
  or _20762_ (_12477_, _12476_, _12475_);
  and _20763_ (_09958_, _12477_, _06444_);
  not _20764_ (_12478_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  nor _20765_ (_12479_, _12461_, _12478_);
  and _20766_ (_12480_, _12461_, word_in[1]);
  nor _20767_ (_12481_, _12480_, _12479_);
  nor _20768_ (_12482_, _12481_, _12455_);
  and _20769_ (_12483_, _12455_, word_in[9]);
  or _20770_ (_12484_, _12483_, _12482_);
  and _20771_ (_12485_, _12484_, _12459_);
  and _20772_ (_12486_, _12458_, _09565_);
  or _20773_ (_12488_, _12486_, _12469_);
  or _20774_ (_12489_, _12488_, _12485_);
  or _20775_ (_12490_, _12473_, word_in[25]);
  and _20776_ (_09960_, _12490_, _12489_);
  or _20777_ (_12491_, _07432_, \oc8051_top_1.oc8051_rom1.data_o [8]);
  not _20778_ (_12492_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nand _20779_ (_12493_, _07432_, _12492_);
  and _20780_ (_12494_, _12493_, _06444_);
  and _20781_ (_09962_, _12494_, _12491_);
  not _20782_ (_12495_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  nor _20783_ (_12496_, _12461_, _12495_);
  and _20784_ (_12497_, _12461_, word_in[2]);
  nor _20785_ (_12498_, _12497_, _12496_);
  nor _20786_ (_12499_, _12498_, _12455_);
  and _20787_ (_12500_, _12455_, word_in[10]);
  or _20788_ (_12501_, _12500_, _12499_);
  and _20789_ (_12502_, _12501_, _12459_);
  and _20790_ (_12503_, _12458_, _10099_);
  or _20791_ (_12504_, _12503_, _12469_);
  or _20792_ (_12505_, _12504_, _12502_);
  or _20793_ (_12506_, _12473_, word_in[26]);
  and _20794_ (_09964_, _12506_, _12505_);
  and _20795_ (_12507_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and _20796_ (_12508_, _12223_, \oc8051_top_1.oc8051_rom1.data_o [22]);
  or _20797_ (_12509_, _12508_, _12507_);
  and _20798_ (_09967_, _12509_, _06444_);
  not _20799_ (_12510_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  nor _20800_ (_12511_, _12461_, _12510_);
  and _20801_ (_12512_, _12461_, word_in[3]);
  nor _20802_ (_12513_, _12512_, _12511_);
  nor _20803_ (_12514_, _12513_, _12455_);
  and _20804_ (_12515_, _12455_, word_in[11]);
  or _20805_ (_12516_, _12515_, _12514_);
  and _20806_ (_12517_, _12516_, _12459_);
  and _20807_ (_12518_, _12458_, _10116_);
  or _20808_ (_12519_, _12518_, _12469_);
  or _20809_ (_12520_, _12519_, _12517_);
  or _20810_ (_12521_, _12473_, word_in[27]);
  and _20811_ (_09969_, _12521_, _12520_);
  or _20812_ (_12522_, _07432_, \oc8051_top_1.oc8051_rom1.data_o [18]);
  nand _20813_ (_12523_, _07432_, _10712_);
  and _20814_ (_12524_, _12523_, _06444_);
  and _20815_ (_09972_, _12524_, _12522_);
  and _20816_ (_12525_, _12461_, word_in[4]);
  not _20817_ (_12526_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  nor _20818_ (_12527_, _12461_, _12526_);
  nor _20819_ (_12528_, _12527_, _12525_);
  nor _20820_ (_12529_, _12528_, _12455_);
  and _20821_ (_12530_, _12455_, word_in[12]);
  or _20822_ (_12531_, _12530_, _12529_);
  and _20823_ (_12532_, _12531_, _12459_);
  and _20824_ (_12533_, _12458_, _10020_);
  or _20825_ (_12534_, _12533_, _12469_);
  or _20826_ (_12535_, _12534_, _12532_);
  or _20827_ (_12536_, _12473_, word_in[28]);
  and _20828_ (_09974_, _12536_, _12535_);
  not _20829_ (_12537_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  nor _20830_ (_12538_, _12461_, _12537_);
  and _20831_ (_12539_, _12461_, word_in[5]);
  nor _20832_ (_12540_, _12539_, _12538_);
  nor _20833_ (_12541_, _12540_, _12455_);
  and _20834_ (_12542_, _12455_, word_in[13]);
  or _20835_ (_12543_, _12542_, _12541_);
  and _20836_ (_12544_, _12543_, _12459_);
  and _20837_ (_12545_, _12458_, _10149_);
  or _20838_ (_12546_, _12545_, _12469_);
  or _20839_ (_12547_, _12546_, _12544_);
  or _20840_ (_12548_, _12473_, word_in[29]);
  and _20841_ (_09976_, _12548_, _12547_);
  or _20842_ (_12549_, _07432_, \oc8051_top_1.oc8051_rom1.data_o [28]);
  nand _20843_ (_12550_, _07432_, _10708_);
  and _20844_ (_12551_, _12550_, _06444_);
  and _20845_ (_09979_, _12551_, _12549_);
  not _20846_ (_12552_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  nor _20847_ (_12553_, _12461_, _12552_);
  and _20848_ (_12554_, _12461_, word_in[6]);
  nor _20849_ (_12555_, _12554_, _12553_);
  nor _20850_ (_12556_, _12555_, _12455_);
  and _20851_ (_12557_, _12455_, word_in[14]);
  or _20852_ (_12558_, _12557_, _12556_);
  and _20853_ (_12559_, _12558_, _12459_);
  and _20854_ (_12560_, _12458_, _10154_);
  or _20855_ (_12561_, _12560_, _12469_);
  or _20856_ (_12562_, _12561_, _12559_);
  or _20857_ (_12563_, _12473_, word_in[30]);
  and _20858_ (_09981_, _12563_, _12562_);
  nor _20859_ (_12564_, _12461_, _08680_);
  and _20860_ (_12565_, _12461_, word_in[7]);
  nor _20861_ (_12566_, _12565_, _12564_);
  nor _20862_ (_12567_, _12566_, _12455_);
  and _20863_ (_12568_, _12455_, word_in[15]);
  or _20864_ (_12569_, _12568_, _12567_);
  and _20865_ (_12570_, _12569_, _12459_);
  and _20866_ (_12571_, _12458_, _08886_);
  or _20867_ (_12572_, _12571_, _12469_);
  or _20868_ (_12573_, _12572_, _12570_);
  or _20869_ (_12574_, _12473_, word_in[31]);
  and _20870_ (_09983_, _12574_, _12573_);
  nor _20871_ (_09996_, _11830_, rst);
  and _20872_ (_12575_, _12048_, _08127_);
  and _20873_ (_12576_, _11452_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor _20874_ (_12577_, _12106_, _12033_);
  and _20875_ (_12578_, _12054_, _11726_);
  or _20876_ (_12579_, _12578_, _12577_);
  or _20877_ (_12580_, _12579_, _12576_);
  or _20878_ (_12581_, _12110_, _12109_);
  and _20879_ (_12582_, _12581_, _12209_);
  nor _20880_ (_12583_, _12581_, _12209_);
  or _20881_ (_12584_, _12583_, _12582_);
  and _20882_ (_12585_, _12584_, _12218_);
  nor _20883_ (_12586_, _12585_, _12580_);
  nand _20884_ (_12587_, _12586_, _12023_);
  or _20885_ (_12588_, _12587_, _12575_);
  and _20886_ (_12589_, _10949_, _08483_);
  nor _20887_ (_12590_, _12589_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor _20888_ (_12591_, _12590_, _12226_);
  or _20889_ (_12592_, _12591_, _12023_);
  and _20890_ (_12593_, _12592_, _06444_);
  and _20891_ (_10009_, _12593_, _12588_);
  or _20892_ (_12594_, _12023_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and _20893_ (_12595_, _12594_, _06444_);
  and _20894_ (_12596_, _12048_, _08019_);
  and _20895_ (_12597_, _11452_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and _20896_ (_12598_, _12032_, _12191_);
  and _20897_ (_12600_, _12054_, _11848_);
  or _20898_ (_12601_, _12600_, _12598_);
  or _20899_ (_12602_, _12601_, _12597_);
  or _20900_ (_12603_, _12193_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  not _20901_ (_12604_, _12194_);
  or _20902_ (_12605_, _12045_, _12034_);
  and _20903_ (_12606_, _12605_, _12052_);
  and _20904_ (_12607_, _12606_, _12604_);
  and _20905_ (_12608_, _12607_, _12603_);
  or _20906_ (_12609_, _12608_, _12602_);
  nor _20907_ (_12610_, _12609_, _12596_);
  nand _20908_ (_12611_, _12610_, _12023_);
  and _20909_ (_10012_, _12611_, _12595_);
  and _20910_ (_12612_, _12227_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and _20911_ (_12613_, _12612_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and _20912_ (_12614_, _12613_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and _20913_ (_12615_, _12614_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and _20914_ (_12616_, _12615_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  or _20915_ (_12617_, _12616_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nand _20916_ (_12618_, _12616_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and _20917_ (_12619_, _12618_, _12617_);
  or _20918_ (_12620_, _12619_, _12023_);
  and _20919_ (_12621_, _12620_, _06444_);
  and _20920_ (_12622_, _11452_, _08230_);
  and _20921_ (_12623_, _12026_, _08267_);
  and _20922_ (_12624_, _11650_, _12032_);
  and _20923_ (_12625_, _12047_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  or _20924_ (_12626_, _12625_, _12624_);
  or _20925_ (_12627_, _12626_, _12623_);
  or _20926_ (_12628_, _12627_, _12622_);
  and _20927_ (_12629_, _12079_, _08376_);
  and _20928_ (_12630_, _07429_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  and _20929_ (_12631_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and _20930_ (_12632_, _07254_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  not _20931_ (_12633_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor _20932_ (_12634_, _07241_, _12633_);
  nor _20933_ (_12635_, _12634_, _12632_);
  and _20934_ (_12636_, _07248_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and _20935_ (_12637_, _07238_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor _20936_ (_12638_, _12637_, _12636_);
  and _20937_ (_12639_, _12638_, _12635_);
  and _20938_ (_12640_, _07246_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and _20939_ (_12641_, _07251_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor _20940_ (_12643_, _12641_, _12640_);
  and _20941_ (_12644_, _12643_, _12639_);
  nor _20942_ (_12645_, _12644_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _20943_ (_12646_, _12645_, _12631_);
  nor _20944_ (_12647_, _12646_, _07429_);
  nor _20945_ (_12648_, _12647_, _12630_);
  and _20946_ (_12649_, _12648_, _12038_);
  nor _20947_ (_12650_, _12649_, _12629_);
  and _20948_ (_12651_, _12650_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor _20949_ (_12652_, _12650_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor _20950_ (_12653_, _12652_, _12651_);
  or _20951_ (_12654_, _12212_, _12084_);
  and _20952_ (_12655_, _12654_, _12653_);
  or _20953_ (_12656_, _12655_, _12651_);
  or _20954_ (_12657_, _12656_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  or _20955_ (_12658_, _12657_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  or _20956_ (_12659_, _12658_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  or _20957_ (_12660_, _12659_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nand _20958_ (_12661_, _12660_, _12650_);
  not _20959_ (_12662_, _12650_);
  and _20960_ (_12663_, \oc8051_top_1.oc8051_memory_interface1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and _20961_ (_12664_, _12663_, _12656_);
  and _20962_ (_12665_, _12664_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  nand _20963_ (_12666_, _12665_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nand _20964_ (_12667_, _12666_, _12662_);
  nand _20965_ (_12668_, _12667_, _12661_);
  nand _20966_ (_12669_, _12668_, _08150_);
  or _20967_ (_12670_, _12668_, _08150_);
  and _20968_ (_12671_, _12670_, _12669_);
  and _20969_ (_12672_, _12671_, _12218_);
  or _20970_ (_12673_, _12672_, _12628_);
  and _20971_ (_12674_, \oc8051_top_1.oc8051_memory_interface1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and _20972_ (_12675_, \oc8051_top_1.oc8051_memory_interface1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and _20973_ (_12676_, _12675_, _12674_);
  and _20974_ (_12677_, \oc8051_top_1.oc8051_memory_interface1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and _20975_ (_12678_, \oc8051_top_1.oc8051_memory_interface1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and _20976_ (_12679_, _12678_, _12663_);
  and _20977_ (_12680_, _12679_, _12677_);
  and _20978_ (_12681_, _12680_, _12676_);
  and _20979_ (_12682_, _12681_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _20980_ (_12683_, _12682_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor _20981_ (_12684_, _12682_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor _20982_ (_12685_, _12684_, _12683_);
  nand _20983_ (_12686_, _12685_, _12054_);
  nand _20984_ (_12687_, _12686_, _12023_);
  or _20985_ (_12688_, _12687_, _12673_);
  and _20986_ (_10017_, _12688_, _12621_);
  or _20987_ (_12689_, _10963_, _10957_);
  and _20988_ (_12690_, _12689_, _10964_);
  or _20989_ (_12691_, _12690_, _08374_);
  or _20990_ (_12692_, _08373_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and _20991_ (_12693_, _12692_, _10894_);
  and _20992_ (_12694_, _12693_, _12691_);
  and _20993_ (_12695_, _10976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  or _20994_ (_10025_, _12695_, _12694_);
  nor _20995_ (_12696_, _10947_, _10933_);
  nor _20996_ (_12697_, _12696_, _10948_);
  or _20997_ (_12698_, _12697_, _08374_);
  or _20998_ (_12699_, _08373_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and _20999_ (_12700_, _12699_, _10894_);
  and _21000_ (_12701_, _12700_, _12698_);
  and _21001_ (_12702_, _10976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  or _21002_ (_10029_, _12702_, _12701_);
  and _21003_ (_12703_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _06444_);
  not _21004_ (_12704_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  nor _21005_ (_12705_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  nor _21006_ (_12706_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and _21007_ (_12707_, _12706_, _12705_);
  not _21008_ (_12708_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  nor _21009_ (_12709_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and _21010_ (_12710_, _12709_, _12708_);
  and _21011_ (_12711_, _12710_, _12707_);
  and _21012_ (_12712_, _12711_, _12704_);
  and _21013_ (_12713_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _06444_);
  and _21014_ (_12714_, _12713_, _12712_);
  or _21015_ (_10037_, _12714_, _12703_);
  and _21016_ (_12715_, _09554_, _08859_);
  and _21017_ (_12716_, _08878_, word_in[0]);
  not _21018_ (_12717_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  nor _21019_ (_12718_, _08878_, _12717_);
  nor _21020_ (_12719_, _12718_, _12716_);
  nor _21021_ (_12720_, _12719_, _08871_);
  and _21022_ (_12721_, _08871_, word_in[8]);
  or _21023_ (_12722_, _12721_, _12720_);
  and _21024_ (_12723_, _12722_, _08868_);
  and _21025_ (_12724_, _09837_, _08867_);
  or _21026_ (_12725_, _12724_, _12723_);
  and _21027_ (_12726_, _12725_, _08862_);
  or _21028_ (_14572_, _12726_, _12715_);
  nor _21029_ (_10040_, _11725_, rst);
  and _21030_ (_12727_, _11261_, _08859_);
  and _21031_ (_12728_, _08878_, word_in[1]);
  not _21032_ (_12729_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  nor _21033_ (_12730_, _08878_, _12729_);
  nor _21034_ (_12731_, _12730_, _12728_);
  nor _21035_ (_12732_, _12731_, _08871_);
  and _21036_ (_12733_, _08871_, word_in[9]);
  or _21037_ (_12734_, _12733_, _12732_);
  and _21038_ (_12735_, _12734_, _08868_);
  and _21039_ (_12736_, _09565_, _08867_);
  or _21040_ (_12737_, _12736_, _12735_);
  and _21041_ (_12738_, _12737_, _08862_);
  or _21042_ (_14573_, _12738_, _12727_);
  and _21043_ (_12739_, _09582_, _08859_);
  and _21044_ (_12740_, _08878_, word_in[2]);
  not _21045_ (_12741_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  nor _21046_ (_12742_, _08878_, _12741_);
  nor _21047_ (_12743_, _12742_, _12740_);
  nor _21048_ (_12744_, _12743_, _08871_);
  and _21049_ (_12745_, _08871_, word_in[10]);
  or _21050_ (_12746_, _12745_, _12744_);
  and _21051_ (_12747_, _12746_, _08868_);
  and _21052_ (_12748_, _10099_, _08867_);
  or _21053_ (_12750_, _12748_, _12747_);
  and _21054_ (_12751_, _12750_, _08862_);
  or _21055_ (_14574_, _12751_, _12739_);
  and _21056_ (_12753_, _08878_, word_in[3]);
  not _21057_ (_12754_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  nor _21058_ (_12755_, _08878_, _12754_);
  nor _21059_ (_12756_, _12755_, _12753_);
  nor _21060_ (_12757_, _12756_, _08871_);
  and _21061_ (_12758_, _08871_, word_in[11]);
  or _21062_ (_12759_, _12758_, _12757_);
  and _21063_ (_12760_, _12759_, _08868_);
  and _21064_ (_12761_, _10116_, _08867_);
  or _21065_ (_12762_, _12761_, _12760_);
  and _21066_ (_12763_, _12762_, _08862_);
  and _21067_ (_12764_, _08859_, word_in[27]);
  or _21068_ (_14575_, _12764_, _12763_);
  and _21069_ (_12765_, _08878_, word_in[4]);
  not _21070_ (_12766_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  nor _21071_ (_12767_, _08878_, _12766_);
  nor _21072_ (_12768_, _12767_, _12765_);
  nor _21073_ (_12770_, _12768_, _08871_);
  and _21074_ (_12771_, _08871_, word_in[12]);
  or _21075_ (_12772_, _12771_, _12770_);
  and _21076_ (_12773_, _12772_, _08868_);
  and _21077_ (_12774_, _10020_, _08867_);
  or _21078_ (_12775_, _12774_, _12773_);
  and _21079_ (_12776_, _12775_, _08862_);
  and _21080_ (_12777_, _08859_, word_in[28]);
  or _21081_ (_14576_, _12777_, _12776_);
  and _21082_ (_12778_, _08878_, word_in[5]);
  not _21083_ (_12779_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  nor _21084_ (_12780_, _08878_, _12779_);
  nor _21085_ (_12781_, _12780_, _12778_);
  nor _21086_ (_12782_, _12781_, _08871_);
  and _21087_ (_12783_, _08871_, word_in[13]);
  or _21088_ (_12784_, _12783_, _12782_);
  and _21089_ (_12785_, _12784_, _08868_);
  and _21090_ (_12786_, _10149_, _08867_);
  or _21091_ (_12787_, _12786_, _12785_);
  and _21092_ (_12788_, _12787_, _08862_);
  and _21093_ (_12789_, _08859_, word_in[29]);
  or _21094_ (_14577_, _12789_, _12788_);
  and _21095_ (_12790_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], _08478_);
  and _21096_ (_12791_, \oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or _21097_ (_12792_, _12791_, _12790_);
  and _21098_ (_10053_, _12792_, _06444_);
  and _21099_ (_12793_, _08878_, word_in[6]);
  not _21100_ (_12794_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  nor _21101_ (_12795_, _08878_, _12794_);
  nor _21102_ (_12796_, _12795_, _12793_);
  nor _21103_ (_12797_, _12796_, _08871_);
  and _21104_ (_12798_, _08871_, word_in[14]);
  or _21105_ (_12799_, _12798_, _12797_);
  and _21106_ (_12800_, _12799_, _08868_);
  and _21107_ (_12801_, _10154_, _08867_);
  or _21108_ (_12802_, _12801_, _12800_);
  and _21109_ (_12803_, _12802_, _08862_);
  and _21110_ (_12804_, _08859_, word_in[30]);
  or _21111_ (_14578_, _12804_, _12803_);
  and _21112_ (_12805_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  nor _21113_ (_12806_, _07432_, _11044_);
  or _21114_ (_12807_, _12806_, _12805_);
  and _21115_ (_10345_, _12807_, _06444_);
  or _21116_ (_12808_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  nand _21117_ (_12809_, _07432_, _11220_);
  and _21118_ (_12810_, _12809_, _06444_);
  and _21119_ (_10354_, _12810_, _12808_);
  and _21120_ (_12811_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  not _21121_ (_12812_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor _21122_ (_12813_, _07432_, _12812_);
  or _21123_ (_12814_, _12813_, _12811_);
  and _21124_ (_10357_, _12814_, _06444_);
  or _21125_ (_12815_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  nand _21126_ (_12816_, _07432_, _12137_);
  and _21127_ (_12817_, _12816_, _06444_);
  and _21128_ (_10362_, _12817_, _12815_);
  or _21129_ (_12818_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  nand _21130_ (_12819_, _07432_, _10728_);
  and _21131_ (_12820_, _12819_, _06444_);
  and _21132_ (_10364_, _12820_, _12818_);
  nor _21133_ (_12821_, _06299_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  nor _21134_ (_12822_, _12821_, _08473_);
  and _21135_ (_10468_, _12822_, _06443_);
  and _21136_ (_10560_, t2_i, _06444_);
  not _21137_ (_12823_, _07159_);
  and _21138_ (_12824_, _09331_, _12823_);
  or _21139_ (_12825_, _12824_, _07158_);
  and _21140_ (_12826_, _12825_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  nand _21141_ (_12827_, _06439_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  nor _21142_ (_12828_, _12827_, _07415_);
  and _21143_ (_12829_, _07416_, _06439_);
  not _21144_ (_12830_, _12829_);
  nor _21145_ (_12831_, _12830_, _11589_);
  or _21146_ (_12832_, _12831_, _12828_);
  or _21147_ (_12833_, _12832_, _12826_);
  and _21148_ (_10727_, _12833_, _06444_);
  not _21149_ (_12834_, _12824_);
  nor _21150_ (_12835_, _07156_, _12834_);
  nand _21151_ (_12836_, _07415_, _06439_);
  or _21152_ (_12837_, _12836_, _12835_);
  and _21153_ (_12838_, _12837_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  nand _21154_ (_12839_, _06439_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  nor _21155_ (_12840_, _12839_, _07418_);
  nor _21156_ (_12841_, _09526_, _07158_);
  and _21157_ (_12842_, _12841_, _07044_);
  or _21158_ (_12843_, _12842_, _12840_);
  or _21159_ (_12844_, _12843_, _12838_);
  and _21160_ (_10802_, _12844_, _06444_);
  and _21161_ (_12845_, _08064_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  not _21162_ (_12846_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nor _21163_ (_12847_, _08064_, _12846_);
  or _21164_ (_12848_, _12847_, _12845_);
  and _21165_ (_10809_, _12848_, _06444_);
  nor _21166_ (_12849_, _11589_, _06449_);
  and _21167_ (_12850_, _06449_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  or _21168_ (_12851_, _12850_, _12849_);
  and _21169_ (_10905_, _12851_, _06444_);
  or _21170_ (_12852_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  nand _21171_ (_12853_, _07432_, _12092_);
  and _21172_ (_12854_, _12853_, _06444_);
  and _21173_ (_10922_, _12854_, _12852_);
  and _21174_ (_12855_, _08558_, word_in[0]);
  nand _21175_ (_12856_, _08480_, _11230_);
  or _21176_ (_12857_, _08480_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and _21177_ (_12858_, _12857_, _12856_);
  and _21178_ (_12859_, _12858_, _08506_);
  nand _21179_ (_12860_, _08480_, _12347_);
  or _21180_ (_12861_, _08480_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  and _21181_ (_12862_, _12861_, _12860_);
  and _21182_ (_12863_, _12862_, _08503_);
  nand _21183_ (_12865_, _08480_, _10608_);
  or _21184_ (_12866_, _08480_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  and _21185_ (_12867_, _12866_, _12865_);
  and _21186_ (_12868_, _12867_, _08523_);
  or _21187_ (_12869_, _12868_, _12863_);
  or _21188_ (_12871_, _12869_, _12859_);
  nand _21189_ (_12872_, _08480_, _12717_);
  or _21190_ (_12873_, _08480_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and _21191_ (_12874_, _12873_, _12872_);
  and _21192_ (_12875_, _12874_, _08513_);
  or _21193_ (_12876_, _12875_, _08532_);
  or _21194_ (_12877_, _12876_, _12871_);
  nand _21195_ (_12878_, _08480_, _09941_);
  or _21196_ (_12879_, _08480_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  and _21197_ (_12880_, _12879_, _12878_);
  and _21198_ (_12881_, _12880_, _08506_);
  nand _21199_ (_12882_, _08480_, _09697_);
  or _21200_ (_12883_, _08480_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  and _21201_ (_12884_, _12883_, _12882_);
  and _21202_ (_12885_, _12884_, _08523_);
  nand _21203_ (_12886_, _08480_, _10183_);
  or _21204_ (_12887_, _08480_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  and _21205_ (_12888_, _12887_, _12886_);
  and _21206_ (_12890_, _12888_, _08503_);
  or _21207_ (_12891_, _12890_, _12885_);
  or _21208_ (_12892_, _12891_, _12881_);
  nand _21209_ (_12893_, _08480_, _10396_);
  or _21210_ (_12894_, _08480_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  and _21211_ (_12895_, _12894_, _12893_);
  and _21212_ (_12896_, _12895_, _08513_);
  or _21213_ (_12897_, _12896_, _08489_);
  or _21214_ (_12898_, _12897_, _12892_);
  and _21215_ (_12899_, _12898_, _12877_);
  and _21216_ (_12900_, _12899_, _08557_);
  or _21217_ (\oc8051_symbolic_cxrom1.cxrom_data_out [0], _12900_, _12855_);
  and _21218_ (_12901_, _08558_, word_in[1]);
  nand _21219_ (_12902_, _08480_, _10624_);
  or _21220_ (_12903_, _08480_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  and _21221_ (_12904_, _12903_, _12902_);
  and _21222_ (_12905_, _12904_, _08523_);
  nand _21223_ (_12906_, _08480_, _11249_);
  or _21224_ (_12907_, _08480_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  and _21225_ (_12908_, _12907_, _12906_);
  and _21226_ (_12909_, _12908_, _08506_);
  nand _21227_ (_12910_, _08480_, _12365_);
  or _21228_ (_12911_, _08480_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  and _21229_ (_12912_, _12911_, _12910_);
  and _21230_ (_12913_, _12912_, _08503_);
  or _21231_ (_12914_, _12913_, _12909_);
  or _21232_ (_12915_, _12914_, _12905_);
  nand _21233_ (_12916_, _08480_, _12729_);
  or _21234_ (_12917_, _08480_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  and _21235_ (_12918_, _12917_, _12916_);
  and _21236_ (_12919_, _12918_, _08513_);
  or _21237_ (_12920_, _12919_, _08532_);
  or _21238_ (_12921_, _12920_, _12915_);
  nand _21239_ (_12922_, _08480_, _09720_);
  or _21240_ (_12923_, _08480_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  and _21241_ (_12924_, _12923_, _12922_);
  and _21242_ (_12925_, _12924_, _08523_);
  nand _21243_ (_12926_, _08480_, _09963_);
  or _21244_ (_12927_, _08480_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  and _21245_ (_12928_, _12927_, _12926_);
  and _21246_ (_12929_, _12928_, _08506_);
  nand _21247_ (_12930_, _08480_, _10197_);
  or _21248_ (_12931_, _08480_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  and _21249_ (_12932_, _12931_, _12930_);
  and _21250_ (_12933_, _12932_, _08503_);
  or _21251_ (_12934_, _12933_, _12929_);
  or _21252_ (_12935_, _12934_, _12925_);
  nand _21253_ (_12936_, _08480_, _10406_);
  or _21254_ (_12937_, _08480_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  and _21255_ (_12938_, _12937_, _12936_);
  and _21256_ (_12939_, _12938_, _08513_);
  or _21257_ (_12940_, _12939_, _08489_);
  or _21258_ (_12941_, _12940_, _12935_);
  and _21259_ (_12942_, _12941_, _12921_);
  and _21260_ (_12943_, _12942_, _08557_);
  or _21261_ (\oc8051_symbolic_cxrom1.cxrom_data_out [1], _12943_, _12901_);
  and _21262_ (_12944_, _08558_, word_in[2]);
  nand _21263_ (_12945_, _08480_, _10636_);
  or _21264_ (_12946_, _08480_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  and _21265_ (_12947_, _12946_, _12945_);
  and _21266_ (_12948_, _12947_, _08523_);
  nand _21267_ (_12949_, _08480_, _11267_);
  or _21268_ (_12950_, _08480_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  and _21269_ (_12951_, _12950_, _12949_);
  and _21270_ (_12952_, _12951_, _08506_);
  nand _21271_ (_12953_, _08480_, _12378_);
  or _21272_ (_12954_, _08480_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  and _21273_ (_12955_, _12954_, _12953_);
  and _21274_ (_12956_, _12955_, _08503_);
  or _21275_ (_12957_, _12956_, _12952_);
  or _21276_ (_12958_, _12957_, _12948_);
  nand _21277_ (_12959_, _08480_, _12741_);
  or _21278_ (_12960_, _08480_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  and _21279_ (_12961_, _12960_, _12959_);
  and _21280_ (_12962_, _12961_, _08513_);
  or _21281_ (_12963_, _12962_, _08532_);
  or _21282_ (_12964_, _12963_, _12958_);
  nand _21283_ (_12965_, _08480_, _09734_);
  or _21284_ (_12966_, _08480_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  and _21285_ (_12967_, _12966_, _12965_);
  and _21286_ (_12968_, _12967_, _08523_);
  nand _21287_ (_12969_, _08480_, _09985_);
  or _21288_ (_12970_, _08480_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  and _21289_ (_12971_, _12970_, _12969_);
  and _21290_ (_12972_, _12971_, _08506_);
  nand _21291_ (_12973_, _08480_, _10209_);
  or _21292_ (_12974_, _08480_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  and _21293_ (_12975_, _12974_, _12973_);
  and _21294_ (_12976_, _12975_, _08503_);
  or _21295_ (_12977_, _12976_, _12972_);
  or _21296_ (_12978_, _12977_, _12968_);
  nand _21297_ (_12979_, _08480_, _10420_);
  or _21298_ (_12980_, _08480_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  and _21299_ (_12981_, _12980_, _12979_);
  and _21300_ (_12982_, _12981_, _08513_);
  or _21301_ (_12983_, _12982_, _08489_);
  or _21302_ (_12984_, _12983_, _12978_);
  and _21303_ (_12985_, _12984_, _12964_);
  and _21304_ (_12986_, _12985_, _08557_);
  or _21305_ (\oc8051_symbolic_cxrom1.cxrom_data_out [2], _12986_, _12944_);
  and _21306_ (_12987_, _08558_, word_in[3]);
  nand _21307_ (_12988_, _08480_, _10649_);
  or _21308_ (_12989_, _08480_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  and _21309_ (_12990_, _12989_, _12988_);
  and _21310_ (_12991_, _12990_, _08523_);
  nand _21311_ (_12992_, _08480_, _11279_);
  or _21312_ (_12993_, _08480_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  and _21313_ (_12994_, _12993_, _12992_);
  and _21314_ (_12995_, _12994_, _08506_);
  nand _21315_ (_12996_, _08480_, _12391_);
  or _21316_ (_12997_, _08480_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  and _21317_ (_12998_, _12997_, _12996_);
  and _21318_ (_12999_, _12998_, _08503_);
  or _21319_ (_13000_, _12999_, _12995_);
  or _21320_ (_13001_, _13000_, _12991_);
  nand _21321_ (_13002_, _08480_, _12754_);
  or _21322_ (_13003_, _08480_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  and _21323_ (_13004_, _13003_, _13002_);
  and _21324_ (_13005_, _13004_, _08513_);
  or _21325_ (_13006_, _13005_, _08532_);
  or _21326_ (_13007_, _13006_, _13001_);
  nand _21327_ (_13008_, _08480_, _09749_);
  or _21328_ (_13009_, _08480_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  and _21329_ (_13010_, _13009_, _13008_);
  and _21330_ (_13012_, _13010_, _08523_);
  nand _21331_ (_13013_, _08480_, _09998_);
  or _21332_ (_13014_, _08480_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  and _21333_ (_13015_, _13014_, _13013_);
  and _21334_ (_13016_, _13015_, _08506_);
  nand _21335_ (_13017_, _08480_, _10221_);
  or _21336_ (_13018_, _08480_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  and _21337_ (_13019_, _13018_, _13017_);
  and _21338_ (_13020_, _13019_, _08503_);
  or _21339_ (_13021_, _13020_, _13016_);
  or _21340_ (_13022_, _13021_, _13012_);
  nand _21341_ (_13024_, _08480_, _10431_);
  or _21342_ (_13025_, _08480_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  and _21343_ (_13026_, _13025_, _13024_);
  and _21344_ (_13027_, _13026_, _08513_);
  or _21345_ (_13028_, _13027_, _08489_);
  or _21346_ (_13029_, _13028_, _13022_);
  and _21347_ (_13030_, _13029_, _13007_);
  and _21348_ (_13031_, _13030_, _08557_);
  or _21349_ (\oc8051_symbolic_cxrom1.cxrom_data_out [3], _13031_, _12987_);
  and _21350_ (_13032_, _08558_, word_in[4]);
  nand _21351_ (_13033_, _08480_, _10660_);
  or _21352_ (_13034_, _08480_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  and _21353_ (_13035_, _13034_, _13033_);
  and _21354_ (_13036_, _13035_, _08523_);
  nand _21355_ (_13037_, _08480_, _11292_);
  or _21356_ (_13039_, _08480_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  and _21357_ (_13040_, _13039_, _13037_);
  and _21358_ (_13041_, _13040_, _08506_);
  nand _21359_ (_13042_, _08480_, _12403_);
  or _21360_ (_13043_, _08480_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  and _21361_ (_13044_, _13043_, _13042_);
  and _21362_ (_13045_, _13044_, _08503_);
  or _21363_ (_13047_, _13045_, _13041_);
  or _21364_ (_13048_, _13047_, _13036_);
  nand _21365_ (_13049_, _08480_, _12766_);
  or _21366_ (_13051_, _08480_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  and _21367_ (_13052_, _13051_, _13049_);
  and _21368_ (_13053_, _13052_, _08513_);
  or _21369_ (_13054_, _13053_, _08532_);
  or _21370_ (_13055_, _13054_, _13048_);
  nand _21371_ (_13056_, _08480_, _09761_);
  or _21372_ (_13057_, _08480_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  and _21373_ (_13058_, _13057_, _13056_);
  and _21374_ (_13059_, _13058_, _08523_);
  nand _21375_ (_13060_, _08480_, _10011_);
  or _21376_ (_13061_, _08480_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  and _21377_ (_13062_, _13061_, _13060_);
  and _21378_ (_13063_, _13062_, _08506_);
  nand _21379_ (_13064_, _08480_, _10233_);
  or _21380_ (_13065_, _08480_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  and _21381_ (_13066_, _13065_, _13064_);
  and _21382_ (_13067_, _13066_, _08503_);
  or _21383_ (_13068_, _13067_, _13063_);
  or _21384_ (_13069_, _13068_, _13059_);
  nand _21385_ (_13070_, _08480_, _10443_);
  or _21386_ (_13071_, _08480_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  and _21387_ (_13072_, _13071_, _13070_);
  and _21388_ (_13073_, _13072_, _08513_);
  or _21389_ (_13074_, _13073_, _08489_);
  or _21390_ (_13075_, _13074_, _13069_);
  and _21391_ (_13076_, _13075_, _13055_);
  and _21392_ (_13077_, _13076_, _08557_);
  or _21393_ (\oc8051_symbolic_cxrom1.cxrom_data_out [4], _13077_, _13032_);
  and _21394_ (_13079_, _08558_, word_in[5]);
  nand _21395_ (_13080_, _08480_, _10672_);
  or _21396_ (_13081_, _08480_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  and _21397_ (_13082_, _13081_, _13080_);
  and _21398_ (_13083_, _13082_, _08523_);
  nand _21399_ (_13084_, _08480_, _11305_);
  or _21400_ (_13085_, _08480_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  and _21401_ (_13086_, _13085_, _13084_);
  and _21402_ (_13087_, _13086_, _08506_);
  nand _21403_ (_13088_, _08480_, _12416_);
  or _21404_ (_13089_, _08480_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  and _21405_ (_13090_, _13089_, _13088_);
  and _21406_ (_13091_, _13090_, _08503_);
  or _21407_ (_13092_, _13091_, _13087_);
  or _21408_ (_13093_, _13092_, _13083_);
  nand _21409_ (_13094_, _08480_, _12779_);
  or _21410_ (_13095_, _08480_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  and _21411_ (_13096_, _13095_, _13094_);
  and _21412_ (_13097_, _13096_, _08513_);
  or _21413_ (_13098_, _13097_, _08532_);
  or _21414_ (_13099_, _13098_, _13093_);
  nand _21415_ (_13100_, _08480_, _09775_);
  or _21416_ (_13101_, _08480_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  and _21417_ (_13102_, _13101_, _13100_);
  and _21418_ (_13103_, _13102_, _08523_);
  nand _21419_ (_13104_, _08480_, _10027_);
  or _21420_ (_13105_, _08480_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  and _21421_ (_13106_, _13105_, _13104_);
  and _21422_ (_13107_, _13106_, _08506_);
  nand _21423_ (_13109_, _08480_, _10245_);
  or _21424_ (_13110_, _08480_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  and _21425_ (_13111_, _13110_, _13109_);
  and _21426_ (_13112_, _13111_, _08503_);
  or _21427_ (_13113_, _13112_, _13107_);
  or _21428_ (_13114_, _13113_, _13103_);
  nand _21429_ (_13115_, _08480_, _10454_);
  or _21430_ (_13116_, _08480_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  and _21431_ (_13117_, _13116_, _13115_);
  and _21432_ (_13118_, _13117_, _08513_);
  or _21433_ (_13119_, _13118_, _08489_);
  or _21434_ (_13120_, _13119_, _13114_);
  and _21435_ (_13121_, _13120_, _13099_);
  and _21436_ (_13122_, _13121_, _08557_);
  or _21437_ (\oc8051_symbolic_cxrom1.cxrom_data_out [5], _13122_, _13079_);
  and _21438_ (_13123_, _08558_, word_in[6]);
  nand _21439_ (_13124_, _08480_, _11318_);
  or _21440_ (_13125_, _08480_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  and _21441_ (_13126_, _13125_, _13124_);
  and _21442_ (_13127_, _13126_, _08506_);
  nand _21443_ (_13128_, _08480_, _12429_);
  or _21444_ (_13129_, _08480_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  and _21445_ (_13130_, _13129_, _13128_);
  and _21446_ (_13131_, _13130_, _08503_);
  nand _21447_ (_13132_, _08480_, _10685_);
  or _21448_ (_13133_, _08480_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  and _21449_ (_13134_, _13133_, _13132_);
  and _21450_ (_13135_, _13134_, _08523_);
  or _21451_ (_13136_, _13135_, _13131_);
  or _21452_ (_13137_, _13136_, _13127_);
  nand _21453_ (_13139_, _08480_, _12794_);
  or _21454_ (_13140_, _08480_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  and _21455_ (_13141_, _13140_, _13139_);
  and _21456_ (_13142_, _13141_, _08513_);
  or _21457_ (_13143_, _13142_, _08532_);
  or _21458_ (_13144_, _13143_, _13137_);
  nand _21459_ (_13145_, _08480_, _10042_);
  or _21460_ (_13146_, _08480_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  and _21461_ (_13147_, _13146_, _13145_);
  and _21462_ (_13149_, _13147_, _08506_);
  nand _21463_ (_13151_, _08480_, _09792_);
  or _21464_ (_13152_, _08480_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  and _21465_ (_13153_, _13152_, _13151_);
  and _21466_ (_13154_, _13153_, _08523_);
  nand _21467_ (_13155_, _08480_, _10258_);
  or _21468_ (_13156_, _08480_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  and _21469_ (_13157_, _13156_, _13155_);
  and _21470_ (_13158_, _13157_, _08503_);
  or _21471_ (_13159_, _13158_, _13154_);
  or _21472_ (_13160_, _13159_, _13149_);
  nand _21473_ (_13162_, _08480_, _10469_);
  or _21474_ (_13163_, _08480_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  and _21475_ (_13164_, _13163_, _13162_);
  and _21476_ (_13165_, _13164_, _08513_);
  or _21477_ (_13166_, _13165_, _08489_);
  or _21478_ (_13167_, _13166_, _13160_);
  and _21479_ (_13168_, _13167_, _13144_);
  and _21480_ (_13169_, _13168_, _08557_);
  or _21481_ (\oc8051_symbolic_cxrom1.cxrom_data_out [6], _13169_, _13123_);
  and _21482_ (_13170_, _08664_, word_in[8]);
  nand _21483_ (_13171_, _08480_, _10998_);
  or _21484_ (_13172_, _08480_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and _21485_ (_13173_, _13172_, _13171_);
  and _21486_ (_13174_, _13173_, _08666_);
  nand _21487_ (_13175_, _08480_, _10504_);
  or _21488_ (_13176_, _08480_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  and _21489_ (_13177_, _13176_, _13175_);
  and _21490_ (_13178_, _13177_, _08665_);
  or _21491_ (_13179_, _13178_, _13174_);
  and _21492_ (_13180_, _13179_, _08623_);
  nand _21493_ (_13181_, _08480_, _12460_);
  or _21494_ (_13182_, _08480_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  and _21495_ (_13183_, _13182_, _13181_);
  and _21496_ (_13184_, _13183_, _08666_);
  nand _21497_ (_13185_, _08480_, _12240_);
  or _21498_ (_13186_, _08480_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  and _21499_ (_13187_, _13186_, _13185_);
  and _21500_ (_13188_, _13187_, _08665_);
  or _21501_ (_13189_, _13188_, _13184_);
  and _21502_ (_13190_, _13189_, _08679_);
  nand _21503_ (_13191_, _08480_, _10290_);
  or _21504_ (_13192_, _08480_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  and _21505_ (_13193_, _13192_, _13191_);
  and _21506_ (_13194_, _13193_, _08666_);
  nand _21507_ (_13195_, _08480_, _10068_);
  or _21508_ (_13196_, _08480_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  and _21509_ (_13197_, _13196_, _13195_);
  and _21510_ (_13198_, _13197_, _08665_);
  or _21511_ (_13199_, _13198_, _13194_);
  and _21512_ (_13200_, _13199_, _08708_);
  nand _21513_ (_13201_, _08480_, _09821_);
  or _21514_ (_13202_, _08480_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  and _21515_ (_13203_, _13202_, _13201_);
  and _21516_ (_13204_, _13203_, _08666_);
  and _21517_ (_13205_, _08480_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  nor _21518_ (_13206_, _08480_, _09697_);
  or _21519_ (_13207_, _13206_, _13205_);
  and _21520_ (_13208_, _13207_, _08665_);
  or _21521_ (_13209_, _13208_, _13204_);
  and _21522_ (_13210_, _13209_, _08626_);
  or _21523_ (_13211_, _13210_, _13200_);
  or _21524_ (_13212_, _13211_, _13190_);
  nor _21525_ (_13213_, _13212_, _13180_);
  nor _21526_ (_13214_, _13213_, _08664_);
  or _21527_ (\oc8051_symbolic_cxrom1.cxrom_data_out [8], _13214_, _13170_);
  and _21528_ (_13215_, _08664_, word_in[9]);
  nand _21529_ (_13216_, _08480_, _11019_);
  or _21530_ (_13217_, _08480_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  and _21531_ (_13218_, _13217_, _13216_);
  and _21532_ (_13219_, _13218_, _08666_);
  nand _21533_ (_13220_, _08480_, _10522_);
  or _21534_ (_13221_, _08480_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  and _21535_ (_13222_, _13221_, _13220_);
  and _21536_ (_13223_, _13222_, _08665_);
  or _21537_ (_13224_, _13223_, _13219_);
  and _21538_ (_13225_, _13224_, _08623_);
  nand _21539_ (_13226_, _08480_, _12478_);
  or _21540_ (_13227_, _08480_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  and _21541_ (_13228_, _13227_, _13226_);
  and _21542_ (_13229_, _13228_, _08666_);
  nand _21543_ (_13230_, _08480_, _12254_);
  or _21544_ (_13231_, _08480_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  and _21545_ (_13232_, _13231_, _13230_);
  and _21546_ (_13233_, _13232_, _08665_);
  or _21547_ (_13234_, _13233_, _13229_);
  and _21548_ (_13235_, _13234_, _08679_);
  nand _21549_ (_13236_, _08480_, _10301_);
  or _21550_ (_13237_, _08480_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  and _21551_ (_13238_, _13237_, _13236_);
  and _21552_ (_13239_, _13238_, _08666_);
  nand _21553_ (_13240_, _08480_, _10087_);
  or _21554_ (_13241_, _08480_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  and _21555_ (_13242_, _13241_, _13240_);
  and _21556_ (_13243_, _13242_, _08665_);
  or _21557_ (_13244_, _13243_, _13239_);
  and _21558_ (_13245_, _13244_, _08708_);
  nand _21559_ (_13246_, _08480_, _09843_);
  or _21560_ (_13247_, _08480_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  and _21561_ (_13248_, _13247_, _13246_);
  and _21562_ (_13249_, _13248_, _08666_);
  nand _21563_ (_13250_, _08480_, _09556_);
  or _21564_ (_13251_, _08480_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  and _21565_ (_13252_, _13251_, _13250_);
  and _21566_ (_13253_, _13252_, _08665_);
  or _21567_ (_13254_, _13253_, _13249_);
  and _21568_ (_13255_, _13254_, _08626_);
  or _21569_ (_13256_, _13255_, _13245_);
  or _21570_ (_13257_, _13256_, _13235_);
  nor _21571_ (_13258_, _13257_, _13225_);
  nor _21572_ (_13259_, _13258_, _08664_);
  or _21573_ (\oc8051_symbolic_cxrom1.cxrom_data_out [9], _13259_, _13215_);
  and _21574_ (_13260_, _08664_, word_in[10]);
  nand _21575_ (_13261_, _08480_, _11032_);
  or _21576_ (_13262_, _08480_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  and _21577_ (_13263_, _13262_, _13261_);
  and _21578_ (_13264_, _13263_, _08666_);
  nand _21579_ (_13265_, _08480_, _10534_);
  or _21580_ (_13266_, _08480_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  and _21581_ (_13267_, _13266_, _13265_);
  and _21582_ (_13268_, _13267_, _08665_);
  or _21583_ (_13269_, _13268_, _13264_);
  and _21584_ (_13270_, _13269_, _08623_);
  nand _21585_ (_13271_, _08480_, _12495_);
  or _21586_ (_13272_, _08480_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  and _21587_ (_13273_, _13272_, _13271_);
  and _21588_ (_13274_, _13273_, _08666_);
  nand _21589_ (_13275_, _08480_, _12267_);
  or _21590_ (_13276_, _08480_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  and _21591_ (_13277_, _13276_, _13275_);
  and _21592_ (_13278_, _13277_, _08665_);
  or _21593_ (_13279_, _13278_, _13274_);
  and _21594_ (_13280_, _13279_, _08679_);
  nand _21595_ (_13281_, _08480_, _10313_);
  or _21596_ (_13282_, _08480_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  and _21597_ (_13283_, _13282_, _13281_);
  and _21598_ (_13284_, _13283_, _08666_);
  nand _21599_ (_13285_, _08480_, _10101_);
  or _21600_ (_13286_, _08480_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  and _21601_ (_13287_, _13286_, _13285_);
  and _21602_ (_13288_, _13287_, _08665_);
  or _21603_ (_13289_, _13288_, _13284_);
  and _21604_ (_13290_, _13289_, _08708_);
  nand _21605_ (_13291_, _08480_, _09857_);
  or _21606_ (_13292_, _08480_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  and _21607_ (_13293_, _13292_, _13291_);
  and _21608_ (_13294_, _13293_, _08666_);
  and _21609_ (_13295_, _08480_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  nor _21610_ (_13296_, _08480_, _09734_);
  or _21611_ (_13297_, _13296_, _13295_);
  and _21612_ (_13298_, _13297_, _08665_);
  or _21613_ (_13299_, _13298_, _13294_);
  and _21614_ (_13301_, _13299_, _08626_);
  or _21615_ (_13302_, _13301_, _13290_);
  or _21616_ (_13303_, _13302_, _13280_);
  nor _21617_ (_13304_, _13303_, _13270_);
  nor _21618_ (_13305_, _13304_, _08664_);
  or _21619_ (\oc8051_symbolic_cxrom1.cxrom_data_out [10], _13305_, _13260_);
  and _21620_ (_13306_, _08664_, word_in[11]);
  nand _21621_ (_13307_, _08480_, _11047_);
  or _21622_ (_13308_, _08480_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  and _21623_ (_13309_, _13308_, _13307_);
  and _21624_ (_13310_, _13309_, _08666_);
  nand _21625_ (_13311_, _08480_, _10546_);
  or _21626_ (_13312_, _08480_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  and _21627_ (_13313_, _13312_, _13311_);
  and _21628_ (_13314_, _13313_, _08665_);
  or _21629_ (_13315_, _13314_, _13310_);
  and _21630_ (_13316_, _13315_, _08623_);
  nand _21631_ (_13317_, _08480_, _12510_);
  or _21632_ (_13318_, _08480_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  and _21633_ (_13319_, _13318_, _13317_);
  and _21634_ (_13320_, _13319_, _08666_);
  nand _21635_ (_13321_, _08480_, _12280_);
  or _21636_ (_13322_, _08480_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  and _21637_ (_13323_, _13322_, _13321_);
  and _21638_ (_13324_, _13323_, _08665_);
  or _21639_ (_13325_, _13324_, _13320_);
  and _21640_ (_13326_, _13325_, _08679_);
  nand _21641_ (_13327_, _08480_, _10325_);
  or _21642_ (_13328_, _08480_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  and _21643_ (_13329_, _13328_, _13327_);
  and _21644_ (_13330_, _13329_, _08666_);
  nand _21645_ (_13331_, _08480_, _10118_);
  or _21646_ (_13332_, _08480_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  and _21647_ (_13333_, _13332_, _13331_);
  and _21648_ (_13334_, _13333_, _08665_);
  or _21649_ (_13335_, _13334_, _13330_);
  and _21650_ (_13336_, _13335_, _08708_);
  nand _21651_ (_13337_, _08480_, _09871_);
  or _21652_ (_13338_, _08480_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  and _21653_ (_13340_, _13338_, _13337_);
  and _21654_ (_13341_, _13340_, _08666_);
  and _21655_ (_13342_, _08480_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  nor _21656_ (_13343_, _08480_, _09749_);
  or _21657_ (_13344_, _13343_, _13342_);
  and _21658_ (_13345_, _13344_, _08665_);
  or _21659_ (_13346_, _13345_, _13341_);
  and _21660_ (_13347_, _13346_, _08626_);
  or _21661_ (_13348_, _13347_, _13336_);
  or _21662_ (_13349_, _13348_, _13326_);
  nor _21663_ (_13350_, _13349_, _13316_);
  nor _21664_ (_13351_, _13350_, _08664_);
  or _21665_ (\oc8051_symbolic_cxrom1.cxrom_data_out [11], _13351_, _13306_);
  and _21666_ (_13352_, _08664_, word_in[12]);
  nand _21667_ (_13353_, _08480_, _11059_);
  or _21668_ (_13354_, _08480_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  and _21669_ (_13355_, _13354_, _13353_);
  and _21670_ (_13356_, _13355_, _08666_);
  nand _21671_ (_13357_, _08480_, _10558_);
  or _21672_ (_13358_, _08480_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  and _21673_ (_13359_, _13358_, _13357_);
  and _21674_ (_13360_, _13359_, _08665_);
  or _21675_ (_13361_, _13360_, _13356_);
  and _21676_ (_13362_, _13361_, _08623_);
  nand _21677_ (_13363_, _08480_, _09889_);
  or _21678_ (_13365_, _08480_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  and _21679_ (_13366_, _13365_, _13363_);
  and _21680_ (_13367_, _13366_, _08666_);
  and _21681_ (_13368_, _08480_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  nor _21682_ (_13369_, _08480_, _09761_);
  or _21683_ (_13370_, _13369_, _13368_);
  and _21684_ (_13371_, _13370_, _08665_);
  or _21685_ (_13372_, _13371_, _13367_);
  and _21686_ (_13373_, _13372_, _08626_);
  nand _21687_ (_13374_, _08480_, _10337_);
  or _21688_ (_13375_, _08480_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  and _21689_ (_13376_, _13375_, _13374_);
  and _21690_ (_13377_, _13376_, _08666_);
  nand _21691_ (_13378_, _08480_, _10129_);
  or _21692_ (_13379_, _08480_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  and _21693_ (_13380_, _13379_, _13378_);
  and _21694_ (_13381_, _13380_, _08665_);
  or _21695_ (_13382_, _13381_, _13377_);
  and _21696_ (_13383_, _13382_, _08708_);
  or _21697_ (_13384_, _13383_, _13373_);
  nand _21698_ (_13385_, _08480_, _12526_);
  or _21699_ (_13386_, _08480_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  and _21700_ (_13388_, _13386_, _13385_);
  and _21701_ (_13389_, _13388_, _08666_);
  nand _21702_ (_13390_, _08480_, _12292_);
  or _21703_ (_13391_, _08480_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  and _21704_ (_13392_, _13391_, _13390_);
  and _21705_ (_13393_, _13392_, _08665_);
  or _21706_ (_13394_, _13393_, _13389_);
  and _21707_ (_13395_, _13394_, _08679_);
  or _21708_ (_13396_, _13395_, _13384_);
  nor _21709_ (_13397_, _13396_, _13362_);
  nor _21710_ (_13398_, _13397_, _08664_);
  or _21711_ (\oc8051_symbolic_cxrom1.cxrom_data_out [12], _13398_, _13352_);
  and _21712_ (_13399_, _08664_, word_in[13]);
  nand _21713_ (_13400_, _08480_, _11071_);
  or _21714_ (_13401_, _08480_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  and _21715_ (_13402_, _13401_, _13400_);
  and _21716_ (_13403_, _13402_, _08666_);
  nand _21717_ (_13404_, _08480_, _10571_);
  or _21718_ (_13405_, _08480_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  and _21719_ (_13406_, _13405_, _13404_);
  and _21720_ (_13407_, _13406_, _08665_);
  or _21721_ (_13408_, _13407_, _13403_);
  and _21722_ (_13409_, _13408_, _08623_);
  and _21723_ (_13410_, _08480_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  nor _21724_ (_13411_, _08480_, _10027_);
  or _21725_ (_13412_, _13411_, _13410_);
  and _21726_ (_13413_, _13412_, _08666_);
  and _21727_ (_13414_, _08480_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  nor _21728_ (_13415_, _08480_, _09775_);
  or _21729_ (_13416_, _13415_, _13414_);
  and _21730_ (_13417_, _13416_, _08665_);
  or _21731_ (_13418_, _13417_, _13413_);
  and _21732_ (_13419_, _13418_, _08626_);
  nand _21733_ (_13420_, _08480_, _10350_);
  or _21734_ (_13421_, _08480_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  and _21735_ (_13423_, _13421_, _13420_);
  and _21736_ (_13424_, _13423_, _08666_);
  nand _21737_ (_13425_, _08480_, _10141_);
  or _21738_ (_13426_, _08480_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  and _21739_ (_13427_, _13426_, _13425_);
  and _21740_ (_13428_, _13427_, _08665_);
  or _21741_ (_13429_, _13428_, _13424_);
  and _21742_ (_13430_, _13429_, _08708_);
  or _21743_ (_13431_, _13430_, _13419_);
  nand _21744_ (_13432_, _08480_, _12537_);
  or _21745_ (_13433_, _08480_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  and _21746_ (_13434_, _13433_, _13432_);
  and _21747_ (_13435_, _13434_, _08666_);
  nand _21748_ (_13436_, _08480_, _12303_);
  or _21749_ (_13437_, _08480_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  and _21750_ (_13438_, _13437_, _13436_);
  and _21751_ (_13439_, _13438_, _08665_);
  or _21752_ (_13440_, _13439_, _13435_);
  and _21753_ (_13441_, _13440_, _08679_);
  or _21754_ (_13442_, _13441_, _13431_);
  nor _21755_ (_13443_, _13442_, _13409_);
  nor _21756_ (_13444_, _13443_, _08664_);
  or _21757_ (\oc8051_symbolic_cxrom1.cxrom_data_out [13], _13444_, _13399_);
  and _21758_ (_13445_, _08664_, word_in[14]);
  nand _21759_ (_13446_, _08480_, _11084_);
  or _21760_ (_13447_, _08480_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  and _21761_ (_13448_, _13447_, _13446_);
  and _21762_ (_13449_, _13448_, _08666_);
  nand _21763_ (_13450_, _08480_, _10583_);
  or _21764_ (_13451_, _08480_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  and _21765_ (_13452_, _13451_, _13450_);
  and _21766_ (_13453_, _13452_, _08665_);
  or _21767_ (_13454_, _13453_, _13449_);
  and _21768_ (_13455_, _13454_, _08623_);
  nand _21769_ (_13456_, _08480_, _12552_);
  or _21770_ (_13457_, _08480_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  and _21771_ (_13458_, _13457_, _13456_);
  and _21772_ (_13459_, _13458_, _08666_);
  nand _21773_ (_13460_, _08480_, _12318_);
  or _21774_ (_13461_, _08480_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  and _21775_ (_13462_, _13461_, _13460_);
  and _21776_ (_13463_, _13462_, _08665_);
  or _21777_ (_13464_, _13463_, _13459_);
  and _21778_ (_13465_, _13464_, _08679_);
  nand _21779_ (_13466_, _08480_, _10366_);
  or _21780_ (_13467_, _08480_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  and _21781_ (_13468_, _13467_, _13466_);
  and _21782_ (_13469_, _13468_, _08666_);
  nand _21783_ (_13470_, _08480_, _10156_);
  or _21784_ (_13471_, _08480_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  and _21785_ (_13472_, _13471_, _13470_);
  and _21786_ (_13473_, _13472_, _08665_);
  or _21787_ (_13474_, _13473_, _13469_);
  and _21788_ (_13475_, _13474_, _08708_);
  nand _21789_ (_13476_, _08480_, _09915_);
  or _21790_ (_13477_, _08480_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  and _21791_ (_13478_, _13477_, _13476_);
  and _21792_ (_13479_, _13478_, _08666_);
  and _21793_ (_13480_, _08480_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  nor _21794_ (_13481_, _08480_, _09792_);
  or _21795_ (_13482_, _13481_, _13480_);
  and _21796_ (_13483_, _13482_, _08665_);
  or _21797_ (_13484_, _13483_, _13479_);
  and _21798_ (_13485_, _13484_, _08626_);
  or _21799_ (_13486_, _13485_, _13475_);
  or _21800_ (_13487_, _13486_, _13465_);
  nor _21801_ (_13488_, _13487_, _13455_);
  nor _21802_ (_13489_, _13488_, _08664_);
  or _21803_ (\oc8051_symbolic_cxrom1.cxrom_data_out [14], _13489_, _13445_);
  and _21804_ (_13490_, _08769_, word_in[16]);
  and _21805_ (_13491_, _12888_, _08506_);
  and _21806_ (_13492_, _12884_, _08513_);
  or _21807_ (_13493_, _13492_, _13491_);
  and _21808_ (_13494_, _12895_, _08503_);
  and _21809_ (_13495_, _12880_, _08523_);
  or _21810_ (_13496_, _13495_, _13494_);
  or _21811_ (_13497_, _13496_, _13493_);
  or _21812_ (_13498_, _13497_, _08731_);
  and _21813_ (_13499_, _12862_, _08506_);
  and _21814_ (_13500_, _12867_, _08513_);
  or _21815_ (_13501_, _13500_, _13499_);
  and _21816_ (_13502_, _12874_, _08503_);
  and _21817_ (_13503_, _12858_, _08523_);
  or _21818_ (_13504_, _13503_, _13502_);
  or _21819_ (_13505_, _13504_, _13501_);
  or _21820_ (_13506_, _13505_, _08770_);
  nand _21821_ (_13507_, _13506_, _13498_);
  nor _21822_ (_13508_, _13507_, _08769_);
  or _21823_ (\oc8051_symbolic_cxrom1.cxrom_data_out [16], _13508_, _13490_);
  and _21824_ (_13509_, _08769_, word_in[17]);
  and _21825_ (_13510_, _12924_, _08513_);
  and _21826_ (_13511_, _12938_, _08503_);
  or _21827_ (_13512_, _13511_, _13510_);
  and _21828_ (_13513_, _12932_, _08506_);
  and _21829_ (_13514_, _12928_, _08523_);
  or _21830_ (_13515_, _13514_, _13513_);
  or _21831_ (_13516_, _13515_, _13512_);
  or _21832_ (_13517_, _13516_, _08731_);
  and _21833_ (_13518_, _12912_, _08506_);
  and _21834_ (_13520_, _12904_, _08513_);
  or _21835_ (_13521_, _13520_, _13518_);
  and _21836_ (_13522_, _12918_, _08503_);
  and _21837_ (_13523_, _12908_, _08523_);
  or _21838_ (_13524_, _13523_, _13522_);
  or _21839_ (_13526_, _13524_, _13521_);
  or _21840_ (_13527_, _13526_, _08770_);
  nand _21841_ (_13528_, _13527_, _13517_);
  nor _21842_ (_13529_, _13528_, _08769_);
  or _21843_ (\oc8051_symbolic_cxrom1.cxrom_data_out [17], _13529_, _13509_);
  and _21844_ (_13530_, _08769_, word_in[18]);
  and _21845_ (_13531_, _12975_, _08506_);
  and _21846_ (_13532_, _12967_, _08513_);
  or _21847_ (_13533_, _13532_, _13531_);
  and _21848_ (_13534_, _12981_, _08503_);
  and _21849_ (_13535_, _12971_, _08523_);
  or _21850_ (_13536_, _13535_, _13534_);
  or _21851_ (_13537_, _13536_, _13533_);
  or _21852_ (_13538_, _13537_, _08731_);
  and _21853_ (_13539_, _12955_, _08506_);
  and _21854_ (_13540_, _12947_, _08513_);
  or _21855_ (_13541_, _13540_, _13539_);
  and _21856_ (_13542_, _12961_, _08503_);
  and _21857_ (_13543_, _12951_, _08523_);
  or _21858_ (_13544_, _13543_, _13542_);
  or _21859_ (_13545_, _13544_, _13541_);
  or _21860_ (_13546_, _13545_, _08770_);
  nand _21861_ (_13547_, _13546_, _13538_);
  nor _21862_ (_13549_, _13547_, _08769_);
  or _21863_ (\oc8051_symbolic_cxrom1.cxrom_data_out [18], _13549_, _13530_);
  and _21864_ (_13550_, _08769_, word_in[19]);
  and _21865_ (_13552_, _13010_, _08513_);
  and _21866_ (_13553_, _13026_, _08503_);
  or _21867_ (_13554_, _13553_, _13552_);
  and _21868_ (_13555_, _13019_, _08506_);
  and _21869_ (_13556_, _13015_, _08523_);
  or _21870_ (_13557_, _13556_, _13555_);
  or _21871_ (_13558_, _13557_, _13554_);
  or _21872_ (_13559_, _13558_, _08731_);
  and _21873_ (_13560_, _12998_, _08506_);
  and _21874_ (_13561_, _12990_, _08513_);
  or _21875_ (_13562_, _13561_, _13560_);
  and _21876_ (_13563_, _13004_, _08503_);
  and _21877_ (_13564_, _12994_, _08523_);
  or _21878_ (_13565_, _13564_, _13563_);
  or _21879_ (_13566_, _13565_, _13562_);
  or _21880_ (_13567_, _13566_, _08770_);
  nand _21881_ (_13568_, _13567_, _13559_);
  nor _21882_ (_13569_, _13568_, _08769_);
  or _21883_ (\oc8051_symbolic_cxrom1.cxrom_data_out [19], _13569_, _13550_);
  and _21884_ (_13570_, _08769_, word_in[20]);
  and _21885_ (_13571_, _13058_, _08513_);
  and _21886_ (_13572_, _13072_, _08503_);
  or _21887_ (_13573_, _13572_, _13571_);
  and _21888_ (_13574_, _13066_, _08506_);
  and _21889_ (_13575_, _13062_, _08523_);
  or _21890_ (_13576_, _13575_, _13574_);
  or _21891_ (_13577_, _13576_, _13573_);
  or _21892_ (_13578_, _13577_, _08731_);
  and _21893_ (_13579_, _13035_, _08513_);
  and _21894_ (_13580_, _13052_, _08503_);
  or _21895_ (_13581_, _13580_, _13579_);
  and _21896_ (_13582_, _13044_, _08506_);
  and _21897_ (_13583_, _13040_, _08523_);
  or _21898_ (_13584_, _13583_, _13582_);
  or _21899_ (_13585_, _13584_, _13581_);
  or _21900_ (_13586_, _13585_, _08770_);
  nand _21901_ (_13587_, _13586_, _13578_);
  nor _21902_ (_13588_, _13587_, _08769_);
  or _21903_ (\oc8051_symbolic_cxrom1.cxrom_data_out [20], _13588_, _13570_);
  and _21904_ (_13590_, _08769_, word_in[21]);
  and _21905_ (_13591_, _13102_, _08513_);
  and _21906_ (_13592_, _13117_, _08503_);
  or _21907_ (_13593_, _13592_, _13591_);
  and _21908_ (_13594_, _13111_, _08506_);
  and _21909_ (_13595_, _13106_, _08523_);
  or _21910_ (_13597_, _13595_, _13594_);
  or _21911_ (_13598_, _13597_, _13593_);
  or _21912_ (_13599_, _13598_, _08731_);
  and _21913_ (_13600_, _13082_, _08513_);
  and _21914_ (_13601_, _13096_, _08503_);
  or _21915_ (_13602_, _13601_, _13600_);
  and _21916_ (_13603_, _13090_, _08506_);
  and _21917_ (_13604_, _13086_, _08523_);
  or _21918_ (_13605_, _13604_, _13603_);
  or _21919_ (_13606_, _13605_, _13602_);
  or _21920_ (_13607_, _13606_, _08770_);
  nand _21921_ (_13608_, _13607_, _13599_);
  nor _21922_ (_13609_, _13608_, _08769_);
  or _21923_ (\oc8051_symbolic_cxrom1.cxrom_data_out [21], _13609_, _13590_);
  and _21924_ (_13610_, _08769_, word_in[22]);
  and _21925_ (_13611_, _13157_, _08506_);
  and _21926_ (_13612_, _13153_, _08513_);
  or _21927_ (_13613_, _13612_, _13611_);
  and _21928_ (_13614_, _13164_, _08503_);
  and _21929_ (_13615_, _13147_, _08523_);
  or _21930_ (_13616_, _13615_, _13614_);
  or _21931_ (_13617_, _13616_, _13613_);
  or _21932_ (_13618_, _13617_, _08731_);
  and _21933_ (_13619_, _13130_, _08506_);
  and _21934_ (_13620_, _13134_, _08513_);
  or _21935_ (_13621_, _13620_, _13619_);
  and _21936_ (_13622_, _13141_, _08503_);
  and _21937_ (_13623_, _13126_, _08523_);
  or _21938_ (_13624_, _13623_, _13622_);
  or _21939_ (_13625_, _13624_, _13621_);
  or _21940_ (_13626_, _13625_, _08770_);
  nand _21941_ (_13627_, _13626_, _13618_);
  nor _21942_ (_13628_, _13627_, _08769_);
  or _21943_ (\oc8051_symbolic_cxrom1.cxrom_data_out [22], _13628_, _13610_);
  and _21944_ (_13629_, _08828_, word_in[24]);
  and _21945_ (_13630_, _13207_, _08666_);
  and _21946_ (_13631_, _13203_, _08665_);
  or _21947_ (_13632_, _13631_, _13630_);
  and _21948_ (_13633_, _13632_, _08814_);
  and _21949_ (_13635_, _13177_, _08666_);
  and _21950_ (_13636_, _13173_, _08665_);
  or _21951_ (_13638_, _13636_, _13635_);
  and _21952_ (_13639_, _13638_, _08800_);
  and _21953_ (_13640_, _13197_, _08666_);
  and _21954_ (_13641_, _13193_, _08665_);
  or _21955_ (_13642_, _13641_, _13640_);
  and _21956_ (_13643_, _13642_, _08837_);
  and _21957_ (_13644_, _13187_, _08666_);
  and _21958_ (_13645_, _13183_, _08665_);
  or _21959_ (_13646_, _13645_, _13644_);
  and _21960_ (_13647_, _13646_, _08842_);
  or _21961_ (_13648_, _13647_, _13643_);
  or _21962_ (_13649_, _13648_, _13639_);
  nor _21963_ (_13650_, _13649_, _13633_);
  nor _21964_ (_13651_, _13650_, _08828_);
  or _21965_ (\oc8051_symbolic_cxrom1.cxrom_data_out [24], _13651_, _13629_);
  and _21966_ (_13652_, _08828_, word_in[25]);
  and _21967_ (_13653_, _13222_, _08666_);
  and _21968_ (_13654_, _13218_, _08665_);
  or _21969_ (_13655_, _13654_, _13653_);
  and _21970_ (_13656_, _13655_, _08800_);
  and _21971_ (_13657_, _13252_, _08666_);
  and _21972_ (_13658_, _13248_, _08665_);
  or _21973_ (_13659_, _13658_, _13657_);
  and _21974_ (_13660_, _13659_, _08814_);
  and _21975_ (_13662_, _13242_, _08666_);
  and _21976_ (_13663_, _13238_, _08665_);
  or _21977_ (_13664_, _13663_, _13662_);
  and _21978_ (_13666_, _13664_, _08837_);
  and _21979_ (_13667_, _13232_, _08666_);
  and _21980_ (_13668_, _13228_, _08665_);
  or _21981_ (_13669_, _13668_, _13667_);
  and _21982_ (_13670_, _13669_, _08842_);
  or _21983_ (_13671_, _13670_, _13666_);
  or _21984_ (_13672_, _13671_, _13660_);
  nor _21985_ (_13673_, _13672_, _13656_);
  nor _21986_ (_13674_, _13673_, _08828_);
  or _21987_ (\oc8051_symbolic_cxrom1.cxrom_data_out [25], _13674_, _13652_);
  and _21988_ (_13676_, _08828_, word_in[26]);
  and _21989_ (_13677_, _13297_, _08666_);
  and _21990_ (_13678_, _13293_, _08665_);
  or _21991_ (_13679_, _13678_, _13677_);
  and _21992_ (_13680_, _13679_, _08814_);
  and _21993_ (_13681_, _13267_, _08666_);
  and _21994_ (_13682_, _13263_, _08665_);
  or _21995_ (_13683_, _13682_, _13681_);
  and _21996_ (_13684_, _13683_, _08800_);
  and _21997_ (_13685_, _13287_, _08666_);
  and _21998_ (_13686_, _13283_, _08665_);
  or _21999_ (_13687_, _13686_, _13685_);
  and _22000_ (_13688_, _13687_, _08837_);
  and _22001_ (_13689_, _13277_, _08666_);
  and _22002_ (_13691_, _13273_, _08665_);
  or _22003_ (_13692_, _13691_, _13689_);
  and _22004_ (_13694_, _13692_, _08842_);
  or _22005_ (_13695_, _13694_, _13688_);
  or _22006_ (_13696_, _13695_, _13684_);
  nor _22007_ (_13697_, _13696_, _13680_);
  nor _22008_ (_13698_, _13697_, _08828_);
  or _22009_ (\oc8051_symbolic_cxrom1.cxrom_data_out [26], _13698_, _13676_);
  and _22010_ (_13699_, _08828_, word_in[27]);
  and _22011_ (_13700_, _13313_, _08666_);
  and _22012_ (_13701_, _13309_, _08665_);
  or _22013_ (_13702_, _13701_, _13700_);
  and _22014_ (_13703_, _13702_, _08800_);
  and _22015_ (_13704_, _13344_, _08666_);
  and _22016_ (_13705_, _13340_, _08665_);
  or _22017_ (_13706_, _13705_, _13704_);
  and _22018_ (_13707_, _13706_, _08814_);
  and _22019_ (_13708_, _13333_, _08666_);
  and _22020_ (_13709_, _13329_, _08665_);
  or _22021_ (_13710_, _13709_, _13708_);
  and _22022_ (_13711_, _13710_, _08837_);
  and _22023_ (_13712_, _13323_, _08666_);
  and _22024_ (_13713_, _13319_, _08665_);
  or _22025_ (_13715_, _13713_, _13712_);
  and _22026_ (_13716_, _13715_, _08842_);
  or _22027_ (_13717_, _13716_, _13711_);
  or _22028_ (_13718_, _13717_, _13707_);
  nor _22029_ (_13719_, _13718_, _13703_);
  nor _22030_ (_13720_, _13719_, _08828_);
  or _22031_ (\oc8051_symbolic_cxrom1.cxrom_data_out [27], _13720_, _13699_);
  and _22032_ (_13722_, _08828_, word_in[28]);
  and _22033_ (_13723_, _13359_, _08666_);
  and _22034_ (_13724_, _13355_, _08665_);
  or _22035_ (_13725_, _13724_, _13723_);
  and _22036_ (_13726_, _13725_, _08800_);
  and _22037_ (_13728_, _13370_, _08666_);
  and _22038_ (_13729_, _13366_, _08665_);
  or _22039_ (_13730_, _13729_, _13728_);
  and _22040_ (_13731_, _13730_, _08814_);
  and _22041_ (_13732_, _13380_, _08666_);
  and _22042_ (_13733_, _13376_, _08665_);
  or _22043_ (_13734_, _13733_, _13732_);
  and _22044_ (_13735_, _13734_, _08837_);
  and _22045_ (_13736_, _13392_, _08666_);
  and _22046_ (_13737_, _13388_, _08665_);
  or _22047_ (_13738_, _13737_, _13736_);
  and _22048_ (_13740_, _13738_, _08842_);
  or _22049_ (_13741_, _13740_, _13735_);
  or _22050_ (_13743_, _13741_, _13731_);
  nor _22051_ (_13744_, _13743_, _13726_);
  nor _22052_ (_13746_, _13744_, _08828_);
  or _22053_ (\oc8051_symbolic_cxrom1.cxrom_data_out [28], _13746_, _13722_);
  and _22054_ (_13748_, _08828_, word_in[29]);
  and _22055_ (_13749_, _13406_, _08666_);
  and _22056_ (_13750_, _13402_, _08665_);
  or _22057_ (_13751_, _13750_, _13749_);
  and _22058_ (_13752_, _13751_, _08800_);
  and _22059_ (_13753_, _13416_, _08666_);
  and _22060_ (_13755_, _13412_, _08665_);
  or _22061_ (_13756_, _13755_, _13753_);
  and _22062_ (_13757_, _13756_, _08814_);
  and _22063_ (_13758_, _13427_, _08666_);
  and _22064_ (_13759_, _13423_, _08665_);
  or _22065_ (_13760_, _13759_, _13758_);
  and _22066_ (_13761_, _13760_, _08837_);
  and _22067_ (_13762_, _13438_, _08666_);
  and _22068_ (_13763_, _13434_, _08665_);
  or _22069_ (_13764_, _13763_, _13762_);
  and _22070_ (_13765_, _13764_, _08842_);
  or _22071_ (_13766_, _13765_, _13761_);
  or _22072_ (_13767_, _13766_, _13757_);
  nor _22073_ (_13768_, _13767_, _13752_);
  nor _22074_ (_13769_, _13768_, _08828_);
  or _22075_ (\oc8051_symbolic_cxrom1.cxrom_data_out [29], _13769_, _13748_);
  and _22076_ (_13770_, _08828_, word_in[30]);
  and _22077_ (_13771_, _13482_, _08666_);
  and _22078_ (_13772_, _13478_, _08665_);
  or _22079_ (_13773_, _13772_, _13771_);
  and _22080_ (_13774_, _13773_, _08814_);
  and _22081_ (_13775_, _13452_, _08666_);
  and _22082_ (_13776_, _13448_, _08665_);
  or _22083_ (_13777_, _13776_, _13775_);
  and _22084_ (_13778_, _13777_, _08800_);
  and _22085_ (_13779_, _13472_, _08666_);
  and _22086_ (_13780_, _13468_, _08665_);
  or _22087_ (_13781_, _13780_, _13779_);
  and _22088_ (_13782_, _13781_, _08837_);
  and _22089_ (_13784_, _13462_, _08666_);
  and _22090_ (_13785_, _13458_, _08665_);
  or _22091_ (_13786_, _13785_, _13784_);
  and _22092_ (_13787_, _13786_, _08842_);
  or _22093_ (_13788_, _13787_, _13782_);
  or _22094_ (_13789_, _13788_, _13778_);
  nor _22095_ (_13790_, _13789_, _13774_);
  nor _22096_ (_13791_, _13790_, _08828_);
  or _22097_ (\oc8051_symbolic_cxrom1.cxrom_data_out [30], _13791_, _13770_);
  and _22098_ (_11141_, _07987_, _06444_);
  and _22099_ (_11154_, _09095_, _06444_);
  and _22100_ (_11159_, _07927_, _06444_);
  nor _22101_ (_13792_, _07602_, _07606_);
  and _22102_ (_13793_, _07602_, _07606_);
  or _22103_ (_13794_, _13793_, _13792_);
  and _22104_ (_11176_, _13794_, _06444_);
  and _22105_ (_11198_, _08097_, _06444_);
  and _22106_ (_11214_, _08205_, _06444_);
  and _22107_ (_11219_, _09196_, _06444_);
  and _22108_ (_11222_, _09275_, _06444_);
  and _22109_ (_11239_, _08284_, _06444_);
  and _22110_ (_11248_, _07635_, _06444_);
  and _22111_ (_11252_, _07628_, _06444_);
  and _22112_ (_11298_, _08163_, _06444_);
  and _22113_ (_11304_, _08246_, _06444_);
  and _22114_ (_11308_, _08332_, _06444_);
  and _22115_ (_13795_, _08064_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  not _22116_ (_13796_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _22117_ (_13797_, _08064_, _13796_);
  or _22118_ (_13798_, _13797_, _13795_);
  and _22119_ (_11397_, _13798_, _06444_);
  or _22120_ (_13799_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  nand _22121_ (_13800_, _07432_, _11718_);
  and _22122_ (_13801_, _13800_, _06444_);
  and _22123_ (_11462_, _13801_, _13799_);
  and _22124_ (_13802_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  and _22125_ (_13803_, _12223_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  or _22126_ (_13804_, _13803_, _13802_);
  and _22127_ (_11506_, _13804_, _06444_);
  and _22128_ (_13806_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor _22129_ (_13807_, _07432_, _11016_);
  or _22130_ (_13808_, _13807_, _13806_);
  and _22131_ (_11748_, _13808_, _06444_);
  or _22132_ (_13809_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  nand _22133_ (_13810_, _07432_, _11194_);
  and _22134_ (_13811_, _13810_, _06444_);
  and _22135_ (_11752_, _13811_, _13809_);
  or _22136_ (_13812_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  nand _22137_ (_13813_, _07432_, _12171_);
  and _22138_ (_13814_, _13813_, _06444_);
  and _22139_ (_11768_, _13814_, _13812_);
  or _22140_ (_13815_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  nand _22141_ (_13816_, _07432_, _09662_);
  and _22142_ (_13817_, _13816_, _06444_);
  and _22143_ (_11783_, _13817_, _13815_);
  nand _22144_ (_13818_, _11589_, _10112_);
  or _22145_ (_13819_, _10112_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  and _22146_ (_13820_, _13819_, _06444_);
  and _22147_ (_11806_, _13820_, _13818_);
  or _22148_ (_13821_, _09339_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  or _22149_ (_13822_, _09467_, _09373_);
  and _22150_ (_11894_, _13822_, _13821_);
  and _22151_ (_11898_, _07765_, _06444_);
  and _22152_ (_11913_, _08278_, _06444_);
  nor _22153_ (_11916_, _09092_, rst);
  nor _22154_ (_13823_, _07190_, _06666_);
  and _22155_ (_13824_, _07190_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  or _22156_ (_13825_, _13824_, _13823_);
  and _22157_ (_11956_, _13825_, _06444_);
  nand _22158_ (_13826_, _08474_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  or _22159_ (_13827_, _08474_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  and _22160_ (_13828_, _13827_, _13826_);
  and _22161_ (_11985_, _13828_, _06443_);
  and _22162_ (_13830_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor _22163_ (_13832_, _07432_, _12492_);
  or _22164_ (_13833_, _13832_, _13830_);
  and _22165_ (_11988_, _13833_, _06444_);
  and _22166_ (_13835_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans , \oc8051_top_1.oc8051_sfr1.pres_ow );
  and _22167_ (_13836_, _13835_, _06295_);
  nor _22168_ (_13837_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  nor _22169_ (_13838_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  and _22170_ (_13840_, _13838_, _13837_);
  nor _22171_ (_13841_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  nor _22172_ (_13842_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  nor _22173_ (_13843_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  and _22174_ (_13845_, _13843_, _13842_);
  and _22175_ (_13846_, _13845_, _13841_);
  and _22176_ (_13847_, _13846_, _13840_);
  and _22177_ (_13848_, _13847_, _13836_);
  not _22178_ (_13849_, _13836_);
  nand _22179_ (_13850_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  nor _22180_ (_13851_, _13850_, _06298_);
  nor _22181_ (_13852_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  nor _22182_ (_13853_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  and _22183_ (_13854_, _13853_, _13852_);
  not _22184_ (_13855_, _13854_);
  nor _22185_ (_13856_, _13855_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  nand _22186_ (_13857_, _13856_, _13847_);
  nand _22187_ (_13858_, _13855_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  nand _22188_ (_13859_, _13858_, _13857_);
  and _22189_ (_13860_, _13859_, _06298_);
  or _22190_ (_13861_, _13860_, _13851_);
  and _22191_ (_13862_, _13861_, _13849_);
  or _22192_ (_13863_, _13862_, _13848_);
  and _22193_ (_11992_, _13863_, _06443_);
  and _22194_ (_13864_, _06440_, _06382_);
  and _22195_ (_13865_, _13864_, _06434_);
  not _22196_ (_13866_, _06297_);
  or _22197_ (_13867_, _13857_, _13866_);
  nand _22198_ (_13868_, _13867_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  nor _22199_ (_13869_, _13868_, _13848_);
  or _22200_ (_13870_, _13869_, _13865_);
  and _22201_ (_12000_, _13870_, _06444_);
  not _22202_ (_13871_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  and _22203_ (_13872_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  not _22204_ (_13873_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and _22205_ (_13874_, _07382_, _13873_);
  not _22206_ (_13875_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  nor _22207_ (_13876_, _13875_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  or _22208_ (_13877_, _13876_, _13874_);
  nor _22209_ (_13878_, _13877_, _13872_);
  nand _22210_ (_13879_, _13878_, _13871_);
  nor _22211_ (_13880_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nor _22212_ (_13881_, _13880_, _13878_);
  nand _22213_ (_13882_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nand _22214_ (_13883_, _13882_, _13881_);
  and _22215_ (_13884_, _13883_, _06444_);
  and _22216_ (_12007_, _13884_, _13879_);
  and _22217_ (_12010_, _13881_, _06444_);
  and _22218_ (_13885_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  not _22219_ (_13886_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor _22220_ (_13887_, _07432_, _13886_);
  or _22221_ (_13888_, _13887_, _13885_);
  and _22222_ (_12027_, _13888_, _06444_);
  and _22223_ (_13889_, _07214_, _06933_);
  and _22224_ (_13890_, _13889_, _07402_);
  or _22225_ (_13891_, _13890_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  and _22226_ (_13892_, _13891_, _06444_);
  and _22227_ (_13893_, _08978_, _06933_);
  nand _22228_ (_13894_, _13893_, _06978_);
  and _22229_ (_12036_, _13894_, _13892_);
  and _22230_ (_13895_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  not _22231_ (_13896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor _22232_ (_13898_, _07432_, _13896_);
  or _22233_ (_13899_, _13898_, _13895_);
  and _22234_ (_12049_, _13899_, _06444_);
  nor _22235_ (_13900_, _06394_, _06336_);
  and _22236_ (_13901_, _07401_, _06676_);
  and _22237_ (_13902_, _13901_, _13900_);
  and _22238_ (_13903_, _13902_, _06933_);
  nand _22239_ (_13904_, _13903_, _06930_);
  or _22240_ (_13905_, _13903_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  and _22241_ (_13906_, _06945_, _06382_);
  not _22242_ (_13907_, _13906_);
  and _22243_ (_13908_, _13907_, _13905_);
  and _22244_ (_13909_, _13908_, _13904_);
  nor _22245_ (_13910_, _13907_, _06978_);
  or _22246_ (_13911_, _13910_, _13909_);
  and _22247_ (_12053_, _13911_, _06444_);
  and _22248_ (_12057_, _08078_, _06444_);
  and _22249_ (_13912_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  not _22250_ (_13913_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and _22251_ (_13914_, _07382_, _13913_);
  or _22252_ (_13915_, _13914_, _13876_);
  nor _22253_ (_13916_, _13915_, _13912_);
  or _22254_ (_13917_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  nand _22255_ (_13918_, _13917_, _06444_);
  nor _22256_ (_12083_, _13918_, _13916_);
  nor _22257_ (_12089_, _07381_, rst);
  not _22258_ (_13919_, rxd_i);
  nand _22259_ (_13920_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r , _13919_);
  nand _22260_ (_13921_, _13920_, _09353_);
  or _22261_ (_13922_, _09354_, _09343_);
  and _22262_ (_13923_, _13922_, _13921_);
  not _22263_ (_13924_, _09340_);
  nand _22264_ (_13926_, _09427_, _13924_);
  or _22265_ (_13927_, _13926_, _13923_);
  and _22266_ (_12133_, _13927_, _09373_);
  and _22267_ (_13929_, _09678_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and _22268_ (_13930_, _13929_, _09345_);
  and _22269_ (_13931_, _09677_, _13930_);
  not _22270_ (_13932_, _09344_);
  nor _22271_ (_13933_, _13929_, _13932_);
  or _22272_ (_13934_, _13933_, _09675_);
  and _22273_ (_13935_, _13934_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  or _22274_ (_13936_, _13935_, _13931_);
  and _22275_ (_12140_, _13936_, _06444_);
  and _22276_ (_13937_, _09679_, _09346_);
  and _22277_ (_13938_, _09677_, _13937_);
  nand _22278_ (_13939_, _13938_, _13919_);
  or _22279_ (_13940_, _13938_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  and _22280_ (_13941_, _13940_, _06444_);
  and _22281_ (_12143_, _13941_, _13939_);
  not _22282_ (_13942_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r );
  nor _22283_ (_13943_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , _09355_);
  not _22284_ (_13944_, _13943_);
  nor _22285_ (_13945_, _06295_, _09339_);
  and _22286_ (_13946_, _13945_, _13944_);
  and _22287_ (_13947_, _13946_, _13932_);
  nor _22288_ (_13948_, _13947_, _13942_);
  and _22289_ (_13949_, _13947_, rxd_i);
  or _22290_ (_13950_, _13949_, rst);
  or _22291_ (_12153_, _13950_, _13948_);
  or _22292_ (_13951_, _09351_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  or _22293_ (_13952_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _22294_ (_13953_, _13952_, _06295_);
  or _22295_ (_13954_, _13953_, _09344_);
  nand _22296_ (_13955_, _13954_, _13951_);
  nand _22297_ (_12159_, _13955_, _09373_);
  and _22298_ (_13956_, _09328_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  and _22299_ (_13957_, _06439_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  and _22300_ (_13958_, _13957_, _09332_);
  and _22301_ (_13959_, _07425_, _07359_);
  or _22302_ (_13960_, _13959_, _13958_);
  or _22303_ (_13961_, _13960_, _13956_);
  and _22304_ (_12259_, _13961_, _06444_);
  nand _22305_ (_13962_, _07613_, _07602_);
  or _22306_ (_13963_, _07602_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  and _22307_ (_13964_, _13963_, _06444_);
  and _22308_ (_12304_, _13964_, _13962_);
  and _22309_ (_12317_, _08990_, _06444_);
  and _22310_ (_13967_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  not _22311_ (_13968_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nor _22312_ (_13969_, _07432_, _13968_);
  or _22313_ (_13970_, _13969_, _13967_);
  and _22314_ (_12334_, _13970_, _06444_);
  or _22315_ (_13971_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  nand _22316_ (_13972_, _07432_, _11838_);
  and _22317_ (_13973_, _13972_, _06444_);
  and _22318_ (_12341_, _13973_, _13971_);
  nand _22319_ (_13975_, _12829_, _10494_);
  or _22320_ (_13976_, _12829_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  and _22321_ (_13977_, _13976_, _06444_);
  and _22322_ (_12351_, _13977_, _13975_);
  and _22323_ (_13979_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  not _22324_ (_13980_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nor _22325_ (_13982_, _07432_, _13980_);
  or _22326_ (_13983_, _13982_, _13979_);
  and _22327_ (_12356_, _13983_, _06444_);
  and _22328_ (_13984_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  not _22329_ (_13985_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nor _22330_ (_13986_, _07432_, _13985_);
  or _22331_ (_13987_, _13986_, _13984_);
  and _22332_ (_12375_, _13987_, _06444_);
  and _22333_ (_13989_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  not _22334_ (_13990_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  nor _22335_ (_13992_, _07432_, _13990_);
  or _22336_ (_13993_, _13992_, _13989_);
  and _22337_ (_12380_, _13993_, _06444_);
  and _22338_ (_13994_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  and _22339_ (_13995_, _12223_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  or _22340_ (_13997_, _13995_, _13994_);
  and _22341_ (_12407_, _13997_, _06444_);
  and _22342_ (_13998_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  not _22343_ (_13999_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nor _22344_ (_14001_, _07432_, _13999_);
  or _22345_ (_14002_, _14001_, _13998_);
  and _22346_ (_12409_, _14002_, _06444_);
  and _22347_ (_14003_, _07425_, _07378_);
  and _22348_ (_14004_, _07153_, _07271_);
  or _22349_ (_14005_, _14004_, _07420_);
  and _22350_ (_14006_, _14005_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  or _22351_ (_14007_, _14006_, _14003_);
  and _22352_ (_12465_, _14007_, _06444_);
  and _22353_ (_14008_, _07190_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  nor _22354_ (_14010_, _07190_, _06978_);
  or _22355_ (_14011_, _14010_, _14008_);
  and _22356_ (_12599_, _14011_, _06444_);
  nor _22357_ (_14013_, _12830_, _06666_);
  not _22358_ (_14014_, _07415_);
  or _22359_ (_14015_, _12825_, _14014_);
  and _22360_ (_14016_, _14015_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  or _22361_ (_14017_, _14016_, _14013_);
  and _22362_ (_12642_, _14017_, _06444_);
  and _22363_ (_14018_, _07046_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  nor _22364_ (_14019_, _07300_, _07046_);
  or _22365_ (_14020_, _14019_, _14018_);
  and _22366_ (_12752_, _14020_, _06444_);
  and _22367_ (_14022_, _07070_, _06448_);
  and _22368_ (_14024_, _06449_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  or _22369_ (_14025_, _14024_, _14022_);
  and _22370_ (_12864_, _14025_, _06444_);
  and _22371_ (_14027_, _09373_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  or _22372_ (_12870_, _14027_, _09425_);
  and _22373_ (_12889_, _06444_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  and _22374_ (_14028_, _09373_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  or _22375_ (_13011_, _14028_, _09418_);
  or _22376_ (_14029_, _09431_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  or _22377_ (_14030_, _14029_, _13932_);
  and _22378_ (_14031_, _14030_, _09430_);
  or _22379_ (_14033_, _14031_, rxd_i);
  and _22380_ (_14034_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1], rxd_i);
  nor _22381_ (_14035_, _14034_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0]);
  and _22382_ (_14036_, _14035_, _09349_);
  and _22383_ (_14038_, _14036_, _09344_);
  nor _22384_ (_14039_, _14038_, _09360_);
  and _22385_ (_14041_, _14039_, _14033_);
  or _22386_ (_14042_, _14041_, _09339_);
  nor _22387_ (_14043_, _09351_, _09339_);
  or _22388_ (_14044_, _14043_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  and _22389_ (_14045_, _14044_, _06444_);
  and _22390_ (_13023_, _14045_, _14042_);
  and _22391_ (_14046_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  nor _22392_ (_14048_, _07432_, _12452_);
  or _22393_ (_14049_, _14048_, _14046_);
  and _22394_ (_13038_, _14049_, _06444_);
  and _22395_ (_13046_, _06444_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  and _22396_ (_13050_, _07586_, _06444_);
  and _22397_ (_14050_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  not _22398_ (_14051_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor _22399_ (_14052_, _07432_, _14051_);
  or _22400_ (_14053_, _14052_, _14050_);
  and _22401_ (_13078_, _14053_, _06444_);
  and _22402_ (_14054_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  not _22403_ (_14056_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nor _22404_ (_14057_, _07432_, _14056_);
  or _22405_ (_14058_, _14057_, _14054_);
  and _22406_ (_13108_, _14058_, _06444_);
  and _22407_ (_14059_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  not _22408_ (_14060_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor _22409_ (_14061_, _07432_, _14060_);
  or _22410_ (_14062_, _14061_, _14059_);
  and _22411_ (_13138_, _14062_, _06444_);
  nor _22412_ (_14063_, _11589_, _09146_);
  and _22413_ (_14064_, _09146_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  or _22414_ (_14065_, _14064_, _14063_);
  or _22415_ (_14066_, _14065_, _07158_);
  or _22416_ (_14067_, _06439_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  and _22417_ (_14068_, _14067_, _06444_);
  and _22418_ (_13148_, _14068_, _14066_);
  and _22419_ (_14069_, _07154_, _06439_);
  not _22420_ (_14070_, _14069_);
  and _22421_ (_14071_, _14070_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  nor _22422_ (_14072_, _14070_, _11589_);
  or _22423_ (_14074_, _14072_, _14071_);
  and _22424_ (_13161_, _14074_, _06444_);
  nand _22425_ (_14075_, _10112_, _07188_);
  or _22426_ (_14076_, _10112_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  and _22427_ (_14077_, _14076_, _06444_);
  and _22428_ (_13300_, _14077_, _14075_);
  nor _22429_ (_14078_, _11919_, _11703_);
  and _22430_ (_14079_, _11861_, _11809_);
  and _22431_ (_14080_, _14079_, _14078_);
  and _22432_ (_14081_, _11669_, _11741_);
  nor _22433_ (_14082_, _11630_, _11782_);
  and _22434_ (_14083_, _14082_, _14081_);
  and _22435_ (_14084_, _14083_, _14080_);
  not _22436_ (_14085_, _11703_);
  and _22437_ (_14086_, _11919_, _14085_);
  and _22438_ (_14087_, _14079_, _14086_);
  and _22439_ (_14088_, _14083_, _14087_);
  nor _22440_ (_14089_, _14088_, _14084_);
  not _22441_ (_14090_, _11861_);
  nor _22442_ (_14091_, _14090_, _11809_);
  and _22443_ (_14092_, _14091_, _14086_);
  and _22444_ (_14093_, _14083_, _14092_);
  and _22445_ (_14094_, _14090_, _11809_);
  and _22446_ (_14095_, _14094_, _14078_);
  and _22447_ (_14096_, _14083_, _14095_);
  nor _22448_ (_14097_, _14096_, _14093_);
  and _22449_ (_14098_, _14097_, _14089_);
  not _22450_ (_14099_, _11782_);
  nor _22451_ (_14100_, _11630_, _14099_);
  and _22452_ (_14101_, _14081_, _14100_);
  and _22453_ (_14102_, _14087_, _14101_);
  nor _22454_ (_14103_, _11861_, _11809_);
  and _22455_ (_14104_, _14086_, _14103_);
  and _22456_ (_14105_, _14083_, _14104_);
  nor _22457_ (_14106_, _14105_, _14102_);
  not _22458_ (_14107_, _11741_);
  and _22459_ (_14108_, _14100_, _14107_);
  and _22460_ (_14109_, _14108_, _11669_);
  and _22461_ (_14110_, _14109_, _14087_);
  not _22462_ (_14111_, _11669_);
  and _22463_ (_14112_, _14108_, _14111_);
  not _22464_ (_14113_, _11919_);
  and _22465_ (_14114_, _14103_, _14113_);
  and _22466_ (_14115_, _14114_, _11703_);
  and _22467_ (_14116_, _14115_, _14112_);
  nor _22468_ (_14117_, _14116_, _14110_);
  and _22469_ (_14118_, _14117_, _14106_);
  and _22470_ (_14119_, _14118_, _14098_);
  and _22471_ (_14120_, _14104_, _14101_);
  and _22472_ (_14121_, _14094_, _14086_);
  and _22473_ (_14122_, _14121_, _14101_);
  nor _22474_ (_14123_, _14122_, _14120_);
  and _22475_ (_14124_, _14095_, _14101_);
  and _22476_ (_14125_, _14092_, _14101_);
  nor _22477_ (_14126_, _14125_, _14124_);
  and _22478_ (_14127_, _14126_, _14123_);
  and _22479_ (_14128_, _14100_, _11741_);
  and _22480_ (_14129_, _14128_, _14111_);
  and _22481_ (_14130_, _14129_, _14121_);
  and _22482_ (_14131_, _14129_, _14087_);
  nor _22483_ (_14132_, _14131_, _14130_);
  and _22484_ (_14133_, _14080_, _14101_);
  and _22485_ (_14134_, _14115_, _14101_);
  nor _22486_ (_14135_, _14134_, _14133_);
  and _22487_ (_14136_, _14135_, _14132_);
  and _22488_ (_14137_, _14136_, _14127_);
  and _22489_ (_14138_, _14137_, _14119_);
  and _22490_ (_14139_, _11919_, _11703_);
  and _22491_ (_14140_, _14139_, _14079_);
  and _22492_ (_14141_, _14140_, _14111_);
  and _22493_ (_14142_, _14082_, _11741_);
  and _22494_ (_14143_, _14142_, _14141_);
  and _22495_ (_14144_, _14082_, _14107_);
  and _22496_ (_14145_, _14140_, _11669_);
  and _22497_ (_14146_, _14145_, _14144_);
  nor _22498_ (_14147_, _14146_, _14143_);
  nand _22499_ (_14148_, _14140_, _14100_);
  and _22500_ (_14149_, _14139_, _14101_);
  and _22501_ (_14150_, _14149_, _14091_);
  and _22502_ (_14151_, _14139_, _14103_);
  and _22503_ (_14152_, _14151_, _14101_);
  nor _22504_ (_14153_, _14152_, _14150_);
  and _22505_ (_14154_, _14144_, _14141_);
  and _22506_ (_14155_, _14139_, _14094_);
  and _22507_ (_14156_, _14155_, _14101_);
  nor _22508_ (_14157_, _14156_, _14154_);
  and _22509_ (_14158_, _14157_, _14153_);
  and _22510_ (_14159_, _14158_, _14148_);
  and _22511_ (_14160_, _14159_, _14147_);
  nand _22512_ (_14161_, _14160_, _14138_);
  and _22513_ (_14162_, _14143_, _12008_);
  and _22514_ (_14163_, _14149_, _14103_);
  and _22515_ (_14164_, _14163_, _08975_);
  nor _22516_ (_14165_, _14164_, _14162_);
  nor _22517_ (_14166_, _14165_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not _22518_ (_14167_, _14166_);
  not _22519_ (_14168_, _06676_);
  nor _22520_ (_14169_, _14114_, _14168_);
  nand _22521_ (_14170_, _14169_, _11789_);
  nand _22522_ (_14171_, _14146_, _08025_);
  and _22523_ (_14172_, _14171_, _14170_);
  and _22524_ (_14173_, _14172_, _11928_);
  and _22525_ (_14174_, _14173_, _14167_);
  nand _22526_ (_14175_, _14174_, _14161_);
  and _22527_ (_14176_, _14175_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  and _22528_ (_14178_, _14150_, _08975_);
  and _22529_ (_14179_, _14088_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  and _22530_ (_14181_, _14084_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  or _22531_ (_14183_, _14181_, _14179_);
  and _22532_ (_14184_, _14096_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  and _22533_ (_14185_, _14093_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  or _22534_ (_14186_, _14185_, _14184_);
  or _22535_ (_14187_, _14186_, _14183_);
  and _22536_ (_14188_, _14102_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and _22537_ (_14189_, _14105_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  or _22538_ (_14190_, _14189_, _14188_);
  and _22539_ (_14191_, _14110_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and _22540_ (_14192_, _14116_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  or _22541_ (_14193_, _14192_, _14191_);
  or _22542_ (_14194_, _14193_, _14190_);
  or _22543_ (_14195_, _14194_, _14187_);
  and _22544_ (_14196_, _14120_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and _22545_ (_14198_, _14122_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  or _22546_ (_14199_, _14198_, _14196_);
  and _22547_ (_14200_, _14124_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and _22548_ (_14201_, _14125_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  or _22549_ (_14202_, _14201_, _14200_);
  or _22550_ (_14203_, _14202_, _14199_);
  and _22551_ (_14204_, _14130_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  and _22552_ (_14205_, _14131_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  or _22553_ (_14206_, _14205_, _14204_);
  and _22554_ (_14208_, _14133_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and _22555_ (_14209_, _14134_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  or _22556_ (_14210_, _14209_, _14208_);
  or _22557_ (_14211_, _14210_, _14206_);
  or _22558_ (_14212_, _14211_, _14203_);
  or _22559_ (_14213_, _14212_, _14195_);
  and _22560_ (_14214_, _14146_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and _22561_ (_14215_, _14143_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  or _22562_ (_14216_, _14215_, _14214_);
  and _22563_ (_14217_, _14154_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and _22564_ (_14218_, _14156_, _11775_);
  or _22565_ (_14219_, _14218_, _14217_);
  and _22566_ (_14220_, _14150_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and _22567_ (_14221_, _14152_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or _22568_ (_14222_, _14221_, _14220_);
  or _22569_ (_14223_, _14222_, _14219_);
  and _22570_ (_14224_, _14140_, _14101_);
  and _22571_ (_14225_, _11437_, _11965_);
  or _22572_ (_14226_, _14225_, _11513_);
  nor _22573_ (_14227_, _14226_, _11512_);
  and _22574_ (_14228_, _11528_, _11374_);
  not _22575_ (_14229_, _14228_);
  nor _22576_ (_14230_, _11536_, _11428_);
  and _22577_ (_14231_, _14230_, _14229_);
  and _22578_ (_14232_, _11493_, _11430_);
  nor _22579_ (_14233_, _14232_, _11524_);
  and _22580_ (_14234_, _11519_, _11374_);
  nor _22581_ (_14235_, _14234_, _11503_);
  and _22582_ (_14236_, _14235_, _14233_);
  nor _22583_ (_14237_, _11352_, _11372_);
  and _22584_ (_14238_, _14237_, _11364_);
  and _22585_ (_14239_, _11976_, _11412_);
  and _22586_ (_14240_, _11407_, _11406_);
  or _22587_ (_14241_, _14240_, _14239_);
  nor _22588_ (_14242_, _14241_, _14238_);
  and _22589_ (_14243_, _14242_, _14236_);
  and _22590_ (_14244_, _14243_, _14231_);
  and _22591_ (_14245_, _14244_, _11499_);
  and _22592_ (_14246_, _14245_, _14227_);
  nor _22593_ (_14247_, _14246_, _11343_);
  or _22594_ (_14248_, _14247_, p0_in[6]);
  not _22595_ (_14249_, _14247_);
  or _22596_ (_14250_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and _22597_ (_14251_, _14250_, _14248_);
  and _22598_ (_14252_, _14251_, _14224_);
  and _22599_ (_14253_, _14129_, _14140_);
  or _22600_ (_14254_, _14247_, p1_in[6]);
  or _22601_ (_14255_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and _22602_ (_14256_, _14255_, _14254_);
  and _22603_ (_14258_, _14256_, _14253_);
  or _22604_ (_14259_, _14258_, _14252_);
  and _22605_ (_14260_, _14112_, _14140_);
  or _22606_ (_14261_, _14247_, p3_in[6]);
  or _22607_ (_14262_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and _22608_ (_14263_, _14262_, _14261_);
  and _22609_ (_14264_, _14263_, _14260_);
  and _22610_ (_14265_, _14109_, _14140_);
  or _22611_ (_14266_, _14247_, p2_in[6]);
  or _22612_ (_14267_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and _22613_ (_14268_, _14267_, _14266_);
  and _22614_ (_14269_, _14268_, _14265_);
  or _22615_ (_14270_, _14269_, _14264_);
  or _22616_ (_14271_, _14270_, _14259_);
  or _22617_ (_14272_, _14271_, _14223_);
  or _22618_ (_14273_, _14272_, _14216_);
  or _22619_ (_14274_, _14273_, _14213_);
  and _22620_ (_14275_, _14274_, _14174_);
  or _22621_ (_14276_, _14275_, _14178_);
  or _22622_ (_14277_, _14276_, _14176_);
  nand _22623_ (_14278_, _14178_, _09045_);
  and _22624_ (_14279_, _14278_, _06444_);
  and _22625_ (_13364_, _14279_, _14277_);
  and _22626_ (_14280_, _07189_, _07070_);
  and _22627_ (_14281_, _10497_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  or _22628_ (_14282_, _14281_, _14280_);
  and _22629_ (_13387_, _14282_, _06444_);
  and _22630_ (_13422_, _07757_, _06444_);
  and _22631_ (_14283_, _14175_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  and _22632_ (_14284_, _14088_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and _22633_ (_14285_, _14084_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or _22634_ (_14286_, _14285_, _14284_);
  and _22635_ (_14287_, _14096_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and _22636_ (_14288_, _14093_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  or _22637_ (_14289_, _14288_, _14287_);
  or _22638_ (_14290_, _14289_, _14286_);
  and _22639_ (_14291_, _14102_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and _22640_ (_14292_, _14105_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  or _22641_ (_14293_, _14292_, _14291_);
  and _22642_ (_14294_, _14110_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and _22643_ (_14296_, _14116_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  or _22644_ (_14297_, _14296_, _14294_);
  or _22645_ (_14298_, _14297_, _14293_);
  or _22646_ (_14299_, _14298_, _14290_);
  and _22647_ (_14300_, _14120_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  and _22648_ (_14301_, _14122_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  or _22649_ (_14302_, _14301_, _14300_);
  and _22650_ (_14303_, _14125_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  and _22651_ (_14304_, _14124_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or _22652_ (_14305_, _14304_, _14303_);
  or _22653_ (_14306_, _14305_, _14302_);
  and _22654_ (_14307_, _14131_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  and _22655_ (_14308_, _14130_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  or _22656_ (_14309_, _14308_, _14307_);
  and _22657_ (_14310_, _14133_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and _22658_ (_14311_, _14134_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  or _22659_ (_14312_, _14311_, _14310_);
  or _22660_ (_14313_, _14312_, _14309_);
  or _22661_ (_14314_, _14313_, _14306_);
  or _22662_ (_14315_, _14314_, _14299_);
  and _22663_ (_14316_, _14154_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and _22664_ (_14317_, _14156_, _11700_);
  or _22665_ (_14318_, _14317_, _14316_);
  and _22666_ (_14319_, _14150_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and _22667_ (_14320_, _14152_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or _22668_ (_14321_, _14320_, _14319_);
  or _22669_ (_14322_, _14321_, _14318_);
  or _22670_ (_14323_, _14247_, p0_in[3]);
  or _22671_ (_14324_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and _22672_ (_14325_, _14324_, _14323_);
  and _22673_ (_14326_, _14325_, _14224_);
  or _22674_ (_14327_, _14247_, p1_in[3]);
  or _22675_ (_14328_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and _22676_ (_14329_, _14328_, _14327_);
  and _22677_ (_14330_, _14329_, _14253_);
  or _22678_ (_14331_, _14330_, _14326_);
  or _22679_ (_14332_, _14247_, p2_in[3]);
  or _22680_ (_14333_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and _22681_ (_14334_, _14333_, _14332_);
  and _22682_ (_14335_, _14334_, _14265_);
  or _22683_ (_14336_, _14247_, p3_in[3]);
  or _22684_ (_14337_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and _22685_ (_14338_, _14337_, _14336_);
  and _22686_ (_14339_, _14338_, _14260_);
  or _22687_ (_14340_, _14339_, _14335_);
  or _22688_ (_14341_, _14340_, _14331_);
  or _22689_ (_14342_, _14341_, _14322_);
  and _22690_ (_14343_, _14143_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and _22691_ (_14344_, _14146_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or _22692_ (_14345_, _14344_, _14343_);
  or _22693_ (_14347_, _14345_, _14342_);
  or _22694_ (_14349_, _14347_, _14315_);
  and _22695_ (_14350_, _14349_, _14174_);
  or _22696_ (_14351_, _14350_, _14178_);
  or _22697_ (_14352_, _14351_, _14283_);
  not _22698_ (_14353_, _14178_);
  or _22699_ (_14354_, _14353_, _08308_);
  and _22700_ (_14355_, _14354_, _06444_);
  and _22701_ (_13519_, _14355_, _14352_);
  and _22702_ (_14357_, _14175_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  and _22703_ (_14358_, _14084_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and _22704_ (_14359_, _14088_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or _22705_ (_14360_, _14359_, _14358_);
  and _22706_ (_14361_, _14096_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and _22707_ (_14362_, _14093_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  or _22708_ (_14363_, _14362_, _14361_);
  or _22709_ (_14364_, _14363_, _14360_);
  and _22710_ (_14366_, _14102_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and _22711_ (_14367_, _14105_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  or _22712_ (_14368_, _14367_, _14366_);
  and _22713_ (_14369_, _14110_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and _22714_ (_14370_, _14116_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or _22715_ (_14371_, _14370_, _14369_);
  or _22716_ (_14372_, _14371_, _14368_);
  or _22717_ (_14373_, _14372_, _14364_);
  and _22718_ (_14374_, _14122_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and _22719_ (_14375_, _14120_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  or _22720_ (_14376_, _14375_, _14374_);
  and _22721_ (_14377_, _14125_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  and _22722_ (_14378_, _14124_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  or _22723_ (_14379_, _14378_, _14377_);
  or _22724_ (_14380_, _14379_, _14376_);
  and _22725_ (_14381_, _14131_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  and _22726_ (_14382_, _14130_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  or _22727_ (_14383_, _14382_, _14381_);
  and _22728_ (_14384_, _14133_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _22729_ (_14385_, _14134_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  or _22730_ (_14386_, _14385_, _14384_);
  or _22731_ (_14387_, _14386_, _14383_);
  or _22732_ (_14388_, _14387_, _14380_);
  or _22733_ (_14389_, _14388_, _14373_);
  and _22734_ (_14390_, _14146_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and _22735_ (_14391_, _14143_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or _22736_ (_14393_, _14391_, _14390_);
  and _22737_ (_14394_, _14150_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and _22738_ (_14395_, _14152_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or _22739_ (_14396_, _14395_, _14394_);
  and _22740_ (_14397_, _14154_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and _22741_ (_14398_, _14156_, _11914_);
  or _22742_ (_14399_, _14398_, _14397_);
  or _22743_ (_14400_, _14399_, _14396_);
  or _22744_ (_14401_, _14247_, p2_in[2]);
  or _22745_ (_14402_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and _22746_ (_14403_, _14402_, _14401_);
  and _22747_ (_14404_, _14403_, _14265_);
  or _22748_ (_14405_, _14247_, p3_in[2]);
  or _22749_ (_14406_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and _22750_ (_14407_, _14406_, _14405_);
  and _22751_ (_14408_, _14407_, _14260_);
  or _22752_ (_14409_, _14408_, _14404_);
  or _22753_ (_14410_, _14247_, p0_in[2]);
  or _22754_ (_14411_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and _22755_ (_14412_, _14411_, _14410_);
  and _22756_ (_14413_, _14412_, _14224_);
  or _22757_ (_14414_, _14247_, p1_in[2]);
  or _22758_ (_14415_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and _22759_ (_14417_, _14415_, _14414_);
  and _22760_ (_14418_, _14417_, _14253_);
  or _22761_ (_14419_, _14418_, _14413_);
  or _22762_ (_14420_, _14419_, _14409_);
  or _22763_ (_14421_, _14420_, _14400_);
  or _22764_ (_14422_, _14421_, _14393_);
  or _22765_ (_14423_, _14422_, _14389_);
  and _22766_ (_14424_, _14423_, _14174_);
  or _22767_ (_14425_, _14424_, _14178_);
  or _22768_ (_14426_, _14425_, _14357_);
  nand _22769_ (_14427_, _14178_, _09138_);
  and _22770_ (_14428_, _14427_, _06444_);
  and _22771_ (_13525_, _14428_, _14426_);
  and _22772_ (_14429_, _14175_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  and _22773_ (_14430_, _14084_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and _22774_ (_14431_, _14088_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or _22775_ (_14432_, _14431_, _14430_);
  and _22776_ (_14433_, _14096_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and _22777_ (_14434_, _14093_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  or _22778_ (_14435_, _14434_, _14433_);
  or _22779_ (_14436_, _14435_, _14432_);
  and _22780_ (_14437_, _14102_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  and _22781_ (_14438_, _14105_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  or _22782_ (_14439_, _14438_, _14437_);
  and _22783_ (_14440_, _14110_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and _22784_ (_14441_, _14116_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  or _22785_ (_14442_, _14441_, _14440_);
  or _22786_ (_14443_, _14442_, _14439_);
  or _22787_ (_14444_, _14443_, _14436_);
  and _22788_ (_14445_, _14120_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  and _22789_ (_14446_, _14122_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  or _22790_ (_14447_, _14446_, _14445_);
  and _22791_ (_14448_, _14125_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and _22792_ (_14449_, _14124_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  or _22793_ (_14450_, _14449_, _14448_);
  or _22794_ (_14451_, _14450_, _14447_);
  and _22795_ (_14452_, _14131_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  and _22796_ (_14453_, _14130_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  or _22797_ (_14454_, _14453_, _14452_);
  and _22798_ (_14455_, _14133_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and _22799_ (_14456_, _14134_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  or _22800_ (_14457_, _14456_, _14455_);
  or _22801_ (_14458_, _14457_, _14454_);
  or _22802_ (_14459_, _14458_, _14451_);
  or _22803_ (_14460_, _14459_, _14444_);
  and _22804_ (_14461_, _14154_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and _22805_ (_14462_, _14156_, _11803_);
  or _22806_ (_14463_, _14462_, _14461_);
  and _22807_ (_14464_, _14150_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and _22808_ (_14465_, _14152_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or _22809_ (_14466_, _14465_, _14464_);
  or _22810_ (_14467_, _14466_, _14463_);
  or _22811_ (_14468_, _14247_, p3_in[1]);
  or _22812_ (_14469_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and _22813_ (_14470_, _14469_, _14468_);
  and _22814_ (_14471_, _14470_, _14260_);
  or _22815_ (_14472_, _14247_, p2_in[1]);
  or _22816_ (_14473_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and _22817_ (_14474_, _14473_, _14472_);
  and _22818_ (_14475_, _14474_, _14265_);
  or _22819_ (_14476_, _14475_, _14471_);
  or _22820_ (_14477_, _14247_, p0_in[1]);
  or _22821_ (_14478_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and _22822_ (_14479_, _14478_, _14477_);
  and _22823_ (_14480_, _14479_, _14224_);
  or _22824_ (_14481_, _14247_, p1_in[1]);
  or _22825_ (_14482_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and _22826_ (_14483_, _14482_, _14481_);
  and _22827_ (_14484_, _14483_, _14253_);
  or _22828_ (_14485_, _14484_, _14480_);
  or _22829_ (_14486_, _14485_, _14476_);
  or _22830_ (_14487_, _14486_, _14467_);
  and _22831_ (_14488_, _14146_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and _22832_ (_14489_, _14143_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  or _22833_ (_14490_, _14489_, _14488_);
  or _22834_ (_14491_, _14490_, _14487_);
  or _22835_ (_14492_, _14491_, _14460_);
  and _22836_ (_14493_, _14492_, _14174_);
  or _22837_ (_14494_, _14493_, _14178_);
  or _22838_ (_14495_, _14494_, _14429_);
  nor _22839_ (_14496_, _14178_, rst);
  and _22840_ (_14497_, _07959_, _06444_);
  or _22841_ (_14498_, _14497_, _14496_);
  and _22842_ (_13548_, _14498_, _14495_);
  nor _22843_ (_14499_, _07300_, _06449_);
  and _22844_ (_14500_, _06449_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  or _22845_ (_14501_, _14500_, _14499_);
  and _22846_ (_13551_, _14501_, _06444_);
  or _22847_ (_14502_, _11137_, _08980_);
  or _22848_ (_14503_, _08982_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and _22849_ (_14504_, _14503_, _06444_);
  and _22850_ (_13589_, _14504_, _14502_);
  and _22851_ (_14505_, _11137_, _09157_);
  and _22852_ (_14506_, _09158_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or _22853_ (_14507_, _14506_, _08975_);
  or _22854_ (_14508_, _14507_, _14505_);
  or _22855_ (_14509_, _11177_, _09208_);
  and _22856_ (_14510_, _14509_, _06444_);
  and _22857_ (_13596_, _14510_, _14508_);
  and _22858_ (_14511_, _07402_, _06434_);
  and _22859_ (_14512_, _14511_, _06440_);
  nand _22860_ (_14513_, _14512_, _11589_);
  or _22861_ (_14514_, _14512_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and _22862_ (_14516_, _14514_, _06444_);
  and _22863_ (_13634_, _14516_, _14513_);
  nand _22864_ (_14517_, _14512_, _07069_);
  or _22865_ (_14518_, _14512_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _22866_ (_14519_, _14518_, _06444_);
  and _22867_ (_13637_, _14519_, _14517_);
  or _22868_ (_14520_, _14512_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  and _22869_ (_14521_, _14520_, _06444_);
  nand _22870_ (_14523_, _14512_, _07300_);
  and _22871_ (_13661_, _14523_, _14521_);
  or _22872_ (_14525_, _14512_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and _22873_ (_14526_, _14525_, _06444_);
  nand _22874_ (_14527_, _14512_, _07188_);
  and _22875_ (_13665_, _14527_, _14526_);
  not _22876_ (_14528_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  nor _22877_ (_14529_, _14512_, _14528_);
  and _22878_ (_14530_, _14512_, _09527_);
  or _22879_ (_14531_, _14530_, _14529_);
  and _22880_ (_13675_, _14531_, _06444_);
  and _22881_ (_14532_, _07402_, _06984_);
  nand _22882_ (_14533_, _14532_, _06666_);
  and _22883_ (_14534_, _14528_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  not _22884_ (_14535_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _22885_ (_14536_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _14535_);
  or _22886_ (_14537_, _14536_, _14534_);
  not _22887_ (_14538_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _22888_ (_14539_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and _22889_ (_14540_, _14539_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _22890_ (_14541_, _14540_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  not _22891_ (_14542_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and _22892_ (_14543_, _14542_, \oc8051_top_1.oc8051_sfr1.pres_ow );
  not _22893_ (_14545_, t0_i);
  and _22894_ (_14546_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and _22895_ (_14547_, _14546_, _14545_);
  or _22896_ (_14548_, _14547_, _14543_);
  and _22897_ (_14549_, _14548_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and _22898_ (_14550_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and _22899_ (_14551_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  and _22900_ (_14552_, _14551_, _14550_);
  and _22901_ (_14553_, _14552_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and _22902_ (_14554_, _14553_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and _22903_ (_00001_, _14554_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and _22904_ (_00002_, _00001_, _14549_);
  and _22905_ (_00003_, _00002_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and _22906_ (_00004_, _00003_, _14541_);
  and _22907_ (_00005_, _00004_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _22908_ (_00006_, _00005_, _14535_);
  nor _22909_ (_00007_, _00006_, _14538_);
  and _22910_ (_00008_, _00006_, _14538_);
  or _22911_ (_00009_, _00008_, _00007_);
  and _22912_ (_00010_, _00009_, _14537_);
  and _22913_ (_00011_, \oc8051_top_1.oc8051_sfr1.pres_ow , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and _22914_ (_00012_, _00011_, _14541_);
  and _22915_ (_00013_, _00012_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or _22916_ (_00014_, _00013_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _22917_ (_00015_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _22918_ (_00016_, _00013_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  not _22919_ (_00017_, _00016_);
  and _22920_ (_00018_, _00017_, _00015_);
  and _22921_ (_00019_, _00018_, _00014_);
  and _22922_ (_00020_, _14549_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and _22923_ (_00021_, _00020_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and _22924_ (_00022_, _00021_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  and _22925_ (_00023_, _00022_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  and _22926_ (_00024_, _00023_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and _22927_ (_00025_, _00024_, _14541_);
  and _22928_ (_00026_, _00025_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or _22929_ (_00027_, _00026_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nor _22930_ (_00028_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  not _22931_ (_00029_, _00028_);
  and _22932_ (_00030_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _22933_ (_00031_, _00030_, _14541_);
  and _22934_ (_00032_, _00031_, _00024_);
  nor _22935_ (_00033_, _00032_, _00029_);
  and _22936_ (_00034_, _00033_, _00027_);
  or _22937_ (_00035_, _00034_, _00019_);
  or _22938_ (_00036_, _00035_, _00010_);
  or _22939_ (_00037_, _00036_, _14532_);
  and _22940_ (_00039_, _09483_, _07402_);
  not _22941_ (_00040_, _00039_);
  and _22942_ (_00041_, _00040_, _00037_);
  and _22943_ (_00042_, _00041_, _14533_);
  and _22944_ (_00043_, _00039_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  or _22945_ (_00044_, _00043_, _00042_);
  and _22946_ (_13690_, _00044_, _06444_);
  nand _22947_ (_00045_, _14532_, _10494_);
  and _22948_ (_00046_, _00032_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or _22949_ (_00047_, _00032_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nand _22950_ (_00048_, _00047_, _00028_);
  nor _22951_ (_00049_, _00048_, _00046_);
  and _22952_ (_00050_, _00031_, _00003_);
  or _22953_ (_00051_, _00050_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and _22954_ (_00052_, _00050_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  not _22955_ (_00053_, _00052_);
  and _22956_ (_00054_, _00053_, _14536_);
  and _22957_ (_00055_, _00054_, _00051_);
  and _22958_ (_00057_, _00016_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or _22959_ (_00058_, _00057_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nand _22960_ (_00059_, _00057_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and _22961_ (_00060_, _00059_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _22962_ (_00062_, _00060_, _00058_);
  or _22963_ (_00063_, _00062_, _00055_);
  or _22964_ (_00065_, _00063_, _00049_);
  or _22965_ (_00067_, _00065_, _14532_);
  and _22966_ (_00068_, _00067_, _00040_);
  and _22967_ (_00069_, _00068_, _00045_);
  and _22968_ (_00070_, _00039_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or _22969_ (_00071_, _00070_, _00069_);
  and _22970_ (_13693_, _00071_, _06444_);
  nand _22971_ (_00072_, _14532_, _09526_);
  or _22972_ (_00073_, _00024_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and _22973_ (_00074_, _00024_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nor _22974_ (_00075_, _00074_, _00029_);
  and _22975_ (_00076_, _00075_, _00073_);
  not _22976_ (_00077_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and _22977_ (_00078_, _00003_, _14535_);
  and _22978_ (_00079_, _00078_, _00077_);
  nor _22979_ (_00080_, _00078_, _00077_);
  or _22980_ (_00081_, _00080_, _00079_);
  and _22981_ (_00083_, _00081_, _14537_);
  and _22982_ (_00084_, _00011_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or _22983_ (_00086_, _00011_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand _22984_ (_00087_, _00086_, _00015_);
  nor _22985_ (_00089_, _00087_, _00084_);
  or _22986_ (_00090_, _00089_, _00083_);
  or _22987_ (_00091_, _00090_, _00076_);
  or _22988_ (_00092_, _00091_, _14532_);
  and _22989_ (_00093_, _00092_, _00072_);
  or _22990_ (_00094_, _00093_, _00039_);
  nand _22991_ (_00095_, _00039_, _00077_);
  and _22992_ (_00096_, _00095_, _06444_);
  and _22993_ (_13714_, _00096_, _00094_);
  nand _22994_ (_00097_, _00039_, _10494_);
  or _22995_ (_00098_, _00028_, _14532_);
  and _22996_ (_00099_, _00098_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and _22997_ (_00100_, _00024_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  or _22998_ (_00101_, _00100_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  nor _22999_ (_00102_, _00028_, _00002_);
  and _23000_ (_00103_, _00102_, _00101_);
  and _23001_ (_00104_, _14534_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and _23002_ (_00105_, _00104_, _00003_);
  nor _23003_ (_00106_, _00105_, _00103_);
  nor _23004_ (_00107_, _00106_, _14532_);
  or _23005_ (_00108_, _00107_, _00099_);
  or _23006_ (_00109_, _00108_, _00039_);
  and _23007_ (_00110_, _00109_, _06444_);
  and _23008_ (_13721_, _00110_, _00097_);
  nand _23009_ (_00111_, _00039_, _06666_);
  and _23010_ (_00112_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and _23011_ (_00113_, _00112_, _14549_);
  and _23012_ (_00114_, _00113_, _14553_);
  and _23013_ (_00115_, _14534_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and _23014_ (_00116_, _00115_, _00114_);
  nand _23015_ (_00117_, _00116_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nor _23016_ (_00118_, _00028_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  nand _23017_ (_00119_, _00118_, _00024_);
  and _23018_ (_00120_, _00119_, _00117_);
  nor _23019_ (_00121_, _00120_, _14532_);
  not _23020_ (_00122_, _00024_);
  or _23021_ (_00123_, _00098_, _00122_);
  and _23022_ (_00124_, _00123_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  or _23023_ (_00125_, _00124_, _00121_);
  or _23024_ (_00126_, _00125_, _00039_);
  and _23025_ (_00127_, _00126_, _06444_);
  and _23026_ (_13727_, _00127_, _00111_);
  nand _23027_ (_00128_, _14532_, _11589_);
  and _23028_ (_00129_, _00003_, _14539_);
  or _23029_ (_00130_, _00129_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nand _23030_ (_00131_, _00129_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _23031_ (_00132_, _00131_, _14536_);
  and _23032_ (_00133_, _00132_, _00130_);
  not _23033_ (_00134_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _23034_ (_00135_, _14553_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and _23035_ (_00136_, _14549_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and _23036_ (_00137_, _00136_, _00135_);
  and _23037_ (_00138_, _00137_, _00134_);
  nor _23038_ (_00139_, _00137_, _00134_);
  or _23039_ (_00140_, _00139_, _00138_);
  and _23040_ (_00141_, _00140_, _00028_);
  and _23041_ (_00142_, _00011_, _14539_);
  and _23042_ (_00144_, _00142_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  nand _23043_ (_00146_, _00144_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  or _23044_ (_00148_, _00144_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _23045_ (_00150_, _00148_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _23046_ (_00152_, _00150_, _00146_);
  or _23047_ (_00154_, _00152_, _00141_);
  or _23048_ (_00155_, _00154_, _00133_);
  or _23049_ (_00156_, _00155_, _14532_);
  and _23050_ (_00157_, _00156_, _00040_);
  and _23051_ (_00158_, _00157_, _00128_);
  and _23052_ (_00159_, _00039_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  or _23053_ (_00160_, _00159_, _00158_);
  and _23054_ (_13739_, _00160_, _06444_);
  nand _23055_ (_00161_, _14532_, _07188_);
  nor _23056_ (_00163_, _00025_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nor _23057_ (_00165_, _00163_, _00026_);
  and _23058_ (_00167_, _00165_, _00028_);
  or _23059_ (_00168_, _00004_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  not _23060_ (_00170_, _00005_);
  and _23061_ (_00171_, _00170_, _14536_);
  and _23062_ (_00173_, _00171_, _00168_);
  and _23063_ (_00174_, _14534_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nor _23064_ (_00175_, _00012_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nor _23065_ (_00176_, _00175_, _00013_);
  and _23066_ (_00178_, _00176_, _00015_);
  or _23067_ (_00179_, _00178_, _00174_);
  or _23068_ (_00180_, _00179_, _00173_);
  or _23069_ (_00181_, _00180_, _00167_);
  or _23070_ (_00182_, _00181_, _14532_);
  and _23071_ (_00183_, _00182_, _00040_);
  and _23072_ (_00184_, _00183_, _00161_);
  and _23073_ (_00185_, _00039_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or _23074_ (_00186_, _00185_, _00184_);
  and _23075_ (_13742_, _00186_, _06444_);
  nand _23076_ (_00187_, _14532_, _07300_);
  and _23077_ (_00188_, _00024_, _14540_);
  or _23078_ (_00190_, _00188_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  nor _23079_ (_00192_, _00025_, _00029_);
  and _23080_ (_00193_, _00192_, _00190_);
  and _23081_ (_00194_, _00078_, _14540_);
  or _23082_ (_00195_, _00194_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  not _23083_ (_00196_, _00004_);
  or _23084_ (_00197_, _00196_, _14534_);
  and _23085_ (_00198_, _00197_, _14537_);
  and _23086_ (_00199_, _00198_, _00195_);
  and _23087_ (_00200_, _00011_, _14540_);
  or _23088_ (_00201_, _00200_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  not _23089_ (_00202_, _00012_);
  and _23090_ (_00203_, _00015_, _00202_);
  and _23091_ (_00204_, _00203_, _00201_);
  or _23092_ (_00206_, _00204_, _00199_);
  or _23093_ (_00207_, _00206_, _00193_);
  or _23094_ (_00208_, _00207_, _14532_);
  and _23095_ (_00209_, _00208_, _00040_);
  and _23096_ (_00210_, _00209_, _00187_);
  and _23097_ (_00212_, _00039_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  or _23098_ (_00213_, _00212_, _00210_);
  and _23099_ (_13745_, _00213_, _06444_);
  not _23100_ (_00214_, _00074_);
  nor _23101_ (_00215_, _00214_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and _23102_ (_00216_, _00214_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  or _23103_ (_00217_, _00216_, _00215_);
  and _23104_ (_00218_, _00217_, _00028_);
  or _23105_ (_00219_, _00084_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  not _23106_ (_00220_, _00142_);
  and _23107_ (_00221_, _00015_, _00220_);
  and _23108_ (_00222_, _00221_, _00219_);
  and _23109_ (_00223_, _00003_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and _23110_ (_00224_, _00223_, _14535_);
  or _23111_ (_00225_, _00224_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  not _23112_ (_00226_, _00129_);
  and _23113_ (_00227_, _00226_, _14536_);
  or _23114_ (_00228_, _00227_, _14534_);
  and _23115_ (_00229_, _00228_, _00225_);
  or _23116_ (_00230_, _00229_, _00222_);
  or _23117_ (_00231_, _00230_, _00218_);
  or _23118_ (_00232_, _00231_, _14532_);
  nand _23119_ (_00233_, _14532_, _07069_);
  and _23120_ (_00234_, _00233_, _00040_);
  and _23121_ (_00235_, _00234_, _00232_);
  and _23122_ (_00236_, _00039_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  or _23123_ (_00237_, _00236_, _00235_);
  and _23124_ (_13747_, _00237_, _06444_);
  nor _23125_ (_00238_, _06430_, _06418_);
  and _23126_ (_00240_, _00238_, _06406_);
  and _23127_ (_00241_, _13902_, _00240_);
  nand _23128_ (_00242_, _00241_, _06930_);
  or _23129_ (_00243_, _00241_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  and _23130_ (_00244_, _00243_, _13907_);
  and _23131_ (_00245_, _00244_, _00242_);
  nor _23132_ (_00246_, _13907_, _10494_);
  or _23133_ (_00248_, _00246_, _00245_);
  and _23134_ (_13754_, _00248_, _06444_);
  and _23135_ (_00249_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and _23136_ (_00250_, _12223_, \oc8051_top_1.oc8051_rom1.data_o [25]);
  or _23137_ (_00251_, _00250_, _00249_);
  and _23138_ (_13783_, _00251_, _06444_);
  and _23139_ (_00253_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and _23140_ (_00254_, _12223_, \oc8051_top_1.oc8051_rom1.data_o [27]);
  or _23141_ (_00255_, _00254_, _00253_);
  and _23142_ (_13805_, _00255_, _06444_);
  nor _23143_ (_00257_, _00022_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  nor _23144_ (_00258_, _00257_, _00023_);
  and _23145_ (_00259_, _00116_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  nor _23146_ (_00260_, _00259_, _00258_);
  nor _23147_ (_00261_, _00260_, _14532_);
  and _23148_ (_00262_, _14532_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  or _23149_ (_00263_, _00262_, _00261_);
  and _23150_ (_00264_, _00263_, _00040_);
  nor _23151_ (_00265_, _00040_, _07300_);
  or _23152_ (_00266_, _00265_, _00264_);
  and _23153_ (_13829_, _00266_, _06444_);
  nand _23154_ (_00267_, _00039_, _07188_);
  nor _23155_ (_00268_, _00023_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  nor _23156_ (_00269_, _00268_, _00024_);
  and _23157_ (_00270_, _00174_, _00003_);
  nor _23158_ (_00271_, _00270_, _00269_);
  nor _23159_ (_00273_, _00271_, _14532_);
  and _23160_ (_00275_, _14532_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  or _23161_ (_00277_, _00275_, _00273_);
  or _23162_ (_00279_, _00277_, _00039_);
  and _23163_ (_00281_, _00279_, _06444_);
  and _23164_ (_13831_, _00281_, _00267_);
  nor _23165_ (_00283_, _00021_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  nor _23166_ (_00284_, _00283_, _00022_);
  and _23167_ (_00285_, _00116_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nor _23168_ (_00286_, _00285_, _00284_);
  nor _23169_ (_00288_, _00286_, _14532_);
  and _23170_ (_00289_, _14532_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  or _23171_ (_00290_, _00289_, _00288_);
  and _23172_ (_00291_, _00290_, _00040_);
  nor _23173_ (_00292_, _00040_, _11589_);
  or _23174_ (_00293_, _00292_, _00291_);
  and _23175_ (_13834_, _00293_, _06444_);
  or _23176_ (_00294_, _14512_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and _23177_ (_00296_, _00294_, _06444_);
  nand _23178_ (_00297_, _14512_, _10494_);
  and _23179_ (_13839_, _00297_, _00296_);
  or _23180_ (_00298_, _14512_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and _23181_ (_00300_, _00298_, _06444_);
  nand _23182_ (_00301_, _14512_, _06666_);
  and _23183_ (_13844_, _00301_, _00300_);
  and _23184_ (_00302_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and _23185_ (_00303_, _12223_, \oc8051_top_1.oc8051_rom1.data_o [26]);
  or _23186_ (_00304_, _00303_, _00302_);
  and _23187_ (_13897_, _00304_, _06444_);
  nor _23188_ (_00305_, _14549_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  nor _23189_ (_00306_, _00305_, _00020_);
  and _23190_ (_00307_, _00116_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nor _23191_ (_00308_, _00307_, _00306_);
  nor _23192_ (_00309_, _00308_, _14532_);
  and _23193_ (_00310_, _14532_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  or _23194_ (_00311_, _00310_, _00309_);
  and _23195_ (_00312_, _00311_, _00040_);
  and _23196_ (_00313_, _00039_, _09527_);
  or _23197_ (_00314_, _00313_, _00312_);
  and _23198_ (_13925_, _00314_, _06444_);
  nor _23199_ (_00315_, _00020_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  nor _23200_ (_00316_, _00315_, _00021_);
  and _23201_ (_00317_, _00116_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nor _23202_ (_00318_, _00317_, _00316_);
  nor _23203_ (_00319_, _00318_, _14532_);
  and _23204_ (_00320_, _14532_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  or _23205_ (_00321_, _00320_, _00319_);
  and _23206_ (_00322_, _00321_, _00040_);
  nor _23207_ (_00323_, _00040_, _07069_);
  or _23208_ (_00324_, _00323_, _00322_);
  and _23209_ (_13928_, _00324_, _06444_);
  and _23210_ (_00325_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and _23211_ (_00327_, _12223_, \oc8051_top_1.oc8051_rom1.data_o [31]);
  or _23212_ (_00328_, _00327_, _00325_);
  and _23213_ (_13965_, _00328_, _06444_);
  nor _23214_ (_00329_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , rst);
  and _23215_ (_13966_, _00329_, \oc8051_top_1.oc8051_memory_interface1.int_ack_buff );
  and _23216_ (_00330_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and _23217_ (_00332_, _12223_, \oc8051_top_1.oc8051_rom1.data_o [24]);
  or _23218_ (_00333_, _00332_, _00330_);
  and _23219_ (_13974_, _00333_, _06444_);
  and _23220_ (_00334_, _07402_, _06988_);
  nand _23221_ (_00335_, _00334_, _10494_);
  not _23222_ (_00336_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and _23223_ (_00337_, _00336_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  not _23224_ (_00338_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and _23225_ (_00340_, _00338_, \oc8051_top_1.oc8051_sfr1.pres_ow );
  not _23226_ (_00341_, t1_i);
  and _23227_ (_00343_, _00341_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and _23228_ (_00344_, _00343_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff );
  or _23229_ (_00346_, _00344_, _00340_);
  and _23230_ (_00347_, _00346_, _00337_);
  and _23231_ (_00348_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and _23232_ (_00349_, _00348_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and _23233_ (_00351_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and _23234_ (_00352_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  and _23235_ (_00353_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  and _23236_ (_00354_, _00353_, _00352_);
  and _23237_ (_00355_, _00354_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and _23238_ (_00356_, _00355_, _00351_);
  and _23239_ (_00357_, _00356_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and _23240_ (_00358_, _00357_, _00349_);
  and _23241_ (_00359_, _00358_, _00347_);
  or _23242_ (_00360_, _00359_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nor _23243_ (_00361_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  not _23244_ (_00362_, _00361_);
  and _23245_ (_00363_, _00359_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nor _23246_ (_00364_, _00363_, _00362_);
  not _23247_ (_00365_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and _23248_ (_00366_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _00365_);
  and _23249_ (_00367_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and _23250_ (_00369_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and _23251_ (_00370_, _00369_, _00367_);
  and _23252_ (_00372_, _00370_, _00354_);
  and _23253_ (_00373_, _00372_, _00351_);
  and _23254_ (_00374_, _00373_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and _23255_ (_00375_, _00374_, _00347_);
  and _23256_ (_00376_, _00375_, _00349_);
  nand _23257_ (_00377_, _00376_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and _23258_ (_00378_, _00377_, _00366_);
  or _23259_ (_00379_, _00378_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and _23260_ (_00380_, _00367_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and _23261_ (_00381_, _00366_, _00380_);
  or _23262_ (_00382_, _00381_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and _23263_ (_00383_, _00382_, _00379_);
  or _23264_ (_00384_, _00383_, _00364_);
  and _23265_ (_00385_, _00384_, _00360_);
  or _23266_ (_00386_, _00385_, _00334_);
  and _23267_ (_00387_, _09478_, _07402_);
  not _23268_ (_00388_, _00387_);
  and _23269_ (_00389_, _00388_, _00386_);
  and _23270_ (_00390_, _00389_, _00335_);
  and _23271_ (_00391_, _00387_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  or _23272_ (_00392_, _00391_, _00390_);
  and _23273_ (_13978_, _00392_, _06444_);
  nand _23274_ (_00393_, _00334_, _06666_);
  not _23275_ (_00394_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  not _23276_ (_00395_, _00366_);
  nor _23277_ (_00396_, _00375_, _00395_);
  not _23278_ (_00397_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and _23279_ (_00398_, _00361_, _00397_);
  and _23280_ (_00399_, _00355_, _00347_);
  and _23281_ (_00400_, _00399_, _00351_);
  nor _23282_ (_00401_, _00362_, _00400_);
  nor _23283_ (_00402_, _00401_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  not _23284_ (_00403_, _00402_);
  nor _23285_ (_00404_, _00403_, _00398_);
  not _23286_ (_00405_, _00404_);
  or _23287_ (_00406_, _00405_, _00396_);
  not _23288_ (_00407_, _00406_);
  and _23289_ (_00408_, _00407_, _00348_);
  nor _23290_ (_00409_, _00408_, _00394_);
  and _23291_ (_00410_, _00408_, _00394_);
  or _23292_ (_00411_, _00410_, _00409_);
  or _23293_ (_00412_, _00411_, _00334_);
  and _23294_ (_00413_, _00412_, _00388_);
  and _23295_ (_00414_, _00413_, _00393_);
  and _23296_ (_00415_, _00387_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  or _23297_ (_00416_, _00415_, _00414_);
  and _23298_ (_13981_, _00416_, _06444_);
  nand _23299_ (_00417_, _00334_, _07300_);
  nor _23300_ (_00418_, _00406_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and _23301_ (_00419_, _00406_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or _23302_ (_00420_, _00419_, _00418_);
  or _23303_ (_00421_, _00420_, _00334_);
  and _23304_ (_00422_, _00421_, _00388_);
  and _23305_ (_00423_, _00422_, _00417_);
  and _23306_ (_00424_, _00387_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or _23307_ (_00425_, _00424_, _00423_);
  and _23308_ (_13988_, _00425_, _06444_);
  nand _23309_ (_00426_, _00334_, _07188_);
  not _23310_ (_00427_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and _23311_ (_00428_, _00407_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nor _23312_ (_00429_, _00428_, _00427_);
  and _23313_ (_00430_, _00428_, _00427_);
  or _23314_ (_00431_, _00430_, _00429_);
  or _23315_ (_00432_, _00431_, _00334_);
  and _23316_ (_00433_, _00432_, _00426_);
  or _23317_ (_00435_, _00433_, _00387_);
  nand _23318_ (_00436_, _00387_, _00427_);
  and _23319_ (_00437_, _00436_, _06444_);
  and _23320_ (_13991_, _00437_, _00435_);
  nand _23321_ (_00438_, _00334_, _07069_);
  and _23322_ (_00439_, _00399_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and _23323_ (_00440_, _00439_, _00380_);
  nor _23324_ (_00441_, _00440_, _00395_);
  or _23325_ (_00442_, _00441_, _00403_);
  and _23326_ (_00443_, _00442_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and _23327_ (_00444_, _00439_, _00401_);
  nor _23328_ (_00445_, _00395_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and _23329_ (_00446_, _00445_, _00440_);
  or _23330_ (_00448_, _00446_, _00444_);
  or _23331_ (_00449_, _00448_, _00443_);
  or _23332_ (_00450_, _00449_, _00334_);
  and _23333_ (_00451_, _00450_, _00438_);
  or _23334_ (_00452_, _00451_, _00387_);
  or _23335_ (_00453_, _00388_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and _23336_ (_00454_, _00453_, _06444_);
  and _23337_ (_13996_, _00454_, _00452_);
  nand _23338_ (_00455_, _00334_, _11589_);
  and _23339_ (_00456_, _00406_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and _23340_ (_00457_, _00366_, _00397_);
  and _23341_ (_00458_, _00457_, _00380_);
  or _23342_ (_00459_, _00458_, _00398_);
  and _23343_ (_00460_, _00459_, _00400_);
  or _23344_ (_00461_, _00460_, _00456_);
  or _23345_ (_00462_, _00461_, _00334_);
  and _23346_ (_00463_, _00462_, _00455_);
  or _23347_ (_00464_, _00463_, _00387_);
  nand _23348_ (_00465_, _00387_, _00397_);
  and _23349_ (_00466_, _00465_, _06444_);
  and _23350_ (_14000_, _00466_, _00464_);
  not _23351_ (_00467_, \oc8051_top_1.oc8051_sfr1.prescaler [2]);
  and _23352_ (_00468_, \oc8051_top_1.oc8051_sfr1.prescaler [0], \oc8051_top_1.oc8051_sfr1.prescaler [1]);
  and _23353_ (_00469_, _00468_, _00467_);
  and _23354_ (_00470_, _00469_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  nor _23355_ (_00472_, _00468_, _00467_);
  or _23356_ (_00473_, _00472_, _00469_);
  nand _23357_ (_00474_, _00473_, _06444_);
  nor _23358_ (_14009_, _00474_, _00470_);
  or _23359_ (_00476_, \oc8051_top_1.oc8051_sfr1.prescaler [0], \oc8051_top_1.oc8051_sfr1.prescaler [1]);
  nor _23360_ (_00477_, _00468_, rst);
  and _23361_ (_14012_, _00477_, _00476_);
  and _23362_ (_00478_, _00399_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  nor _23363_ (_00479_, _00399_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  nor _23364_ (_00480_, _00479_, _00478_);
  nor _23365_ (_00481_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _00365_);
  nor _23366_ (_00482_, _00481_, _00366_);
  nor _23367_ (_00483_, _00482_, _00334_);
  and _23368_ (_00484_, _00483_, _00480_);
  not _23369_ (_00485_, _00483_);
  and _23370_ (_00486_, _00485_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and _23371_ (_00487_, _00380_, _00399_);
  and _23372_ (_00488_, _00481_, _00487_);
  nand _23373_ (_00489_, _00488_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  nor _23374_ (_00490_, _00489_, _00334_);
  or _23375_ (_00491_, _00490_, _00486_);
  or _23376_ (_00492_, _00491_, _00484_);
  and _23377_ (_00493_, _00492_, _00388_);
  nor _23378_ (_00494_, _00388_, _06666_);
  or _23379_ (_00495_, _00494_, _00493_);
  and _23380_ (_14021_, _00495_, _06444_);
  nand _23381_ (_00496_, _00387_, _10494_);
  and _23382_ (_00497_, _00478_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nor _23383_ (_00498_, _00478_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nor _23384_ (_00499_, _00498_, _00497_);
  and _23385_ (_00500_, _00499_, _00483_);
  and _23386_ (_00502_, _00485_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nand _23387_ (_00503_, _00488_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nor _23388_ (_00505_, _00503_, _00334_);
  or _23389_ (_00506_, _00505_, _00502_);
  or _23390_ (_00507_, _00506_, _00500_);
  or _23391_ (_00508_, _00507_, _00387_);
  and _23392_ (_00510_, _00508_, _06444_);
  and _23393_ (_14023_, _00510_, _00496_);
  and _23394_ (_00511_, _00347_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and _23395_ (_00512_, _00511_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  and _23396_ (_00513_, _00512_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  and _23397_ (_00514_, _00513_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nor _23398_ (_00515_, _00514_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  nor _23399_ (_00516_, _00515_, _00399_);
  and _23400_ (_00517_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  nor _23401_ (_00518_, _00517_, _00334_);
  and _23402_ (_00519_, _00518_, _00516_);
  not _23403_ (_00520_, _00518_);
  and _23404_ (_00521_, _00520_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and _23405_ (_00522_, _00481_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nand _23406_ (_00523_, _00522_, _00487_);
  nor _23407_ (_00524_, _00523_, _00334_);
  or _23408_ (_00525_, _00524_, _00521_);
  or _23409_ (_00526_, _00525_, _00519_);
  and _23410_ (_00527_, _00526_, _00388_);
  nor _23411_ (_00528_, _00388_, _07188_);
  or _23412_ (_00529_, _00528_, _00527_);
  and _23413_ (_14026_, _00529_, _06444_);
  nor _23414_ (_00530_, _00512_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  or _23415_ (_00531_, _00530_, _00513_);
  nand _23416_ (_00532_, _00531_, _00518_);
  or _23417_ (_00533_, _00518_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  and _23418_ (_00534_, _00533_, _00532_);
  and _23419_ (_00535_, _00497_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and _23420_ (_00536_, _00481_, _00535_);
  nand _23421_ (_00537_, _00536_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nor _23422_ (_00538_, _00537_, _00334_);
  or _23423_ (_00539_, _00538_, _00387_);
  or _23424_ (_00540_, _00539_, _00534_);
  nand _23425_ (_00541_, _00387_, _11589_);
  and _23426_ (_00542_, _00541_, _06444_);
  and _23427_ (_14032_, _00542_, _00540_);
  and _23428_ (_00543_, _00520_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nand _23429_ (_00545_, _00536_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nor _23430_ (_00546_, _00545_, _00334_);
  or _23431_ (_00547_, _00546_, _00543_);
  nor _23432_ (_00548_, _00513_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nor _23433_ (_00549_, _00548_, _00514_);
  and _23434_ (_00551_, _00549_, _00518_);
  or _23435_ (_00552_, _00551_, _00387_);
  or _23436_ (_00553_, _00552_, _00547_);
  nand _23437_ (_00554_, _00387_, _07300_);
  and _23438_ (_00555_, _00554_, _06444_);
  and _23439_ (_14037_, _00555_, _00553_);
  nor _23440_ (_00556_, _00511_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  or _23441_ (_00557_, _00556_, _00512_);
  nand _23442_ (_00558_, _00557_, _00518_);
  or _23443_ (_00559_, _00518_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  and _23444_ (_00560_, _00559_, _00558_);
  nand _23445_ (_00561_, _00536_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nor _23446_ (_00562_, _00561_, _00334_);
  or _23447_ (_00563_, _00562_, _00387_);
  or _23448_ (_00564_, _00563_, _00560_);
  nand _23449_ (_00565_, _00387_, _07069_);
  and _23450_ (_00566_, _00565_, _06444_);
  and _23451_ (_14040_, _00566_, _00564_);
  or _23452_ (_00567_, _00388_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and _23453_ (_00568_, _00567_, _06444_);
  or _23454_ (_00570_, _00399_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  nor _23455_ (_00571_, _00439_, _00362_);
  and _23456_ (_00573_, _00571_, _00570_);
  or _23457_ (_00574_, _00487_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and _23458_ (_00575_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  or _23459_ (_00576_, _00575_, _00441_);
  and _23460_ (_00577_, _00576_, _00574_);
  nor _23461_ (_00578_, _00577_, _00573_);
  nor _23462_ (_00579_, _00578_, _00334_);
  and _23463_ (_00580_, _00334_, _09527_);
  or _23464_ (_00581_, _00580_, _00579_);
  or _23465_ (_00582_, _00581_, _00387_);
  and _23466_ (_14047_, _00582_, _00568_);
  and _23467_ (_00583_, _08064_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  not _23468_ (_00584_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nor _23469_ (_00585_, _08064_, _00584_);
  or _23470_ (_00586_, _00585_, _00583_);
  and _23471_ (_14073_, _00586_, _06444_);
  nor _23472_ (_14177_, _11630_, rst);
  and _23473_ (_00587_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  and _23474_ (_00588_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and _23475_ (_00589_, _00588_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor _23476_ (_00590_, _00588_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor _23477_ (_00591_, _00590_, _00589_);
  or _23478_ (_00592_, _00591_, _00587_);
  and _23479_ (_14180_, _00592_, _06444_);
  not _23480_ (_00593_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  nor _23481_ (_00594_, _00587_, _00593_);
  nor _23482_ (_00595_, _00594_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and _23483_ (_00596_, _00594_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  or _23484_ (_00597_, _00596_, _00595_);
  nor _23485_ (_14182_, _00597_, rst);
  and _23486_ (_00598_, _00587_, _00593_);
  nor _23487_ (_00599_, _00598_, _00594_);
  and _23488_ (_14197_, _00599_, _06444_);
  and _23489_ (_00600_, _08064_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  not _23490_ (_00601_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  nor _23491_ (_00602_, _08064_, _00601_);
  or _23492_ (_00603_, _00602_, _00600_);
  and _23493_ (_14207_, _00603_, _06444_);
  and _23494_ (_00604_, _12011_, _08030_);
  and _23495_ (_00605_, _00604_, _07401_);
  and _23496_ (_00606_, _00605_, _06933_);
  nand _23497_ (_00607_, _00606_, _06930_);
  or _23498_ (_00609_, _00606_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and _23499_ (_00610_, _00609_, _06674_);
  and _23500_ (_00611_, _00610_, _00607_);
  and _23501_ (_00612_, _07150_, _06382_);
  nand _23502_ (_00613_, _00612_, _06978_);
  or _23503_ (_00614_, _00612_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and _23504_ (_00615_, _00614_, _06440_);
  and _23505_ (_00616_, _00615_, _00613_);
  and _23506_ (_00617_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  or _23507_ (_00618_, _00617_, rst);
  or _23508_ (_00619_, _00618_, _00616_);
  or _23509_ (_14346_, _00619_, _00611_);
  and _23510_ (_00620_, _08064_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  not _23511_ (_00621_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor _23512_ (_00622_, _08064_, _00621_);
  or _23513_ (_00623_, _00622_, _00620_);
  and _23514_ (_14348_, _00623_, _06444_);
  nand _23515_ (_00624_, _10112_, _06978_);
  or _23516_ (_00625_, _10112_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  and _23517_ (_00626_, _00625_, _06444_);
  and _23518_ (_14356_, _00626_, _00624_);
  and _23519_ (_00627_, _09373_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  or _23520_ (_14365_, _00627_, _09368_);
  and _23521_ (_00628_, _00520_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  or _23522_ (_00630_, _00347_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nor _23523_ (_00631_, _00511_, _00517_);
  and _23524_ (_00632_, _00631_, _00630_);
  and _23525_ (_00633_, _00481_, _00440_);
  nor _23526_ (_00634_, _00633_, _00632_);
  nor _23527_ (_00635_, _00634_, _00334_);
  or _23528_ (_00636_, _00635_, _00387_);
  or _23529_ (_00637_, _00636_, _00628_);
  nand _23530_ (_00638_, _00387_, _09526_);
  and _23531_ (_00639_, _00638_, _06444_);
  and _23532_ (_14392_, _00639_, _00637_);
  and _23533_ (_00640_, _07402_, _06394_);
  and _23534_ (_00641_, _00640_, _06933_);
  nand _23535_ (_00642_, _00641_, _06930_);
  or _23536_ (_00643_, _00641_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and _23537_ (_00644_, _00643_, _06674_);
  and _23538_ (_00645_, _00644_, _00642_);
  and _23539_ (_00646_, _07402_, _07150_);
  nand _23540_ (_00647_, _00646_, _06978_);
  or _23541_ (_00648_, _00646_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and _23542_ (_00649_, _00648_, _06440_);
  and _23543_ (_00651_, _00649_, _00647_);
  and _23544_ (_00652_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  or _23545_ (_00653_, _00652_, rst);
  or _23546_ (_00654_, _00653_, _00651_);
  or _23547_ (_14416_, _00654_, _00645_);
  nand _23548_ (_00656_, _10112_, _07069_);
  or _23549_ (_00657_, _10112_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  and _23550_ (_00658_, _00657_, _06444_);
  and _23551_ (_14515_, _00658_, _00656_);
  and _23552_ (_00659_, _08064_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  not _23553_ (_00660_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  nor _23554_ (_00661_, _08064_, _00660_);
  or _23555_ (_00662_, _00661_, _00659_);
  and _23556_ (_14522_, _00662_, _06444_);
  or _23557_ (_00663_, _08064_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  not _23558_ (_00664_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nand _23559_ (_00665_, _08064_, _00664_);
  and _23560_ (_00666_, _00665_, _06444_);
  and _23561_ (_14524_, _00666_, _00663_);
  and _23562_ (_00667_, _09373_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  or _23563_ (_14544_, _00667_, _09376_);
  and _23564_ (_00668_, _08912_, _06676_);
  and _23565_ (_00669_, _00668_, _13900_);
  and _23566_ (_00670_, _00669_, _00240_);
  nand _23567_ (_00672_, _00670_, _06930_);
  or _23568_ (_00673_, _00670_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  nor _23569_ (_00674_, _06350_, _06336_);
  and _23570_ (_00675_, _00674_, _06381_);
  and _23571_ (_00677_, _00675_, _13889_);
  not _23572_ (_00678_, _00677_);
  and _23573_ (_00679_, _00678_, _00673_);
  and _23574_ (_00680_, _00679_, _00672_);
  nor _23575_ (_00681_, _00678_, _10494_);
  or _23576_ (_00682_, _00681_, _00680_);
  and _23577_ (_00038_, _00682_, _06444_);
  and _23578_ (_00683_, _00669_, _06987_);
  nand _23579_ (_00684_, _00683_, _06930_);
  or _23580_ (_00685_, _00683_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and _23581_ (_00686_, _00685_, _00678_);
  and _23582_ (_00687_, _00686_, _00684_);
  nor _23583_ (_00689_, _00678_, _06666_);
  or _23584_ (_00690_, _00689_, _00687_);
  and _23585_ (_00056_, _00690_, _06444_);
  and _23586_ (_00692_, _06430_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  or _23587_ (_00693_, _00692_, _08233_);
  and _23588_ (_00694_, _00693_, _00669_);
  not _23589_ (_00696_, _00669_);
  nor _23590_ (_00697_, _06982_, _06430_);
  or _23591_ (_00698_, _00697_, _00696_);
  and _23592_ (_00699_, _00698_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  or _23593_ (_00700_, _00699_, _00677_);
  or _23594_ (_00702_, _00700_, _00694_);
  nand _23595_ (_00703_, _00677_, _07188_);
  and _23596_ (_00704_, _00703_, _06444_);
  and _23597_ (_00061_, _00704_, _00702_);
  and _23598_ (_00705_, _00669_, _08310_);
  nand _23599_ (_00706_, _00705_, _06930_);
  or _23600_ (_00707_, _00705_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and _23601_ (_00708_, _00707_, _00678_);
  and _23602_ (_00709_, _00708_, _00706_);
  nor _23603_ (_00710_, _00678_, _07300_);
  or _23604_ (_00711_, _00710_, _00709_);
  and _23605_ (_00064_, _00711_, _06444_);
  not _23606_ (_00712_, _08977_);
  nor _23607_ (_00713_, _00712_, _06930_);
  and _23608_ (_00714_, _06431_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or _23609_ (_00715_, _00714_, _00713_);
  and _23610_ (_00716_, _00715_, _00669_);
  or _23611_ (_00717_, _06932_, _06931_);
  or _23612_ (_00718_, _00696_, _00717_);
  and _23613_ (_00719_, _00718_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or _23614_ (_00720_, _00719_, _00677_);
  or _23615_ (_00721_, _00720_, _00716_);
  nand _23616_ (_00722_, _00677_, _11589_);
  and _23617_ (_00723_, _00722_, _06444_);
  and _23618_ (_00066_, _00723_, _00721_);
  and _23619_ (_00725_, _00669_, _06432_);
  nand _23620_ (_00726_, _00725_, _06930_);
  or _23621_ (_00727_, _00725_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and _23622_ (_00728_, _00727_, _00678_);
  and _23623_ (_00729_, _00728_, _00726_);
  nor _23624_ (_00730_, _00678_, _07069_);
  or _23625_ (_00731_, _00730_, _00729_);
  and _23626_ (_00082_, _00731_, _06444_);
  and _23627_ (_00732_, _00669_, _06942_);
  nand _23628_ (_00733_, _00732_, _06930_);
  or _23629_ (_00734_, _00732_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and _23630_ (_00735_, _00734_, _00678_);
  and _23631_ (_00736_, _00735_, _00733_);
  and _23632_ (_00737_, _00677_, _09527_);
  or _23633_ (_00738_, _00737_, _00736_);
  and _23634_ (_00085_, _00738_, _06444_);
  or _23635_ (_00739_, _07432_, \oc8051_top_1.oc8051_rom1.data_o [30]);
  nand _23636_ (_00740_, _07432_, _07434_);
  and _23637_ (_00741_, _00740_, _06444_);
  and _23638_ (_00088_, _00741_, _00739_);
  and _23639_ (_00742_, _00668_, _06670_);
  and _23640_ (_00743_, _00742_, _08310_);
  nand _23641_ (_00744_, _00743_, _06930_);
  or _23642_ (_00745_, _00743_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and _23643_ (_00746_, _08912_, _06945_);
  and _23644_ (_00747_, _00746_, _06940_);
  not _23645_ (_00748_, _00747_);
  and _23646_ (_00749_, _00748_, _00745_);
  and _23647_ (_00750_, _00749_, _00744_);
  nor _23648_ (_00751_, _00748_, _07300_);
  or _23649_ (_00752_, _00751_, _00750_);
  and _23650_ (_00143_, _00752_, _06444_);
  and _23651_ (_00753_, _00742_, _00240_);
  nand _23652_ (_00754_, _00753_, _06930_);
  or _23653_ (_00755_, _00753_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and _23654_ (_00756_, _00755_, _00748_);
  and _23655_ (_00757_, _00756_, _00754_);
  nor _23656_ (_00758_, _00748_, _10494_);
  or _23657_ (_00759_, _00758_, _00757_);
  and _23658_ (_00145_, _00759_, _06444_);
  and _23659_ (_00760_, _00742_, _06987_);
  nand _23660_ (_00761_, _00760_, _06930_);
  or _23661_ (_00762_, _00760_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and _23662_ (_00763_, _00762_, _00748_);
  and _23663_ (_00764_, _00763_, _00761_);
  nor _23664_ (_00765_, _00748_, _06666_);
  or _23665_ (_00766_, _00765_, _00764_);
  and _23666_ (_00147_, _00766_, _06444_);
  and _23667_ (_00767_, _06430_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  or _23668_ (_00768_, _00767_, _08233_);
  and _23669_ (_00769_, _00768_, _00742_);
  not _23670_ (_00770_, _00742_);
  or _23671_ (_00771_, _00770_, _00697_);
  and _23672_ (_00772_, _00771_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  or _23673_ (_00773_, _00772_, _00747_);
  or _23674_ (_00774_, _00773_, _00769_);
  nand _23675_ (_00775_, _00747_, _07188_);
  and _23676_ (_00776_, _00775_, _06444_);
  and _23677_ (_00149_, _00776_, _00774_);
  and _23678_ (_00777_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], _08478_);
  and _23679_ (_00778_, \oc8051_top_1.oc8051_memory_interface1.istb_t , \oc8051_top_1.oc8051_rom1.data_o [2]);
  or _23680_ (_00779_, _00778_, _00777_);
  and _23681_ (_00151_, _00779_, _06444_);
  and _23682_ (_00780_, _06431_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or _23683_ (_00781_, _00780_, _00713_);
  and _23684_ (_00782_, _00781_, _00742_);
  or _23685_ (_00783_, _00770_, _00717_);
  and _23686_ (_00784_, _00783_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or _23687_ (_00785_, _00784_, _00747_);
  or _23688_ (_00786_, _00785_, _00782_);
  nand _23689_ (_00787_, _00747_, _11589_);
  and _23690_ (_00788_, _00787_, _06444_);
  and _23691_ (_00153_, _00788_, _00786_);
  and _23692_ (_00789_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], _08478_);
  and _23693_ (_00790_, \oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or _23694_ (_00791_, _00790_, _00789_);
  and _23695_ (_00162_, _00791_, _06444_);
  and _23696_ (_00792_, _08478_, \oc8051_top_1.oc8051_memory_interface1.cdata [5]);
  and _23697_ (_00793_, \oc8051_top_1.oc8051_memory_interface1.istb_t , \oc8051_top_1.oc8051_rom1.data_o [5]);
  or _23698_ (_00794_, _00793_, _00792_);
  and _23699_ (_00164_, _00794_, _06444_);
  and _23700_ (_00795_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], _08478_);
  and _23701_ (_00796_, \oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or _23702_ (_00797_, _00796_, _00795_);
  and _23703_ (_00166_, _00797_, _06444_);
  and _23704_ (_00798_, _00742_, _06432_);
  nand _23705_ (_00799_, _00798_, _06930_);
  or _23706_ (_00800_, _00798_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and _23707_ (_00801_, _00800_, _00748_);
  and _23708_ (_00802_, _00801_, _00799_);
  nor _23709_ (_00803_, _00748_, _07069_);
  or _23710_ (_00804_, _00803_, _00802_);
  and _23711_ (_00169_, _00804_, _06444_);
  and _23712_ (_00805_, _00742_, _06942_);
  nand _23713_ (_00806_, _00805_, _06930_);
  or _23714_ (_00807_, _00805_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and _23715_ (_00808_, _00807_, _00748_);
  and _23716_ (_00809_, _00808_, _00806_);
  and _23717_ (_00810_, _00747_, _09527_);
  or _23718_ (_00811_, _00810_, _00809_);
  and _23719_ (_00172_, _00811_, _06444_);
  and _23720_ (_00812_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], _08478_);
  and _23721_ (_00813_, \oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or _23722_ (_00814_, _00813_, _00812_);
  and _23723_ (_00177_, _00814_, _06444_);
  and _23724_ (_00815_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], _08478_);
  and _23725_ (_00816_, \oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or _23726_ (_00817_, _00816_, _00815_);
  and _23727_ (_00189_, _00817_, _06444_);
  and _23728_ (_00818_, _13901_, _06670_);
  and _23729_ (_00819_, _00818_, _06983_);
  nand _23730_ (_00820_, _00819_, _06930_);
  or _23731_ (_00821_, _00819_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and _23732_ (_00822_, _00821_, _07408_);
  and _23733_ (_00823_, _00822_, _00820_);
  nor _23734_ (_00824_, _07408_, _07188_);
  or _23735_ (_00825_, _00824_, _00823_);
  and _23736_ (_00191_, _00825_, _06444_);
  and _23737_ (_00826_, _00818_, _08977_);
  nand _23738_ (_00827_, _00826_, _06930_);
  or _23739_ (_00828_, _00826_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and _23740_ (_00829_, _00828_, _07408_);
  and _23741_ (_00830_, _00829_, _00827_);
  nor _23742_ (_00831_, _11589_, _07408_);
  or _23743_ (_00832_, _00831_, _00830_);
  and _23744_ (_00205_, _00832_, _06444_);
  and _23745_ (_00833_, _00818_, _06942_);
  or _23746_ (_00834_, _00833_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and _23747_ (_00835_, _00834_, _07408_);
  nand _23748_ (_00836_, _00833_, _06930_);
  and _23749_ (_00837_, _00836_, _00835_);
  and _23750_ (_00838_, _09527_, _07407_);
  or _23751_ (_00839_, _00838_, _00837_);
  and _23752_ (_00211_, _00839_, _06444_);
  and _23753_ (_00840_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _23754_ (_00841_, _00840_, _09452_);
  and _23755_ (_00239_, _00841_, _06444_);
  nor _23756_ (_00842_, _13916_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or _23757_ (_00843_, _00842_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  nand _23758_ (_00844_, _00842_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  and _23759_ (_00845_, _00844_, _06444_);
  and _23760_ (_00247_, _00845_, _00843_);
  nand _23761_ (_00846_, _07199_, _07195_);
  and _23762_ (_00847_, _07199_, _07108_);
  or _23763_ (_00848_, _00847_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0]);
  and _23764_ (_00849_, _00848_, _06444_);
  and _23765_ (_00252_, _00849_, _00846_);
  nor _23766_ (_00850_, _07073_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nand _23767_ (_00851_, _00850_, _07195_);
  and _23768_ (_00852_, _00850_, _07108_);
  or _23769_ (_00853_, _00852_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0]);
  and _23770_ (_00854_, _00853_, _06444_);
  and _23771_ (_00256_, _00854_, _00851_);
  not _23772_ (_00855_, _11452_);
  and _23773_ (_00856_, _12023_, _00855_);
  and _23774_ (_00272_, _00856_, _06444_);
  or _23775_ (_00857_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and _23776_ (_00858_, _00857_, _07120_);
  or _23777_ (_00859_, _00858_, _07126_);
  and _23778_ (_00860_, _07111_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or _23779_ (_00861_, _00860_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and _23780_ (_00862_, _07113_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _23781_ (_00863_, _00862_, _07116_);
  and _23782_ (_00864_, _00863_, _00861_);
  nand _23783_ (_00865_, _07394_, _07116_);
  nand _23784_ (_00866_, _00865_, _07125_);
  or _23785_ (_00867_, _00866_, _00864_);
  and _23786_ (_00868_, _00867_, _00859_);
  and _23787_ (_00869_, _07394_, _07119_);
  or _23788_ (_00870_, _00869_, _07130_);
  or _23789_ (_00871_, _00870_, _00868_);
  or _23790_ (_00872_, _07131_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and _23791_ (_00873_, _00872_, _00871_);
  and _23792_ (_00874_, _00873_, _07134_);
  and _23793_ (_00875_, _00857_, _07085_);
  or _23794_ (_00876_, _00875_, _07091_);
  and _23795_ (_00877_, _07095_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or _23796_ (_00878_, _00877_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  nor _23797_ (_00879_, _07101_, _07077_);
  nor _23798_ (_00880_, _00879_, _07104_);
  and _23799_ (_00881_, _00880_, _00878_);
  nand _23800_ (_00882_, _07394_, _07104_);
  nand _23801_ (_00883_, _00882_, _07090_);
  or _23802_ (_00884_, _00883_, _00881_);
  and _23803_ (_00885_, _00884_, _00876_);
  and _23804_ (_00886_, _07394_, _07084_);
  or _23805_ (_00887_, _00886_, _00885_);
  and _23806_ (_00888_, _00887_, _07108_);
  or _23807_ (_00889_, _00888_, _07073_);
  or _23808_ (_00890_, _00889_, _00874_);
  or _23809_ (_00891_, _07075_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and _23810_ (_00892_, _00891_, _06444_);
  and _23811_ (_00274_, _00892_, _00890_);
  or _23812_ (_00893_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  or _23813_ (_00894_, _00893_, _07085_);
  not _23814_ (_00895_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  or _23815_ (_00896_, _00877_, _00895_);
  nand _23816_ (_00897_, _00896_, _00880_);
  or _23817_ (_00898_, _07385_, _07105_);
  and _23818_ (_00899_, _00898_, _00897_);
  or _23819_ (_00900_, _00899_, _07089_);
  not _23820_ (_00901_, _07087_);
  not _23821_ (_00902_, _07089_);
  or _23822_ (_00903_, _00893_, _00902_);
  and _23823_ (_00904_, _00903_, _00901_);
  and _23824_ (_00905_, _00904_, _00900_);
  and _23825_ (_00906_, _07385_, _07087_);
  or _23826_ (_00907_, _00906_, _07084_);
  or _23827_ (_00908_, _00907_, _00905_);
  and _23828_ (_00909_, _00908_, _00894_);
  or _23829_ (_00910_, _00909_, _07134_);
  or _23830_ (_00911_, _00893_, _07120_);
  or _23831_ (_00912_, _00860_, _00895_);
  nand _23832_ (_00913_, _00912_, _00863_);
  or _23833_ (_00914_, _07385_, _07117_);
  and _23834_ (_00915_, _00914_, _00913_);
  or _23835_ (_00916_, _00915_, _07124_);
  not _23836_ (_00917_, _07122_);
  not _23837_ (_00918_, _07124_);
  or _23838_ (_00919_, _00893_, _00918_);
  and _23839_ (_00920_, _00919_, _00917_);
  and _23840_ (_00921_, _00920_, _00916_);
  and _23841_ (_00922_, _07385_, _07122_);
  or _23842_ (_00923_, _00922_, _07119_);
  or _23843_ (_00924_, _00923_, _00921_);
  and _23844_ (_00925_, _00924_, _00911_);
  or _23845_ (_00926_, _00925_, _07196_);
  and _23846_ (_00927_, _00926_, _00910_);
  or _23847_ (_00928_, _00927_, _07073_);
  nor _23848_ (_00929_, _07132_, _07073_);
  or _23849_ (_00930_, _00929_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  and _23850_ (_00931_, _00930_, _06444_);
  and _23851_ (_00276_, _00931_, _00928_);
  or _23852_ (_00932_, _00589_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  and _23853_ (_00278_, _00932_, _06444_);
  and _23854_ (_00933_, _06442_, _06444_);
  and _23855_ (_00934_, _00933_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  and _23856_ (_00935_, _13854_, _06298_);
  nor _23857_ (_00936_, _00935_, _13836_);
  and _23858_ (_00937_, _00936_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  and _23859_ (_00938_, _00937_, _06443_);
  or _23860_ (_00280_, _00938_, _00934_);
  nor _23861_ (_00282_, _12648_, rst);
  and _23862_ (_00287_, _11576_, _06444_);
  or _23863_ (_00939_, _07077_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and _23864_ (_00940_, _00939_, _07120_);
  or _23865_ (_00941_, _00940_, _07126_);
  and _23866_ (_00942_, _07111_, _07077_);
  or _23867_ (_00943_, _00942_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and _23868_ (_00944_, _07113_, _07077_);
  nor _23869_ (_00945_, _00944_, _07116_);
  and _23870_ (_00946_, _00945_, _00943_);
  nand _23871_ (_00947_, _07393_, _07116_);
  nand _23872_ (_00948_, _00947_, _07125_);
  or _23873_ (_00949_, _00948_, _00946_);
  and _23874_ (_00950_, _00949_, _00941_);
  and _23875_ (_00951_, _07393_, _07119_);
  or _23876_ (_00952_, _00951_, _07130_);
  or _23877_ (_00953_, _00952_, _00950_);
  or _23878_ (_00954_, _07131_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and _23879_ (_00955_, _00954_, _00953_);
  and _23880_ (_00956_, _00955_, _07134_);
  and _23881_ (_00957_, _00939_, _07085_);
  or _23882_ (_00958_, _00957_, _07091_);
  and _23883_ (_00959_, _07393_, _07104_);
  nor _23884_ (_00960_, _07101_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _23885_ (_00961_, _00960_, _07104_);
  and _23886_ (_00962_, _07095_, _07077_);
  or _23887_ (_00963_, _00962_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  nand _23888_ (_00964_, _00963_, _00961_);
  nand _23889_ (_00965_, _00964_, _07090_);
  or _23890_ (_00966_, _00965_, _00959_);
  and _23891_ (_00967_, _00966_, _00958_);
  and _23892_ (_00968_, _07393_, _07084_);
  or _23893_ (_00969_, _00968_, _00967_);
  and _23894_ (_00970_, _00969_, _07108_);
  or _23895_ (_00971_, _00970_, _00956_);
  or _23896_ (_00972_, _00971_, _07073_);
  or _23897_ (_00973_, _07075_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and _23898_ (_00974_, _00973_, _06444_);
  and _23899_ (_00295_, _00974_, _00972_);
  or _23900_ (_00975_, _07077_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  or _23901_ (_00977_, _00975_, _07120_);
  or _23902_ (_00978_, _07384_, _00917_);
  not _23903_ (_00979_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  or _23904_ (_00980_, _00942_, _00979_);
  nand _23905_ (_00981_, _00980_, _00945_);
  or _23906_ (_00982_, _07384_, _07117_);
  and _23907_ (_00983_, _00982_, _00918_);
  and _23908_ (_00984_, _00983_, _00981_);
  and _23909_ (_00985_, _00975_, _07124_);
  or _23910_ (_00986_, _00985_, _07122_);
  or _23911_ (_00987_, _00986_, _00984_);
  and _23912_ (_00988_, _00987_, _00978_);
  or _23913_ (_00989_, _00988_, _07119_);
  and _23914_ (_00990_, _00989_, _00977_);
  or _23915_ (_00991_, _00990_, _07196_);
  or _23916_ (_00992_, _00975_, _07085_);
  or _23917_ (_00993_, _00962_, _00979_);
  nand _23918_ (_00994_, _00993_, _00961_);
  or _23919_ (_00995_, _07384_, _07105_);
  and _23920_ (_00996_, _00995_, _00994_);
  or _23921_ (_00997_, _00996_, _07089_);
  or _23922_ (_00998_, _00975_, _00902_);
  and _23923_ (_01000_, _00998_, _00901_);
  and _23924_ (_01001_, _01000_, _00997_);
  and _23925_ (_01002_, _07384_, _07087_);
  or _23926_ (_01003_, _01002_, _07084_);
  or _23927_ (_01004_, _01003_, _01001_);
  and _23928_ (_01005_, _01004_, _00992_);
  or _23929_ (_01006_, _01005_, _07134_);
  and _23930_ (_01007_, _01006_, _00991_);
  or _23931_ (_01008_, _01007_, _07073_);
  or _23932_ (_01009_, _00929_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  and _23933_ (_01010_, _01009_, _06444_);
  and _23934_ (_00299_, _01010_, _01008_);
  nor _23935_ (_01011_, _07108_, _07073_);
  or _23936_ (_01012_, _01011_, _07077_);
  nand _23937_ (_01013_, _00850_, _07132_);
  and _23938_ (_01014_, _01013_, _06444_);
  and _23939_ (_00326_, _01014_, _01012_);
  and _23940_ (_01015_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _06444_);
  and _23941_ (_00331_, _01015_, _07073_);
  nand _23942_ (_01016_, _07127_, _07203_);
  nor _23943_ (_01017_, _01016_, _07108_);
  and _23944_ (_01018_, _07073_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  or _23945_ (_01019_, _07104_, _07073_);
  nor _23946_ (_01020_, _01019_, _07082_);
  not _23947_ (_01021_, _07091_);
  nor _23948_ (_01022_, _07102_, _01021_);
  and _23949_ (_01023_, _01022_, _01020_);
  or _23950_ (_01024_, _01023_, _01018_);
  or _23951_ (_01025_, _01024_, _01017_);
  and _23952_ (_00339_, _01025_, _06444_);
  or _23953_ (_01026_, _07124_, _07116_);
  and _23954_ (_01027_, _07114_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or _23955_ (_01028_, _01027_, _01026_);
  and _23956_ (_01029_, _01028_, _00917_);
  and _23957_ (_01030_, _07195_, _07120_);
  and _23958_ (_01031_, _01030_, _01029_);
  or _23959_ (_01032_, _07104_, _07089_);
  and _23960_ (_01033_, _07102_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or _23961_ (_01034_, _01033_, _01032_);
  and _23962_ (_01035_, _01034_, _00901_);
  and _23963_ (_01036_, _07108_, _07085_);
  and _23964_ (_01037_, _01036_, _01035_);
  or _23965_ (_01038_, _01037_, _07073_);
  or _23966_ (_01039_, _01038_, _01031_);
  or _23967_ (_01040_, _07075_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and _23968_ (_01041_, _01040_, _06444_);
  and _23969_ (_00342_, _01041_, _01039_);
  nor _23970_ (_01042_, _07111_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nor _23971_ (_01043_, _01042_, _07113_);
  or _23972_ (_01044_, _01043_, _07116_);
  and _23973_ (_01045_, _01044_, _00918_);
  or _23974_ (_01046_, _01045_, _07122_);
  and _23975_ (_01047_, _01046_, _01030_);
  or _23976_ (_01048_, _07095_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and _23977_ (_01049_, _01048_, _07101_);
  or _23978_ (_01050_, _01049_, _07104_);
  and _23979_ (_01051_, _01050_, _00902_);
  or _23980_ (_01052_, _01051_, _07087_);
  and _23981_ (_01053_, _01052_, _01036_);
  or _23982_ (_01054_, _01053_, _07073_);
  or _23983_ (_01055_, _01054_, _01047_);
  or _23984_ (_01056_, _07075_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and _23985_ (_01057_, _01056_, _06444_);
  and _23986_ (_00345_, _01057_, _01055_);
  and _23987_ (_00350_, _12703_, _07073_);
  and _23988_ (_01058_, _07073_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  or _23989_ (_01059_, _01058_, _00929_);
  and _23990_ (_00368_, _01059_, _06444_);
  and _23991_ (_01060_, _07073_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  or _23992_ (_01061_, _01060_, _00929_);
  and _23993_ (_00371_, _01061_, _06444_);
  and _23994_ (_01062_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and _23995_ (_01063_, _12223_, \oc8051_top_1.oc8051_rom1.data_o [29]);
  or _23996_ (_01064_, _01063_, _01062_);
  and _23997_ (_00434_, _01064_, _06444_);
  and _23998_ (_01065_, _08064_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  not _23999_ (_01066_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor _24000_ (_01067_, _08064_, _01066_);
  or _24001_ (_01068_, _01067_, _01065_);
  and _24002_ (_00447_, _01068_, _06444_);
  and _24003_ (_01069_, _12825_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  nand _24004_ (_01070_, _06439_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  nor _24005_ (_01071_, _01070_, _07415_);
  and _24006_ (_01072_, _12829_, _07070_);
  or _24007_ (_01073_, _01072_, _01071_);
  or _24008_ (_01074_, _01073_, _01069_);
  and _24009_ (_00471_, _01074_, _06444_);
  or _24010_ (_01075_, _08064_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  not _24011_ (_01076_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  nand _24012_ (_01077_, _08064_, _01076_);
  and _24013_ (_01078_, _01077_, _06444_);
  and _24014_ (_00475_, _01078_, _01075_);
  and _24015_ (_01079_, _00604_, _08912_);
  and _24016_ (_01080_, _01079_, _06933_);
  nand _24017_ (_01081_, _01080_, _06930_);
  or _24018_ (_01082_, _01080_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and _24019_ (_01083_, _01082_, _06674_);
  and _24020_ (_01084_, _01083_, _01081_);
  and _24021_ (_01085_, _00674_, _07150_);
  and _24022_ (_01086_, _01085_, _06381_);
  not _24023_ (_01087_, _01086_);
  nor _24024_ (_01088_, _01087_, _06978_);
  and _24025_ (_01089_, _01087_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or _24026_ (_01090_, _01089_, _01088_);
  and _24027_ (_01091_, _01090_, _06440_);
  and _24028_ (_01092_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or _24029_ (_01093_, _01092_, rst);
  or _24030_ (_01094_, _01093_, _01091_);
  or _24031_ (_00501_, _01094_, _01084_);
  and _24032_ (_01095_, _14070_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  nor _24033_ (_01096_, _14070_, _07188_);
  or _24034_ (_01097_, _01096_, _01095_);
  and _24035_ (_00504_, _01097_, _06444_);
  nor _24036_ (_01098_, _12830_, _07300_);
  nor _24037_ (_01099_, _07415_, _07158_);
  or _24038_ (_01100_, _01099_, _12825_);
  and _24039_ (_01101_, _01100_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  or _24040_ (_01102_, _01101_, _01098_);
  and _24041_ (_00509_, _01102_, _06444_);
  and _24042_ (_01103_, _09373_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  or _24043_ (_00544_, _01103_, _09383_);
  and _24044_ (_01104_, _09373_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  or _24045_ (_00550_, _01104_, _09390_);
  or _24046_ (_01105_, _08064_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  not _24047_ (_01106_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  nand _24048_ (_01107_, _08064_, _01106_);
  and _24049_ (_01108_, _01107_, _06444_);
  and _24050_ (_00569_, _01108_, _01105_);
  and _24051_ (_01109_, _08064_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  not _24052_ (_01110_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  nor _24053_ (_01111_, _08064_, _01110_);
  or _24054_ (_01112_, _01111_, _01109_);
  and _24055_ (_00572_, _01112_, _06444_);
  nor _24056_ (_00608_, _11688_, rst);
  nor _24057_ (_01113_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and _24058_ (_01114_, _01113_, _06296_);
  and _24059_ (_01115_, _01114_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  not _24060_ (_01116_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  nor _24061_ (_01117_, _01114_, _01116_);
  or _24062_ (_01118_, _01117_, _01115_);
  or _24063_ (_01119_, _01118_, _13902_);
  or _24064_ (_01120_, _08977_, _01116_);
  nand _24065_ (_01121_, _01120_, _13902_);
  or _24066_ (_01122_, _01121_, _00713_);
  and _24067_ (_01123_, _01122_, _01119_);
  or _24068_ (_01124_, _01123_, _13906_);
  nand _24069_ (_01125_, _13906_, _11589_);
  and _24070_ (_01126_, _01125_, _06444_);
  and _24071_ (_00629_, _01126_, _01124_);
  and _24072_ (_01127_, _08064_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  not _24073_ (_01128_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nor _24074_ (_01129_, _08064_, _01128_);
  or _24075_ (_01130_, _01129_, _01127_);
  and _24076_ (_00650_, _01130_, _06444_);
  and _24077_ (_01131_, _10891_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  or _24078_ (_01132_, _10882_, _07236_);
  nand _24079_ (_01133_, _10882_, _07236_);
  and _24080_ (_01134_, _01133_, _01132_);
  nand _24081_ (_01135_, _01134_, _01131_);
  or _24082_ (_01136_, _01134_, _01131_);
  and _24083_ (_01137_, _01136_, _01135_);
  or _24084_ (_01138_, _01137_, _07429_);
  or _24085_ (_01139_, _07230_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and _24086_ (_01140_, _01139_, _10894_);
  and _24087_ (_00655_, _01140_, _01138_);
  or _24088_ (_01141_, _08064_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  not _24089_ (_01142_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nand _24090_ (_01143_, _08064_, _01142_);
  and _24091_ (_01144_, _01143_, _06444_);
  and _24092_ (_00671_, _01144_, _01141_);
  and _24093_ (_01146_, _08064_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  nor _24094_ (_01147_, _08064_, _01142_);
  or _24095_ (_01148_, _01147_, _01146_);
  and _24096_ (_00676_, _01148_, _06444_);
  or _24097_ (_01149_, _08064_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  not _24098_ (_01150_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nand _24099_ (_01151_, _08064_, _01150_);
  and _24100_ (_01152_, _01151_, _06444_);
  and _24101_ (_00688_, _01152_, _01149_);
  and _24102_ (_01153_, _08064_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  not _24103_ (_01154_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor _24104_ (_01155_, _08064_, _01154_);
  or _24105_ (_01156_, _01155_, _01153_);
  and _24106_ (_00691_, _01156_, _06444_);
  and _24107_ (_01158_, _13902_, _06987_);
  nand _24108_ (_01160_, _01158_, _06930_);
  or _24109_ (_01161_, _01158_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  and _24110_ (_01162_, _01161_, _13907_);
  and _24111_ (_01163_, _01162_, _01160_);
  nor _24112_ (_01165_, _13907_, _06666_);
  or _24113_ (_01166_, _01165_, _01163_);
  and _24114_ (_00695_, _01166_, _06444_);
  and _24115_ (_01167_, _13902_, _06983_);
  nand _24116_ (_01168_, _01167_, _06930_);
  or _24117_ (_01169_, _01167_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and _24118_ (_01170_, _01169_, _13907_);
  and _24119_ (_01171_, _01170_, _01168_);
  nor _24120_ (_01172_, _13907_, _07188_);
  or _24121_ (_01173_, _01172_, _01171_);
  and _24122_ (_00701_, _01173_, _06444_);
  or _24123_ (_01174_, _07432_, \oc8051_top_1.oc8051_rom1.data_o [14]);
  nand _24124_ (_01175_, _07432_, _13985_);
  and _24125_ (_01176_, _01175_, _06444_);
  and _24126_ (_00724_, _01176_, _01174_);
  and _24127_ (_01177_, _12712_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  or _24128_ (_01178_, _01177_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and _24129_ (_00976_, _01178_, _06444_);
  and _24130_ (_01179_, _12712_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  or _24131_ (_01180_, _01179_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  and _24132_ (_00999_, _01180_, _06444_);
  nor _24133_ (_01181_, _06978_, _06449_);
  and _24134_ (_01182_, _06449_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  or _24135_ (_01184_, _01182_, _01181_);
  and _24136_ (_01157_, _01184_, _06444_);
  and _24137_ (_01185_, _13902_, _08310_);
  nand _24138_ (_01186_, _01185_, _06930_);
  or _24139_ (_01187_, _01185_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  and _24140_ (_01188_, _01187_, _13907_);
  and _24141_ (_01189_, _01188_, _01186_);
  nor _24142_ (_01190_, _13907_, _07300_);
  or _24143_ (_01191_, _01190_, _01189_);
  and _24144_ (_01159_, _01191_, _06444_);
  and _24145_ (_01192_, _14175_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  and _24146_ (_01193_, _14088_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and _24147_ (_01194_, _14084_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or _24148_ (_01195_, _01194_, _01193_);
  and _24149_ (_01196_, _14093_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and _24150_ (_01197_, _14096_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or _24151_ (_01198_, _01197_, _01196_);
  or _24152_ (_01199_, _01198_, _01195_);
  and _24153_ (_01200_, _14102_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and _24154_ (_01201_, _14105_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  or _24155_ (_01202_, _01201_, _01200_);
  and _24156_ (_01203_, _14110_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and _24157_ (_01204_, _14116_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  or _24158_ (_01205_, _01204_, _01203_);
  or _24159_ (_01206_, _01205_, _01202_);
  or _24160_ (_01207_, _01206_, _01199_);
  and _24161_ (_01208_, _14120_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and _24162_ (_01209_, _14122_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  or _24163_ (_01210_, _01209_, _01208_);
  and _24164_ (_01211_, _14124_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and _24165_ (_01212_, _14125_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  or _24166_ (_01213_, _01212_, _01211_);
  or _24167_ (_01214_, _01213_, _01210_);
  and _24168_ (_01215_, _14131_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  and _24169_ (_01216_, _14130_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  or _24170_ (_01217_, _01216_, _01215_);
  and _24171_ (_01219_, _14133_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _24172_ (_01220_, _14134_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  or _24173_ (_01221_, _01220_, _01219_);
  or _24174_ (_01222_, _01221_, _01217_);
  or _24175_ (_01223_, _01222_, _01214_);
  or _24176_ (_01224_, _01223_, _01207_);
  and _24177_ (_01225_, _14154_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  not _24178_ (_01226_, _11734_);
  and _24179_ (_01227_, _14156_, _01226_);
  or _24180_ (_01228_, _01227_, _01225_);
  and _24181_ (_01229_, _14150_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and _24182_ (_01230_, _14152_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or _24183_ (_01231_, _01230_, _01229_);
  or _24184_ (_01232_, _01231_, _01228_);
  or _24185_ (_01233_, _14247_, p3_in[5]);
  or _24186_ (_01234_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and _24187_ (_01235_, _01234_, _01233_);
  and _24188_ (_01236_, _01235_, _14260_);
  or _24189_ (_01237_, _14247_, p2_in[5]);
  or _24190_ (_01238_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and _24191_ (_01239_, _01238_, _01237_);
  and _24192_ (_01240_, _01239_, _14265_);
  or _24193_ (_01241_, _01240_, _01236_);
  or _24194_ (_01242_, _14247_, p0_in[5]);
  or _24195_ (_01243_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and _24196_ (_01244_, _01243_, _01242_);
  and _24197_ (_01245_, _01244_, _14224_);
  or _24198_ (_01246_, _14247_, p1_in[5]);
  or _24199_ (_01248_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and _24200_ (_01249_, _01248_, _01246_);
  and _24201_ (_01250_, _01249_, _14253_);
  or _24202_ (_01251_, _01250_, _01245_);
  or _24203_ (_01252_, _01251_, _01241_);
  or _24204_ (_01253_, _01252_, _01232_);
  and _24205_ (_01254_, _14146_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and _24206_ (_01255_, _14143_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  or _24207_ (_01256_, _01255_, _01254_);
  or _24208_ (_01257_, _01256_, _01253_);
  or _24209_ (_01258_, _01257_, _01224_);
  and _24210_ (_01259_, _01258_, _14174_);
  or _24211_ (_01260_, _01259_, _14178_);
  or _24212_ (_01261_, _01260_, _01192_);
  or _24213_ (_01262_, _14353_, _08127_);
  and _24214_ (_01263_, _01262_, _06444_);
  and _24215_ (_01164_, _01263_, _01261_);
  nor _24216_ (_01264_, _11589_, _07190_);
  and _24217_ (_01265_, _10497_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  or _24218_ (_01266_, _01265_, _01264_);
  and _24219_ (_01183_, _01266_, _06444_);
  and _24220_ (_01267_, _06449_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  and _24221_ (_01268_, _12841_, _06447_);
  or _24222_ (_01269_, _01268_, _01267_);
  and _24223_ (_01218_, _01269_, _06444_);
  and _24224_ (_01270_, _07414_, _06439_);
  or _24225_ (_01271_, _01270_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  nand _24226_ (_01272_, _01270_, _09526_);
  and _24227_ (_01273_, _01272_, _06444_);
  and _24228_ (_01247_, _01273_, _01271_);
  or _24229_ (_01274_, _08064_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  not _24230_ (_01275_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  nand _24231_ (_01276_, _08064_, _01275_);
  and _24232_ (_01277_, _01276_, _06444_);
  and _24233_ (_01378_, _01277_, _01274_);
  and _24234_ (_01278_, _08064_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  not _24235_ (_01279_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _24236_ (_01280_, _08064_, _01279_);
  or _24237_ (_01281_, _01280_, _01278_);
  and _24238_ (_01394_, _01281_, _06444_);
  nor _24239_ (_01282_, _14070_, _07300_);
  and _24240_ (_01283_, _14070_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  or _24241_ (_01284_, _01283_, _01282_);
  and _24242_ (_01641_, _01284_, _06444_);
  nor _24243_ (_01285_, \oc8051_top_1.oc8051_decoder1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  and _24244_ (_01286_, _01285_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  not _24245_ (_01287_, _01286_);
  or _24246_ (_01288_, _01287_, _08308_);
  or _24247_ (_01289_, _01286_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3]);
  and _24248_ (_01290_, _01289_, _06444_);
  and _24249_ (_01650_, _01290_, _01288_);
  and _24250_ (_01291_, _12711_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  or _24251_ (_01292_, _01291_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  and _24252_ (_01676_, _01292_, _06444_);
  and _24253_ (_01293_, _12712_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  or _24254_ (_01294_, _01293_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  and _24255_ (_01679_, _01294_, _06444_);
  and _24256_ (_01295_, _12712_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  or _24257_ (_01296_, _01295_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and _24258_ (_01684_, _01296_, _06444_);
  nand _24259_ (_01297_, _01286_, _09138_);
  or _24260_ (_01298_, _01286_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2]);
  and _24261_ (_01299_, _01298_, _06444_);
  and _24262_ (_01697_, _01299_, _01297_);
  not _24263_ (_01300_, _06432_);
  nor _24264_ (_01301_, _06930_, _01300_);
  nand _24265_ (_01302_, _01300_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  nand _24266_ (_01303_, _01302_, _13902_);
  or _24267_ (_01304_, _01303_, _01301_);
  or _24268_ (_01305_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  or _24269_ (_01306_, _01305_, _13902_);
  and _24270_ (_01307_, _01306_, _01304_);
  or _24271_ (_01308_, _01307_, _13906_);
  nand _24272_ (_01309_, _13906_, _07069_);
  and _24273_ (_01310_, _01309_, _06444_);
  and _24274_ (_01700_, _01310_, _01308_);
  not _24275_ (_01311_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  or _24276_ (_01312_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _01311_);
  or _24277_ (_01313_, _01312_, _06295_);
  and _24278_ (_01314_, _01313_, _01113_);
  or _24279_ (_01315_, _01314_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or _24280_ (_01316_, _01315_, _13902_);
  nand _24281_ (_01317_, _08021_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  nand _24282_ (_01318_, _01317_, _13902_);
  or _24283_ (_01319_, _01318_, _08022_);
  and _24284_ (_01320_, _01319_, _01316_);
  or _24285_ (_01321_, _01320_, _13906_);
  nand _24286_ (_01322_, _13906_, _09526_);
  and _24287_ (_01323_, _01322_, _06444_);
  and _24288_ (_01702_, _01323_, _01321_);
  and _24289_ (_01324_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and _24290_ (_01325_, _12223_, \oc8051_top_1.oc8051_rom1.data_o [17]);
  or _24291_ (_01326_, _01325_, _01324_);
  and _24292_ (_01708_, _01326_, _06444_);
  and _24293_ (_01327_, _12712_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  or _24294_ (_01328_, _01327_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and _24295_ (_01716_, _01328_, _06444_);
  and _24296_ (_01329_, _14070_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  nor _24297_ (_01330_, _14070_, _10494_);
  or _24298_ (_01331_, _01330_, _01329_);
  and _24299_ (_01734_, _01331_, _06444_);
  or _24300_ (_01332_, _01287_, _07959_);
  or _24301_ (_01333_, _01286_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1]);
  and _24302_ (_01334_, _01333_, _06444_);
  and _24303_ (_01752_, _01334_, _01332_);
  or _24304_ (_01335_, _01287_, _08019_);
  or _24305_ (_01336_, _01286_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  and _24306_ (_01337_, _01336_, _06444_);
  and _24307_ (_01786_, _01337_, _01335_);
  and _24308_ (_01338_, _08064_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor _24309_ (_01339_, _08064_, _00664_);
  or _24310_ (_01340_, _01339_, _01338_);
  and _24311_ (_01790_, _01340_, _06444_);
  and _24312_ (_01341_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and _24313_ (_01343_, _12223_, \oc8051_top_1.oc8051_rom1.data_o [16]);
  or _24314_ (_01344_, _01343_, _01341_);
  and _24315_ (_01803_, _01344_, _06444_);
  nor _24316_ (_01806_, \oc8051_top_1.oc8051_sfr1.prescaler [0], rst);
  and _24317_ (_01345_, _08230_, _06444_);
  or _24318_ (_01346_, _01345_, _14496_);
  and _24319_ (_01347_, _14175_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  and _24320_ (_01348_, _14084_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and _24321_ (_01349_, _14088_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  or _24322_ (_01350_, _01349_, _01348_);
  and _24323_ (_01351_, _14093_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and _24324_ (_01352_, _14096_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or _24325_ (_01353_, _01352_, _01351_);
  or _24326_ (_01354_, _01353_, _01350_);
  and _24327_ (_01355_, _14102_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and _24328_ (_01356_, _14105_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  or _24329_ (_01357_, _01356_, _01355_);
  and _24330_ (_01358_, _14110_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  and _24331_ (_01359_, _14116_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  or _24332_ (_01360_, _01359_, _01358_);
  or _24333_ (_01361_, _01360_, _01357_);
  or _24334_ (_01362_, _01361_, _01354_);
  and _24335_ (_01363_, _14120_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and _24336_ (_01364_, _14122_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  or _24337_ (_01365_, _01364_, _01363_);
  and _24338_ (_01366_, _14125_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and _24339_ (_01367_, _14124_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  or _24340_ (_01368_, _01367_, _01366_);
  or _24341_ (_01369_, _01368_, _01365_);
  and _24342_ (_01370_, _14131_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and _24343_ (_01371_, _14130_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  or _24344_ (_01372_, _01371_, _01370_);
  and _24345_ (_01373_, _14133_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _24346_ (_01374_, _14134_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  or _24347_ (_01375_, _01374_, _01373_);
  or _24348_ (_01376_, _01375_, _01372_);
  or _24349_ (_01377_, _01376_, _01369_);
  or _24350_ (_01379_, _01377_, _01362_);
  and _24351_ (_01380_, _14150_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and _24352_ (_01381_, _14152_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or _24353_ (_01382_, _01381_, _01380_);
  and _24354_ (_01383_, _14154_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and _24355_ (_01384_, _14156_, _11664_);
  or _24356_ (_01385_, _01384_, _01383_);
  or _24357_ (_01386_, _01385_, _01382_);
  or _24358_ (_01387_, _14247_, p0_in[4]);
  or _24359_ (_01388_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and _24360_ (_01389_, _01388_, _01387_);
  and _24361_ (_01390_, _01389_, _14224_);
  or _24362_ (_01391_, _14247_, p1_in[4]);
  or _24363_ (_01392_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and _24364_ (_01393_, _01392_, _01391_);
  and _24365_ (_01395_, _01393_, _14253_);
  or _24366_ (_01396_, _01395_, _01390_);
  or _24367_ (_01397_, _14247_, p3_in[4]);
  or _24368_ (_01398_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and _24369_ (_01399_, _01398_, _01397_);
  and _24370_ (_01400_, _01399_, _14260_);
  or _24371_ (_01401_, _14247_, p2_in[4]);
  or _24372_ (_01402_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and _24373_ (_01403_, _01402_, _01401_);
  and _24374_ (_01404_, _01403_, _14265_);
  or _24375_ (_01405_, _01404_, _01400_);
  or _24376_ (_01406_, _01405_, _01396_);
  or _24377_ (_01407_, _01406_, _01386_);
  and _24378_ (_01408_, _14143_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and _24379_ (_01409_, _14146_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or _24380_ (_01410_, _01409_, _01408_);
  or _24381_ (_01411_, _01410_, _01407_);
  or _24382_ (_01412_, _01411_, _01379_);
  and _24383_ (_01413_, _01412_, _14174_);
  or _24384_ (_01414_, _01413_, _14178_);
  or _24385_ (_01415_, _01414_, _01347_);
  and _24386_ (_01808_, _01415_, _01346_);
  and _24387_ (_01416_, _08019_, _06444_);
  or _24388_ (_01417_, _01416_, _14496_);
  and _24389_ (_01418_, _14096_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and _24390_ (_01419_, _14093_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  or _24391_ (_01420_, _01419_, _01418_);
  and _24392_ (_01421_, _14088_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and _24393_ (_01422_, _14084_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  or _24394_ (_01423_, _01422_, _01421_);
  or _24395_ (_01424_, _01423_, _01420_);
  and _24396_ (_01425_, _14102_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and _24397_ (_01426_, _14105_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  or _24398_ (_01427_, _01426_, _01425_);
  and _24399_ (_01428_, _14110_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and _24400_ (_01429_, _14116_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  or _24401_ (_01430_, _01429_, _01428_);
  or _24402_ (_01431_, _01430_, _01427_);
  or _24403_ (_01432_, _01431_, _01424_);
  and _24404_ (_01433_, _14124_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and _24405_ (_01434_, _14125_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  or _24406_ (_01435_, _01434_, _01433_);
  and _24407_ (_01436_, _14122_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and _24408_ (_01437_, _14120_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  or _24409_ (_01438_, _01437_, _01436_);
  or _24410_ (_01439_, _01438_, _01435_);
  and _24411_ (_01440_, _14131_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  and _24412_ (_01441_, _14130_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  or _24413_ (_01442_, _01441_, _01440_);
  and _24414_ (_01443_, _14133_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and _24415_ (_01444_, _14134_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  or _24416_ (_01445_, _01444_, _01443_);
  or _24417_ (_01446_, _01445_, _01442_);
  or _24418_ (_01447_, _01446_, _01439_);
  or _24419_ (_01448_, _01447_, _01432_);
  and _24420_ (_01449_, _14154_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  and _24421_ (_01450_, _14156_, _11858_);
  or _24422_ (_01451_, _01450_, _01449_);
  and _24423_ (_01452_, _14150_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and _24424_ (_01453_, _14152_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or _24425_ (_01454_, _01453_, _01452_);
  or _24426_ (_01455_, _01454_, _01451_);
  or _24427_ (_01456_, _14247_, p3_in[0]);
  or _24428_ (_01457_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and _24429_ (_01458_, _01457_, _01456_);
  and _24430_ (_01459_, _01458_, _14260_);
  or _24431_ (_01460_, _14247_, p2_in[0]);
  or _24432_ (_01461_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and _24433_ (_01462_, _01461_, _01460_);
  and _24434_ (_01463_, _01462_, _14265_);
  or _24435_ (_01464_, _01463_, _01459_);
  or _24436_ (_01465_, _14247_, p0_in[0]);
  or _24437_ (_01466_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  and _24438_ (_01467_, _01466_, _01465_);
  and _24439_ (_01468_, _01467_, _14224_);
  or _24440_ (_01469_, _14247_, p1_in[0]);
  or _24441_ (_01470_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and _24442_ (_01471_, _01470_, _01469_);
  and _24443_ (_01472_, _01471_, _14253_);
  or _24444_ (_01473_, _01472_, _01468_);
  or _24445_ (_01474_, _01473_, _01464_);
  or _24446_ (_01475_, _01474_, _01455_);
  or _24447_ (_01476_, _08269_, _08196_);
  nand _24448_ (_01477_, _08269_, _08196_);
  nand _24449_ (_01478_, _01477_, _01476_);
  or _24450_ (_01479_, _09045_, _07652_);
  not _24451_ (_01480_, _00240_);
  nor _24452_ (_01481_, _01480_, _06930_);
  nor _24453_ (_01482_, _00240_, _06736_);
  nor _24454_ (_01483_, _01482_, _01481_);
  nor _24455_ (_01484_, _01483_, _08028_);
  and _24456_ (_01485_, _08036_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or _24457_ (_01486_, _01485_, _07439_);
  nor _24458_ (_01487_, _01486_, _01484_);
  nand _24459_ (_01488_, _01487_, _01479_);
  and _24460_ (_01489_, _09201_, _07439_);
  not _24461_ (_01490_, _01489_);
  and _24462_ (_01491_, _01490_, _01488_);
  or _24463_ (_01492_, _01491_, _11179_);
  nand _24464_ (_01493_, _01491_, _11179_);
  and _24465_ (_01494_, _01493_, _01492_);
  nand _24466_ (_01495_, _01494_, _01478_);
  or _24467_ (_01496_, _01494_, _01478_);
  and _24468_ (_01497_, _01496_, _01495_);
  or _24469_ (_01498_, _08063_, _07976_);
  nand _24470_ (_01499_, _08063_, _07976_);
  nand _24471_ (_01500_, _01499_, _01498_);
  or _24472_ (_01501_, _09138_, _07652_);
  nor _24473_ (_01502_, _08977_, _06782_);
  nor _24474_ (_01503_, _01502_, _00713_);
  nor _24475_ (_01504_, _01503_, _08028_);
  and _24476_ (_01505_, _08036_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or _24477_ (_01506_, _01505_, _07439_);
  nor _24478_ (_01507_, _01506_, _01504_);
  and _24479_ (_01508_, _01507_, _01501_);
  and _24480_ (_01509_, _09280_, _07439_);
  or _24481_ (_01510_, _01509_, _01508_);
  nand _24482_ (_01511_, _01510_, _08344_);
  or _24483_ (_01512_, _01510_, _08344_);
  and _24484_ (_01513_, _01512_, _01511_);
  nand _24485_ (_01514_, _01513_, _01500_);
  or _24486_ (_01515_, _01513_, _01500_);
  and _24487_ (_01516_, _01515_, _01514_);
  nor _24488_ (_01517_, _01516_, _01497_);
  and _24489_ (_01518_, _01516_, _01497_);
  or _24490_ (_01519_, _01518_, _01517_);
  and _24491_ (_01520_, _01519_, _14143_);
  and _24492_ (_01521_, _14146_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or _24493_ (_01522_, _01521_, _01520_);
  or _24494_ (_01523_, _01522_, _01475_);
  or _24495_ (_01524_, _01523_, _01448_);
  and _24496_ (_01525_, _01524_, _14174_);
  and _24497_ (_01526_, _14175_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  or _24498_ (_01527_, _01526_, _14178_);
  or _24499_ (_01528_, _01527_, _01525_);
  and _24500_ (_01810_, _01528_, _01417_);
  not _24501_ (_01529_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  not _24502_ (_01530_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and _24503_ (_01531_, _10967_, _01530_);
  and _24504_ (_01532_, _01531_, _01529_);
  nor _24505_ (_01533_, _01531_, _01529_);
  nor _24506_ (_01534_, _01533_, _01532_);
  not _24507_ (_01535_, _01534_);
  nor _24508_ (_01536_, _10967_, _01530_);
  or _24509_ (_01537_, _01536_, _01531_);
  and _24510_ (_01538_, _01537_, _10970_);
  and _24511_ (_01539_, _01538_, _01535_);
  nor _24512_ (_01540_, _01538_, _01535_);
  nor _24513_ (_01541_, _01540_, _01539_);
  or _24514_ (_01542_, _01541_, _08374_);
  or _24515_ (_01543_, _08373_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _24516_ (_01544_, _01543_, _10894_);
  and _24517_ (_01545_, _01544_, _01542_);
  and _24518_ (_01546_, _10976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  or _24519_ (_01846_, _01546_, _01545_);
  not _24520_ (_01547_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  not _24521_ (_01548_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  not _24522_ (_01549_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and _24523_ (_01550_, _01532_, _01549_);
  and _24524_ (_01551_, _01550_, _01548_);
  nor _24525_ (_01552_, _01551_, _01547_);
  and _24526_ (_01553_, _01551_, _01547_);
  nor _24527_ (_01554_, _01553_, _01552_);
  not _24528_ (_01555_, _01554_);
  nor _24529_ (_01556_, _01550_, _01548_);
  or _24530_ (_01557_, _01556_, _01551_);
  nor _24531_ (_01558_, _01532_, _01549_);
  nor _24532_ (_01559_, _01558_, _01550_);
  not _24533_ (_01561_, _01559_);
  and _24534_ (_01562_, _01561_, _01539_);
  and _24535_ (_01563_, _01562_, _01557_);
  and _24536_ (_01564_, _01563_, _01555_);
  nor _24537_ (_01565_, _01563_, _01555_);
  nor _24538_ (_01566_, _01565_, _01564_);
  or _24539_ (_01567_, _01566_, _08374_);
  or _24540_ (_01568_, _08373_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and _24541_ (_01569_, _01568_, _10894_);
  and _24542_ (_01570_, _01569_, _01567_);
  and _24543_ (_01571_, _10976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or _24544_ (_01849_, _01571_, _01570_);
  nor _24545_ (_01572_, _01562_, _01557_);
  nor _24546_ (_01573_, _01572_, _01563_);
  or _24547_ (_01574_, _01573_, _08374_);
  or _24548_ (_01575_, _08373_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and _24549_ (_01576_, _01575_, _10894_);
  and _24550_ (_01577_, _01576_, _01574_);
  and _24551_ (_01578_, _10976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or _24552_ (_01854_, _01578_, _01577_);
  and _24553_ (_01579_, _08064_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  not _24554_ (_01580_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nor _24555_ (_01581_, _08064_, _01580_);
  or _24556_ (_01582_, _01581_, _01579_);
  and _24557_ (_01974_, _01582_, _06444_);
  and _24558_ (_01583_, _10976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor _24559_ (_01584_, _01561_, _01539_);
  nor _24560_ (_01585_, _01584_, _01562_);
  or _24561_ (_01586_, _01585_, _08374_);
  or _24562_ (_01587_, _08373_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _24563_ (_01588_, _01587_, _10894_);
  and _24564_ (_01589_, _01588_, _01586_);
  or _24565_ (_02013_, _01589_, _01583_);
  and _24566_ (_01590_, _08064_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  not _24567_ (_01591_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nor _24568_ (_01592_, _08064_, _01591_);
  or _24569_ (_01593_, _01592_, _01590_);
  and _24570_ (_02042_, _01593_, _06444_);
  nor _24571_ (_01594_, _01537_, _10970_);
  nor _24572_ (_01595_, _01594_, _01538_);
  or _24573_ (_01596_, _01595_, _08374_);
  or _24574_ (_01597_, _08373_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and _24575_ (_01598_, _01597_, _10894_);
  and _24576_ (_01599_, _01598_, _01596_);
  and _24577_ (_01600_, _10976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  or _24578_ (_02046_, _01600_, _01599_);
  and _24579_ (_01601_, _08064_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  not _24580_ (_01602_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nor _24581_ (_01603_, _08064_, _01602_);
  or _24582_ (_01604_, _01603_, _01601_);
  and _24583_ (_02090_, _01604_, _06444_);
  and _24584_ (_01605_, _07425_, _11568_);
  and _24585_ (_01606_, _09328_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  and _24586_ (_01607_, _06439_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  and _24587_ (_01608_, _01607_, _09332_);
  or _24588_ (_01609_, _01608_, _01606_);
  or _24589_ (_01610_, _01609_, _01605_);
  and _24590_ (_02146_, _01610_, _06444_);
  or _24591_ (_01611_, _13890_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  and _24592_ (_01612_, _01611_, _06444_);
  nand _24593_ (_01613_, _13893_, _06666_);
  and _24594_ (_02191_, _01613_, _01612_);
  or _24595_ (_01614_, _13890_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  and _24596_ (_01615_, _01614_, _06444_);
  nand _24597_ (_01616_, _13893_, _10494_);
  and _24598_ (_02204_, _01616_, _01615_);
  or _24599_ (_01617_, _09675_, _09347_);
  or _24600_ (_01618_, _09677_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and _24601_ (_01619_, _01618_, _06444_);
  and _24602_ (_02236_, _01619_, _01617_);
  or _24603_ (_01620_, _13931_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0]);
  nand _24604_ (_01621_, _13931_, _13919_);
  and _24605_ (_01622_, _01621_, _06444_);
  and _24606_ (_02250_, _01622_, _01620_);
  and _24607_ (_01623_, _06449_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  nor _24608_ (_01624_, _10494_, _06449_);
  or _24609_ (_01625_, _01624_, _01623_);
  and _24610_ (_02266_, _01625_, _06444_);
  nor _24611_ (_01626_, _07188_, _09146_);
  and _24612_ (_01627_, _09146_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  or _24613_ (_01628_, _01627_, _07158_);
  or _24614_ (_01629_, _01628_, _01626_);
  or _24615_ (_01630_, _06439_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  and _24616_ (_01631_, _01630_, _06444_);
  and _24617_ (_02269_, _01631_, _01629_);
  or _24618_ (_01632_, _13890_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  and _24619_ (_01633_, _01632_, _06444_);
  nand _24620_ (_01634_, _13893_, _07188_);
  and _24621_ (_02313_, _01634_, _01633_);
  and _24622_ (_02560_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _06444_);
  or _24623_ (_01635_, _07432_, \oc8051_top_1.oc8051_rom1.data_o [15]);
  nand _24624_ (_01636_, _07432_, _13980_);
  and _24625_ (_01637_, _01636_, _06444_);
  and _24626_ (_02566_, _01637_, _01635_);
  or _24627_ (_01638_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  nand _24628_ (_01639_, _07432_, _12633_);
  and _24629_ (_01640_, _01639_, _06444_);
  and _24630_ (_02583_, _01640_, _01638_);
  or _24631_ (_01642_, _13890_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  and _24632_ (_01643_, _01642_, _06444_);
  nand _24633_ (_01644_, _13893_, _07300_);
  and _24634_ (_02632_, _01644_, _01643_);
  and _24635_ (_01645_, _09527_, _07148_);
  and _24636_ (_01646_, _07190_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  or _24637_ (_01647_, _01646_, _01645_);
  or _24638_ (_01648_, _06439_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  and _24639_ (_01649_, _01648_, _06444_);
  and _24640_ (_02645_, _01649_, _01647_);
  or _24641_ (_01651_, _14512_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and _24642_ (_01652_, _01651_, _06444_);
  nand _24643_ (_01653_, _14512_, _06978_);
  and _24644_ (_02649_, _01653_, _01652_);
  nand _24645_ (_01654_, _14532_, _06978_);
  or _24646_ (_01655_, _00046_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand _24647_ (_01656_, _01655_, _00028_);
  and _24648_ (_01657_, _00046_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nor _24649_ (_01658_, _01657_, _01656_);
  and _24650_ (_01659_, _00016_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and _24651_ (_01660_, _01659_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or _24652_ (_01661_, _01659_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand _24653_ (_01662_, _01661_, _00015_);
  nor _24654_ (_01663_, _01662_, _01660_);
  and _24655_ (_01664_, _00052_, _14535_);
  or _24656_ (_01665_, _01664_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand _24657_ (_01666_, _01664_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and _24658_ (_01667_, _01666_, _01665_);
  and _24659_ (_01668_, _01667_, _14537_);
  or _24660_ (_01669_, _01668_, _01663_);
  or _24661_ (_01670_, _01669_, _01658_);
  or _24662_ (_01671_, _01670_, _14532_);
  and _24663_ (_01672_, _01671_, _00040_);
  and _24664_ (_01673_, _01672_, _01654_);
  and _24665_ (_01674_, _00039_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or _24666_ (_01675_, _01674_, _01673_);
  and _24667_ (_02652_, _01675_, _06444_);
  not _24668_ (_01677_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 );
  nor _24669_ (_01678_, _00011_, _01677_);
  or _24670_ (_01680_, _01678_, _01660_);
  and _24671_ (_01681_, _01680_, _00015_);
  not _24672_ (_01682_, _14532_);
  nor _24673_ (_01683_, _00039_, rst);
  and _24674_ (_01685_, _01683_, _01682_);
  and _24675_ (_02658_, _01685_, _01681_);
  nand _24676_ (_01686_, _00039_, _06978_);
  not _24677_ (_01687_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and _24678_ (_01688_, _00029_, _00002_);
  and _24679_ (_01689_, _01688_, _01682_);
  nor _24680_ (_01690_, _01689_, _01687_);
  and _24681_ (_01691_, _01689_, _01687_);
  or _24682_ (_01692_, _01691_, _01690_);
  and _24683_ (_01693_, _00115_, _00002_);
  nand _24684_ (_01694_, _01693_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nor _24685_ (_01695_, _01694_, _14532_);
  or _24686_ (_01696_, _01695_, _01692_);
  or _24687_ (_01698_, _01696_, _00039_);
  and _24688_ (_01699_, _01698_, _06444_);
  and _24689_ (_02661_, _01699_, _01686_);
  not _24690_ (_01701_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  nor _24691_ (_01703_, _14549_, _01701_);
  or _24692_ (_01704_, _01703_, _01657_);
  and _24693_ (_01705_, _01704_, _00028_);
  and _24694_ (_01706_, _00052_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or _24695_ (_01707_, _01706_, _01703_);
  and _24696_ (_01709_, _01707_, _14536_);
  or _24697_ (_01710_, _01703_, _00003_);
  and _24698_ (_01711_, _01710_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  or _24699_ (_01712_, _01711_, _01709_);
  or _24700_ (_01713_, _01712_, _01705_);
  and _24701_ (_02664_, _01713_, _01685_);
  and _24702_ (_01714_, _00517_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  not _24703_ (_01715_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  nor _24704_ (_01717_, _00347_, _01715_);
  and _24705_ (_01718_, _01717_, _00481_);
  or _24706_ (_01719_, _01718_, _01714_);
  and _24707_ (_01720_, _00347_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and _24708_ (_01721_, _01720_, _00349_);
  and _24709_ (_01722_, _01721_, _00374_);
  and _24710_ (_01723_, _01722_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  or _24711_ (_01724_, _01723_, _01717_);
  and _24712_ (_01725_, _01724_, _00366_);
  or _24713_ (_01726_, _01725_, _01719_);
  and _24714_ (_01727_, _00363_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  or _24715_ (_01728_, _01727_, _01717_);
  and _24716_ (_01729_, _01728_, _00361_);
  or _24717_ (_01730_, _01729_, _00536_);
  or _24718_ (_01731_, _01730_, _01726_);
  and _24719_ (_01732_, _01731_, _06444_);
  nand _24720_ (_01733_, _01732_, _00388_);
  nor _24721_ (_02666_, _01733_, _00334_);
  and _24722_ (_02670_, t0_i, _06444_);
  nand _24723_ (_01735_, _00334_, _06978_);
  or _24724_ (_01736_, _00363_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor _24725_ (_01737_, _01727_, _00362_);
  and _24726_ (_01738_, _01737_, _01736_);
  and _24727_ (_01739_, _00379_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  or _24728_ (_01740_, _00377_, _00395_);
  nor _24729_ (_01741_, _01740_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  or _24730_ (_01742_, _01741_, _01739_);
  or _24731_ (_01743_, _01742_, _01738_);
  or _24732_ (_01744_, _01743_, _00334_);
  and _24733_ (_01745_, _01744_, _00388_);
  and _24734_ (_01746_, _01745_, _01735_);
  and _24735_ (_01747_, _00387_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  or _24736_ (_01748_, _01747_, _01746_);
  and _24737_ (_02673_, _01748_, _06444_);
  nand _24738_ (_01749_, _00387_, _06978_);
  nor _24739_ (_01750_, _00497_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  nor _24740_ (_01751_, _01750_, _00487_);
  and _24741_ (_01753_, _01751_, _00483_);
  and _24742_ (_01754_, _00485_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  nand _24743_ (_01755_, _00488_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor _24744_ (_01756_, _01755_, _00334_);
  or _24745_ (_01757_, _01756_, _01754_);
  or _24746_ (_01758_, _01757_, _01753_);
  or _24747_ (_01759_, _01758_, _00387_);
  and _24748_ (_01760_, _01759_, _06444_);
  and _24749_ (_02676_, _01760_, _01749_);
  and _24750_ (_02679_, t1_i, _06444_);
  nand _24751_ (_01761_, _12829_, _06978_);
  or _24752_ (_01762_, _12829_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  and _24753_ (_01763_, _01762_, _06444_);
  and _24754_ (_02763_, _01763_, _01761_);
  and _24755_ (_01764_, _01079_, _06432_);
  nand _24756_ (_01765_, _01764_, _06930_);
  or _24757_ (_01766_, _01764_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and _24758_ (_01767_, _01766_, _06674_);
  and _24759_ (_01768_, _01767_, _01765_);
  nor _24760_ (_01769_, _01087_, _07069_);
  and _24761_ (_01770_, _01087_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or _24762_ (_01771_, _01770_, _01769_);
  and _24763_ (_01772_, _01771_, _06440_);
  and _24764_ (_01773_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or _24765_ (_01774_, _01773_, rst);
  or _24766_ (_01775_, _01774_, _01772_);
  or _24767_ (_02879_, _01775_, _01768_);
  and _24768_ (_01776_, _01079_, _06987_);
  nand _24769_ (_01777_, _01776_, _06930_);
  or _24770_ (_01778_, _01776_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and _24771_ (_01779_, _01778_, _06674_);
  and _24772_ (_01780_, _01779_, _01777_);
  nor _24773_ (_01781_, _01087_, _06666_);
  and _24774_ (_01782_, _01087_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or _24775_ (_01783_, _01782_, _01781_);
  and _24776_ (_01784_, _01783_, _06440_);
  and _24777_ (_01785_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or _24778_ (_01787_, _01785_, rst);
  or _24779_ (_01788_, _01787_, _01784_);
  or _24780_ (_02881_, _01788_, _01780_);
  and _24781_ (_01789_, _08913_, _06432_);
  nand _24782_ (_01791_, _01789_, _06930_);
  or _24783_ (_01792_, _01789_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and _24784_ (_01793_, _01792_, _06674_);
  and _24785_ (_01794_, _01793_, _01791_);
  and _24786_ (_01795_, _08919_, _07070_);
  and _24787_ (_01796_, _08920_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or _24788_ (_01797_, _01796_, _01795_);
  and _24789_ (_01798_, _01797_, _06440_);
  and _24790_ (_01799_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or _24791_ (_01800_, _01799_, rst);
  or _24792_ (_01801_, _01800_, _01798_);
  or _24793_ (_02883_, _01801_, _01794_);
  and _24794_ (_01802_, _08913_, _06987_);
  nand _24795_ (_01804_, _01802_, _06930_);
  or _24796_ (_01805_, _01802_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and _24797_ (_01807_, _01805_, _06674_);
  and _24798_ (_01809_, _01807_, _01804_);
  nor _24799_ (_01811_, _08920_, _06666_);
  and _24800_ (_01812_, _08920_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or _24801_ (_01813_, _01812_, _01811_);
  and _24802_ (_01814_, _01813_, _06440_);
  and _24803_ (_01815_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or _24804_ (_01816_, _01815_, rst);
  or _24805_ (_01817_, _01816_, _01814_);
  or _24806_ (_02886_, _01817_, _01809_);
  and _24807_ (_01818_, _00605_, _08977_);
  nand _24808_ (_01819_, _01818_, _06930_);
  or _24809_ (_01820_, _01818_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and _24810_ (_01821_, _01820_, _06674_);
  and _24811_ (_01822_, _01821_, _01819_);
  nand _24812_ (_01823_, _11589_, _00612_);
  or _24813_ (_01824_, _00612_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and _24814_ (_01825_, _01824_, _06440_);
  and _24815_ (_01826_, _01825_, _01823_);
  and _24816_ (_01827_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  or _24817_ (_01828_, _01827_, rst);
  or _24818_ (_01829_, _01828_, _01826_);
  or _24819_ (_02888_, _01829_, _01822_);
  and _24820_ (_01830_, _00640_, _06987_);
  nand _24821_ (_01831_, _01830_, _06930_);
  or _24822_ (_01832_, _01830_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and _24823_ (_01833_, _01832_, _06674_);
  and _24824_ (_01834_, _01833_, _01831_);
  nand _24825_ (_01835_, _00646_, _06666_);
  or _24826_ (_01836_, _00646_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and _24827_ (_01837_, _01836_, _06440_);
  and _24828_ (_01838_, _01837_, _01835_);
  and _24829_ (_01839_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  or _24830_ (_01840_, _01839_, rst);
  or _24831_ (_01841_, _01840_, _01838_);
  or _24832_ (_02890_, _01841_, _01834_);
  and _24833_ (_01842_, _07402_, _07043_);
  nand _24834_ (_01843_, _01842_, _06930_);
  or _24835_ (_01844_, _01842_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and _24836_ (_01845_, _01844_, _06674_);
  and _24837_ (_01847_, _01845_, _01843_);
  nand _24838_ (_01848_, _00646_, _07069_);
  or _24839_ (_01850_, _00646_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and _24840_ (_01851_, _01850_, _06440_);
  and _24841_ (_01852_, _01851_, _01848_);
  and _24842_ (_01853_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  or _24843_ (_01855_, _01853_, rst);
  or _24844_ (_01856_, _01855_, _01852_);
  or _24845_ (_02893_, _01856_, _01847_);
  and _24846_ (_01857_, _08064_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor _24847_ (_01858_, _08064_, _01150_);
  or _24848_ (_01859_, _01858_, _01857_);
  and _24849_ (_02898_, _01859_, _06444_);
  and _24850_ (_01860_, _06934_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or _24851_ (_01861_, _01860_, _06935_);
  and _24852_ (_01862_, _01861_, _12012_);
  nand _24853_ (_01863_, _12008_, _06930_);
  nor _24854_ (_01864_, _12008_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor _24855_ (_01865_, _01864_, _12012_);
  and _24856_ (_01866_, _01865_, _01863_);
  or _24857_ (_01867_, _01866_, _07218_);
  or _24858_ (_01868_, _01867_, _01862_);
  nand _24859_ (_01869_, _07218_, _06978_);
  and _24860_ (_01870_, _01869_, _06444_);
  and _24861_ (_02905_, _01870_, _01868_);
  and _24862_ (_01871_, _08064_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  not _24863_ (_01872_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nor _24864_ (_01873_, _08064_, _01872_);
  or _24865_ (_01874_, _01873_, _01871_);
  and _24866_ (_02908_, _01874_, _06444_);
  and _24867_ (_01875_, _01079_, _06942_);
  nand _24868_ (_01876_, _01875_, _06930_);
  or _24869_ (_01877_, _01875_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and _24870_ (_01878_, _01877_, _06674_);
  and _24871_ (_01879_, _01878_, _01876_);
  and _24872_ (_01880_, _01086_, _09527_);
  and _24873_ (_01881_, _01087_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  or _24874_ (_01882_, _01881_, _01880_);
  and _24875_ (_01883_, _01882_, _06440_);
  and _24876_ (_01884_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  or _24877_ (_01885_, _01884_, rst);
  or _24878_ (_01886_, _01885_, _01883_);
  or _24879_ (_02914_, _01886_, _01879_);
  and _24880_ (_01887_, _01079_, _08310_);
  nand _24881_ (_01888_, _01887_, _06930_);
  or _24882_ (_01889_, _01887_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and _24883_ (_01890_, _01889_, _06674_);
  and _24884_ (_01891_, _01890_, _01888_);
  nor _24885_ (_01892_, _01087_, _07300_);
  and _24886_ (_01893_, _01087_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or _24887_ (_01894_, _01893_, _01892_);
  and _24888_ (_01895_, _01894_, _06440_);
  and _24889_ (_01896_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or _24890_ (_01897_, _01896_, rst);
  or _24891_ (_01898_, _01897_, _01895_);
  or _24892_ (_02916_, _01898_, _01891_);
  and _24893_ (_01899_, _00605_, _00240_);
  nand _24894_ (_01900_, _01899_, _06930_);
  or _24895_ (_01901_, _01899_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and _24896_ (_01902_, _01901_, _06674_);
  and _24897_ (_01903_, _01902_, _01900_);
  nand _24898_ (_01904_, _10494_, _00612_);
  or _24899_ (_01905_, _00612_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and _24900_ (_01906_, _01905_, _06440_);
  and _24901_ (_01907_, _01906_, _01904_);
  and _24902_ (_01908_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  or _24903_ (_01909_, _01908_, rst);
  or _24904_ (_01910_, _01909_, _01907_);
  or _24905_ (_02919_, _01910_, _01903_);
  nand _24906_ (_01911_, _00612_, _06930_);
  or _24907_ (_01912_, _00612_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and _24908_ (_01913_, _01912_, _06674_);
  and _24909_ (_01914_, _01913_, _01911_);
  nand _24910_ (_01915_, _09526_, _00612_);
  and _24911_ (_01916_, _01915_, _06440_);
  and _24912_ (_01917_, _01916_, _01912_);
  and _24913_ (_01918_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  or _24914_ (_01919_, _01918_, rst);
  or _24915_ (_01920_, _01919_, _01917_);
  or _24916_ (_02921_, _01920_, _01914_);
  nand _24917_ (_01921_, _00646_, _06930_);
  or _24918_ (_01922_, _00646_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  and _24919_ (_01923_, _01922_, _06674_);
  and _24920_ (_01924_, _01923_, _01921_);
  nand _24921_ (_01925_, _09526_, _00646_);
  and _24922_ (_01926_, _01922_, _06440_);
  and _24923_ (_01927_, _01926_, _01925_);
  and _24924_ (_01928_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  or _24925_ (_01929_, _01928_, rst);
  or _24926_ (_01930_, _01929_, _01927_);
  or _24927_ (_02924_, _01930_, _01924_);
  and _24928_ (_01931_, _00640_, _08310_);
  nand _24929_ (_01932_, _01931_, _06930_);
  or _24930_ (_01933_, _01931_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and _24931_ (_01934_, _01933_, _06674_);
  and _24932_ (_01935_, _01934_, _01932_);
  nand _24933_ (_01937_, _00646_, _07300_);
  or _24934_ (_01938_, _00646_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and _24935_ (_01939_, _01938_, _06440_);
  and _24936_ (_01940_, _01939_, _01937_);
  and _24937_ (_01941_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or _24938_ (_01942_, _01941_, rst);
  or _24939_ (_01943_, _01942_, _01940_);
  or _24940_ (_02926_, _01943_, _01935_);
  and _24941_ (_01944_, _08064_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor _24942_ (_01945_, _08064_, _01076_);
  or _24943_ (_01946_, _01945_, _01944_);
  and _24944_ (_02945_, _01946_, _06444_);
  nand _24945_ (_01947_, _12829_, _09526_);
  or _24946_ (_01948_, _12829_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  and _24947_ (_01949_, _01948_, _01947_);
  and _24948_ (_03036_, _01949_, _06444_);
  and _24949_ (_01950_, _00605_, _06987_);
  nand _24950_ (_01951_, _01950_, _06930_);
  or _24951_ (_01952_, _01950_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and _24952_ (_01953_, _01952_, _06674_);
  and _24953_ (_01954_, _01953_, _01951_);
  nand _24954_ (_01955_, _00612_, _06666_);
  or _24955_ (_01956_, _00612_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and _24956_ (_01957_, _01956_, _06440_);
  and _24957_ (_01958_, _01957_, _01955_);
  and _24958_ (_01959_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  or _24959_ (_01960_, _01959_, rst);
  or _24960_ (_01961_, _01960_, _01958_);
  or _24961_ (_03040_, _01961_, _01954_);
  and _24962_ (_01962_, _00605_, _06983_);
  nand _24963_ (_01963_, _01962_, _06930_);
  or _24964_ (_01964_, _01962_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and _24965_ (_01965_, _01964_, _06674_);
  and _24966_ (_01966_, _01965_, _01963_);
  nand _24967_ (_01967_, _00612_, _07188_);
  or _24968_ (_01968_, _00612_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and _24969_ (_01969_, _01968_, _06440_);
  and _24970_ (_01970_, _01969_, _01967_);
  and _24971_ (_01971_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  or _24972_ (_01972_, _01971_, rst);
  or _24973_ (_01973_, _01972_, _01970_);
  or _24974_ (_03042_, _01973_, _01966_);
  and _24975_ (_01975_, _08913_, _06983_);
  nand _24976_ (_01976_, _01975_, _06930_);
  or _24977_ (_01977_, _01975_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and _24978_ (_01978_, _01977_, _06674_);
  and _24979_ (_01979_, _01978_, _01976_);
  nor _24980_ (_01980_, _08920_, _07188_);
  and _24981_ (_01981_, _08920_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or _24982_ (_01982_, _01981_, _01980_);
  and _24983_ (_01983_, _01982_, _06440_);
  and _24984_ (_01984_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or _24985_ (_01985_, _01984_, rst);
  or _24986_ (_01986_, _01985_, _01983_);
  or _24987_ (_03044_, _01986_, _01979_);
  and _24988_ (_01987_, _08913_, _08310_);
  nand _24989_ (_01988_, _01987_, _06930_);
  or _24990_ (_01989_, _01987_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and _24991_ (_01990_, _01989_, _06674_);
  and _24992_ (_01991_, _01990_, _01988_);
  nor _24993_ (_01992_, _08920_, _07300_);
  and _24994_ (_01993_, _08920_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or _24995_ (_01994_, _01993_, _01992_);
  and _24996_ (_01995_, _01994_, _06440_);
  and _24997_ (_01996_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or _24998_ (_01997_, _01996_, rst);
  or _24999_ (_01998_, _01997_, _01995_);
  or _25000_ (_03046_, _01998_, _01991_);
  nand _25001_ (_01999_, _13890_, _11589_);
  or _25002_ (_02000_, _13890_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  and _25003_ (_02001_, _02000_, _06444_);
  and _25004_ (_03049_, _02001_, _01999_);
  nand _25005_ (_02002_, _13890_, _07069_);
  or _25006_ (_02003_, _13890_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  and _25007_ (_02004_, _02003_, _06444_);
  and _25008_ (_03061_, _02004_, _02002_);
  and _25009_ (_02005_, _00640_, _00240_);
  nand _25010_ (_02006_, _02005_, _06930_);
  or _25011_ (_02007_, _02005_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and _25012_ (_02008_, _02007_, _06674_);
  and _25013_ (_02009_, _02008_, _02006_);
  nand _25014_ (_02010_, _10494_, _00646_);
  or _25015_ (_02011_, _00646_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and _25016_ (_02012_, _02011_, _06440_);
  and _25017_ (_02014_, _02012_, _02010_);
  and _25018_ (_02015_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  or _25019_ (_02016_, _02015_, rst);
  or _25020_ (_02017_, _02016_, _02014_);
  or _25021_ (_03070_, _02017_, _02009_);
  and _25022_ (_02018_, _00640_, _06983_);
  nand _25023_ (_02019_, _02018_, _06930_);
  or _25024_ (_02020_, _02018_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and _25025_ (_02021_, _02020_, _06674_);
  and _25026_ (_02022_, _02021_, _02019_);
  nand _25027_ (_02023_, _00646_, _07188_);
  or _25028_ (_02024_, _00646_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and _25029_ (_02025_, _02024_, _06440_);
  and _25030_ (_02026_, _02025_, _02023_);
  and _25031_ (_02027_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or _25032_ (_02028_, _02027_, rst);
  or _25033_ (_02029_, _02028_, _02026_);
  or _25034_ (_03072_, _02029_, _02022_);
  not _25035_ (_02030_, _00640_);
  or _25036_ (_02031_, _02030_, _00717_);
  and _25037_ (_02032_, _02031_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and _25038_ (_02033_, _06431_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or _25039_ (_02034_, _02033_, _00713_);
  and _25040_ (_02035_, _02034_, _00640_);
  or _25041_ (_02036_, _02035_, _02032_);
  and _25042_ (_02037_, _02036_, _06674_);
  nand _25043_ (_02038_, _11589_, _00646_);
  or _25044_ (_02039_, _00646_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and _25045_ (_02040_, _02039_, _06440_);
  and _25046_ (_02041_, _02040_, _02038_);
  and _25047_ (_02043_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or _25048_ (_02044_, _02043_, rst);
  or _25049_ (_02045_, _02044_, _02041_);
  or _25050_ (_03074_, _02045_, _02037_);
  and _25051_ (_02047_, _00605_, _08310_);
  nand _25052_ (_02048_, _02047_, _06930_);
  or _25053_ (_02049_, _02047_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and _25054_ (_02050_, _02049_, _06674_);
  and _25055_ (_02051_, _02050_, _02048_);
  nand _25056_ (_02052_, _00612_, _07300_);
  or _25057_ (_02053_, _00612_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and _25058_ (_02054_, _02053_, _06440_);
  and _25059_ (_02055_, _02054_, _02052_);
  and _25060_ (_02056_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or _25061_ (_02057_, _02056_, rst);
  or _25062_ (_02058_, _02057_, _02055_);
  or _25063_ (_03076_, _02058_, _02051_);
  and _25064_ (_02059_, _08913_, _00240_);
  nand _25065_ (_02060_, _02059_, _06930_);
  or _25066_ (_02061_, _02059_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and _25067_ (_02062_, _02061_, _06674_);
  and _25068_ (_02063_, _02062_, _02060_);
  nor _25069_ (_02064_, _10494_, _08920_);
  and _25070_ (_02065_, _08920_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or _25071_ (_02066_, _02065_, _02064_);
  and _25072_ (_02067_, _02066_, _06440_);
  and _25073_ (_02068_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or _25074_ (_02069_, _02068_, rst);
  or _25075_ (_02070_, _02069_, _02067_);
  or _25076_ (_03078_, _02070_, _02063_);
  and _25077_ (_02071_, _00605_, _06432_);
  nand _25078_ (_02072_, _02071_, _06930_);
  or _25079_ (_02073_, _02071_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and _25080_ (_02074_, _02073_, _06674_);
  and _25081_ (_02075_, _02074_, _02072_);
  or _25082_ (_02076_, _00612_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  nand _25083_ (_02077_, _00612_, _07069_);
  and _25084_ (_02078_, _02077_, _06440_);
  and _25085_ (_02079_, _02078_, _02076_);
  and _25086_ (_02080_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  or _25087_ (_02081_, _02080_, rst);
  or _25088_ (_02082_, _02081_, _02079_);
  or _25089_ (_03080_, _02082_, _02075_);
  and _25090_ (_02083_, _08913_, _08977_);
  nand _25091_ (_02084_, _02083_, _06930_);
  or _25092_ (_02085_, _02083_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and _25093_ (_02086_, _02085_, _06674_);
  and _25094_ (_02087_, _02086_, _02084_);
  nor _25095_ (_02088_, _11589_, _08920_);
  and _25096_ (_02089_, _08920_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or _25097_ (_02091_, _02089_, _02088_);
  and _25098_ (_02092_, _02091_, _06440_);
  and _25099_ (_02093_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or _25100_ (_02094_, _02093_, rst);
  or _25101_ (_02095_, _02094_, _02092_);
  or _25102_ (_03081_, _02095_, _02087_);
  nand _25103_ (_02096_, _08919_, _06930_);
  or _25104_ (_02097_, _08919_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and _25105_ (_02098_, _02097_, _06674_);
  and _25106_ (_02099_, _02098_, _02096_);
  and _25107_ (_02100_, _09527_, _08919_);
  and _25108_ (_02101_, _08920_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  or _25109_ (_02102_, _02101_, _02100_);
  and _25110_ (_02103_, _02102_, _06440_);
  and _25111_ (_02104_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  or _25112_ (_02105_, _02104_, rst);
  or _25113_ (_02106_, _02105_, _02103_);
  or _25114_ (_03084_, _02106_, _02099_);
  and _25115_ (_02107_, _01079_, _00240_);
  nand _25116_ (_02108_, _02107_, _06930_);
  or _25117_ (_02109_, _02107_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and _25118_ (_02110_, _02109_, _06674_);
  and _25119_ (_02111_, _02110_, _02108_);
  nor _25120_ (_02112_, _01087_, _10494_);
  and _25121_ (_02113_, _01087_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or _25122_ (_02114_, _02113_, _02112_);
  and _25123_ (_02115_, _02114_, _06440_);
  and _25124_ (_02116_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or _25125_ (_02117_, _02116_, rst);
  or _25126_ (_02118_, _02117_, _02115_);
  or _25127_ (_03086_, _02118_, _02111_);
  and _25128_ (_02119_, _01079_, _06983_);
  nand _25129_ (_02120_, _02119_, _06930_);
  or _25130_ (_02121_, _02119_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and _25131_ (_02122_, _02121_, _06674_);
  and _25132_ (_02123_, _02122_, _02120_);
  nor _25133_ (_02124_, _01087_, _07188_);
  and _25134_ (_02125_, _01087_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or _25135_ (_02126_, _02125_, _02124_);
  and _25136_ (_02127_, _02126_, _06440_);
  and _25137_ (_02128_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or _25138_ (_02129_, _02128_, rst);
  or _25139_ (_02130_, _02129_, _02127_);
  or _25140_ (_03088_, _02130_, _02123_);
  and _25141_ (_02131_, _01079_, _08977_);
  nand _25142_ (_02132_, _02131_, _06930_);
  or _25143_ (_02133_, _02131_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and _25144_ (_02134_, _02133_, _06674_);
  and _25145_ (_02135_, _02134_, _02132_);
  nor _25146_ (_02136_, _01087_, _11589_);
  and _25147_ (_02137_, _01087_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or _25148_ (_02138_, _02137_, _02136_);
  and _25149_ (_02139_, _02138_, _06440_);
  and _25150_ (_02140_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or _25151_ (_02141_, _02140_, rst);
  or _25152_ (_02142_, _02141_, _02139_);
  or _25153_ (_03091_, _02142_, _02135_);
  nand _25154_ (_02143_, _13890_, _09526_);
  or _25155_ (_02144_, _13890_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  and _25156_ (_02145_, _02144_, _06444_);
  and _25157_ (_03118_, _02145_, _02143_);
  and _25158_ (_03132_, _01286_, _06444_);
  and _25159_ (_03406_, \oc8051_top_1.oc8051_memory_interface1.istb_t , _06444_);
  and _25160_ (_02147_, _03406_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or _25161_ (_03144_, _02147_, _03132_);
  or _25162_ (_02148_, _07432_, \oc8051_top_1.oc8051_rom1.data_o [13]);
  nand _25163_ (_02149_, _07432_, _13990_);
  and _25164_ (_02150_, _02149_, _06444_);
  and _25165_ (_03147_, _02150_, _02148_);
  nand _25166_ (_02151_, _07226_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _25167_ (_03150_, _02151_, _06444_);
  and _25168_ (_03196_, _00287_, _11574_);
  and _25169_ (_03293_, _07982_, _06444_);
  nor _25170_ (_02152_, _07432_, _07429_);
  nand _25171_ (_02153_, _01135_, _01132_);
  and _25172_ (_02154_, _02153_, _07230_);
  and _25173_ (_02155_, _02154_, _07235_);
  nor _25174_ (_02156_, _02154_, _07235_);
  nor _25175_ (_02157_, _02156_, _02155_);
  nor _25176_ (_02158_, _02157_, _02152_);
  and _25177_ (_02159_, _07240_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and _25178_ (_02160_, _02159_, _02152_);
  and _25179_ (_02161_, _02160_, _10890_);
  or _25180_ (_02162_, _02161_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _25181_ (_02163_, _02162_, _02158_);
  and _25182_ (_03295_, _02163_, _06444_);
  and _25183_ (_03300_, _11622_, _06444_);
  and _25184_ (_02164_, _12712_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  or _25185_ (_02165_, _02164_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  and _25186_ (_03304_, _02165_, _06444_);
  and _25187_ (_03307_, _01491_, _06444_);
  not _25188_ (_02166_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  nand _25189_ (_02167_, _07230_, _02166_);
  nand _25190_ (_02168_, _02167_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nand _25191_ (_02169_, _02168_, _12712_);
  and _25192_ (_03309_, _02169_, _06444_);
  and _25193_ (_02170_, _14070_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  and _25194_ (_02171_, _12841_, _07154_);
  or _25195_ (_02172_, _02171_, _02170_);
  and _25196_ (_03321_, _02172_, _06444_);
  nor _25197_ (_02173_, _12830_, _07188_);
  and _25198_ (_02174_, _01100_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  or _25199_ (_02175_, _02174_, _02173_);
  and _25200_ (_03325_, _02175_, _06444_);
  and _25201_ (_03331_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , _06444_);
  and _25202_ (_02176_, _07046_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  nor _25203_ (_02177_, _07188_, _07046_);
  or _25204_ (_02178_, _02177_, _02176_);
  and _25205_ (_03344_, _02178_, _06444_);
  nor _25206_ (_03350_, _01510_, rst);
  nor _25207_ (_02179_, _10946_, _10944_);
  nor _25208_ (_02180_, _02179_, _10947_);
  or _25209_ (_02181_, _02180_, _08374_);
  or _25210_ (_02182_, _08373_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and _25211_ (_02183_, _02182_, _10894_);
  and _25212_ (_02184_, _02183_, _02181_);
  and _25213_ (_02185_, _10976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  or _25214_ (_03355_, _02185_, _02184_);
  and _25215_ (_02186_, _14069_, _07070_);
  and _25216_ (_02187_, _14070_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  or _25217_ (_02188_, _02187_, _02186_);
  and _25218_ (_03357_, _02188_, _06444_);
  or _25219_ (_02189_, _10942_, _10940_);
  and _25220_ (_02190_, _02189_, _10943_);
  or _25221_ (_02192_, _02190_, _08374_);
  or _25222_ (_02193_, _08373_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and _25223_ (_02194_, _02193_, _10894_);
  and _25224_ (_02195_, _02194_, _02192_);
  and _25225_ (_02196_, _10976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or _25226_ (_03360_, _02196_, _02195_);
  nor _25227_ (_02197_, _10939_, _10891_);
  nor _25228_ (_02198_, _02197_, _10940_);
  or _25229_ (_02199_, _02198_, _08374_);
  or _25230_ (_02200_, _08373_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and _25231_ (_02201_, _02200_, _10894_);
  and _25232_ (_02202_, _02201_, _02199_);
  and _25233_ (_02203_, _10976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  or _25234_ (_03385_, _02203_, _02202_);
  not _25235_ (_02205_, _00599_);
  and _25236_ (_02206_, _02205_, _00597_);
  and _25237_ (_02207_, _00278_, _00592_);
  and _25238_ (_03398_, _02207_, _02206_);
  and _25239_ (_02208_, \oc8051_top_1.oc8051_memory_interface1.cdata [7], _08478_);
  and _25240_ (_02209_, \oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or _25241_ (_02210_, _02209_, _02208_);
  and _25242_ (_03414_, _02210_, _06444_);
  and _25243_ (_02211_, _11763_, _07425_);
  and _25244_ (_02212_, _09328_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  and _25245_ (_02213_, _06439_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  and _25246_ (_02214_, _02213_, _09332_);
  or _25247_ (_02215_, _02214_, _02212_);
  or _25248_ (_02216_, _02215_, _02211_);
  and _25249_ (_03425_, _02216_, _06444_);
  and _25250_ (_02217_, _08421_, _08356_);
  and _25251_ (_02218_, _02217_, _08453_);
  and _25252_ (_02219_, _08437_, _08405_);
  and _25253_ (_02220_, _02219_, _08468_);
  and _25254_ (_02221_, _07231_, _06444_);
  and _25255_ (_02222_, _02221_, _08388_);
  and _25256_ (_02223_, _02222_, _07259_);
  and _25257_ (_02224_, _02223_, _02220_);
  and _25258_ (_03428_, _02224_, _02218_);
  nor _25259_ (_02225_, _14070_, _06666_);
  and _25260_ (_02226_, _14070_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  or _25261_ (_02227_, _02226_, _02225_);
  and _25262_ (_03429_, _02227_, _06444_);
  or _25263_ (_02228_, _07432_, \oc8051_top_1.oc8051_rom1.data_o [19]);
  nand _25264_ (_02229_, _07432_, _11264_);
  and _25265_ (_02230_, _02229_, _06444_);
  and _25266_ (_03460_, _02230_, _02228_);
  and _25267_ (_02231_, _13934_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and _25268_ (_02232_, _09678_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and _25269_ (_02233_, _02232_, _13933_);
  or _25270_ (_02234_, _02233_, _02231_);
  and _25271_ (_03483_, _02234_, _06444_);
  and _25272_ (_02235_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and _25273_ (_02237_, _12223_, \oc8051_top_1.oc8051_rom1.data_o [21]);
  or _25274_ (_02238_, _02237_, _02235_);
  and _25275_ (_03495_, _02238_, _06444_);
  and _25276_ (_02239_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and _25277_ (_02240_, _12223_, \oc8051_top_1.oc8051_rom1.data_o [20]);
  or _25278_ (_02241_, _02240_, _02239_);
  and _25279_ (_03502_, _02241_, _06444_);
  not _25280_ (_02242_, _00850_);
  or _25281_ (_02243_, _02242_, _07198_);
  and _25282_ (_02244_, _00850_, _07208_);
  and _25283_ (_02245_, _02244_, _07206_);
  or _25284_ (_02246_, _02245_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  and _25285_ (_02247_, _02246_, _06444_);
  and _25286_ (_03515_, _02247_, _02243_);
  nor _25287_ (_03523_, _11570_, rst);
  nor _25288_ (_03532_, _07222_, rst);
  and _25289_ (_02248_, _11443_, _11385_);
  and _25290_ (_02249_, _11408_, _11394_);
  or _25291_ (_02251_, _02249_, _11483_);
  or _25292_ (_02252_, _02251_, _02248_);
  and _25293_ (_02253_, _11394_, _11523_);
  and _25294_ (_02254_, _11394_, _11493_);
  and _25295_ (_02255_, _11394_, _11458_);
  or _25296_ (_02256_, _02255_, _02254_);
  or _25297_ (_02257_, _02256_, _02253_);
  or _25298_ (_02258_, _11519_, _11394_);
  and _25299_ (_02259_, _02258_, _11418_);
  and _25300_ (_02260_, _11426_, _11355_);
  or _25301_ (_02261_, _02260_, _02259_);
  or _25302_ (_02262_, _02261_, _02257_);
  and _25303_ (_02263_, _11433_, _11965_);
  and _25304_ (_02264_, _11443_, _11965_);
  or _25305_ (_02265_, _02264_, _02263_);
  or _25306_ (_02267_, _02265_, _11379_);
  and _25307_ (_02268_, _11370_, _11423_);
  and _25308_ (_02270_, _11528_, _11418_);
  or _25309_ (_02271_, _14240_, _02270_);
  or _25310_ (_02272_, _02271_, _02268_);
  or _25311_ (_02273_, _02272_, _02267_);
  or _25312_ (_02274_, _02273_, _02262_);
  and _25313_ (_02275_, _11431_, _11965_);
  and _25314_ (_02276_, _11407_, _11976_);
  and _25315_ (_02277_, _11431_, _11526_);
  or _25316_ (_02278_, _02277_, _02276_);
  and _25317_ (_02279_, _11370_, _11976_);
  or _25318_ (_02280_, _02279_, _11439_);
  or _25319_ (_02281_, _02280_, _02278_);
  or _25320_ (_02282_, _02281_, _02275_);
  and _25321_ (_02283_, _11394_, _11475_);
  or _25322_ (_02284_, _02283_, _14234_);
  and _25323_ (_02285_, _11519_, _11407_);
  or _25324_ (_02286_, _02285_, _11537_);
  or _25325_ (_02287_, _02286_, _02284_);
  or _25326_ (_02288_, _14225_, _14228_);
  or _25327_ (_02289_, _02288_, _02287_);
  or _25328_ (_02290_, _02289_, _02282_);
  or _25329_ (_02291_, _02290_, _02274_);
  or _25330_ (_02292_, _02291_, _02252_);
  and _25331_ (_02293_, _02292_, _07230_);
  and _25332_ (_02294_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  not _25333_ (_02295_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and _25334_ (_02296_, _11453_, _02295_);
  and _25335_ (_02297_, _11370_, _11355_);
  nor _25336_ (_02298_, _11385_, _11354_);
  not _25337_ (_02299_, _02298_);
  and _25338_ (_02300_, _02299_, _11419_);
  nor _25339_ (_02301_, _02300_, _02297_);
  not _25340_ (_02302_, _02301_);
  and _25341_ (_02303_, _02302_, _02296_);
  or _25342_ (_02304_, _02303_, _02294_);
  or _25343_ (_02305_, _02304_, _02293_);
  and _25344_ (_03537_, _02305_, _06444_);
  and _25345_ (_02306_, _06444_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and _25346_ (_02307_, _02306_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  or _25347_ (_02308_, _11394_, _11526_);
  and _25348_ (_02309_, _02308_, _11486_);
  and _25349_ (_02310_, _11528_, _11373_);
  or _25350_ (_02311_, _02310_, _11442_);
  or _25351_ (_02312_, _02311_, _11424_);
  or _25352_ (_02314_, _02312_, _02309_);
  not _25353_ (_02315_, _11430_);
  or _25354_ (_02316_, _11995_, _02315_);
  nand _25355_ (_02317_, _02316_, _11505_);
  or _25356_ (_02318_, _02317_, _02314_);
  or _25357_ (_02319_, _02318_, _02252_);
  or _25358_ (_02320_, _02264_, _14225_);
  or _25359_ (_02321_, _02320_, _02263_);
  and _25360_ (_02322_, _02321_, _07311_);
  and _25361_ (_02323_, _11519_, _11411_);
  or _25362_ (_02324_, _14234_, _02323_);
  and _25363_ (_02325_, _11395_, _11355_);
  or _25364_ (_02326_, _11419_, _11431_);
  and _25365_ (_02327_, _02326_, _11394_);
  or _25366_ (_02328_, _02327_, _02325_);
  or _25367_ (_02329_, _02328_, _02324_);
  or _25368_ (_02330_, _02329_, _02322_);
  or _25369_ (_02331_, _02330_, _02319_);
  and _25370_ (_02332_, _07230_, _06444_);
  and _25371_ (_02333_, _02332_, _02331_);
  or _25372_ (_03545_, _02333_, _02307_);
  and _25373_ (_02334_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or _25374_ (_02335_, _02334_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and _25375_ (_02336_, _06870_, _06847_);
  and _25376_ (_02337_, _06838_, _06680_);
  nand _25377_ (_02338_, _06640_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nand _25378_ (_02339_, _02338_, _02334_);
  or _25379_ (_02340_, _02339_, _02337_);
  or _25380_ (_02341_, _02340_, _02336_);
  and _25381_ (_02342_, _02341_, _02335_);
  or _25382_ (_02343_, _02342_, _12012_);
  or _25383_ (_02344_, _00240_, _08294_);
  nand _25384_ (_02345_, _02344_, _12012_);
  or _25385_ (_02346_, _02345_, _01481_);
  and _25386_ (_02347_, _02346_, _02343_);
  or _25387_ (_02348_, _02347_, _07218_);
  nand _25388_ (_02349_, _10494_, _07218_);
  and _25389_ (_02350_, _02349_, _06444_);
  and _25390_ (_03547_, _02350_, _02348_);
  and _25391_ (_02351_, _11459_, _11389_);
  not _25392_ (_02352_, _11399_);
  and _25393_ (_02353_, _02352_, _02296_);
  and _25394_ (_02354_, _11934_, _11347_);
  and _25395_ (_02355_, _11933_, _11347_);
  or _25396_ (_02356_, _02355_, _02354_);
  and _25397_ (_02357_, _02356_, _11389_);
  or _25398_ (_02358_, _02357_, _02353_);
  or _25399_ (_02359_, _02358_, _02351_);
  and _25400_ (_02360_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _25401_ (_02361_, _11524_, _11494_);
  or _25402_ (_02362_, _02361_, _11509_);
  not _25403_ (_02363_, _11354_);
  nor _25404_ (_02364_, _11995_, _02363_);
  or _25405_ (_02365_, _02364_, _02354_);
  or _25406_ (_02366_, _02365_, _02362_);
  and _25407_ (_02367_, _11482_, _11347_);
  and _25408_ (_02368_, _02367_, _11417_);
  or _25409_ (_02369_, _11534_, _11504_);
  or _25410_ (_02370_, _02369_, _02368_);
  nor _25411_ (_02371_, _11495_, _11413_);
  nand _25412_ (_02372_, _02371_, _11492_);
  or _25413_ (_02373_, _02372_, _02370_);
  or _25414_ (_02374_, _02373_, _02366_);
  not _25415_ (_02375_, _11513_);
  nand _25416_ (_02376_, _02375_, _11416_);
  and _25417_ (_02377_, _11519_, _11370_);
  or _25418_ (_02378_, _02377_, _02355_);
  or _25419_ (_02379_, _02378_, _02376_);
  or _25420_ (_02380_, _02379_, _02374_);
  and _25421_ (_02381_, _02380_, _07230_);
  or _25422_ (_02382_, _02381_, _02360_);
  or _25423_ (_02383_, _02382_, _02359_);
  and _25424_ (_03554_, _02383_, _06444_);
  and _25425_ (_02384_, _11423_, _11417_);
  or _25426_ (_02385_, _11529_, _11428_);
  or _25427_ (_02386_, _02385_, _02384_);
  and _25428_ (_02387_, _11413_, _11376_);
  or _25429_ (_02388_, _02387_, _11442_);
  or _25430_ (_02389_, _02388_, _02356_);
  or _25431_ (_02390_, _02389_, _02386_);
  and _25432_ (_02391_, _02390_, _07230_);
  and _25433_ (_02392_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _25434_ (_02393_, _02392_, _02358_);
  or _25435_ (_02394_, _02393_, _02391_);
  and _25436_ (_03573_, _02394_, _06444_);
  nand _25437_ (_02395_, _01480_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  nand _25438_ (_02396_, _02395_, _06678_);
  or _25439_ (_02397_, _02396_, _01481_);
  and _25440_ (_02398_, _07015_, _06981_);
  or _25441_ (_02399_, _02398_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or _25442_ (_02400_, _02399_, _06678_);
  and _25443_ (_02401_, _02400_, _02397_);
  or _25444_ (_02402_, _02401_, _06946_);
  nand _25445_ (_02403_, _10494_, _06946_);
  and _25446_ (_02404_, _02403_, _06444_);
  and _25447_ (_03597_, _02404_, _02402_);
  and _25448_ (_02405_, _07147_, _06440_);
  and _25449_ (_02406_, _02405_, _06941_);
  and _25450_ (_02407_, _06987_, _06678_);
  nand _25451_ (_02408_, _02407_, _06930_);
  or _25452_ (_02409_, _02407_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and _25453_ (_02410_, _02409_, _02408_);
  or _25454_ (_02411_, _02410_, _02406_);
  nand _25455_ (_02412_, _06946_, _06666_);
  and _25456_ (_02413_, _02412_, _06444_);
  and _25457_ (_03599_, _02413_, _02411_);
  and _25458_ (_02414_, _06983_, _06678_);
  nand _25459_ (_02415_, _02414_, _06930_);
  not _25460_ (_02416_, _06946_);
  or _25461_ (_02417_, _02414_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and _25462_ (_02418_, _02417_, _02416_);
  and _25463_ (_02419_, _02418_, _02415_);
  nor _25464_ (_02420_, _07188_, _02416_);
  or _25465_ (_02421_, _02420_, _02419_);
  and _25466_ (_03606_, _02421_, _06444_);
  and _25467_ (_02422_, _10976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor _25468_ (_02423_, _10956_, _10920_);
  nor _25469_ (_02424_, _02423_, _10957_);
  or _25470_ (_02425_, _02424_, _08374_);
  or _25471_ (_02426_, _08373_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and _25472_ (_02427_, _02426_, _10894_);
  and _25473_ (_02428_, _02427_, _02425_);
  or _25474_ (_03621_, _02428_, _02422_);
  nor _25475_ (_03623_, _11402_, rst);
  nand _25476_ (_02429_, _02332_, _11418_);
  or _25477_ (_03625_, _02429_, _02298_);
  and _25478_ (_02430_, _10839_, _10751_);
  and _25479_ (_02431_, _02430_, _10836_);
  and _25480_ (_02432_, _10850_, _10746_);
  and _25481_ (_02433_, _10874_, _10836_);
  or _25482_ (_02434_, _02433_, _02432_);
  or _25483_ (_02435_, _02434_, _02431_);
  nor _25484_ (_02436_, _10884_, _10848_);
  nand _25485_ (_02437_, _02436_, _10786_);
  or _25486_ (_02438_, _02437_, _02435_);
  nand _25487_ (_02439_, _10822_, _10776_);
  or _25488_ (_02440_, _02439_, _02438_);
  and _25489_ (_02441_, _10820_, _10753_);
  and _25490_ (_02442_, _10743_, _08425_);
  and _25491_ (_02443_, _10739_, _08457_);
  and _25492_ (_02444_, _10770_, _02443_);
  or _25493_ (_02445_, _02444_, _02442_);
  or _25494_ (_02446_, _02445_, _02441_);
  or _25495_ (_02447_, _10831_, _10826_);
  and _25496_ (_02448_, _10799_, _10753_);
  and _25497_ (_02449_, _02448_, _10812_);
  and _25498_ (_02450_, _10736_, _10812_);
  and _25499_ (_02451_, _10782_, _02450_);
  and _25500_ (_02452_, _10736_, _10741_);
  and _25501_ (_02453_, _10850_, _02452_);
  or _25502_ (_02454_, _02453_, _02451_);
  or _25503_ (_02455_, _02454_, _02449_);
  or _25504_ (_02456_, _02455_, _02447_);
  or _25505_ (_02457_, _02456_, _02446_);
  or _25506_ (_02458_, _02457_, _02440_);
  and _25507_ (_02459_, _02458_, _07231_);
  and _25508_ (_02460_, _07228_, _06308_);
  and _25509_ (_02461_, _02460_, _11386_);
  nor _25510_ (_02462_, _02461_, _02295_);
  or _25511_ (_02463_, _02462_, rst);
  or _25512_ (_03627_, _02463_, _02459_);
  not _25513_ (_02464_, _07229_);
  or _25514_ (_02465_, _08360_, _02464_);
  or _25515_ (_02466_, _07229_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and _25516_ (_02467_, _02466_, _06444_);
  and _25517_ (_03630_, _02467_, _02465_);
  and _25518_ (_02468_, _02306_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and _25519_ (_02469_, _11490_, _11355_);
  or _25520_ (_02470_, _02469_, _11986_);
  and _25521_ (_02471_, _11419_, _11394_);
  and _25522_ (_02472_, _11493_, _11354_);
  or _25523_ (_02473_, _02472_, _02471_);
  or _25524_ (_02474_, _02473_, _02470_);
  or _25525_ (_02475_, _11491_, _12040_);
  or _25526_ (_02476_, _02475_, _02325_);
  nor _25527_ (_02477_, _02476_, _02474_);
  nand _25528_ (_02478_, _02477_, _11461_);
  and _25529_ (_02479_, _02478_, _02332_);
  or _25530_ (_03632_, _02479_, _02468_);
  or _25531_ (_02480_, _02248_, _11379_);
  and _25532_ (_02481_, _11519_, _11412_);
  or _25533_ (_02482_, _02481_, _11442_);
  and _25534_ (_02483_, _11490_, _11965_);
  or _25535_ (_02484_, _02483_, _02482_);
  or _25536_ (_02485_, _02484_, _02480_);
  and _25537_ (_02486_, _02485_, _07230_);
  and _25538_ (_02487_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _25539_ (_02488_, _02487_, _02353_);
  or _25540_ (_02489_, _02488_, _02486_);
  and _25541_ (_03634_, _02489_, _06444_);
  and _25542_ (_02490_, _02306_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and _25543_ (_02491_, _11443_, _11394_);
  not _25544_ (_02492_, _11429_);
  and _25545_ (_02493_, _11427_, _11526_);
  or _25546_ (_02494_, _02493_, _14239_);
  or _25547_ (_02495_, _02494_, _02492_);
  or _25548_ (_02496_, _02495_, _02491_);
  and _25549_ (_02497_, _11965_, _11458_);
  or _25550_ (_02498_, _02361_, _02253_);
  or _25551_ (_02499_, _02498_, _02497_);
  or _25552_ (_02500_, _02480_, _02309_);
  or _25553_ (_02501_, _02500_, _02499_);
  or _25554_ (_02502_, _02501_, _02496_);
  and _25555_ (_02503_, _02502_, _02332_);
  or _25556_ (_03637_, _02503_, _02490_);
  and _25557_ (_02504_, _12012_, _06987_);
  nand _25558_ (_02505_, _02504_, _06930_);
  or _25559_ (_02506_, _02504_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and _25560_ (_02507_, _02506_, _07219_);
  and _25561_ (_02508_, _02507_, _02505_);
  nor _25562_ (_02509_, _07219_, _06666_);
  or _25563_ (_02510_, _02509_, _02508_);
  and _25564_ (_03640_, _02510_, _06444_);
  and _25565_ (_02511_, _07029_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and _25566_ (_02512_, _02511_, _07026_);
  and _25567_ (_02513_, _07011_, _06994_);
  or _25568_ (_02514_, _02513_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  nand _25569_ (_02515_, _07011_, _06995_);
  and _25570_ (_02516_, _02515_, _02514_);
  or _25571_ (_02517_, _02516_, _02512_);
  and _25572_ (_02518_, _02517_, _07035_);
  and _25573_ (_02519_, _07017_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  or _25574_ (_02520_, _02519_, _06985_);
  or _25575_ (_02521_, _02520_, _02518_);
  nand _25576_ (_02522_, _07188_, _06985_);
  and _25577_ (_02523_, _02522_, _09503_);
  and _25578_ (_02524_, _02523_, _02521_);
  and _25579_ (_02525_, _06989_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or _25580_ (_02526_, _02525_, _02524_);
  and _25581_ (_03644_, _02526_, _06444_);
  and _25582_ (_02527_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and _25583_ (_02528_, _11534_, _07230_);
  or _25584_ (_02529_, _02528_, _02527_);
  or _25585_ (_02530_, _02529_, _02353_);
  and _25586_ (_03646_, _02530_, _06444_);
  or _25587_ (_02531_, _02356_, _02325_);
  and _25588_ (_02532_, _02531_, _11342_);
  or _25589_ (_02533_, _02303_, \oc8051_top_1.oc8051_sfr1.wait_data );
  or _25590_ (_02534_, _02533_, _02357_);
  or _25591_ (_02535_, _02534_, _02532_);
  or _25592_ (_02536_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2], _06308_);
  and _25593_ (_02537_, _02536_, _06444_);
  and _25594_ (_03648_, _02537_, _02535_);
  not _25595_ (_02538_, _06985_);
  and _25596_ (_02539_, _07017_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and _25597_ (_02540_, _07011_, _06993_);
  nor _25598_ (_02541_, _02540_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  nor _25599_ (_02542_, _02541_, _02513_);
  and _25600_ (_02543_, _07029_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and _25601_ (_02544_, _02543_, _07026_);
  or _25602_ (_02545_, _02544_, _02542_);
  and _25603_ (_02546_, _02545_, _07035_);
  or _25604_ (_02547_, _02546_, _02539_);
  and _25605_ (_02548_, _02547_, _02538_);
  nor _25606_ (_02549_, _07300_, _02538_);
  or _25607_ (_02550_, _02549_, _06989_);
  or _25608_ (_02551_, _02550_, _02548_);
  or _25609_ (_02552_, _09503_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and _25610_ (_02553_, _02552_, _06444_);
  and _25611_ (_03651_, _02553_, _02551_);
  and _25612_ (_02554_, _02306_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  or _25613_ (_02555_, _11412_, _11427_);
  and _25614_ (_02556_, _02555_, _11976_);
  or _25615_ (_02557_, _11379_, _11494_);
  or _25616_ (_02558_, _02557_, _02556_);
  or _25617_ (_02559_, _02481_, _11504_);
  or _25618_ (_02561_, _11533_, _11489_);
  or _25619_ (_02562_, _02561_, _02559_);
  or _25620_ (_02563_, _02472_, _02497_);
  and _25621_ (_02564_, _11490_, _11406_);
  and _25622_ (_02565_, _11406_, _11458_);
  or _25623_ (_02567_, _02565_, _02564_);
  or _25624_ (_02568_, _02567_, _02563_);
  or _25625_ (_02569_, _02568_, _02562_);
  or _25626_ (_02570_, _02569_, _02558_);
  and _25627_ (_02571_, _02570_, _02332_);
  or _25628_ (_03653_, _02571_, _02554_);
  and _25629_ (_02572_, _02306_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  not _25630_ (_02573_, _11478_);
  or _25631_ (_02574_, _02249_, _02573_);
  or _25632_ (_02575_, _02311_, _02260_);
  or _25633_ (_02576_, _02575_, _02494_);
  nor _25634_ (_02577_, _02576_, _02574_);
  and _25635_ (_02578_, _02577_, _11488_);
  or _25636_ (_02579_, _02483_, _02263_);
  nor _25637_ (_02580_, _02579_, _02324_);
  nand _25638_ (_02581_, _02580_, _11484_);
  nor _25639_ (_02582_, _02581_, _02499_);
  and _25640_ (_02584_, _02582_, _14230_);
  nand _25641_ (_02585_, _02584_, _02578_);
  and _25642_ (_02586_, _02585_, _02332_);
  or _25643_ (_03656_, _02586_, _02572_);
  or _25644_ (_02587_, _02275_, _02268_);
  or _25645_ (_02588_, _02280_, _02277_);
  or _25646_ (_02589_, _02588_, _02587_);
  or _25647_ (_02590_, _02264_, _02352_);
  or _25648_ (_02591_, _02590_, _02589_);
  and _25649_ (_02592_, _02591_, _02332_);
  nor _25650_ (_02593_, _11399_, _11342_);
  and _25651_ (_02594_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _25652_ (_02595_, _02594_, _02593_);
  and _25653_ (_02596_, _02595_, _06444_);
  or _25654_ (_03658_, _02596_, _02592_);
  and _25655_ (_02597_, _11976_, _11417_);
  or _25656_ (_02598_, _02597_, _02355_);
  and _25657_ (_02599_, _11519_, _11369_);
  or _25658_ (_02600_, _02599_, _02482_);
  or _25659_ (_02601_, _02600_, _02598_);
  or _25660_ (_02602_, _02601_, _02376_);
  or _25661_ (_02603_, _02494_, _02386_);
  or _25662_ (_02604_, _02603_, _02602_);
  or _25663_ (_02605_, _02604_, _02374_);
  and _25664_ (_02606_, _02605_, _07230_);
  and _25665_ (_02607_, \oc8051_top_1.oc8051_decoder1.wr , \oc8051_top_1.oc8051_sfr1.wait_data );
  or _25666_ (_02608_, _02607_, _02359_);
  or _25667_ (_02609_, _02608_, _02606_);
  and _25668_ (_03660_, _02609_, _06444_);
  and _25669_ (_02610_, _07017_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and _25670_ (_02611_, _07011_, _06992_);
  nor _25671_ (_02612_, _02611_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  nor _25672_ (_02613_, _02612_, _02540_);
  and _25673_ (_02614_, _07029_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and _25674_ (_02615_, _02614_, _07026_);
  or _25675_ (_02616_, _02615_, _02613_);
  and _25676_ (_02617_, _02616_, _07035_);
  or _25677_ (_02618_, _02617_, _02610_);
  and _25678_ (_02619_, _02618_, _02538_);
  nor _25679_ (_02620_, _11589_, _02538_);
  or _25680_ (_02621_, _02620_, _06989_);
  or _25681_ (_02622_, _02621_, _02619_);
  or _25682_ (_02623_, _09503_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and _25683_ (_02624_, _02623_, _06444_);
  and _25684_ (_03663_, _02624_, _02622_);
  and _25685_ (_02625_, _07011_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  nor _25686_ (_02626_, _02625_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  nor _25687_ (_02627_, _02626_, _02611_);
  and _25688_ (_02628_, _07029_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and _25689_ (_02629_, _02628_, _07026_);
  or _25690_ (_02630_, _02629_, _02627_);
  and _25691_ (_02631_, _02630_, _07035_);
  and _25692_ (_02633_, _07017_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  or _25693_ (_02634_, _02633_, _06985_);
  or _25694_ (_02635_, _02634_, _02631_);
  nand _25695_ (_02636_, _07069_, _06985_);
  and _25696_ (_02637_, _02636_, _09503_);
  and _25697_ (_02638_, _02637_, _02635_);
  and _25698_ (_02639_, _06989_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  or _25699_ (_02640_, _02639_, _02638_);
  and _25700_ (_03667_, _02640_, _06444_);
  and _25701_ (_02641_, _10976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor _25702_ (_02642_, _10955_, _10925_);
  nor _25703_ (_02643_, _02642_, _10956_);
  or _25704_ (_02644_, _02643_, _08374_);
  or _25705_ (_02646_, _08373_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and _25706_ (_02647_, _02646_, _10894_);
  and _25707_ (_02648_, _02647_, _02644_);
  or _25708_ (_03669_, _02648_, _02641_);
  nand _25709_ (_02650_, _01085_, _07216_);
  or _25710_ (_02651_, _02650_, _08230_);
  not _25711_ (_02653_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nand _25712_ (_02654_, _02650_, _02653_);
  and _25713_ (_02655_, _02654_, _06440_);
  and _25714_ (_02656_, _02655_, _02651_);
  nor _25715_ (_02657_, _06673_, _02653_);
  and _25716_ (_02659_, _00604_, _07963_);
  and _25717_ (_02660_, _02659_, _06983_);
  nand _25718_ (_02662_, _02660_, _06930_);
  or _25719_ (_02663_, _02660_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and _25720_ (_02665_, _02663_, _06674_);
  and _25721_ (_02667_, _02665_, _02662_);
  or _25722_ (_02668_, _02667_, _02657_);
  or _25723_ (_02669_, _02668_, _02656_);
  and _25724_ (_03678_, _02669_, _06444_);
  and _25725_ (_02671_, _07029_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  nand _25726_ (_02672_, _02671_, _07006_);
  nand _25727_ (_02674_, _02672_, _02625_);
  or _25728_ (_02675_, _07011_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and _25729_ (_02677_, _02675_, _07035_);
  and _25730_ (_02678_, _02677_, _02674_);
  and _25731_ (_02680_, _07017_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  or _25732_ (_02681_, _02680_, _06985_);
  or _25733_ (_02682_, _02681_, _02678_);
  nand _25734_ (_02683_, _09526_, _06985_);
  and _25735_ (_02684_, _02683_, _09503_);
  and _25736_ (_02685_, _02684_, _02682_);
  and _25737_ (_02686_, _06989_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  or _25738_ (_02687_, _02686_, _02685_);
  and _25739_ (_03685_, _02687_, _06444_);
  not _25740_ (_02688_, _02332_);
  or _25741_ (_03688_, _02688_, _02301_);
  or _25742_ (_02689_, _07432_, \oc8051_top_1.oc8051_rom1.data_o [7]);
  nand _25743_ (_02690_, _07432_, _13886_);
  and _25744_ (_02691_, _02690_, _06444_);
  and _25745_ (_03692_, _02691_, _02689_);
  or _25746_ (_02692_, _07432_, \oc8051_top_1.oc8051_rom1.data_o [6]);
  nand _25747_ (_02693_, _07432_, _13896_);
  and _25748_ (_02694_, _02693_, _06444_);
  and _25749_ (_03700_, _02694_, _02692_);
  or _25750_ (_02695_, _02650_, _08019_);
  not _25751_ (_02696_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nand _25752_ (_02697_, _02650_, _02696_);
  and _25753_ (_02698_, _02697_, _06440_);
  and _25754_ (_02699_, _02698_, _02695_);
  nor _25755_ (_02700_, _06673_, _02696_);
  or _25756_ (_02701_, _02650_, _08232_);
  and _25757_ (_02702_, _02697_, _06674_);
  and _25758_ (_02703_, _02702_, _02701_);
  or _25759_ (_02704_, _02703_, _02700_);
  or _25760_ (_02705_, _02704_, _02699_);
  and _25761_ (_03705_, _02705_, _06444_);
  or _25762_ (_02706_, _02650_, _08127_);
  not _25763_ (_02707_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nand _25764_ (_02708_, _02650_, _02707_);
  and _25765_ (_02709_, _02708_, _06440_);
  and _25766_ (_02710_, _02709_, _02706_);
  nor _25767_ (_02711_, _06673_, _02707_);
  and _25768_ (_02712_, _02659_, _06987_);
  nand _25769_ (_02713_, _02712_, _06930_);
  or _25770_ (_02714_, _02712_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and _25771_ (_02715_, _02714_, _06674_);
  and _25772_ (_02716_, _02715_, _02713_);
  or _25773_ (_02717_, _02716_, _02711_);
  or _25774_ (_02718_, _02717_, _02710_);
  and _25775_ (_03708_, _02718_, _06444_);
  and _25776_ (_02719_, _11418_, _11347_);
  and _25777_ (_02720_, _02719_, _11394_);
  or _25778_ (_02721_, _02720_, _02257_);
  or _25779_ (_02722_, _02471_, _11966_);
  or _25780_ (_02723_, _02722_, _11396_);
  or _25781_ (_02724_, _02723_, _02721_);
  or _25782_ (_02725_, _02249_, _02283_);
  or _25783_ (_02726_, _02598_, _02384_);
  or _25784_ (_02727_, _02726_, _02725_);
  and _25785_ (_02728_, _02263_, _07311_);
  or _25786_ (_02729_, _02728_, _02354_);
  or _25787_ (_02730_, _02729_, _02727_);
  or _25788_ (_02731_, _14225_, _11398_);
  and _25789_ (_02732_, _11456_, _11965_);
  or _25790_ (_02733_, _02297_, _02732_);
  or _25791_ (_02734_, _02733_, _02731_);
  and _25792_ (_02735_, _02367_, _11418_);
  and _25793_ (_02736_, _11437_, _11430_);
  and _25794_ (_02737_, _02275_, _11376_);
  or _25795_ (_02738_, _02737_, _02736_);
  or _25796_ (_02739_, _02738_, _02735_);
  or _25797_ (_02740_, _02739_, _02734_);
  or _25798_ (_02741_, _02740_, _02730_);
  or _25799_ (_02742_, _02279_, _02260_);
  or _25800_ (_02743_, _02742_, _11440_);
  or _25801_ (_02744_, _02743_, _02278_);
  and _25802_ (_02745_, _02483_, _07311_);
  or _25803_ (_02746_, _02264_, _11444_);
  or _25804_ (_02747_, _02746_, _11375_);
  or _25805_ (_02748_, _02747_, _02745_);
  or _25806_ (_02749_, _02748_, _02744_);
  or _25807_ (_02750_, _02749_, _02741_);
  or _25808_ (_02751_, _02750_, _02724_);
  and _25809_ (_02752_, _02751_, _07230_);
  and _25810_ (_02753_, \oc8051_top_1.oc8051_sfr1.wait_data , \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  or _25811_ (_02754_, _02593_, _02303_);
  or _25812_ (_02755_, _02754_, _02753_);
  or _25813_ (_02756_, _02755_, _02752_);
  and _25814_ (_03710_, _02756_, _06444_);
  or _25815_ (_02757_, _10954_, _10929_);
  nor _25816_ (_02758_, _10955_, _08374_);
  and _25817_ (_02759_, _02758_, _02757_);
  and _25818_ (_02760_, _08374_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  or _25819_ (_02761_, _02760_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _25820_ (_02762_, _02761_, _02759_);
  or _25821_ (_02764_, _02166_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and _25822_ (_02765_, _02764_, _06444_);
  and _25823_ (_03712_, _02765_, _02762_);
  and _25824_ (_02766_, _11418_, _11385_);
  nor _25825_ (_02767_, _02766_, _02297_);
  or _25826_ (_03715_, _02767_, _02688_);
  or _25827_ (_02768_, _02448_, \oc8051_top_1.oc8051_decoder1.state [1]);
  or _25828_ (_02769_, _02768_, _02454_);
  and _25829_ (_02770_, _02769_, _02461_);
  nor _25830_ (_02771_, _02460_, _11386_);
  or _25831_ (_02772_, _02771_, rst);
  or _25832_ (_03718_, _02772_, _02770_);
  and _25833_ (_02773_, _10976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nor _25834_ (_02774_, _01553_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and _25835_ (_02775_, _01553_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nor _25836_ (_02776_, _02775_, _02774_);
  not _25837_ (_02777_, _02776_);
  nor _25838_ (_02778_, _02777_, _01564_);
  and _25839_ (_02779_, _02777_, _01564_);
  or _25840_ (_02780_, _02779_, _02778_);
  or _25841_ (_02781_, _02780_, _08374_);
  or _25842_ (_02782_, _08373_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and _25843_ (_02783_, _02782_, _10894_);
  and _25844_ (_02784_, _02783_, _02781_);
  or _25845_ (_03720_, _02784_, _02773_);
  and _25846_ (_02785_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8], \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and _25847_ (_02786_, _12225_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and _25848_ (_02787_, _02786_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and _25849_ (_02788_, _02787_, _02785_);
  and _25850_ (_02789_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11], \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nand _25851_ (_02790_, _02789_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor _25852_ (_02791_, _02790_, _07432_);
  and _25853_ (_02792_, _02791_, _02788_);
  and _25854_ (_02793_, _02792_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and _25855_ (_02794_, _02793_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nand _25856_ (_02795_, _02794_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  or _25857_ (_02796_, _02794_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and _25858_ (_02797_, _02796_, _02795_);
  or _25859_ (_02798_, _02797_, _12023_);
  and _25860_ (_02799_, _02798_, _06444_);
  and _25861_ (_02800_, _11452_, _11137_);
  and _25862_ (_02801_, _12026_, _11177_);
  and _25863_ (_02802_, _12032_, _11625_);
  and _25864_ (_02803_, _12047_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  or _25865_ (_02804_, _02803_, _02802_);
  or _25866_ (_02805_, _02804_, _02801_);
  or _25867_ (_02806_, _02805_, _02800_);
  or _25868_ (_02807_, \oc8051_top_1.oc8051_memory_interface1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  or _25869_ (_02808_, _02807_, _12660_);
  or _25870_ (_02809_, _02808_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand _25871_ (_02810_, _02809_, _12650_);
  or _25872_ (_02811_, _12666_, _08150_);
  or _25873_ (_02812_, _02811_, _08155_);
  or _25874_ (_02813_, _02812_, _09186_);
  nand _25875_ (_02814_, _02813_, _12662_);
  nand _25876_ (_02815_, _02814_, _02810_);
  nand _25877_ (_02816_, _02815_, _11165_);
  or _25878_ (_02817_, _02815_, _11165_);
  and _25879_ (_02818_, _02817_, _12218_);
  and _25880_ (_02819_, _02818_, _02816_);
  or _25881_ (_02820_, _02819_, _02806_);
  and _25882_ (_02821_, _12683_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and _25883_ (_02822_, _02821_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor _25884_ (_02823_, _02822_, _11165_);
  and _25885_ (_02824_, _02822_, _11165_);
  or _25886_ (_02825_, _02824_, _02823_);
  nand _25887_ (_02826_, _02825_, _12054_);
  nand _25888_ (_02827_, _02826_, _12023_);
  or _25889_ (_02828_, _02827_, _02820_);
  and _25890_ (_03733_, _02828_, _02799_);
  or _25891_ (_02829_, _02650_, _12024_);
  not _25892_ (_02830_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  nand _25893_ (_02831_, _02650_, _02830_);
  and _25894_ (_02832_, _02831_, _06440_);
  and _25895_ (_02833_, _02832_, _02829_);
  nor _25896_ (_02834_, _06673_, _02830_);
  and _25897_ (_02835_, _02659_, _00240_);
  nand _25898_ (_02836_, _02835_, _06930_);
  or _25899_ (_02837_, _02835_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and _25900_ (_02838_, _02837_, _06674_);
  and _25901_ (_02839_, _02838_, _02836_);
  or _25902_ (_02840_, _02839_, _02834_);
  or _25903_ (_02841_, _02840_, _02833_);
  and _25904_ (_03737_, _02841_, _06444_);
  and _25905_ (_02842_, _11418_, _11976_);
  or _25906_ (_02843_, _02842_, _11513_);
  or _25907_ (_02844_, _02843_, _11517_);
  and _25908_ (_02845_, _02384_, _11410_);
  or _25909_ (_02846_, _02845_, _11371_);
  or _25910_ (_02847_, _02846_, _02844_);
  and _25911_ (_02848_, _02364_, _07268_);
  or _25912_ (_02849_, _02248_, _11398_);
  or _25913_ (_02850_, _02849_, _02368_);
  or _25914_ (_02851_, _02850_, _02848_);
  or _25915_ (_02852_, _02851_, _02847_);
  or _25916_ (_02853_, _02852_, _02749_);
  or _25917_ (_02854_, _02853_, _02724_);
  and _25918_ (_02855_, _02854_, _07230_);
  and _25919_ (_02856_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _25920_ (_02857_, _02856_, _02754_);
  or _25921_ (_02858_, _02857_, _02855_);
  and _25922_ (_03743_, _02858_, _06444_);
  nor _25923_ (_03747_, _12073_, rst);
  and _25924_ (_03752_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _06444_);
  nand _25925_ (_02859_, _10494_, _09479_);
  not _25926_ (_02860_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  nor _25927_ (_02861_, _09485_, _02860_);
  and _25928_ (_02862_, _09485_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or _25929_ (_02863_, _02862_, _02861_);
  or _25930_ (_02864_, _02863_, _09479_);
  and _25931_ (_02865_, _02864_, _06444_);
  and _25932_ (_03756_, _02865_, _02859_);
  nor _25933_ (_03758_, _11547_, rst);
  nand _25934_ (_02866_, _10112_, _09526_);
  or _25935_ (_02867_, _10112_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  and _25936_ (_02868_, _02867_, _02866_);
  and _25937_ (_03765_, _02868_, _06444_);
  and _25938_ (_02869_, _12012_, _06983_);
  nand _25939_ (_02870_, _02869_, _06930_);
  or _25940_ (_02871_, _02869_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and _25941_ (_02872_, _02871_, _07219_);
  and _25942_ (_02873_, _02872_, _02870_);
  or _25943_ (_02874_, _02873_, _07221_);
  and _25944_ (_03784_, _02874_, _06444_);
  or _25945_ (_02875_, _09485_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  or _25946_ (_02876_, _09486_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and _25947_ (_02877_, _02876_, _02875_);
  or _25948_ (_02878_, _02877_, _09479_);
  nand _25949_ (_02880_, _09479_, _07069_);
  and _25950_ (_02882_, _02880_, _06444_);
  and _25951_ (_03787_, _02882_, _02878_);
  nand _25952_ (_02884_, _09479_, _06666_);
  or _25953_ (_02885_, _09485_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  not _25954_ (_02887_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  nand _25955_ (_02889_, _09485_, _02887_);
  and _25956_ (_02891_, _02889_, _02885_);
  or _25957_ (_02892_, _02891_, _09479_);
  and _25958_ (_02894_, _02892_, _06444_);
  and _25959_ (_03791_, _02894_, _02884_);
  nor _25960_ (_03794_, _11470_, rst);
  nand _25961_ (_02895_, _09479_, _07188_);
  and _25962_ (_02896_, _09485_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and _25963_ (_02897_, _09486_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  or _25964_ (_02899_, _02897_, _02896_);
  or _25965_ (_02900_, _02899_, _09479_);
  and _25966_ (_02901_, _02900_, _06444_);
  and _25967_ (_03797_, _02901_, _02895_);
  and _25968_ (_02902_, _09485_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  not _25969_ (_02903_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  nor _25970_ (_02904_, _09485_, _02903_);
  or _25971_ (_02906_, _02904_, _02902_);
  or _25972_ (_02907_, _02906_, _09479_);
  nand _25973_ (_02909_, _09479_, _07300_);
  and _25974_ (_02910_, _02909_, _06444_);
  and _25975_ (_03800_, _02910_, _02907_);
  nor _25976_ (_03802_, _12106_, rst);
  or _25977_ (_02911_, _02650_, _07959_);
  not _25978_ (_02912_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  nand _25979_ (_02913_, _02650_, _02912_);
  and _25980_ (_02915_, _02913_, _06440_);
  and _25981_ (_02917_, _02915_, _02911_);
  nor _25982_ (_02918_, _06673_, _02912_);
  and _25983_ (_02920_, _02659_, _06432_);
  nand _25984_ (_02922_, _02920_, _06930_);
  or _25985_ (_02923_, _02920_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and _25986_ (_02925_, _02923_, _06674_);
  and _25987_ (_02927_, _02925_, _02922_);
  or _25988_ (_02928_, _02927_, _02918_);
  or _25989_ (_02929_, _02928_, _02917_);
  and _25990_ (_03804_, _02929_, _06444_);
  or _25991_ (_02930_, _02650_, _08308_);
  not _25992_ (_02931_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nand _25993_ (_02932_, _02650_, _02931_);
  and _25994_ (_02933_, _02932_, _06440_);
  and _25995_ (_02934_, _02933_, _02930_);
  nor _25996_ (_02935_, _06673_, _02931_);
  and _25997_ (_02936_, _02659_, _08310_);
  nand _25998_ (_02937_, _02936_, _06930_);
  or _25999_ (_02938_, _02936_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and _26000_ (_02939_, _02938_, _06674_);
  and _26001_ (_02940_, _02939_, _02937_);
  or _26002_ (_02941_, _02940_, _02935_);
  or _26003_ (_02942_, _02941_, _02934_);
  and _26004_ (_03807_, _02942_, _06444_);
  nor _26005_ (_03812_, _12128_, rst);
  and _26006_ (_02943_, _02306_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  or _26007_ (_02944_, _11479_, _11476_);
  or _26008_ (_02946_, _11512_, _11487_);
  or _26009_ (_02947_, _02946_, _02944_);
  or _26010_ (_02948_, _02947_, _02558_);
  and _26011_ (_02949_, _02555_, _11356_);
  or _26012_ (_02950_, _11456_, _11486_);
  and _26013_ (_02951_, _02950_, _11355_);
  or _26014_ (_02952_, _02951_, _02949_);
  or _26015_ (_02953_, _02481_, _02264_);
  or _26016_ (_02954_, _02953_, _02279_);
  or _26017_ (_02955_, _02954_, _02952_);
  or _26018_ (_02956_, _02955_, _02948_);
  and _26019_ (_02957_, _02497_, _07311_);
  or _26020_ (_02958_, _02957_, _02254_);
  or _26021_ (_02959_, _02958_, _11495_);
  or _26022_ (_02960_, _02564_, _02732_);
  and _26023_ (_02961_, _11456_, _11526_);
  and _26024_ (_02962_, _11423_, _11426_);
  or _26025_ (_02963_, _02962_, _02961_);
  or _26026_ (_02964_, _02963_, _02960_);
  or _26027_ (_02965_, _11504_, _11444_);
  or _26028_ (_02966_, _02965_, _11509_);
  or _26029_ (_02967_, _02966_, _02964_);
  or _26030_ (_02968_, _02967_, _02959_);
  or _26031_ (_02969_, _02968_, _02956_);
  and _26032_ (_02970_, _02969_, _02332_);
  or _26033_ (_03816_, _02970_, _02943_);
  and _26034_ (_02971_, _09485_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and _26035_ (_02972_, _09486_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  or _26036_ (_02973_, _02972_, _02971_);
  or _26037_ (_02974_, _02973_, _09479_);
  nand _26038_ (_02975_, _11589_, _09479_);
  and _26039_ (_02976_, _02975_, _06444_);
  and _26040_ (_03821_, _02976_, _02974_);
  not _26041_ (_02977_, _09138_);
  or _26042_ (_02978_, _02650_, _02977_);
  not _26043_ (_02979_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  nand _26044_ (_02980_, _02650_, _02979_);
  and _26045_ (_02981_, _02980_, _06440_);
  and _26046_ (_02982_, _02981_, _02978_);
  nor _26047_ (_02983_, _06673_, _02979_);
  not _26048_ (_02984_, _02659_);
  or _26049_ (_02985_, _02984_, _00717_);
  and _26050_ (_02986_, _02985_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and _26051_ (_02987_, _06431_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or _26052_ (_02988_, _02987_, _00713_);
  and _26053_ (_02989_, _02988_, _02659_);
  or _26054_ (_02990_, _02989_, _02986_);
  and _26055_ (_02991_, _02990_, _06674_);
  or _26056_ (_02992_, _02991_, _02983_);
  or _26057_ (_02993_, _02992_, _02982_);
  and _26058_ (_03824_, _02993_, _06444_);
  and _26059_ (_02994_, _12012_, _08310_);
  or _26060_ (_02995_, _02994_, _07278_);
  nand _26061_ (_02996_, _02994_, _06930_);
  and _26062_ (_02997_, _02996_, _02995_);
  or _26063_ (_02998_, _02997_, _07301_);
  and _26064_ (_03828_, _02998_, _06444_);
  or _26065_ (_02999_, _07263_, _02464_);
  or _26066_ (_03000_, _07229_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and _26067_ (_03001_, _03000_, _06444_);
  and _26068_ (_03831_, _03001_, _02999_);
  or _26069_ (_03002_, _08392_, _02464_);
  or _26070_ (_03003_, _07229_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and _26071_ (_03004_, _03003_, _06444_);
  and _26072_ (_03833_, _03004_, _03002_);
  nand _26073_ (_03005_, _08408_, _07229_);
  or _26074_ (_03006_, _07229_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and _26075_ (_03007_, _03006_, _06444_);
  and _26076_ (_03835_, _03007_, _03005_);
  or _26077_ (_03008_, _08425_, _02464_);
  or _26078_ (_03009_, _07229_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and _26079_ (_03010_, _03009_, _06444_);
  and _26080_ (_03837_, _03010_, _03008_);
  or _26081_ (_03011_, _08441_, _02464_);
  or _26082_ (_03012_, _07229_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and _26083_ (_03013_, _03012_, _06444_);
  and _26084_ (_03839_, _03013_, _03011_);
  or _26085_ (_03014_, _08457_, _02464_);
  or _26086_ (_03015_, _07229_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and _26087_ (_03016_, _03015_, _06444_);
  and _26088_ (_03840_, _03016_, _03014_);
  nor _26089_ (_03017_, _10953_, _10948_);
  nor _26090_ (_03018_, _03017_, _10954_);
  or _26091_ (_03019_, _03018_, _08374_);
  or _26092_ (_03020_, _08373_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _26093_ (_03021_, _03020_, _10894_);
  and _26094_ (_03022_, _03021_, _03019_);
  and _26095_ (_03023_, _10976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or _26096_ (_03842_, _03023_, _03022_);
  nand _26097_ (_03024_, _08472_, _07229_);
  or _26098_ (_03025_, _07229_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and _26099_ (_03026_, _03025_, _06444_);
  and _26100_ (_03851_, _03026_, _03024_);
  or _26101_ (_03027_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or _26102_ (_03028_, _07987_, _07927_);
  or _26103_ (_03029_, _03028_, _09095_);
  or _26104_ (_03030_, _03029_, _08284_);
  or _26105_ (_03031_, _03030_, _08097_);
  or _26106_ (_03032_, _03031_, _08996_);
  and _26107_ (_03033_, _03032_, _07602_);
  or _26108_ (_03034_, _06844_, _06842_);
  not _26109_ (_03035_, _06706_);
  nand _26110_ (_03037_, _06842_, _03035_);
  and _26111_ (_03038_, _03037_, _06680_);
  and _26112_ (_03039_, _03038_, _03034_);
  not _26113_ (_03041_, _06707_);
  nand _26114_ (_03043_, _06877_, _03041_);
  nor _26115_ (_03045_, _06878_, _06848_);
  and _26116_ (_03047_, _03045_, _03043_);
  and _26117_ (_03048_, _06752_, _06482_);
  and _26118_ (_03050_, _03048_, _07578_);
  and _26119_ (_03051_, _03050_, _08167_);
  nand _26120_ (_03052_, _03051_, _07459_);
  nand _26121_ (_03053_, _03052_, \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or _26122_ (_03054_, _03053_, _03047_);
  or _26123_ (_03055_, _03054_, _03039_);
  nor _26124_ (_03056_, _03055_, _08206_);
  nand _26125_ (_03057_, _03056_, _11108_);
  or _26126_ (_03058_, _03057_, _03033_);
  and _26127_ (_03059_, _03058_, _03027_);
  or _26128_ (_03060_, _03059_, _12012_);
  and _26129_ (_03062_, _00712_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or _26130_ (_03063_, _03062_, _00713_);
  or _26131_ (_03064_, _03063_, _12013_);
  and _26132_ (_03065_, _03064_, _03060_);
  or _26133_ (_03066_, _03065_, _07218_);
  nand _26134_ (_03067_, _11589_, _07218_);
  and _26135_ (_03068_, _03067_, _06444_);
  and _26136_ (_03860_, _03068_, _03066_);
  or _26137_ (_03069_, _09485_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  or _26138_ (_03071_, _09486_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and _26139_ (_03073_, _03071_, _03069_);
  or _26140_ (_03075_, _03073_, _09479_);
  nand _26141_ (_03077_, _09526_, _09479_);
  and _26142_ (_03079_, _03077_, _06444_);
  and _26143_ (_03864_, _03079_, _03075_);
  and _26144_ (_03082_, _12012_, _06432_);
  nand _26145_ (_03083_, _03082_, _06930_);
  or _26146_ (_03085_, _03082_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and _26147_ (_03087_, _03085_, _07219_);
  and _26148_ (_03089_, _03087_, _03083_);
  nor _26149_ (_03090_, _07219_, _07069_);
  or _26150_ (_03092_, _03090_, _03089_);
  and _26151_ (_03869_, _03092_, _06444_);
  nand _26152_ (_03093_, _09484_, _07300_);
  and _26153_ (_03094_, _09482_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and _26154_ (_03095_, _09481_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or _26155_ (_03096_, _03095_, _03094_);
  or _26156_ (_03097_, _03096_, _09484_);
  and _26157_ (_03098_, _03097_, _09684_);
  and _26158_ (_03099_, _03098_, _03093_);
  and _26159_ (_03100_, _09479_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  or _26160_ (_03101_, _03100_, _03099_);
  and _26161_ (_03911_, _03101_, _06444_);
  nand _26162_ (_03102_, _10494_, _09484_);
  and _26163_ (_03103_, _09482_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and _26164_ (_03104_, _09481_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  or _26165_ (_03105_, _03104_, _03103_);
  or _26166_ (_03106_, _03105_, _09484_);
  and _26167_ (_03107_, _03106_, _09684_);
  and _26168_ (_03108_, _03107_, _03102_);
  and _26169_ (_03109_, _09479_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  or _26170_ (_03110_, _03109_, _03108_);
  and _26171_ (_03914_, _03110_, _06444_);
  and _26172_ (_03111_, _06430_, _06395_);
  and _26173_ (_03112_, _08976_, _03111_);
  and _26174_ (_03113_, _03112_, _06941_);
  and _26175_ (_03114_, _03113_, _06440_);
  or _26176_ (_03115_, _09481_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  not _26177_ (_03116_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  nand _26178_ (_03117_, _09481_, _03116_);
  nand _26179_ (_03119_, _03117_, _03115_);
  nor _26180_ (_03120_, _03119_, _03114_);
  not _26181_ (_03121_, _03114_);
  nor _26182_ (_03122_, _03121_, _06666_);
  or _26183_ (_03123_, _03122_, _03120_);
  or _26184_ (_03124_, _03123_, _09479_);
  or _26185_ (_03125_, _09684_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and _26186_ (_03126_, _03125_, _06444_);
  and _26187_ (_03917_, _03126_, _03124_);
  nand _26188_ (_03127_, _09484_, _07188_);
  and _26189_ (_03128_, _09482_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and _26190_ (_03129_, _09481_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or _26191_ (_03130_, _03129_, _03128_);
  or _26192_ (_03131_, _03130_, _09484_);
  and _26193_ (_03133_, _03131_, _09684_);
  and _26194_ (_03134_, _03133_, _03127_);
  and _26195_ (_03135_, _09479_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  or _26196_ (_03136_, _03135_, _03134_);
  and _26197_ (_03923_, _03136_, _06444_);
  and _26198_ (_03137_, _09482_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and _26199_ (_03138_, _09481_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  nor _26200_ (_03139_, _03138_, _03137_);
  nor _26201_ (_03140_, _03139_, _03114_);
  nor _26202_ (_03141_, _11589_, _03121_);
  or _26203_ (_03142_, _03141_, _03140_);
  or _26204_ (_03143_, _03142_, _09479_);
  or _26205_ (_03145_, _09684_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and _26206_ (_03146_, _03145_, _06444_);
  and _26207_ (_03935_, _03146_, _03143_);
  and _26208_ (_03148_, _07046_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  nor _26209_ (_03149_, _11589_, _07046_);
  or _26210_ (_03151_, _03149_, _03148_);
  and _26211_ (_03944_, _03151_, _06444_);
  or _26212_ (_03152_, _09481_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  or _26213_ (_03153_, _09482_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and _26214_ (_03154_, _03153_, _03152_);
  or _26215_ (_03155_, _03154_, _09484_);
  nand _26216_ (_03156_, _09484_, _07069_);
  and _26217_ (_03157_, _03156_, _03155_);
  or _26218_ (_03158_, _03157_, _09479_);
  or _26219_ (_03159_, _09684_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and _26220_ (_03160_, _03159_, _06444_);
  and _26221_ (_03958_, _03160_, _03158_);
  nand _26222_ (_03161_, _09526_, _09484_);
  or _26223_ (_03162_, _09481_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  or _26224_ (_03163_, _09482_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and _26225_ (_03164_, _03163_, _03162_);
  or _26226_ (_03165_, _03164_, _09484_);
  and _26227_ (_03166_, _03165_, _03161_);
  or _26228_ (_03167_, _03166_, _09479_);
  or _26229_ (_03168_, _09684_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  and _26230_ (_03169_, _03168_, _06444_);
  and _26231_ (_03962_, _03169_, _03167_);
  and _26232_ (_03170_, _02306_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  or _26233_ (_03171_, _02574_, _11381_);
  or _26234_ (_03172_, _03171_, _02734_);
  and _26235_ (_03173_, _02260_, _11347_);
  or _26236_ (_03174_, _02278_, _11440_);
  or _26237_ (_03175_, _03174_, _03173_);
  or _26238_ (_03176_, _02254_, _11409_);
  or _26239_ (_03177_, _02737_, _02483_);
  or _26240_ (_03178_, _03177_, _03176_);
  or _26241_ (_03179_, _02323_, _11343_);
  or _26242_ (_03180_, _03179_, _11442_);
  nor _26243_ (_03181_, _03180_, _11483_);
  nand _26244_ (_03182_, _03181_, _11514_);
  or _26245_ (_03183_, _03182_, _03178_);
  or _26246_ (_03184_, _03183_, _03175_);
  or _26247_ (_03185_, _03184_, _03172_);
  or _26248_ (_03186_, _11398_, _11342_);
  nor _26249_ (_03187_, rst, \oc8051_top_1.oc8051_sfr1.wait_data );
  and _26250_ (_03188_, _03187_, _03186_);
  and _26251_ (_03189_, _03188_, _03185_);
  or _26252_ (_03981_, _03189_, _03170_);
  nor _26253_ (_03190_, _14070_, _06978_);
  and _26254_ (_03191_, _14070_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  or _26255_ (_03192_, _03191_, _03190_);
  and _26256_ (_03986_, _03192_, _06444_);
  and _26257_ (_03193_, _02306_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  or _26258_ (_03194_, _02276_, _11977_);
  or _26259_ (_03195_, _02483_, _11438_);
  nor _26260_ (_03197_, _03195_, _03194_);
  nand _26261_ (_03198_, _03197_, _14227_);
  and _26262_ (_03199_, _11486_, _11355_);
  or _26263_ (_03200_, _02720_, _11489_);
  or _26264_ (_03201_, _03200_, _03199_);
  or _26265_ (_03202_, _03201_, _02954_);
  or _26266_ (_03203_, _03202_, _03198_);
  nor _26267_ (_03204_, _11479_, _11398_);
  nand _26268_ (_03205_, _03204_, _11445_);
  and _26269_ (_03206_, _11431_, _11355_);
  or _26270_ (_03207_, _02722_, _03206_);
  or _26271_ (_03208_, _03207_, _03205_);
  or _26272_ (_03209_, _03208_, _02495_);
  or _26273_ (_03210_, _03209_, _02499_);
  or _26274_ (_03211_, _03210_, _03203_);
  and _26275_ (_03212_, _03211_, _03188_);
  or _26276_ (_03989_, _03212_, _03193_);
  or _26277_ (_03213_, _11442_, _11428_);
  or _26278_ (_03214_, _03213_, _02276_);
  or _26279_ (_03215_, _03214_, _11438_);
  or _26280_ (_03216_, _03215_, _02494_);
  or _26281_ (_03217_, _03201_, _02498_);
  or _26282_ (_03218_, _03217_, _03216_);
  or _26283_ (_03219_, _02559_, _14226_);
  and _26284_ (_03220_, _02260_, _11360_);
  or _26285_ (_03221_, _03220_, _02946_);
  or _26286_ (_03222_, _03221_, _03219_);
  or _26287_ (_03223_, _03222_, _02959_);
  or _26288_ (_03224_, _03223_, _03218_);
  and _26289_ (_03225_, _03224_, _07230_);
  and _26290_ (_03226_, \oc8051_top_1.oc8051_decoder1.alu_op [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and _26291_ (_03227_, _11396_, _06308_);
  or _26292_ (_03228_, _03227_, _03226_);
  or _26293_ (_03229_, _03228_, _03225_);
  and _26294_ (_03994_, _03229_, _06444_);
  and _26295_ (_03230_, _07046_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  nor _26296_ (_03231_, _07046_, _06666_);
  or _26297_ (_03232_, _03231_, _03230_);
  and _26298_ (_03996_, _03232_, _06444_);
  nor _26299_ (_04000_, _12154_, rst);
  and _26300_ (_03233_, _02306_, \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  or _26301_ (_03234_, _02254_, _02264_);
  or _26302_ (_03235_, _03234_, _02469_);
  nor _26303_ (_03236_, _11533_, _11966_);
  nand _26304_ (_03237_, _03236_, _11978_);
  or _26305_ (_03238_, _03237_, _03235_);
  or _26306_ (_03239_, _02952_, _02947_);
  or _26307_ (_03240_, _03239_, _03238_);
  or _26308_ (_03241_, _03240_, _02589_);
  and _26309_ (_03242_, _03241_, _02332_);
  or _26310_ (_04011_, _03242_, _03233_);
  nor _26311_ (_03243_, _06978_, _09146_);
  and _26312_ (_03244_, _09146_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  or _26313_ (_03245_, _03244_, _07158_);
  or _26314_ (_03246_, _03245_, _03243_);
  or _26315_ (_03247_, _06439_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  and _26316_ (_03248_, _03247_, _06444_);
  and _26317_ (_04025_, _03248_, _03246_);
  or _26318_ (_03249_, _07432_, \oc8051_top_1.oc8051_rom1.data_o [11]);
  nand _26319_ (_03250_, _07432_, _13968_);
  and _26320_ (_03251_, _03250_, _06444_);
  and _26321_ (_04050_, _03251_, _03249_);
  or _26322_ (_03252_, _07432_, \oc8051_top_1.oc8051_rom1.data_o [10]);
  nand _26323_ (_03253_, _07432_, _13999_);
  and _26324_ (_03254_, _03253_, _06444_);
  and _26325_ (_04052_, _03254_, _03252_);
  or _26326_ (_03255_, _07432_, \oc8051_top_1.oc8051_rom1.data_o [9]);
  nand _26327_ (_03256_, _07432_, _12812_);
  and _26328_ (_03257_, _03256_, _06444_);
  and _26329_ (_04057_, _03257_, _03255_);
  and _26330_ (_04074_, _06444_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  and _26331_ (_03258_, _07459_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or _26332_ (_03259_, _07459_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand _26333_ (_03260_, _03259_, _06444_);
  nor _26334_ (_04088_, _03260_, _03258_);
  and _26335_ (_04094_, _08201_, _06444_);
  and _26336_ (_03261_, _09328_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  and _26337_ (_03262_, _11882_, _07151_);
  and _26338_ (_03263_, _09332_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  or _26339_ (_03264_, _03263_, _03262_);
  and _26340_ (_03265_, _03264_, _06439_);
  or _26341_ (_03266_, _03265_, _03261_);
  and _26342_ (_04095_, _03266_, _06444_);
  nand _26343_ (_03267_, _10494_, _10112_);
  or _26344_ (_03268_, _10112_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  and _26345_ (_03269_, _03268_, _06444_);
  and _26346_ (_04105_, _03269_, _03267_);
  nor _26347_ (_03270_, _12615_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor _26348_ (_03271_, _03270_, _12616_);
  or _26349_ (_03272_, _03271_, _12023_);
  and _26350_ (_03273_, _03272_, _06444_);
  not _26351_ (_03274_, _12023_);
  and _26352_ (_03275_, _12659_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  or _26353_ (_03276_, _03275_, _12661_);
  or _26354_ (_03277_, _12665_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _26355_ (_03278_, _03277_, _12666_);
  or _26356_ (_03279_, _03278_, _12650_);
  and _26357_ (_03280_, _03279_, _12218_);
  and _26358_ (_03281_, _03280_, _03276_);
  nor _26359_ (_03282_, _12681_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor _26360_ (_03283_, _03282_, _12682_);
  and _26361_ (_03284_, _03283_, _12054_);
  and _26362_ (_03285_, _11452_, _08308_);
  and _26363_ (_03286_, _12026_, _08342_);
  and _26364_ (_03287_, _11689_, _12032_);
  and _26365_ (_03288_, _12047_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  or _26366_ (_03289_, _03288_, _03287_);
  or _26367_ (_03290_, _03289_, _03286_);
  or _26368_ (_03291_, _03290_, _03285_);
  or _26369_ (_03292_, _03291_, _03284_);
  or _26370_ (_03294_, _03292_, _03281_);
  or _26371_ (_03296_, _03294_, _03274_);
  and _26372_ (_04109_, _03296_, _03273_);
  nor _26373_ (_03297_, _00855_, _09138_);
  not _26374_ (_03298_, _12026_);
  nor _26375_ (_03299_, _03298_, _09280_);
  and _26376_ (_03301_, _11905_, _12032_);
  and _26377_ (_03302_, _12047_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  or _26378_ (_03303_, _03302_, _03301_);
  or _26379_ (_03305_, _03303_, _03299_);
  or _26380_ (_03306_, _03305_, _03297_);
  and _26381_ (_03308_, _12658_, _12650_);
  nor _26382_ (_03310_, _12664_, _12650_);
  or _26383_ (_03311_, _03310_, _03308_);
  nand _26384_ (_03312_, _03311_, _08143_);
  or _26385_ (_03313_, _03311_, _08143_);
  and _26386_ (_03314_, _03313_, _03312_);
  and _26387_ (_03315_, _03314_, _12218_);
  or _26388_ (_03316_, _03315_, _03306_);
  nand _26389_ (_03317_, _12054_, _08360_);
  nand _26390_ (_03318_, _03317_, _12023_);
  or _26391_ (_03319_, _03318_, _03316_);
  nor _26392_ (_03320_, _12614_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor _26393_ (_03322_, _03320_, _12615_);
  or _26394_ (_03323_, _03322_, _12023_);
  and _26395_ (_03324_, _03323_, _06444_);
  and _26396_ (_04113_, _03324_, _03319_);
  and _26397_ (_03326_, _12656_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  or _26398_ (_03327_, _03326_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and _26399_ (_03328_, _03327_, _03310_);
  nand _26400_ (_03329_, _12657_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nand _26401_ (_03330_, _03329_, _12658_);
  and _26402_ (_03332_, _03330_, _12650_);
  or _26403_ (_03333_, _03332_, _03328_);
  and _26404_ (_03334_, _03333_, _12218_);
  nor _26405_ (_03335_, _03298_, _07640_);
  and _26406_ (_03336_, _11452_, _07959_);
  and _26407_ (_03337_, _12032_, _11794_);
  and _26408_ (_03338_, _12054_, _10739_);
  and _26409_ (_03339_, _12047_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  or _26410_ (_03340_, _03339_, _03338_);
  or _26411_ (_03341_, _03340_, _03337_);
  or _26412_ (_03342_, _03341_, _03336_);
  or _26413_ (_03343_, _03342_, _03335_);
  or _26414_ (_03345_, _03343_, _03334_);
  or _26415_ (_03346_, _03345_, _03274_);
  nor _26416_ (_03347_, _12613_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  nor _26417_ (_03348_, _03347_, _12614_);
  or _26418_ (_03349_, _03348_, _12023_);
  and _26419_ (_03351_, _03349_, _06444_);
  and _26420_ (_04123_, _03351_, _03346_);
  and _26421_ (_03352_, _11452_, _08019_);
  and _26422_ (_03353_, _12054_, _08457_);
  nor _26423_ (_03354_, _03298_, _08060_);
  and _26424_ (_03356_, _11848_, _12032_);
  and _26425_ (_03358_, _12047_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  or _26426_ (_03359_, _03358_, _03356_);
  or _26427_ (_03361_, _03359_, _03354_);
  or _26428_ (_03362_, _03361_, _03353_);
  nor _26429_ (_03363_, _03362_, _03352_);
  nand _26430_ (_03364_, _03363_, _12023_);
  nand _26431_ (_03365_, _12656_, _07589_);
  or _26432_ (_03366_, _12656_, _07589_);
  and _26433_ (_03367_, _03366_, _03365_);
  nor _26434_ (_03368_, _03367_, _12650_);
  and _26435_ (_03369_, _03367_, _12650_);
  or _26436_ (_03370_, _03369_, _03368_);
  and _26437_ (_03371_, _03370_, _12606_);
  or _26438_ (_03372_, _03371_, _03364_);
  nor _26439_ (_03373_, _12612_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor _26440_ (_03374_, _03373_, _12613_);
  or _26441_ (_03375_, _03374_, _12023_);
  and _26442_ (_03376_, _03375_, _06444_);
  and _26443_ (_04126_, _03376_, _03372_);
  nor _26444_ (_03377_, _12227_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor _26445_ (_03378_, _03377_, _12612_);
  or _26446_ (_03379_, _03378_, _12023_);
  and _26447_ (_03380_, _03379_, _06444_);
  nor _26448_ (_03381_, _12654_, _12653_);
  nor _26449_ (_03382_, _03381_, _12655_);
  and _26450_ (_03383_, _03382_, _12218_);
  and _26451_ (_03384_, _12048_, _11137_);
  and _26452_ (_03386_, _11452_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor _26453_ (_03387_, _12648_, _12033_);
  and _26454_ (_03388_, _12054_, _11625_);
  or _26455_ (_03389_, _03388_, _03387_);
  or _26456_ (_03390_, _03389_, _03386_);
  or _26457_ (_03391_, _03390_, _03384_);
  nor _26458_ (_03392_, _03391_, _03383_);
  nand _26459_ (_03393_, _03392_, _12023_);
  and _26460_ (_04131_, _03393_, _03380_);
  nor _26461_ (_03394_, _03258_, _07471_);
  and _26462_ (_03395_, _03258_, _07471_);
  or _26463_ (_03396_, _03395_, _03394_);
  and _26464_ (_04192_, _03396_, _06444_);
  and _26465_ (_04195_, _11102_, _06444_);
  and _26466_ (_04203_, _06444_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  or _26467_ (_03397_, _07414_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  nand _26468_ (_03399_, _07069_, _07414_);
  and _26469_ (_03400_, _03399_, _03397_);
  or _26470_ (_03401_, _03400_, _07158_);
  or _26471_ (_03402_, _06439_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  and _26472_ (_03403_, _03402_, _06444_);
  and _26473_ (_04204_, _03403_, _03401_);
  not _26474_ (_03404_, _00936_);
  or _26475_ (_03405_, _03404_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  or _26476_ (_03407_, _00936_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  and _26477_ (_03408_, _03407_, _03405_);
  and _26478_ (_03409_, _03408_, _06443_);
  and _26479_ (_03410_, _06442_, _06296_);
  or _26480_ (_03411_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3], _13875_);
  and _26481_ (_03412_, _03411_, _06444_);
  and _26482_ (_03413_, _03412_, _03410_);
  or _26483_ (_04206_, _03413_, _03409_);
  nor _26484_ (_03415_, _07300_, _09146_);
  and _26485_ (_03416_, _09146_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  or _26486_ (_03417_, _03416_, _07158_);
  or _26487_ (_03418_, _03417_, _03415_);
  or _26488_ (_03419_, _06439_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  and _26489_ (_03420_, _03419_, _06444_);
  and _26490_ (_04208_, _03420_, _03418_);
  nor _26491_ (_03421_, _10494_, _09146_);
  and _26492_ (_03422_, _09146_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  or _26493_ (_03423_, _03422_, _07158_);
  or _26494_ (_03424_, _03423_, _03421_);
  or _26495_ (_03426_, _06439_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  and _26496_ (_03427_, _03426_, _06444_);
  and _26497_ (_04210_, _03427_, _03424_);
  nor _26498_ (_03430_, _14085_, _11669_);
  and _26499_ (_03431_, _03430_, _14142_);
  or _26500_ (_03432_, _01519_, _14113_);
  or _26501_ (_03433_, _11919_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and _26502_ (_03434_, _03433_, _14079_);
  and _26503_ (_03435_, _03434_, _03432_);
  and _26504_ (_03436_, _14113_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and _26505_ (_03437_, _11919_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  or _26506_ (_03438_, _03437_, _03436_);
  and _26507_ (_03439_, _03438_, _14094_);
  or _26508_ (_03440_, _14113_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  or _26509_ (_03441_, _11919_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  and _26510_ (_03442_, _03441_, _14103_);
  and _26511_ (_03443_, _03442_, _03440_);
  or _26512_ (_03444_, _03443_, _03439_);
  or _26513_ (_03445_, _11919_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  or _26514_ (_03446_, _14113_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  and _26515_ (_03447_, _03446_, _14091_);
  and _26516_ (_03448_, _03447_, _03445_);
  or _26517_ (_03449_, _03448_, _03444_);
  or _26518_ (_03450_, _03449_, _03435_);
  and _26519_ (_03451_, _03450_, _03431_);
  nor _26520_ (_03452_, _11919_, _07098_);
  and _26521_ (_03453_, _11919_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  or _26522_ (_03454_, _03453_, _03452_);
  and _26523_ (_03455_, _03454_, _14079_);
  or _26524_ (_03456_, _14113_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  or _26525_ (_03457_, _11919_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and _26526_ (_03458_, _03457_, _14094_);
  and _26527_ (_03459_, _03458_, _03456_);
  or _26528_ (_03461_, _03459_, _03455_);
  and _26529_ (_03462_, _14113_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and _26530_ (_03463_, _11919_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or _26531_ (_03464_, _03463_, _03462_);
  and _26532_ (_03465_, _03464_, _14091_);
  or _26533_ (_03466_, _11919_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  or _26534_ (_03467_, _14113_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and _26535_ (_03468_, _03467_, _14103_);
  and _26536_ (_03469_, _03468_, _03466_);
  or _26537_ (_03470_, _03469_, _03465_);
  or _26538_ (_03471_, _03470_, _03461_);
  and _26539_ (_03472_, _03471_, _14109_);
  or _26540_ (_03473_, _14113_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  or _26541_ (_03474_, _11919_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and _26542_ (_03475_, _03474_, _14079_);
  and _26543_ (_03476_, _03475_, _03473_);
  or _26544_ (_03477_, _14113_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or _26545_ (_03478_, _11919_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and _26546_ (_03479_, _03478_, _14094_);
  and _26547_ (_03480_, _03479_, _03477_);
  or _26548_ (_03481_, _03480_, _03476_);
  and _26549_ (_03482_, _14113_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and _26550_ (_03484_, _11919_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or _26551_ (_03485_, _03484_, _03482_);
  and _26552_ (_03486_, _03485_, _14091_);
  or _26553_ (_03487_, _11919_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or _26554_ (_03488_, _14113_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and _26555_ (_03489_, _03488_, _14103_);
  and _26556_ (_03490_, _03489_, _03487_);
  or _26557_ (_03491_, _03490_, _03486_);
  or _26558_ (_03492_, _03491_, _03481_);
  and _26559_ (_03493_, _03492_, _14101_);
  nor _26560_ (_03494_, _11919_, _07110_);
  and _26561_ (_03496_, _11919_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  or _26562_ (_03497_, _03496_, _03494_);
  and _26563_ (_03498_, _03497_, _14094_);
  nand _26564_ (_03499_, _11919_, _07118_);
  or _26565_ (_03500_, _11919_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and _26566_ (_03501_, _03500_, _14079_);
  and _26567_ (_03503_, _03501_, _03499_);
  or _26568_ (_03504_, _03503_, _03498_);
  or _26569_ (_03505_, _11919_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  nand _26570_ (_03506_, _11919_, _07115_);
  and _26571_ (_03507_, _03506_, _14103_);
  and _26572_ (_03508_, _03507_, _03505_);
  or _26573_ (_03509_, _11919_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  nand _26574_ (_03510_, _11919_, _07123_);
  and _26575_ (_03511_, _03510_, _14091_);
  and _26576_ (_03512_, _03511_, _03509_);
  or _26577_ (_03513_, _03512_, _03508_);
  or _26578_ (_03514_, _03513_, _03504_);
  and _26579_ (_03516_, _03514_, _14112_);
  or _26580_ (_03517_, _03516_, _03493_);
  or _26581_ (_03518_, _03517_, _03472_);
  and _26582_ (_03519_, _03518_, _14085_);
  and _26583_ (_03520_, _14108_, _11703_);
  nor _26584_ (_03521_, _03431_, _03520_);
  nand _26585_ (_03522_, _14144_, _11703_);
  and _26586_ (_03524_, _03522_, _03521_);
  nand _26587_ (_03525_, _14129_, _11703_);
  and _26588_ (_03526_, _14083_, _14085_);
  and _26589_ (_03527_, _14101_, _11703_);
  nand _26590_ (_03528_, _14100_, _14085_);
  nand _26591_ (_03529_, _03528_, \oc8051_top_1.oc8051_sfr1.bit_out );
  or _26592_ (_03530_, _03529_, _03527_);
  nor _26593_ (_03531_, _03530_, _03526_);
  and _26594_ (_03533_, _03531_, _03525_);
  and _26595_ (_03534_, _03533_, _03524_);
  and _26596_ (_03535_, _14103_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  and _26597_ (_03536_, _14079_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  or _26598_ (_03538_, _03536_, _11919_);
  or _26599_ (_03539_, _03538_, _03535_);
  and _26600_ (_03540_, _14103_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  and _26601_ (_03541_, _14079_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or _26602_ (_03542_, _03541_, _14113_);
  or _26603_ (_03543_, _03542_, _03540_);
  and _26604_ (_03544_, _03543_, _03539_);
  or _26605_ (_03546_, _11919_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  nand _26606_ (_03548_, _11919_, _01116_);
  and _26607_ (_03549_, _03548_, _14091_);
  and _26608_ (_03550_, _03549_, _03546_);
  nor _26609_ (_03551_, _11919_, _01311_);
  and _26610_ (_03552_, _11919_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  or _26611_ (_03553_, _03552_, _03551_);
  and _26612_ (_03555_, _03553_, _14094_);
  or _26613_ (_03556_, _03555_, _11703_);
  or _26614_ (_03557_, _03556_, _03550_);
  or _26615_ (_03558_, _03557_, _03544_);
  or _26616_ (_03559_, _14247_, p1_in[7]);
  or _26617_ (_03560_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and _26618_ (_03561_, _03560_, _03559_);
  and _26619_ (_03562_, _03561_, _14103_);
  and _26620_ (_03563_, _14256_, _14091_);
  or _26621_ (_03564_, _03563_, _11919_);
  or _26622_ (_03565_, _03564_, _03562_);
  and _26623_ (_03566_, _14329_, _14103_);
  and _26624_ (_03567_, _14417_, _14091_);
  or _26625_ (_03568_, _03567_, _14113_);
  or _26626_ (_03569_, _03568_, _03566_);
  and _26627_ (_03570_, _03569_, _03565_);
  or _26628_ (_03571_, _01471_, _14113_);
  or _26629_ (_03572_, _01393_, _11919_);
  and _26630_ (_03574_, _03572_, _14079_);
  and _26631_ (_03575_, _03574_, _03571_);
  or _26632_ (_03576_, _14483_, _14113_);
  or _26633_ (_03577_, _01249_, _11919_);
  and _26634_ (_03578_, _03577_, _14094_);
  and _26635_ (_03579_, _03578_, _03576_);
  or _26636_ (_03580_, _03579_, _14085_);
  or _26637_ (_03581_, _03580_, _03575_);
  or _26638_ (_03582_, _03581_, _03570_);
  and _26639_ (_03583_, _03582_, _14129_);
  and _26640_ (_03584_, _03583_, _03558_);
  and _26641_ (_03585_, _11925_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and _26642_ (_03586_, _14079_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and _26643_ (_03587_, _14091_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or _26644_ (_03588_, _03587_, _03586_);
  and _26645_ (_03589_, _14103_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  and _26646_ (_03590_, _14094_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  or _26647_ (_03591_, _03590_, _03589_);
  or _26648_ (_03592_, _03591_, _03588_);
  and _26649_ (_03593_, _03592_, _14113_);
  and _26650_ (_03594_, _14079_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and _26651_ (_03595_, _14091_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or _26652_ (_03596_, _03595_, _03594_);
  and _26653_ (_03598_, _14103_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and _26654_ (_03600_, _14094_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or _26655_ (_03601_, _03600_, _03598_);
  or _26656_ (_03602_, _03601_, _03596_);
  and _26657_ (_03603_, _03602_, _11919_);
  or _26658_ (_03604_, _03603_, _03593_);
  and _26659_ (_03605_, _03604_, _03526_);
  or _26660_ (_03607_, _03605_, _03585_);
  or _26661_ (_03608_, _03607_, _03584_);
  or _26662_ (_03609_, _03608_, _03534_);
  or _26663_ (_03610_, _14474_, _14113_);
  or _26664_ (_03611_, _01239_, _11919_);
  and _26665_ (_03612_, _03611_, _14094_);
  and _26666_ (_03613_, _03612_, _03610_);
  or _26667_ (_03614_, _14268_, _11919_);
  or _26668_ (_03615_, _14403_, _14113_);
  and _26669_ (_03616_, _03615_, _14091_);
  and _26670_ (_03617_, _03616_, _03614_);
  or _26671_ (_03618_, _03617_, _03613_);
  or _26672_ (_03619_, _01462_, _14113_);
  or _26673_ (_03620_, _01403_, _11919_);
  and _26674_ (_03622_, _03620_, _14079_);
  and _26675_ (_03624_, _03622_, _03619_);
  or _26676_ (_03626_, _14334_, _14113_);
  or _26677_ (_03628_, _14247_, p2_in[7]);
  or _26678_ (_03629_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and _26679_ (_03631_, _03629_, _03628_);
  or _26680_ (_03633_, _03631_, _11919_);
  and _26681_ (_03635_, _03633_, _14103_);
  and _26682_ (_03636_, _03635_, _03626_);
  or _26683_ (_03638_, _03636_, _03624_);
  or _26684_ (_03639_, _03638_, _03618_);
  and _26685_ (_03641_, _03639_, _11669_);
  and _26686_ (_03642_, _01399_, _14079_);
  or _26687_ (_03643_, _03642_, _11919_);
  and _26688_ (_03645_, _14263_, _14091_);
  and _26689_ (_03647_, _01235_, _14094_);
  or _26690_ (_03649_, _14247_, p3_in[7]);
  or _26691_ (_03650_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and _26692_ (_03652_, _03650_, _03649_);
  and _26693_ (_03654_, _03652_, _14103_);
  or _26694_ (_03655_, _03654_, _03647_);
  or _26695_ (_03657_, _03655_, _03645_);
  or _26696_ (_03659_, _03657_, _03643_);
  and _26697_ (_03661_, _14470_, _14094_);
  or _26698_ (_03662_, _03661_, _14113_);
  and _26699_ (_03664_, _01458_, _14079_);
  and _26700_ (_03665_, _14338_, _14103_);
  and _26701_ (_03666_, _14407_, _14091_);
  or _26702_ (_03668_, _03666_, _03665_);
  or _26703_ (_03670_, _03668_, _03664_);
  or _26704_ (_03671_, _03670_, _03662_);
  and _26705_ (_03672_, _03671_, _14111_);
  and _26706_ (_03673_, _03672_, _03659_);
  or _26707_ (_03674_, _03673_, _03641_);
  and _26708_ (_03675_, _03674_, _03520_);
  and _26709_ (_03676_, _01389_, _14113_);
  and _26710_ (_03677_, _01467_, _11919_);
  or _26711_ (_03679_, _03677_, _03676_);
  and _26712_ (_03680_, _03679_, _14079_);
  or _26713_ (_03681_, _14479_, _14113_);
  or _26714_ (_03682_, _01244_, _11919_);
  and _26715_ (_03683_, _03682_, _14094_);
  and _26716_ (_03684_, _03683_, _03681_);
  or _26717_ (_03686_, _14412_, _14113_);
  or _26718_ (_03687_, _14251_, _11919_);
  and _26719_ (_03689_, _03687_, _14091_);
  and _26720_ (_03690_, _03689_, _03686_);
  or _26721_ (_03691_, _14325_, _14113_);
  or _26722_ (_03693_, _14247_, p0_in[7]);
  or _26723_ (_03694_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and _26724_ (_03695_, _03694_, _03693_);
  or _26725_ (_03696_, _03695_, _11919_);
  and _26726_ (_03697_, _03696_, _14103_);
  and _26727_ (_03698_, _03697_, _03691_);
  or _26728_ (_03699_, _03698_, _03690_);
  or _26729_ (_03701_, _03699_, _03684_);
  or _26730_ (_03702_, _03701_, _03680_);
  and _26731_ (_03703_, _03702_, _03527_);
  and _26732_ (_03704_, _03430_, _14144_);
  and _26733_ (_03706_, _14094_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and _26734_ (_03707_, _14091_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  or _26735_ (_03709_, _03707_, _03706_);
  and _26736_ (_03711_, _03709_, _14113_);
  and _26737_ (_03713_, _14094_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and _26738_ (_03714_, _14091_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or _26739_ (_03716_, _03714_, _03713_);
  and _26740_ (_03717_, _03716_, _11919_);
  not _26741_ (_03719_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  nor _26742_ (_03721_, _11919_, _03719_);
  and _26743_ (_03722_, _11919_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  or _26744_ (_03723_, _03722_, _03721_);
  and _26745_ (_03724_, _03723_, _14103_);
  nor _26746_ (_03725_, _11919_, _02653_);
  and _26747_ (_03726_, _11919_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  or _26748_ (_03727_, _03726_, _03725_);
  and _26749_ (_03728_, _03727_, _14079_);
  or _26750_ (_03729_, _03728_, _03724_);
  or _26751_ (_03730_, _03729_, _03717_);
  or _26752_ (_03731_, _03730_, _03711_);
  and _26753_ (_03732_, _03731_, _03704_);
  and _26754_ (_03734_, _11703_, _11669_);
  and _26755_ (_03735_, _03734_, _14144_);
  and _26756_ (_03736_, _14094_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and _26757_ (_03738_, _14091_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or _26758_ (_03739_, _03738_, _03736_);
  and _26759_ (_03740_, _14103_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and _26760_ (_03741_, _14079_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or _26761_ (_03742_, _03741_, _03740_);
  or _26762_ (_03744_, _03742_, _03739_);
  and _26763_ (_03745_, _03744_, _11919_);
  and _26764_ (_03746_, _14094_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and _26765_ (_03748_, _14091_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or _26766_ (_03749_, _03748_, _03746_);
  and _26767_ (_03750_, _14103_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and _26768_ (_03751_, _14079_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or _26769_ (_03753_, _03751_, _03750_);
  or _26770_ (_03754_, _03753_, _03749_);
  and _26771_ (_03755_, _03754_, _14113_);
  or _26772_ (_03757_, _03755_, _03745_);
  and _26773_ (_03759_, _03757_, _03735_);
  or _26774_ (_03760_, _03759_, _03732_);
  or _26775_ (_03761_, _03760_, _03703_);
  or _26776_ (_03762_, _03761_, _03675_);
  or _26777_ (_03763_, _03762_, _03609_);
  or _26778_ (_03764_, _03763_, _03519_);
  or _26779_ (_03766_, _03764_, _03451_);
  and _26780_ (_03767_, _03735_, _07646_);
  nor _26781_ (_03768_, _03767_, _11931_);
  nand _26782_ (_03769_, _03585_, _06930_);
  and _26783_ (_03770_, _03769_, _03768_);
  and _26784_ (_03771_, _03770_, _03766_);
  and _26785_ (_03772_, _14103_, _11568_);
  and _26786_ (_03773_, _14091_, _11763_);
  or _26787_ (_03774_, _03773_, _03772_);
  and _26788_ (_03775_, _03774_, _14113_);
  and _26789_ (_03776_, _14103_, _07340_);
  and _26790_ (_03777_, _14091_, _11882_);
  or _26791_ (_03778_, _03777_, _03776_);
  and _26792_ (_03779_, _03778_, _11919_);
  nor _26793_ (_03780_, _11919_, _06666_);
  and _26794_ (_03781_, _11919_, _07070_);
  or _26795_ (_03782_, _03781_, _03780_);
  and _26796_ (_03783_, _03782_, _14094_);
  nor _26797_ (_03785_, _11919_, _07188_);
  and _26798_ (_03786_, _11919_, _09527_);
  or _26799_ (_03788_, _03786_, _03785_);
  and _26800_ (_03789_, _03788_, _14079_);
  or _26801_ (_03790_, _03789_, _03783_);
  or _26802_ (_03792_, _03790_, _03779_);
  nor _26803_ (_03793_, _03792_, _03775_);
  nor _26804_ (_03795_, _03793_, _03768_);
  or _26805_ (_03796_, _03795_, _03771_);
  and _26806_ (_04214_, _03796_, _06444_);
  nor _26807_ (_03798_, _00469_, rst);
  or _26808_ (_03799_, _00468_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  nand _26809_ (_03801_, _00468_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  and _26810_ (_03803_, _03801_, _03799_);
  and _26811_ (_04218_, _03803_, _03798_);
  and _26812_ (_04220_, _00470_, _06444_);
  nor _26813_ (_03805_, _02821_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor _26814_ (_03806_, _03805_, _02822_);
  and _26815_ (_03808_, _03806_, _12054_);
  nor _26816_ (_03809_, _00855_, _09045_);
  nor _26817_ (_03810_, _03298_, _09201_);
  and _26818_ (_03811_, _12032_, _11778_);
  and _26819_ (_03813_, _12047_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or _26820_ (_03814_, _03813_, _03811_);
  or _26821_ (_03815_, _03814_, _03810_);
  or _26822_ (_03817_, _03815_, _03809_);
  or _26823_ (_03818_, _03817_, _03808_);
  and _26824_ (_03819_, _02812_, _12662_);
  and _26825_ (_03820_, _02808_, _12650_);
  or _26826_ (_03822_, _03820_, _03819_);
  nand _26827_ (_03823_, _03822_, _09186_);
  or _26828_ (_03825_, _03822_, _09186_);
  and _26829_ (_03826_, _03825_, _03823_);
  and _26830_ (_03827_, _03826_, _12218_);
  or _26831_ (_03829_, _03827_, _03818_);
  or _26832_ (_03830_, _03829_, _03274_);
  nor _26833_ (_03832_, _02793_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor _26834_ (_03834_, _03832_, _02794_);
  or _26835_ (_03836_, _03834_, _12023_);
  and _26836_ (_03838_, _03836_, _06444_);
  and _26837_ (_04222_, _03838_, _03830_);
  or _26838_ (_03841_, _12683_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  not _26839_ (_03843_, _02821_);
  and _26840_ (_03844_, _03843_, _12054_);
  and _26841_ (_03845_, _03844_, _03841_);
  and _26842_ (_03846_, _11452_, _08127_);
  and _26843_ (_03847_, _12026_, _08194_);
  and _26844_ (_03848_, _11726_, _12032_);
  and _26845_ (_03849_, _12047_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or _26846_ (_03850_, _03849_, _03848_);
  or _26847_ (_03852_, _03850_, _03847_);
  or _26848_ (_03853_, _03852_, _03846_);
  nand _26849_ (_03854_, _12650_, _08150_);
  nor _26850_ (_03855_, _03854_, _12660_);
  nor _26851_ (_03856_, _02811_, _12650_);
  nor _26852_ (_03857_, _03856_, _03855_);
  nand _26853_ (_03858_, _03857_, _08155_);
  or _26854_ (_03859_, _03857_, _08155_);
  and _26855_ (_03861_, _03859_, _03858_);
  and _26856_ (_03862_, _03861_, _12218_);
  or _26857_ (_03863_, _03862_, _03853_);
  or _26858_ (_03865_, _03863_, _03845_);
  or _26859_ (_03866_, _03865_, _03274_);
  nor _26860_ (_03867_, _02792_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor _26861_ (_03868_, _03867_, _02793_);
  or _26862_ (_03870_, _03868_, _12023_);
  and _26863_ (_03871_, _03870_, _06444_);
  and _26864_ (_04226_, _03871_, _03866_);
  or _26865_ (_03872_, _07432_, \oc8051_top_1.oc8051_rom1.data_o [0]);
  nand _26866_ (_03873_, _07432_, _14060_);
  and _26867_ (_03874_, _03873_, _06444_);
  and _26868_ (_04313_, _03874_, _03872_);
  or _26869_ (_03875_, _07432_, \oc8051_top_1.oc8051_rom1.data_o [2]);
  nand _26870_ (_03876_, _07432_, _14051_);
  and _26871_ (_03877_, _03876_, _06444_);
  and _26872_ (_04362_, _03877_, _03875_);
  not _26873_ (_03878_, _11453_);
  and _26874_ (_03879_, _11460_, _03878_);
  nor _26875_ (_03880_, _11533_, _11455_);
  nand _26876_ (_03881_, _03880_, _11492_);
  or _26877_ (_03882_, _03881_, _11509_);
  or _26878_ (_03883_, _03882_, _02947_);
  and _26879_ (_03884_, _03883_, _11342_);
  or _26880_ (_03885_, _03884_, _03879_);
  and _26881_ (_04364_, _03885_, _06444_);
  and _26882_ (_03886_, _14088_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  and _26883_ (_03887_, _14084_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or _26884_ (_03888_, _03887_, _03886_);
  and _26885_ (_03889_, _14096_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  and _26886_ (_03890_, _14093_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  or _26887_ (_03891_, _03890_, _03889_);
  or _26888_ (_03892_, _03891_, _03888_);
  and _26889_ (_03893_, _14102_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and _26890_ (_03894_, _14105_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  or _26891_ (_03895_, _03894_, _03893_);
  and _26892_ (_03896_, _14110_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and _26893_ (_03897_, _14116_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  or _26894_ (_03898_, _03897_, _03896_);
  or _26895_ (_03899_, _03898_, _03895_);
  or _26896_ (_03900_, _03899_, _03892_);
  and _26897_ (_03901_, _14120_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and _26898_ (_03902_, _14122_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  or _26899_ (_03903_, _03902_, _03901_);
  and _26900_ (_03904_, _14124_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and _26901_ (_03905_, _14125_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  or _26902_ (_03906_, _03905_, _03904_);
  or _26903_ (_03907_, _03906_, _03903_);
  and _26904_ (_03908_, _14130_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  and _26905_ (_03909_, _14131_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  or _26906_ (_03910_, _03909_, _03908_);
  and _26907_ (_03912_, _14133_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and _26908_ (_03913_, _14134_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or _26909_ (_03915_, _03913_, _03912_);
  or _26910_ (_03916_, _03915_, _03910_);
  or _26911_ (_03918_, _03916_, _03907_);
  or _26912_ (_03919_, _03918_, _03900_);
  and _26913_ (_03920_, _14154_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and _26914_ (_03921_, _14156_, _11622_);
  or _26915_ (_03922_, _03921_, _03920_);
  and _26916_ (_03924_, _14150_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and _26917_ (_03925_, _14152_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or _26918_ (_03926_, _03925_, _03924_);
  or _26919_ (_03927_, _03926_, _03922_);
  and _26920_ (_03928_, _03631_, _14265_);
  and _26921_ (_03929_, _03652_, _14260_);
  or _26922_ (_03930_, _03929_, _03928_);
  and _26923_ (_03931_, _03695_, _14224_);
  and _26924_ (_03932_, _03561_, _14253_);
  or _26925_ (_03933_, _03932_, _03931_);
  or _26926_ (_03934_, _03933_, _03930_);
  or _26927_ (_03936_, _03934_, _03927_);
  and _26928_ (_03937_, _14143_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  and _26929_ (_03938_, _14146_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or _26930_ (_03939_, _03938_, _03937_);
  or _26931_ (_03940_, _03939_, _03936_);
  or _26932_ (_03941_, _03940_, _03919_);
  and _26933_ (_03942_, _03941_, _14174_);
  and _26934_ (_03943_, _14175_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  or _26935_ (_03945_, _03943_, _03942_);
  or _26936_ (_03946_, _03945_, _14178_);
  or _26937_ (_03947_, _14353_, _11137_);
  and _26938_ (_03948_, _03947_, _06444_);
  and _26939_ (_04366_, _03948_, _03946_);
  or _26940_ (_03949_, _00936_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  or _26941_ (_03950_, _03404_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  and _26942_ (_03951_, _03950_, _03949_);
  or _26943_ (_03952_, _03951_, _06442_);
  and _26944_ (_03953_, _03952_, _06444_);
  nand _26945_ (_03954_, _03410_, _06978_);
  and _26946_ (_04369_, _03954_, _03953_);
  or _26947_ (_03955_, _02650_, _11137_);
  nand _26948_ (_03956_, _02650_, _03719_);
  and _26949_ (_03957_, _03956_, _06440_);
  and _26950_ (_03959_, _03957_, _03955_);
  nor _26951_ (_03960_, _06673_, _03719_);
  and _26952_ (_03961_, _02659_, _06933_);
  nand _26953_ (_03963_, _03961_, _06930_);
  or _26954_ (_03964_, _03961_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and _26955_ (_03965_, _03964_, _06674_);
  and _26956_ (_03966_, _03965_, _03963_);
  or _26957_ (_03967_, _03966_, _03960_);
  or _26958_ (_03968_, _03967_, _03959_);
  and _26959_ (_04377_, _03968_, _06444_);
  or _26960_ (_03969_, _03404_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  or _26961_ (_03970_, _00936_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  and _26962_ (_03971_, _03970_, _03969_);
  and _26963_ (_03972_, _03971_, _06443_);
  nand _26964_ (_03973_, _06978_, _06295_);
  nand _26965_ (_03974_, _10494_, _06296_);
  and _26966_ (_03975_, _03974_, _00933_);
  and _26967_ (_03976_, _03975_, _03973_);
  or _26968_ (_04379_, _03976_, _03972_);
  and _26969_ (_03977_, _06442_, _06295_);
  and _26970_ (_03978_, _03977_, _11763_);
  or _26971_ (_03979_, _00936_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  or _26972_ (_03980_, _03404_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  nand _26973_ (_03982_, _03980_, _03979_);
  nor _26974_ (_03983_, _03982_, _06442_);
  and _26975_ (_03984_, _03410_, _07378_);
  or _26976_ (_03985_, _03984_, _03983_);
  or _26977_ (_03987_, _03985_, _03978_);
  and _26978_ (_04383_, _03987_, _06444_);
  nor _26979_ (_04491_, _11904_, rst);
  nand _26980_ (_03988_, _06406_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  nor _26981_ (_03990_, _03988_, _00238_);
  or _26982_ (_03991_, _03990_, _01481_);
  and _26983_ (_03992_, _03991_, _00818_);
  nand _26984_ (_03993_, _00818_, _06406_);
  and _26985_ (_03995_, _03993_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or _26986_ (_03997_, _03995_, _07407_);
  or _26987_ (_03998_, _03997_, _03992_);
  nand _26988_ (_03999_, _10494_, _07407_);
  and _26989_ (_04001_, _03999_, _06444_);
  and _26990_ (_04530_, _04001_, _03998_);
  or _26991_ (_04002_, _07432_, \oc8051_top_1.oc8051_rom1.data_o [1]);
  nand _26992_ (_04003_, _07432_, _14056_);
  and _26993_ (_04004_, _04003_, _06444_);
  and _26994_ (_04533_, _04004_, _04002_);
  and _26995_ (_04005_, _00742_, _06933_);
  nand _26996_ (_04006_, _04005_, _06930_);
  or _26997_ (_04007_, _04005_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and _26998_ (_04008_, _04007_, _00748_);
  and _26999_ (_04009_, _04008_, _04006_);
  nor _27000_ (_04010_, _00748_, _06978_);
  or _27001_ (_04012_, _04010_, _04009_);
  and _27002_ (_04535_, _04012_, _06444_);
  and _27003_ (_04013_, _00669_, _06933_);
  nand _27004_ (_04014_, _04013_, _06930_);
  or _27005_ (_04015_, _04013_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and _27006_ (_04016_, _04015_, _00678_);
  and _27007_ (_04017_, _04016_, _04014_);
  nor _27008_ (_04018_, _00678_, _06978_);
  or _27009_ (_04019_, _04018_, _04017_);
  and _27010_ (_04538_, _04019_, _06444_);
  and _27011_ (_04020_, _08310_, _06678_);
  nand _27012_ (_04021_, _04020_, _06930_);
  or _27013_ (_04022_, _04020_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and _27014_ (_04023_, _04022_, _02416_);
  and _27015_ (_04024_, _04023_, _04021_);
  nor _27016_ (_04026_, _07300_, _02416_);
  or _27017_ (_04027_, _04026_, _04024_);
  and _27018_ (_04545_, _04027_, _06444_);
  and _27019_ (_04028_, _06431_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or _27020_ (_04029_, _04028_, _00713_);
  and _27021_ (_04030_, _04029_, _06678_);
  not _27022_ (_04031_, _06678_);
  or _27023_ (_04032_, _00717_, _04031_);
  and _27024_ (_04033_, _04032_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or _27025_ (_04034_, _04033_, _06946_);
  or _27026_ (_04035_, _04034_, _04030_);
  nand _27027_ (_04036_, _11589_, _06946_);
  and _27028_ (_04037_, _04036_, _06444_);
  and _27029_ (_04548_, _04037_, _04035_);
  and _27030_ (_04038_, _06678_, _06432_);
  nand _27031_ (_04039_, _04038_, _06930_);
  or _27032_ (_04040_, _04038_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  and _27033_ (_04041_, _04040_, _04039_);
  or _27034_ (_04042_, _04041_, _02406_);
  nand _27035_ (_04043_, _07069_, _06946_);
  and _27036_ (_04044_, _04043_, _06444_);
  and _27037_ (_04551_, _04044_, _04042_);
  and _27038_ (_04045_, _06678_, _06942_);
  nand _27039_ (_04046_, _04045_, _06930_);
  or _27040_ (_04047_, _04045_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and _27041_ (_04048_, _04047_, _04046_);
  or _27042_ (_04049_, _04048_, _02406_);
  nand _27043_ (_04051_, _09526_, _06946_);
  and _27044_ (_04053_, _04051_, _06444_);
  and _27045_ (_04555_, _04053_, _04049_);
  not _27046_ (_04054_, _14174_);
  and _27047_ (_04557_, _14496_, _04054_);
  nor _27048_ (_04055_, _08484_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor _27049_ (_04056_, _04055_, _12589_);
  or _27050_ (_04058_, _04056_, _12023_);
  and _27051_ (_04059_, _12048_, _08230_);
  and _27052_ (_04060_, _11452_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor _27053_ (_04061_, _12128_, _12033_);
  and _27054_ (_04062_, _12054_, _11650_);
  or _27055_ (_04063_, _04062_, _04061_);
  or _27056_ (_04064_, _04063_, _04060_);
  or _27057_ (_04065_, _12207_, _12205_);
  and _27058_ (_04066_, _04065_, _12208_);
  and _27059_ (_04067_, _04066_, _12218_);
  or _27060_ (_04068_, _04067_, _04064_);
  nor _27061_ (_04069_, _04068_, _04059_);
  nand _27062_ (_04070_, _04069_, _12023_);
  and _27063_ (_04071_, _04070_, _06444_);
  and _27064_ (_04562_, _04071_, _04058_);
  or _27065_ (_04072_, _12023_, _08486_);
  and _27066_ (_04073_, _12048_, _08308_);
  and _27067_ (_04075_, _11452_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor _27068_ (_04076_, _12154_, _12033_);
  and _27069_ (_04077_, _12054_, _11689_);
  or _27070_ (_04078_, _04077_, _04076_);
  or _27071_ (_04079_, _04078_, _04075_);
  or _27072_ (_04080_, _12157_, _12158_);
  not _27073_ (_04081_, _04080_);
  nand _27074_ (_04082_, _04081_, _12203_);
  or _27075_ (_04083_, _04081_, _12203_);
  and _27076_ (_04084_, _04083_, _12606_);
  and _27077_ (_04085_, _04084_, _04082_);
  or _27078_ (_04086_, _04085_, _04079_);
  nor _27079_ (_04087_, _04086_, _04073_);
  nand _27080_ (_04089_, _04087_, _12023_);
  and _27081_ (_04090_, _04089_, _06444_);
  and _27082_ (_04564_, _04090_, _04072_);
  and _27083_ (_04091_, _08064_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor _27084_ (_04092_, _08064_, _01106_);
  or _27085_ (_04093_, _04092_, _04091_);
  and _27086_ (_04566_, _04093_, _06444_);
  and _27087_ (_04096_, _03977_, _07378_);
  or _27088_ (_04097_, _03404_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  or _27089_ (_04098_, _00936_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  nand _27090_ (_04099_, _04098_, _04097_);
  nor _27091_ (_04100_, _04099_, _06442_);
  and _27092_ (_04101_, _03410_, _07359_);
  or _27093_ (_04102_, _04101_, _04100_);
  or _27094_ (_04103_, _04102_, _04096_);
  and _27095_ (_04573_, _04103_, _06444_);
  and _27096_ (_04104_, _12048_, _02977_);
  and _27097_ (_04106_, _11452_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and _27098_ (_04107_, _12032_, _12162_);
  and _27099_ (_04108_, _12054_, _11905_);
  or _27100_ (_04110_, _04108_, _04107_);
  or _27101_ (_04111_, _04110_, _04106_);
  nor _27102_ (_04112_, _12201_, _12199_);
  nor _27103_ (_04114_, _04112_, _12202_);
  and _27104_ (_04115_, _04114_, _12218_);
  or _27105_ (_04116_, _04115_, _04111_);
  or _27106_ (_04117_, _04116_, _04104_);
  and _27107_ (_04118_, _04117_, _12023_);
  and _27108_ (_04119_, _03274_, _08499_);
  or _27109_ (_04120_, _04119_, _04118_);
  and _27110_ (_04576_, _04120_, _06444_);
  and _27111_ (_04121_, _03977_, _07359_);
  or _27112_ (_04122_, _00936_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  or _27113_ (_04124_, _03404_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  nand _27114_ (_04125_, _04124_, _04122_);
  nor _27115_ (_04127_, _04125_, _06442_);
  and _27116_ (_04128_, _03410_, _07340_);
  or _27117_ (_04129_, _04128_, _04127_);
  or _27118_ (_04130_, _04129_, _04121_);
  and _27119_ (_04580_, _04130_, _06444_);
  not _27120_ (_04132_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  nor _27121_ (_04133_, _00856_, _04132_);
  and _27122_ (_04134_, _12054_, _11794_);
  and _27123_ (_04135_, _12186_, _12032_);
  or _27124_ (_04136_, _04135_, _04134_);
  or _27125_ (_04137_, _12196_, _12194_);
  and _27126_ (_04138_, _12606_, _12198_);
  and _27127_ (_04139_, _04138_, _04137_);
  or _27128_ (_04140_, _04139_, _04136_);
  and _27129_ (_04141_, _12048_, _07959_);
  or _27130_ (_04142_, _04141_, _04140_);
  and _27131_ (_04143_, _04142_, _12023_);
  or _27132_ (_04144_, _04143_, _04133_);
  and _27133_ (_04582_, _04144_, _06444_);
  and _27134_ (_04145_, _07046_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  nor _27135_ (_04146_, _07046_, _06978_);
  or _27136_ (_04147_, _04146_, _04145_);
  and _27137_ (_04587_, _04147_, _06444_);
  or _27138_ (_04148_, _03404_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  or _27139_ (_04149_, _00936_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  nand _27140_ (_04150_, _04149_, _04148_);
  nor _27141_ (_04151_, _04150_, _06442_);
  and _27142_ (_04152_, _03410_, _11882_);
  or _27143_ (_04153_, _04152_, _04151_);
  and _27144_ (_04154_, _13865_, _06295_);
  and _27145_ (_04155_, _04154_, _07340_);
  or _27146_ (_04156_, _04155_, _04153_);
  and _27147_ (_04590_, _04156_, _06444_);
  and _27148_ (_04157_, _07403_, _07402_);
  nand _27149_ (_04158_, _04157_, _08310_);
  nor _27150_ (_04159_, _04158_, _06930_);
  and _27151_ (_04160_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  nand _27152_ (_04161_, _07387_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  nor _27153_ (_04162_, _07396_, _07076_);
  not _27154_ (_04163_, _04162_);
  or _27155_ (_04164_, _04163_, _07392_);
  or _27156_ (_04165_, _04164_, _04161_);
  and _27157_ (_04166_, _04165_, _04160_);
  and _27158_ (_04167_, _04166_, _04158_);
  or _27159_ (_04168_, _04167_, _07407_);
  or _27160_ (_04169_, _04168_, _04159_);
  nand _27161_ (_04170_, _07407_, _07300_);
  and _27162_ (_04171_, _04170_, _06444_);
  and _27163_ (_04592_, _04171_, _04169_);
  and _27164_ (_04172_, _07011_, _07004_);
  nor _27165_ (_04173_, _04172_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or _27166_ (_04174_, _04173_, _07024_);
  nor _27167_ (_04175_, _07028_, _02860_);
  nand _27168_ (_04176_, _04175_, _07026_);
  and _27169_ (_04177_, _04176_, _04174_);
  nor _27170_ (_04178_, _04177_, _07017_);
  and _27171_ (_04179_, _07017_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  or _27172_ (_04180_, _04179_, _06985_);
  or _27173_ (_04181_, _04180_, _04178_);
  or _27174_ (_04182_, _02538_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  and _27175_ (_04183_, _04182_, _09503_);
  and _27176_ (_04184_, _04183_, _04181_);
  nor _27177_ (_04185_, _10494_, _09503_);
  or _27178_ (_04186_, _04185_, _04184_);
  and _27179_ (_04595_, _04186_, _06444_);
  and _27180_ (_04187_, _07029_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and _27181_ (_04188_, _04187_, _07026_);
  nand _27182_ (_04189_, _07011_, _07003_);
  and _27183_ (_04190_, _04189_, _02887_);
  nor _27184_ (_04191_, _04190_, _04172_);
  or _27185_ (_04193_, _04191_, _07017_);
  or _27186_ (_04194_, _04193_, _04188_);
  or _27187_ (_04196_, _07035_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and _27188_ (_04197_, _04196_, _06990_);
  and _27189_ (_04198_, _04197_, _04194_);
  nor _27190_ (_04199_, _09503_, _06666_);
  and _27191_ (_04200_, _06985_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or _27192_ (_04201_, _04200_, _04199_);
  or _27193_ (_04202_, _04201_, _04198_);
  and _27194_ (_04597_, _04202_, _06444_);
  or _27195_ (_04205_, _04162_, _07392_);
  or _27196_ (_04207_, _04205_, _04161_);
  nand _27197_ (_04209_, _04207_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  nand _27198_ (_04211_, _04209_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and _27199_ (_04212_, _14511_, _06674_);
  or _27200_ (_04213_, _04212_, _04211_);
  and _27201_ (_04215_, _04213_, _07408_);
  nand _27202_ (_04216_, _04212_, _06930_);
  and _27203_ (_04217_, _04216_, _04215_);
  nor _27204_ (_04219_, _07408_, _07069_);
  or _27205_ (_04221_, _04219_, _04217_);
  and _27206_ (_04803_, _04221_, _06444_);
  nand _27207_ (_04806_, _11857_, _06444_);
  nand _27208_ (_04808_, _11802_, _06444_);
  nand _27209_ (_04810_, _11912_, _06444_);
  nor _27210_ (_04812_, _11699_, rst);
  nor _27211_ (_04814_, _11663_, rst);
  nor _27212_ (_04822_, _11734_, rst);
  nor _27213_ (_04824_, _11774_, rst);
  nor _27214_ (_04223_, _01701_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff );
  or _27215_ (_04224_, _04164_, _07388_);
  and _27216_ (_04225_, _04224_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or _27217_ (_04227_, _04225_, _04223_);
  and _27218_ (_04228_, _04157_, _06987_);
  or _27219_ (_04229_, _04228_, _04227_);
  and _27220_ (_04230_, _04229_, _07408_);
  nand _27221_ (_04231_, _04228_, _06930_);
  and _27222_ (_04232_, _04231_, _04230_);
  nor _27223_ (_04233_, _07408_, _06666_);
  or _27224_ (_04234_, _04233_, _04232_);
  and _27225_ (_04826_, _04234_, _06444_);
  and _27226_ (_04235_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and _27227_ (_04236_, _04235_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and _27228_ (_04237_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  and _27229_ (_04238_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  and _27230_ (_04239_, _04238_, _04237_);
  and _27231_ (_04240_, _04239_, _04236_);
  and _27232_ (_04241_, _04240_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  and _27233_ (_04242_, _04241_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  and _27234_ (_04243_, _04242_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  and _27235_ (_04244_, _04243_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  and _27236_ (_04245_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  and _27237_ (_04246_, _04245_, _04244_);
  and _27238_ (_04247_, _04246_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor _27239_ (_04248_, _04246_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor _27240_ (_04249_, _04248_, _04247_);
  nor _27241_ (_04250_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  not _27242_ (_04251_, _04250_);
  and _27243_ (_04252_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and _27244_ (_04253_, _04252_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor _27245_ (_04254_, _04252_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor _27246_ (_04255_, _04254_, _04253_);
  not _27247_ (_04256_, _04255_);
  and _27248_ (_04257_, _04253_, _01279_);
  nor _27249_ (_04258_, _04253_, _01279_);
  nor _27250_ (_04259_, _04258_, _04257_);
  nor _27251_ (_04260_, _04259_, _08481_);
  and _27252_ (_04261_, _04259_, \oc8051_symbolic_cxrom1.regvalid [5]);
  nor _27253_ (_04262_, _04261_, _04260_);
  nor _27254_ (_04263_, _04262_, _04256_);
  and _27255_ (_04264_, _04259_, \oc8051_symbolic_cxrom1.regvalid [1]);
  nor _27256_ (_04265_, _04259_, _08521_);
  nor _27257_ (_04266_, _04265_, _04264_);
  nor _27258_ (_04267_, _04266_, _04255_);
  nor _27259_ (_04268_, _04267_, _04263_);
  nor _27260_ (_04269_, _04268_, _04251_);
  and _27261_ (_04270_, _13796_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  not _27262_ (_04271_, _04270_);
  nor _27263_ (_04272_, _04259_, _08515_);
  and _27264_ (_04273_, _04259_, \oc8051_symbolic_cxrom1.regvalid [7]);
  nor _27265_ (_04274_, _04273_, _04272_);
  nor _27266_ (_04275_, _04274_, _04256_);
  and _27267_ (_04276_, _04259_, \oc8051_symbolic_cxrom1.regvalid [3]);
  not _27268_ (_04277_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor _27269_ (_04278_, _04259_, _04277_);
  nor _27270_ (_04279_, _04278_, _04276_);
  nor _27271_ (_04280_, _04279_, _04255_);
  nor _27272_ (_04281_, _04280_, _04275_);
  nor _27273_ (_04282_, _04281_, _04271_);
  nor _27274_ (_04283_, _04282_, _04269_);
  and _27275_ (_04284_, _04259_, \oc8051_symbolic_cxrom1.regvalid [4]);
  not _27276_ (_04285_, \oc8051_symbolic_cxrom1.regvalid [12]);
  nor _27277_ (_04286_, _04259_, _04285_);
  nor _27278_ (_04287_, _04286_, _04284_);
  nor _27279_ (_04288_, _04287_, _04256_);
  and _27280_ (_04289_, _04259_, \oc8051_symbolic_cxrom1.regvalid [0]);
  not _27281_ (_04290_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor _27282_ (_04291_, _04259_, _04290_);
  nor _27283_ (_04292_, _04291_, _04289_);
  nor _27284_ (_04293_, _04292_, _01154_);
  or _27285_ (_04294_, _04293_, _04288_);
  and _27286_ (_04295_, _04294_, _04252_);
  and _27287_ (_04296_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _12846_);
  not _27288_ (_04297_, _04296_);
  nor _27289_ (_04298_, _04259_, _08546_);
  and _27290_ (_04299_, _04259_, \oc8051_symbolic_cxrom1.regvalid [6]);
  nor _27291_ (_04300_, _04299_, _04298_);
  nor _27292_ (_04301_, _04300_, _04256_);
  and _27293_ (_04302_, _04259_, \oc8051_symbolic_cxrom1.regvalid [2]);
  nor _27294_ (_04303_, _04259_, _09302_);
  nor _27295_ (_04304_, _04303_, _04302_);
  nor _27296_ (_04305_, _04304_, _04255_);
  nor _27297_ (_04306_, _04305_, _04301_);
  nor _27298_ (_04307_, _04306_, _04297_);
  nor _27299_ (_04308_, _04307_, _04295_);
  and _27300_ (_04309_, _04308_, _04283_);
  and _27301_ (_04310_, _04296_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  and _27302_ (_04311_, _04252_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  nor _27303_ (_04312_, _04311_, _04310_);
  and _27304_ (_04314_, _04270_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  and _27305_ (_04315_, _04250_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  nor _27306_ (_04316_, _04315_, _04314_);
  and _27307_ (_04317_, _04316_, _04312_);
  and _27308_ (_04318_, _04317_, _04256_);
  not _27309_ (_04319_, _04259_);
  and _27310_ (_04320_, _04270_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  and _27311_ (_04321_, _04250_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  nor _27312_ (_04322_, _04321_, _04320_);
  and _27313_ (_04323_, _04296_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  and _27314_ (_04324_, _04252_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  nor _27315_ (_04325_, _04324_, _04323_);
  and _27316_ (_04326_, _04325_, _04322_);
  and _27317_ (_04327_, _04326_, _04255_);
  or _27318_ (_04328_, _04327_, _04319_);
  nor _27319_ (_04329_, _04328_, _04318_);
  and _27320_ (_04330_, _04296_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  and _27321_ (_04331_, _04270_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  nor _27322_ (_04332_, _04331_, _04330_);
  and _27323_ (_04333_, _04250_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  and _27324_ (_04334_, _04252_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  nor _27325_ (_04335_, _04334_, _04333_);
  and _27326_ (_04336_, _04335_, _04332_);
  and _27327_ (_04337_, _04336_, _04256_);
  and _27328_ (_04338_, _04296_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  and _27329_ (_04339_, _04252_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  nor _27330_ (_04340_, _04339_, _04338_);
  and _27331_ (_04341_, _04270_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  and _27332_ (_04342_, _04250_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  nor _27333_ (_04343_, _04342_, _04341_);
  and _27334_ (_04344_, _04343_, _04340_);
  and _27335_ (_04345_, _04344_, _04255_);
  or _27336_ (_04346_, _04345_, _04259_);
  nor _27337_ (_04347_, _04346_, _04337_);
  nor _27338_ (_04348_, _04347_, _04329_);
  nor _27339_ (_04349_, _04348_, _04309_);
  and _27340_ (_04350_, _04349_, _04249_);
  nor _27341_ (_04351_, _04349_, _04249_);
  nor _27342_ (_04352_, _04351_, _04350_);
  and _27343_ (_04353_, _04244_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor _27344_ (_04354_, _04353_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  nor _27345_ (_04355_, _04354_, _04246_);
  and _27346_ (_04356_, _04355_, _04349_);
  nor _27347_ (_04357_, _04355_, _04349_);
  nor _27348_ (_04358_, _04244_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor _27349_ (_04359_, _04358_, _04353_);
  and _27350_ (_04360_, _04359_, _04349_);
  nor _27351_ (_04361_, _04243_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  nor _27352_ (_04363_, _04361_, _04244_);
  and _27353_ (_04365_, _04363_, _04349_);
  nor _27354_ (_04367_, _04242_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  nor _27355_ (_04368_, _04367_, _04243_);
  and _27356_ (_04370_, _04368_, _04349_);
  nor _27357_ (_04371_, _04363_, _04349_);
  nor _27358_ (_04372_, _04371_, _04365_);
  nor _27359_ (_04373_, _04368_, _04349_);
  nor _27360_ (_04374_, _04373_, _04370_);
  not _27361_ (_04375_, _04374_);
  nor _27362_ (_04376_, _04241_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  nor _27363_ (_04378_, _04376_, _04242_);
  and _27364_ (_04380_, _04378_, _04349_);
  nor _27365_ (_04381_, _04378_, _04349_);
  nor _27366_ (_04382_, _04240_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor _27367_ (_04384_, _04382_, _04241_);
  and _27368_ (_04385_, _04384_, _04349_);
  and _27369_ (_04386_, _04237_, _04236_);
  and _27370_ (_04387_, _04386_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nor _27371_ (_04388_, _04387_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  nor _27372_ (_04389_, _04388_, _04240_);
  and _27373_ (_04390_, _04389_, _04349_);
  nor _27374_ (_04391_, _04389_, _04349_);
  nor _27375_ (_04392_, _04386_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nor _27376_ (_04393_, _04392_, _04387_);
  and _27377_ (_04394_, _04296_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  and _27378_ (_04395_, _04252_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  nor _27379_ (_04396_, _04395_, _04394_);
  and _27380_ (_04397_, _04270_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  and _27381_ (_04398_, _04250_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  nor _27382_ (_04399_, _04398_, _04397_);
  and _27383_ (_04400_, _04399_, _04396_);
  and _27384_ (_04401_, _04400_, _04256_);
  and _27385_ (_04402_, _04270_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  and _27386_ (_04403_, _04250_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  nor _27387_ (_04404_, _04403_, _04402_);
  and _27388_ (_04405_, _04296_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  and _27389_ (_04406_, _04252_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  nor _27390_ (_04407_, _04406_, _04405_);
  and _27391_ (_04408_, _04407_, _04404_);
  and _27392_ (_04409_, _04408_, _04255_);
  or _27393_ (_04410_, _04409_, _04259_);
  nor _27394_ (_04411_, _04410_, _04401_);
  and _27395_ (_04412_, _04270_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  and _27396_ (_04413_, _04296_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  nor _27397_ (_04414_, _04413_, _04412_);
  and _27398_ (_04415_, _04250_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  and _27399_ (_04416_, _04252_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  nor _27400_ (_04417_, _04416_, _04415_);
  and _27401_ (_04418_, _04417_, _04414_);
  nor _27402_ (_04419_, _04418_, _04255_);
  and _27403_ (_04420_, _04296_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  and _27404_ (_04421_, _04252_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  nor _27405_ (_04422_, _04421_, _04420_);
  and _27406_ (_04423_, _04270_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  and _27407_ (_04424_, _04250_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  nor _27408_ (_04425_, _04424_, _04423_);
  and _27409_ (_04426_, _04425_, _04422_);
  nor _27410_ (_04427_, _04426_, _04256_);
  or _27411_ (_04428_, _04427_, _04419_);
  and _27412_ (_04429_, _04428_, _04259_);
  nor _27413_ (_04430_, _04429_, _04411_);
  nor _27414_ (_04431_, _04430_, _04309_);
  and _27415_ (_04432_, _04431_, _04393_);
  nor _27416_ (_04433_, _04431_, _04393_);
  nor _27417_ (_04434_, _04433_, _04432_);
  not _27418_ (_04435_, _04434_);
  and _27419_ (_04436_, _04236_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nor _27420_ (_04437_, _04436_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  nor _27421_ (_04438_, _04437_, _04386_);
  and _27422_ (_04439_, _04296_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  and _27423_ (_04440_, _04252_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  nor _27424_ (_04441_, _04440_, _04439_);
  and _27425_ (_04442_, _04270_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  and _27426_ (_04443_, _04250_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  nor _27427_ (_04444_, _04443_, _04442_);
  and _27428_ (_04445_, _04444_, _04441_);
  and _27429_ (_04446_, _04445_, _04256_);
  and _27430_ (_04447_, _04296_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  and _27431_ (_04448_, _04252_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  nor _27432_ (_04449_, _04448_, _04447_);
  and _27433_ (_04450_, _04270_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  and _27434_ (_04451_, _04250_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  nor _27435_ (_04452_, _04451_, _04450_);
  and _27436_ (_04453_, _04452_, _04449_);
  and _27437_ (_04454_, _04453_, _04255_);
  or _27438_ (_04455_, _04454_, _04259_);
  nor _27439_ (_04456_, _04455_, _04446_);
  and _27440_ (_04457_, _04270_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  and _27441_ (_04458_, _04296_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  nor _27442_ (_04459_, _04458_, _04457_);
  and _27443_ (_04460_, _04250_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  and _27444_ (_04461_, _04252_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  nor _27445_ (_04462_, _04461_, _04460_);
  and _27446_ (_04463_, _04462_, _04459_);
  nor _27447_ (_04464_, _04463_, _04255_);
  and _27448_ (_04465_, _04296_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  and _27449_ (_04466_, _04252_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  nor _27450_ (_04467_, _04466_, _04465_);
  and _27451_ (_04468_, _04270_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  and _27452_ (_04469_, _04250_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  nor _27453_ (_04470_, _04469_, _04468_);
  and _27454_ (_04471_, _04470_, _04467_);
  nor _27455_ (_04472_, _04471_, _04256_);
  or _27456_ (_04473_, _04472_, _04464_);
  and _27457_ (_04474_, _04473_, _04259_);
  nor _27458_ (_04475_, _04474_, _04456_);
  nor _27459_ (_04476_, _04475_, _04309_);
  and _27460_ (_04477_, _04476_, _04438_);
  nor _27461_ (_04478_, _04476_, _04438_);
  nor _27462_ (_04479_, _04478_, _04477_);
  not _27463_ (_04480_, _04479_);
  nor _27464_ (_04481_, _04236_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nor _27465_ (_04482_, _04481_, _04436_);
  and _27466_ (_04483_, _04296_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  and _27467_ (_04484_, _04252_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  nor _27468_ (_04485_, _04484_, _04483_);
  and _27469_ (_04486_, _04270_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  and _27470_ (_04487_, _04250_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  nor _27471_ (_04488_, _04487_, _04486_);
  and _27472_ (_04489_, _04488_, _04485_);
  and _27473_ (_04490_, _04489_, _04256_);
  and _27474_ (_04492_, _04296_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  and _27475_ (_04493_, _04252_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  nor _27476_ (_04494_, _04493_, _04492_);
  and _27477_ (_04495_, _04270_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  and _27478_ (_04496_, _04250_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  nor _27479_ (_04497_, _04496_, _04495_);
  and _27480_ (_04498_, _04497_, _04494_);
  and _27481_ (_04499_, _04498_, _04255_);
  or _27482_ (_04500_, _04499_, _04319_);
  nor _27483_ (_04501_, _04500_, _04490_);
  and _27484_ (_04502_, _04296_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  and _27485_ (_04503_, _04270_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  nor _27486_ (_04504_, _04503_, _04502_);
  and _27487_ (_04505_, _04250_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  and _27488_ (_04506_, _04252_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  nor _27489_ (_04507_, _04506_, _04505_);
  and _27490_ (_04508_, _04507_, _04504_);
  and _27491_ (_04509_, _04508_, _04256_);
  and _27492_ (_04510_, _04296_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  and _27493_ (_04511_, _04252_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  nor _27494_ (_04512_, _04511_, _04510_);
  and _27495_ (_04513_, _04270_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  and _27496_ (_04514_, _04250_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  nor _27497_ (_04515_, _04514_, _04513_);
  and _27498_ (_04516_, _04515_, _04512_);
  and _27499_ (_04517_, _04516_, _04255_);
  or _27500_ (_04518_, _04517_, _04259_);
  nor _27501_ (_04519_, _04518_, _04509_);
  nor _27502_ (_04520_, _04519_, _04501_);
  nor _27503_ (_04521_, _04520_, _04309_);
  and _27504_ (_04522_, _04521_, _04482_);
  and _27505_ (_04523_, _04235_, _01279_);
  nor _27506_ (_04524_, _04235_, _01279_);
  nor _27507_ (_04525_, _04524_, _04523_);
  not _27508_ (_04526_, _04525_);
  and _27509_ (_04527_, _04296_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  and _27510_ (_04528_, _04252_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  nor _27511_ (_04529_, _04528_, _04527_);
  and _27512_ (_04531_, _04270_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  and _27513_ (_04532_, _04250_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  nor _27514_ (_04534_, _04532_, _04531_);
  and _27515_ (_04536_, _04534_, _04529_);
  and _27516_ (_04537_, _04536_, _04256_);
  and _27517_ (_04539_, _04270_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  and _27518_ (_04540_, _04250_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  nor _27519_ (_04541_, _04540_, _04539_);
  and _27520_ (_04542_, _04296_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  and _27521_ (_04543_, _04252_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  nor _27522_ (_04544_, _04543_, _04542_);
  and _27523_ (_04546_, _04544_, _04541_);
  and _27524_ (_04547_, _04546_, _04255_);
  or _27525_ (_04549_, _04547_, _04319_);
  nor _27526_ (_04550_, _04549_, _04537_);
  and _27527_ (_04552_, _04296_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  and _27528_ (_04553_, _04270_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  nor _27529_ (_04554_, _04553_, _04552_);
  and _27530_ (_04556_, _04250_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  and _27531_ (_04558_, _04252_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  nor _27532_ (_04559_, _04558_, _04556_);
  and _27533_ (_04560_, _04559_, _04554_);
  and _27534_ (_04561_, _04560_, _04256_);
  and _27535_ (_04563_, _04296_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  and _27536_ (_04565_, _04252_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  nor _27537_ (_04567_, _04565_, _04563_);
  and _27538_ (_04568_, _04270_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  and _27539_ (_04569_, _04250_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  nor _27540_ (_04570_, _04569_, _04568_);
  and _27541_ (_04571_, _04570_, _04567_);
  and _27542_ (_04572_, _04571_, _04255_);
  or _27543_ (_04574_, _04572_, _04259_);
  nor _27544_ (_04575_, _04574_, _04561_);
  nor _27545_ (_04577_, _04575_, _04550_);
  nor _27546_ (_04578_, _04577_, _04309_);
  and _27547_ (_04579_, _04578_, _04526_);
  nor _27548_ (_04581_, _04578_, _04526_);
  nor _27549_ (_04583_, _04581_, _04579_);
  not _27550_ (_04584_, _04583_);
  and _27551_ (_04585_, _12846_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and _27552_ (_04586_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _01154_);
  nor _27553_ (_04588_, _04586_, _04585_);
  not _27554_ (_04589_, _04588_);
  and _27555_ (_04591_, _04296_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  and _27556_ (_04593_, _04252_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  nor _27557_ (_04594_, _04593_, _04591_);
  and _27558_ (_04596_, _04270_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  and _27559_ (_04598_, _04250_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  nor _27560_ (_04599_, _04598_, _04596_);
  and _27561_ (_04600_, _04599_, _04594_);
  and _27562_ (_04601_, _04600_, _04256_);
  and _27563_ (_04602_, _04296_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  and _27564_ (_04603_, _04252_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  nor _27565_ (_04604_, _04603_, _04602_);
  and _27566_ (_04605_, _04270_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  and _27567_ (_04606_, _04250_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  nor _27568_ (_04607_, _04606_, _04605_);
  and _27569_ (_04608_, _04607_, _04604_);
  and _27570_ (_04609_, _04608_, _04255_);
  or _27571_ (_04610_, _04609_, _04319_);
  nor _27572_ (_04611_, _04610_, _04601_);
  and _27573_ (_04612_, _04296_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  and _27574_ (_04613_, _04270_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  nor _27575_ (_04614_, _04613_, _04612_);
  and _27576_ (_04615_, _04250_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  and _27577_ (_04616_, _04252_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  nor _27578_ (_04617_, _04616_, _04615_);
  and _27579_ (_04618_, _04617_, _04614_);
  and _27580_ (_04619_, _04618_, _04256_);
  and _27581_ (_04620_, _04296_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  and _27582_ (_04621_, _04252_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  nor _27583_ (_04622_, _04621_, _04620_);
  and _27584_ (_04623_, _04270_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  and _27585_ (_04624_, _04250_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  nor _27586_ (_04625_, _04624_, _04623_);
  and _27587_ (_04626_, _04625_, _04622_);
  and _27588_ (_04627_, _04626_, _04255_);
  or _27589_ (_04628_, _04627_, _04259_);
  nor _27590_ (_04629_, _04628_, _04619_);
  nor _27591_ (_04630_, _04629_, _04611_);
  nor _27592_ (_04631_, _04630_, _04309_);
  and _27593_ (_04632_, _04631_, _04589_);
  and _27594_ (_04633_, _04296_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  and _27595_ (_04634_, _04270_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  nor _27596_ (_04635_, _04634_, _04633_);
  and _27597_ (_04636_, _04250_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  and _27598_ (_04637_, _04252_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  nor _27599_ (_04638_, _04637_, _04636_);
  and _27600_ (_04639_, _04638_, _04635_);
  and _27601_ (_04640_, _04639_, _04256_);
  and _27602_ (_04641_, _04296_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  and _27603_ (_04642_, _04252_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  nor _27604_ (_04643_, _04642_, _04641_);
  and _27605_ (_04644_, _04270_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  and _27606_ (_04645_, _04250_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  nor _27607_ (_04646_, _04645_, _04644_);
  and _27608_ (_04647_, _04646_, _04643_);
  and _27609_ (_04648_, _04647_, _04255_);
  or _27610_ (_04649_, _04648_, _04319_);
  nor _27611_ (_04650_, _04649_, _04640_);
  and _27612_ (_04651_, _04296_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  and _27613_ (_04652_, _04270_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  nor _27614_ (_04653_, _04652_, _04651_);
  and _27615_ (_04654_, _04250_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  and _27616_ (_04655_, _04252_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  nor _27617_ (_04656_, _04655_, _04654_);
  and _27618_ (_04657_, _04656_, _04653_);
  and _27619_ (_04658_, _04657_, _04256_);
  and _27620_ (_04659_, _04270_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  and _27621_ (_04660_, _04250_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  nor _27622_ (_04661_, _04660_, _04659_);
  and _27623_ (_04662_, _04296_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  and _27624_ (_04663_, _04252_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  nor _27625_ (_04664_, _04663_, _04662_);
  and _27626_ (_04665_, _04664_, _04661_);
  and _27627_ (_04666_, _04665_, _04255_);
  or _27628_ (_04667_, _04666_, _04259_);
  nor _27629_ (_04668_, _04667_, _04658_);
  nor _27630_ (_04669_, _04668_, _04650_);
  nor _27631_ (_04670_, _04669_, _04309_);
  and _27632_ (_04671_, _04670_, _12846_);
  and _27633_ (_04672_, _04296_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  and _27634_ (_04673_, _04252_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  nor _27635_ (_04674_, _04673_, _04672_);
  and _27636_ (_04675_, _04270_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  and _27637_ (_04676_, _04250_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  nor _27638_ (_04677_, _04676_, _04675_);
  and _27639_ (_04678_, _04677_, _04674_);
  and _27640_ (_04679_, _04678_, _04256_);
  and _27641_ (_04680_, _04270_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  and _27642_ (_04681_, _04250_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  nor _27643_ (_04682_, _04681_, _04680_);
  and _27644_ (_04683_, _04296_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  and _27645_ (_04684_, _04252_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  nor _27646_ (_04685_, _04684_, _04683_);
  and _27647_ (_04686_, _04685_, _04682_);
  and _27648_ (_04687_, _04686_, _04255_);
  or _27649_ (_04688_, _04687_, _04319_);
  nor _27650_ (_04689_, _04688_, _04679_);
  and _27651_ (_04690_, _04296_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and _27652_ (_04691_, _04252_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  nor _27653_ (_04692_, _04691_, _04690_);
  and _27654_ (_04693_, _04270_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and _27655_ (_04694_, _04250_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  nor _27656_ (_04695_, _04694_, _04693_);
  and _27657_ (_04696_, _04695_, _04692_);
  nor _27658_ (_04697_, _04696_, _04255_);
  and _27659_ (_04698_, _04270_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  and _27660_ (_04699_, _04250_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  nor _27661_ (_04700_, _04699_, _04698_);
  and _27662_ (_04701_, _04296_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and _27663_ (_04702_, _04252_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  nor _27664_ (_04703_, _04702_, _04701_);
  and _27665_ (_04704_, _04703_, _04700_);
  nor _27666_ (_04705_, _04704_, _04256_);
  or _27667_ (_04706_, _04705_, _04697_);
  and _27668_ (_04707_, _04706_, _04319_);
  nor _27669_ (_04708_, _04707_, _04689_);
  nor _27670_ (_04709_, _04708_, _04309_);
  and _27671_ (_04710_, _04709_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _27672_ (_04711_, _04670_, _12846_);
  nor _27673_ (_04712_, _04711_, _04671_);
  and _27674_ (_04713_, _04712_, _04710_);
  nor _27675_ (_04714_, _04713_, _04671_);
  nor _27676_ (_04715_, _04631_, _04589_);
  nor _27677_ (_04716_, _04715_, _04632_);
  not _27678_ (_04717_, _04716_);
  nor _27679_ (_04718_, _04717_, _04714_);
  nor _27680_ (_04719_, _04718_, _04632_);
  nor _27681_ (_04720_, _04719_, _04584_);
  nor _27682_ (_04721_, _04720_, _04579_);
  nor _27683_ (_04722_, _04521_, _04482_);
  nor _27684_ (_04723_, _04722_, _04522_);
  not _27685_ (_04724_, _04723_);
  nor _27686_ (_04725_, _04724_, _04721_);
  nor _27687_ (_04726_, _04725_, _04522_);
  nor _27688_ (_04727_, _04726_, _04480_);
  nor _27689_ (_04728_, _04727_, _04477_);
  nor _27690_ (_04729_, _04728_, _04435_);
  nor _27691_ (_04730_, _04729_, _04432_);
  nor _27692_ (_04731_, _04730_, _04391_);
  or _27693_ (_04732_, _04731_, _04390_);
  nor _27694_ (_04733_, _04384_, _04349_);
  nor _27695_ (_04734_, _04733_, _04385_);
  and _27696_ (_04735_, _04734_, _04732_);
  nor _27697_ (_04736_, _04735_, _04385_);
  nor _27698_ (_04737_, _04736_, _04381_);
  nor _27699_ (_04738_, _04737_, _04380_);
  nor _27700_ (_04739_, _04738_, _04375_);
  and _27701_ (_04740_, _04739_, _04372_);
  or _27702_ (_04741_, _04740_, _04370_);
  nor _27703_ (_04742_, _04741_, _04365_);
  nor _27704_ (_04743_, _04359_, _04349_);
  nor _27705_ (_04744_, _04743_, _04360_);
  not _27706_ (_04745_, _04744_);
  nor _27707_ (_04746_, _04745_, _04742_);
  nor _27708_ (_04747_, _04746_, _04360_);
  nor _27709_ (_04748_, _04747_, _04357_);
  or _27710_ (_04749_, _04748_, _04356_);
  and _27711_ (_04750_, _04749_, _04352_);
  nor _27712_ (_04751_, _04750_, _04350_);
  nor _27713_ (_04752_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  and _27714_ (_04753_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  nor _27715_ (_04754_, _04753_, _04752_);
  nor _27716_ (_04755_, _04754_, _04247_);
  and _27717_ (_04756_, _04754_, _04247_);
  nor _27718_ (_04757_, _04756_, _04755_);
  nor _27719_ (_04758_, _04757_, _04349_);
  and _27720_ (_04759_, _04757_, _04349_);
  nor _27721_ (_04760_, _04759_, _04758_);
  nor _27722_ (_04761_, _04760_, _04751_);
  and _27723_ (_04762_, _04745_, _04742_);
  nor _27724_ (_04763_, _04762_, _04746_);
  nor _27725_ (_04764_, _04763_, _00664_);
  nor _27726_ (_04765_, _04739_, _04370_);
  nand _27727_ (_04766_, _04372_, _01602_);
  or _27728_ (_04767_, _04372_, _01602_);
  and _27729_ (_04768_, _04767_, _04766_);
  not _27730_ (_04769_, _04768_);
  nor _27731_ (_04770_, _04769_, _04765_);
  not _27732_ (_04771_, _04349_);
  nor _27733_ (_04772_, _04378_, _01150_);
  and _27734_ (_04773_, _04378_, _01150_);
  or _27735_ (_04774_, _04773_, _04772_);
  nand _27736_ (_04775_, _04774_, _04771_);
  or _27737_ (_04776_, _04774_, _04771_);
  and _27738_ (_04777_, _04776_, _04775_);
  or _27739_ (_04778_, _04777_, _04736_);
  nand _27740_ (_04779_, _04777_, _04736_);
  and _27741_ (_04780_, _04779_, _04778_);
  nor _27742_ (_04781_, _04734_, _04732_);
  nor _27743_ (_04782_, _04781_, _04735_);
  nor _27744_ (_04783_, _04782_, _01872_);
  and _27745_ (_04784_, _04782_, _01872_);
  nor _27746_ (_04785_, _04390_, _04391_);
  nor _27747_ (_04786_, _04785_, _04730_);
  and _27748_ (_04787_, _04785_, _04730_);
  nor _27749_ (_04788_, _04787_, _04786_);
  and _27750_ (_04789_, _04788_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  nor _27751_ (_04790_, _04788_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  and _27752_ (_04791_, _04728_, _04435_);
  nor _27753_ (_04792_, _04791_, _04729_);
  and _27754_ (_04793_, _04792_, _01106_);
  nor _27755_ (_04794_, _04792_, _01106_);
  and _27756_ (_04795_, _04726_, _04480_);
  nor _27757_ (_04796_, _04795_, _04727_);
  nor _27758_ (_04797_, _04796_, _01128_);
  and _27759_ (_04798_, _04796_, _01128_);
  and _27760_ (_04799_, _04724_, _04721_);
  nor _27761_ (_04800_, _04799_, _04725_);
  nor _27762_ (_04801_, _04800_, _01275_);
  not _27763_ (_04802_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _27764_ (_04804_, _04719_, _04584_);
  nor _27765_ (_04805_, _04804_, _04720_);
  nor _27766_ (_04807_, _04805_, _04802_);
  and _27767_ (_04809_, _04805_, _04802_);
  not _27768_ (_04811_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and _27769_ (_04813_, _04717_, _04714_);
  nor _27770_ (_04815_, _04813_, _04718_);
  and _27771_ (_04816_, _04815_, _04811_);
  and _27772_ (_04817_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _27773_ (_04818_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  or _27774_ (_04819_, _04818_, _04817_);
  not _27775_ (_04820_, _04819_);
  nand _27776_ (_04821_, _04820_, _04709_);
  or _27777_ (_04823_, _04820_, _04709_);
  and _27778_ (_04825_, _04823_, _04821_);
  not _27779_ (_04827_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor _27780_ (_04828_, _04712_, _04710_);
  nor _27781_ (_04829_, _04828_, _04713_);
  nor _27782_ (_04830_, _04829_, _04827_);
  and _27783_ (_04831_, _04829_, _04827_);
  or _27784_ (_04832_, _04831_, _04830_);
  or _27785_ (_04833_, _04832_, _04825_);
  nor _27786_ (_04834_, _04815_, _04811_);
  or _27787_ (_04835_, _04834_, _04833_);
  or _27788_ (_04836_, _04835_, _04816_);
  or _27789_ (_04837_, _04836_, _04809_);
  or _27790_ (_04838_, _04837_, _04807_);
  and _27791_ (_04839_, _04800_, _01275_);
  or _27792_ (_04840_, _04839_, _04838_);
  or _27793_ (_04841_, _04840_, _04801_);
  or _27794_ (_04842_, _04841_, _04798_);
  or _27795_ (_04843_, _04842_, _04797_);
  or _27796_ (_04844_, _04843_, _04794_);
  or _27797_ (_04845_, _04844_, _04793_);
  or _27798_ (_04846_, _04845_, _04790_);
  or _27799_ (_04847_, _04846_, _04789_);
  or _27800_ (_04848_, _04847_, _04784_);
  or _27801_ (_04849_, _04848_, _04783_);
  or _27802_ (_04850_, _04849_, _04780_);
  or _27803_ (_04851_, _04850_, _04770_);
  and _27804_ (_04852_, _04738_, _04375_);
  nor _27805_ (_04853_, _04852_, _04739_);
  nor _27806_ (_04854_, _04853_, _01142_);
  and _27807_ (_04855_, _04769_, _04765_);
  and _27808_ (_04856_, _04853_, _01142_);
  or _27809_ (_04857_, _04856_, _04855_);
  or _27810_ (_04858_, _04857_, _04854_);
  or _27811_ (_04859_, _04858_, _04851_);
  or _27812_ (_04860_, _04859_, _04764_);
  nor _27813_ (_04861_, _04355_, _01591_);
  and _27814_ (_04862_, _04355_, _01591_);
  or _27815_ (_04863_, _04862_, _04861_);
  nand _27816_ (_04864_, _04863_, _04349_);
  or _27817_ (_04865_, _04863_, _04349_);
  and _27818_ (_04866_, _04865_, _04864_);
  and _27819_ (_04867_, _04866_, _04747_);
  and _27820_ (_04868_, _04763_, _00664_);
  nor _27821_ (_04869_, _04866_, _04747_);
  or _27822_ (_04870_, _04869_, _04868_);
  or _27823_ (_04871_, _04870_, _04867_);
  or _27824_ (_04872_, _04871_, _04860_);
  or _27825_ (_04873_, _04872_, _04761_);
  nor _27826_ (_04874_, _04749_, _04352_);
  nor _27827_ (_04875_, _04874_, _04750_);
  nor _27828_ (_04876_, _04875_, _01580_);
  and _27829_ (_04877_, _04760_, _04751_);
  and _27830_ (_04878_, _04875_, _01580_);
  or _27831_ (_04879_, _04878_, _04877_);
  or _27832_ (_04880_, _04879_, _04876_);
  or _27833_ (_04881_, _04880_, _04873_);
  or _27834_ (_04882_, _04802_, \oc8051_symbolic_cxrom1.regvalid [13]);
  or _27835_ (_04883_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [5]);
  and _27836_ (_04884_, _04883_, _04882_);
  and _27837_ (_04885_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], _04811_);
  and _27838_ (_04886_, _04885_, _04884_);
  or _27839_ (_04887_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [9]);
  and _27840_ (_04888_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or _27841_ (_04889_, _04802_, \oc8051_symbolic_cxrom1.regvalid [1]);
  and _27842_ (_04890_, _04889_, _04888_);
  and _27843_ (_04891_, _04890_, _04887_);
  or _27844_ (_04892_, _04891_, _04886_);
  nor _27845_ (_04893_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _27846_ (_04895_, _04893_, _04811_);
  nor _27847_ (_04896_, _04895_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _27848_ (_04897_, _04895_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor _27849_ (_04898_, _04897_, _04896_);
  and _27850_ (_04899_, _04898_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and _27851_ (_04900_, _04893_, _04811_);
  nor _27852_ (_04901_, _04900_, _04895_);
  or _27853_ (_04902_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], _09063_);
  nand _27854_ (_04903_, _04902_, _04901_);
  or _27855_ (_04904_, _04903_, _04899_);
  and _27856_ (_04905_, _04904_, _04827_);
  nand _27857_ (_04906_, _04898_, _04277_);
  or _27858_ (_04907_, _04898_, \oc8051_symbolic_cxrom1.regvalid [3]);
  and _27859_ (_04908_, _04907_, _04906_);
  or _27860_ (_04909_, _04901_, _04908_);
  and _27861_ (_04911_, _04909_, _04905_);
  or _27862_ (_04912_, _04911_, _04892_);
  and _27863_ (_04913_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [8]);
  and _27864_ (_04914_, _04802_, \oc8051_symbolic_cxrom1.regvalid [0]);
  or _27865_ (_04915_, _04914_, _04913_);
  and _27866_ (_04917_, _04915_, _04811_);
  and _27867_ (_04918_, _04802_, \oc8051_symbolic_cxrom1.regvalid [4]);
  and _27868_ (_04919_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [12]);
  or _27869_ (_04920_, _04919_, _04918_);
  and _27870_ (_04921_, _04920_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or _27871_ (_04922_, _04921_, _04917_);
  and _27872_ (_04923_, _04922_, _04827_);
  and _27873_ (_04924_, _04888_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _27874_ (_04925_, _04924_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _27875_ (_04927_, _04924_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor _27876_ (_04928_, _04927_, _04925_);
  or _27877_ (_04929_, _04928_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and _27878_ (_04930_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _27879_ (_04931_, _04930_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor _27880_ (_04932_, _04931_, _04924_);
  and _27881_ (_04933_, _04932_, _04882_);
  and _27882_ (_04934_, _04933_, _04929_);
  or _27883_ (_04936_, _04928_, \oc8051_symbolic_cxrom1.regvalid [1]);
  not _27884_ (_04938_, _04932_);
  nand _27885_ (_04939_, _04928_, _08521_);
  and _27886_ (_04940_, _04939_, _04938_);
  and _27887_ (_04941_, _04940_, _04936_);
  or _27888_ (_04942_, _04941_, _04934_);
  and _27889_ (_04944_, _04942_, _04923_);
  or _27890_ (_04946_, _04928_, \oc8051_symbolic_cxrom1.regvalid [7]);
  or _27891_ (_04947_, _04802_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and _27892_ (_04948_, _04947_, _04932_);
  and _27893_ (_04949_, _04948_, _04946_);
  or _27894_ (_04951_, _04928_, \oc8051_symbolic_cxrom1.regvalid [3]);
  nand _27895_ (_04952_, _04928_, _04277_);
  and _27896_ (_04953_, _04952_, _04938_);
  and _27897_ (_04954_, _04953_, _04951_);
  or _27898_ (_04955_, _04954_, _04949_);
  and _27899_ (_04956_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [14]);
  and _27900_ (_04957_, _04802_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or _27901_ (_04958_, _04957_, _04811_);
  or _27902_ (_04959_, _04958_, _04956_);
  or _27903_ (_04961_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [2]);
  or _27904_ (_04962_, _04802_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and _27905_ (_04963_, _04962_, _04961_);
  or _27906_ (_04964_, _04963_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and _27907_ (_04965_, _04964_, _04959_);
  and _27908_ (_04967_, _04965_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and _27909_ (_04968_, _04920_, _04885_);
  or _27910_ (_04969_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [8]);
  or _27911_ (_04970_, _04802_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and _27912_ (_04971_, _04970_, _04888_);
  and _27913_ (_04972_, _04971_, _04969_);
  or _27914_ (_04973_, _04972_, _04968_);
  and _27915_ (_04974_, _04973_, _04967_);
  and _27916_ (_04975_, _04974_, _04955_);
  or _27917_ (_04976_, _04975_, _04944_);
  not _27918_ (_04977_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  or _27919_ (_04978_, _04973_, _04965_);
  and _27920_ (_04979_, _04978_, _04977_);
  and _27921_ (_04980_, _04979_, _04976_);
  and _27922_ (_04981_, _04980_, _04912_);
  or _27923_ (_04982_, _04827_, \oc8051_symbolic_cxrom1.regvalid [2]);
  or _27924_ (_04983_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_symbolic_cxrom1.regvalid [0]);
  and _27925_ (_04985_, _04983_, _04982_);
  or _27926_ (_04987_, _04985_, _04898_);
  or _27927_ (_04988_, _04827_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or _27928_ (_04989_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_symbolic_cxrom1.regvalid [8]);
  nand _27929_ (_04991_, _04989_, _04988_);
  and _27930_ (_04992_, _04991_, _04898_);
  nor _27931_ (_04993_, _04992_, _04901_);
  and _27932_ (_04994_, _04993_, _04987_);
  and _27933_ (_04995_, _04898_, \oc8051_symbolic_cxrom1.regvalid [12]);
  or _27934_ (_04996_, _04918_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  or _27935_ (_04997_, _04996_, _04995_);
  and _27936_ (_04998_, _04898_, \oc8051_symbolic_cxrom1.regvalid [14]);
  or _27937_ (_04999_, _04957_, _04827_);
  or _27938_ (_05000_, _04999_, _04998_);
  and _27939_ (_05001_, _05000_, _04901_);
  and _27940_ (_05002_, _05001_, _04997_);
  or _27941_ (_05003_, _05002_, _04994_);
  or _27942_ (_05004_, _04928_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or _27943_ (_05005_, _04802_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and _27944_ (_05006_, _05005_, _05004_);
  or _27945_ (_05007_, _05006_, _04938_);
  nand _27946_ (_05008_, _04928_, _09302_);
  or _27947_ (_05009_, _04928_, \oc8051_symbolic_cxrom1.regvalid [2]);
  and _27948_ (_05010_, _05009_, _05008_);
  or _27949_ (_05011_, _05010_, _04932_);
  and _27950_ (_05012_, _05011_, _05007_);
  or _27951_ (_05013_, _05012_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  not _27952_ (_05014_, \oc8051_symbolic_cxrom1.regvalid [0]);
  nor _27953_ (_05015_, _04928_, _05014_);
  and _27954_ (_05016_, _04928_, \oc8051_symbolic_cxrom1.regvalid [8]);
  or _27955_ (_05017_, _05016_, _05015_);
  and _27956_ (_05018_, _05017_, _04938_);
  or _27957_ (_05019_, _04928_, \oc8051_symbolic_cxrom1.regvalid [4]);
  or _27958_ (_05021_, _04802_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and _27959_ (_05022_, _05021_, _04932_);
  and _27960_ (_05023_, _05022_, _05019_);
  or _27961_ (_05024_, _05023_, _04827_);
  or _27962_ (_05025_, _05024_, _05018_);
  or _27963_ (_05026_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [7]);
  and _27964_ (_05027_, _05026_, _04947_);
  or _27965_ (_05028_, _05027_, _04811_);
  or _27966_ (_05029_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [3]);
  or _27967_ (_05030_, _04802_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and _27968_ (_05032_, _05030_, _05029_);
  or _27969_ (_05033_, _05032_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and _27970_ (_05034_, _05033_, _05028_);
  and _27971_ (_05035_, _05034_, _04930_);
  and _27972_ (_05036_, _04827_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  or _27973_ (_05037_, _04884_, _04811_);
  or _27974_ (_05038_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [1]);
  or _27975_ (_05039_, _04802_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and _27976_ (_05040_, _05039_, _05038_);
  or _27977_ (_05041_, _05040_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and _27978_ (_05042_, _05041_, _05037_);
  and _27979_ (_05043_, _05042_, _05036_);
  or _27980_ (_05044_, _05043_, _05035_);
  and _27981_ (_05045_, _05034_, _04827_);
  or _27982_ (_05046_, _05045_, _04892_);
  and _27983_ (_05047_, _05046_, _05044_);
  and _27984_ (_05048_, _05047_, _05025_);
  and _27985_ (_05049_, _05048_, _05013_);
  and _27986_ (_05050_, _05049_, _05003_);
  or _27987_ (_05051_, _05050_, _04981_);
  nor _27988_ (_05052_, _04250_, _01154_);
  and _27989_ (_05053_, _05052_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _27990_ (_05054_, _05052_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _27991_ (_05055_, _05054_, _05053_);
  nand _27992_ (_05056_, _05055_, _08515_);
  nor _27993_ (_05057_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and _27994_ (_05058_, _05057_, _13796_);
  nor _27995_ (_05059_, _05058_, _05052_);
  nor _27996_ (_05060_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [7]);
  not _27997_ (_05061_, _05060_);
  and _27998_ (_05062_, _05061_, _05059_);
  and _27999_ (_05063_, _05062_, _05056_);
  not _28000_ (_05064_, _05059_);
  and _28001_ (_05065_, _05055_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor _28002_ (_05066_, _05055_, _08508_);
  or _28003_ (_05067_, _05066_, _05065_);
  and _28004_ (_05068_, _05067_, _05064_);
  or _28005_ (_05069_, _05068_, _05063_);
  and _28006_ (_05070_, _05069_, _04250_);
  or _28007_ (_05071_, _05055_, \oc8051_symbolic_cxrom1.regvalid [4]);
  and _28008_ (_05072_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _04285_);
  nor _28009_ (_05073_, _05072_, _05064_);
  and _28010_ (_05074_, _05073_, _05071_);
  and _28011_ (_05075_, _05055_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor _28012_ (_05076_, _05055_, _05014_);
  or _28013_ (_05077_, _05076_, _05075_);
  and _28014_ (_05078_, _05077_, _05064_);
  or _28015_ (_05079_, _05078_, _05074_);
  and _28016_ (_05080_, _05079_, _04296_);
  or _28017_ (_05081_, _05080_, _05070_);
  nand _28018_ (_05082_, _05055_, _08546_);
  nor _28019_ (_05083_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [6]);
  not _28020_ (_05084_, _05083_);
  and _28021_ (_05085_, _05084_, _05059_);
  and _28022_ (_05086_, _05085_, _05082_);
  or _28023_ (_05087_, _05055_, \oc8051_symbolic_cxrom1.regvalid [2]);
  nand _28024_ (_05088_, _05055_, _09302_);
  and _28025_ (_05089_, _05088_, _05087_);
  and _28026_ (_05090_, _05089_, _05064_);
  or _28027_ (_05091_, _05090_, _05086_);
  and _28028_ (_05092_, _05091_, _04252_);
  or _28029_ (_05093_, _05055_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and _28030_ (_05094_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _08481_);
  nor _28031_ (_05095_, _05094_, _05064_);
  and _28032_ (_05096_, _05095_, _05093_);
  or _28033_ (_05097_, _05055_, \oc8051_symbolic_cxrom1.regvalid [1]);
  nand _28034_ (_05098_, _05055_, _08521_);
  and _28035_ (_05099_, _05098_, _05064_);
  and _28036_ (_05100_, _05099_, _05097_);
  or _28037_ (_05101_, _05100_, _05096_);
  and _28038_ (_05102_, _05101_, _04270_);
  or _28039_ (_05103_, _05102_, _05092_);
  or _28040_ (_05104_, _05103_, _05081_);
  and _28041_ (_05105_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _08515_);
  nor _28042_ (_05106_, _05105_, _01154_);
  and _28043_ (_05107_, _05106_, _05061_);
  and _28044_ (_05108_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _04277_);
  nor _28045_ (_05109_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [3]);
  nor _28046_ (_05110_, _05109_, _05108_);
  and _28047_ (_05111_, _05110_, _01154_);
  nor _28048_ (_05112_, _05111_, _05107_);
  nor _28049_ (_05113_, _05112_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  not _28050_ (_05114_, _04235_);
  and _28051_ (_05115_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [1]);
  and _28052_ (_05116_, _01279_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor _28053_ (_05117_, _05116_, _05115_);
  nor _28054_ (_05118_, _05117_, _05114_);
  nor _28055_ (_05119_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [5]);
  nor _28056_ (_05120_, _05119_, _05094_);
  and _28057_ (_05121_, _05120_, _04586_);
  nor _28058_ (_05122_, _05121_, _05118_);
  not _28059_ (_05123_, _05122_);
  nor _28060_ (_05124_, _05123_, _05113_);
  nor _28061_ (_05125_, _05124_, _13796_);
  not _28062_ (_05126_, _05125_);
  and _28063_ (_05127_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _08546_);
  nor _28064_ (_05128_, _05127_, _01154_);
  and _28065_ (_05129_, _05128_, _05084_);
  and _28066_ (_05130_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _09302_);
  nor _28067_ (_05131_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [2]);
  nor _28068_ (_05132_, _05131_, _05130_);
  and _28069_ (_05133_, _05132_, _01154_);
  nor _28070_ (_05134_, _05133_, _05129_);
  nor _28071_ (_05135_, _05134_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nor _28072_ (_05136_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [4]);
  nor _28073_ (_05137_, _05136_, _05072_);
  and _28074_ (_05138_, _05137_, _04586_);
  nor _28075_ (_05139_, _05138_, _05135_);
  nor _28076_ (_05140_, _05139_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28077_ (_05141_, _04270_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and _28078_ (_05142_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _05014_);
  nor _28079_ (_05143_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [8]);
  nor _28080_ (_05144_, _05143_, _05142_);
  and _28081_ (_05145_, _05144_, _05141_);
  nor _28082_ (_05146_, _05145_, _05140_);
  and _28083_ (_05147_, _05146_, _05126_);
  and _28084_ (_05148_, _05137_, _04585_);
  nor _28085_ (_05149_, _05148_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28086_ (_05150_, _05134_, _12846_);
  and _28087_ (_05151_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _04290_);
  nor _28088_ (_05152_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [0]);
  nor _28089_ (_05153_, _05152_, _05151_);
  and _28090_ (_05154_, _05153_, _05057_);
  nor _28091_ (_05155_, _05154_, _05150_);
  and _28092_ (_05156_, _05155_, _05149_);
  nor _28093_ (_05157_, _05112_, _12846_);
  nor _28094_ (_05158_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [1]);
  and _28095_ (_05159_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _08521_);
  nor _28096_ (_05160_, _05159_, _05158_);
  and _28097_ (_05161_, _05160_, _05057_);
  and _28098_ (_05162_, _05120_, _04585_);
  or _28099_ (_05163_, _05162_, _13796_);
  or _28100_ (_05164_, _05163_, _05161_);
  nor _28101_ (_05165_, _05164_, _05157_);
  nor _28102_ (_05166_, _05165_, _05156_);
  not _28103_ (_05167_, _08064_);
  nor _28104_ (_05168_, _05167_, first_instr);
  nand _28105_ (_05169_, _05168_, _05166_);
  or _28106_ (_05170_, _05169_, _05147_);
  nor _28107_ (_05171_, _05170_, _04309_);
  and _28108_ (_05172_, _05171_, _05104_);
  and _28109_ (_05173_, _05172_, _05051_);
  nor _28110_ (_05174_, \oc8051_symbolic_cxrom1.regarray[0] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28111_ (_05175_, _09720_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28112_ (_05176_, _05175_, _05174_);
  and _28113_ (_05177_, _05176_, _05057_);
  nor _28114_ (_05178_, _05177_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _28115_ (_05179_, \oc8051_symbolic_cxrom1.regarray[4] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28116_ (_05180_, _10197_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28117_ (_05181_, _05180_, _05179_);
  and _28118_ (_05182_, _05181_, _04585_);
  not _28119_ (_05183_, _05182_);
  nor _28120_ (_05184_, \oc8051_symbolic_cxrom1.regarray[2] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28121_ (_05185_, _09963_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28122_ (_05186_, _05185_, _05184_);
  and _28123_ (_05187_, _05186_, _04586_);
  nor _28124_ (_05188_, \oc8051_symbolic_cxrom1.regarray[6] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28125_ (_05189_, _10406_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28126_ (_05190_, _05189_, _05188_);
  and _28127_ (_05191_, _05190_, _04235_);
  nor _28128_ (_05192_, _05191_, _05187_);
  and _28129_ (_05193_, _05192_, _05183_);
  and _28130_ (_05194_, _05193_, _05178_);
  nor _28131_ (_05195_, \oc8051_symbolic_cxrom1.regarray[8] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28132_ (_05196_, _10624_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28133_ (_05197_, _05196_, _05195_);
  and _28134_ (_05198_, _05197_, _05057_);
  nor _28135_ (_05199_, _05198_, _01279_);
  nor _28136_ (_05200_, \oc8051_symbolic_cxrom1.regarray[12] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28137_ (_05201_, _12365_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28138_ (_05202_, _05201_, _05200_);
  and _28139_ (_05203_, _05202_, _04585_);
  not _28140_ (_05204_, _05203_);
  nor _28141_ (_05205_, \oc8051_symbolic_cxrom1.regarray[10] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28142_ (_05206_, _11249_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28143_ (_05207_, _05206_, _05205_);
  and _28144_ (_05208_, _05207_, _04586_);
  nor _28145_ (_05209_, \oc8051_symbolic_cxrom1.regarray[14] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28146_ (_05210_, _12729_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28147_ (_05211_, _05210_, _05209_);
  and _28148_ (_05212_, _05211_, _04235_);
  nor _28149_ (_05213_, _05212_, _05208_);
  and _28150_ (_05214_, _05213_, _05204_);
  and _28151_ (_05215_, _05214_, _05199_);
  nor _28152_ (_05216_, _05215_, _05194_);
  and _28153_ (_05217_, _05216_, _05166_);
  nor _28154_ (_05218_, \oc8051_symbolic_cxrom1.regarray[0] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28155_ (_05219_, _09697_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28156_ (_05220_, _05219_, _05218_);
  and _28157_ (_05221_, _05220_, _05057_);
  nor _28158_ (_05222_, _05221_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _28159_ (_05223_, \oc8051_symbolic_cxrom1.regarray[4] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28160_ (_05224_, _10183_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28161_ (_05225_, _05224_, _05223_);
  and _28162_ (_05226_, _05225_, _04585_);
  not _28163_ (_05227_, _05226_);
  nor _28164_ (_05228_, \oc8051_symbolic_cxrom1.regarray[2] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28165_ (_05229_, _09941_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28166_ (_05230_, _05229_, _05228_);
  and _28167_ (_05231_, _05230_, _04586_);
  nor _28168_ (_05232_, \oc8051_symbolic_cxrom1.regarray[6] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28169_ (_05233_, _10396_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28170_ (_05234_, _05233_, _05232_);
  and _28171_ (_05235_, _05234_, _04235_);
  nor _28172_ (_05236_, _05235_, _05231_);
  and _28173_ (_05237_, _05236_, _05227_);
  and _28174_ (_05238_, _05237_, _05222_);
  nor _28175_ (_05239_, \oc8051_symbolic_cxrom1.regarray[8] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28176_ (_05240_, _10608_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28177_ (_05241_, _05240_, _05239_);
  and _28178_ (_05242_, _05241_, _05057_);
  nor _28179_ (_05243_, _05242_, _01279_);
  nor _28180_ (_05244_, \oc8051_symbolic_cxrom1.regarray[12] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28181_ (_05245_, _12347_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28182_ (_05246_, _05245_, _05244_);
  and _28183_ (_05247_, _05246_, _04585_);
  not _28184_ (_05248_, _05247_);
  nor _28185_ (_05249_, \oc8051_symbolic_cxrom1.regarray[10] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28186_ (_05250_, _11230_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28187_ (_05251_, _05250_, _05249_);
  and _28188_ (_05252_, _05251_, _04586_);
  nor _28189_ (_05253_, \oc8051_symbolic_cxrom1.regarray[14] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28190_ (_05254_, _12717_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28191_ (_05255_, _05254_, _05253_);
  and _28192_ (_05256_, _05255_, _04235_);
  nor _28193_ (_05257_, _05256_, _05252_);
  and _28194_ (_05258_, _05257_, _05248_);
  and _28195_ (_05259_, _05258_, _05243_);
  nor _28196_ (_05260_, _05259_, _05238_);
  and _28197_ (_05261_, _05260_, _05166_);
  nor _28198_ (_05262_, _05261_, _05217_);
  nor _28199_ (_05263_, \oc8051_symbolic_cxrom1.regarray[0] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28200_ (_05264_, _09775_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28201_ (_05265_, _05264_, _05263_);
  and _28202_ (_05266_, _05265_, _05057_);
  nor _28203_ (_05267_, _05266_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _28204_ (_05268_, \oc8051_symbolic_cxrom1.regarray[4] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28205_ (_05269_, _10245_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28206_ (_05270_, _05269_, _05268_);
  and _28207_ (_05271_, _05270_, _04585_);
  not _28208_ (_05272_, _05271_);
  nor _28209_ (_05273_, \oc8051_symbolic_cxrom1.regarray[2] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28210_ (_05274_, _10027_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28211_ (_05275_, _05274_, _05273_);
  and _28212_ (_05276_, _05275_, _04586_);
  nor _28213_ (_05277_, \oc8051_symbolic_cxrom1.regarray[6] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28214_ (_05278_, _10454_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28215_ (_05279_, _05278_, _05277_);
  and _28216_ (_05280_, _05279_, _04235_);
  nor _28217_ (_05281_, _05280_, _05276_);
  and _28218_ (_05282_, _05281_, _05272_);
  and _28219_ (_05283_, _05282_, _05267_);
  nor _28220_ (_05284_, \oc8051_symbolic_cxrom1.regarray[8] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28221_ (_05285_, _10672_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28222_ (_05286_, _05285_, _05284_);
  and _28223_ (_05287_, _05286_, _05057_);
  nor _28224_ (_05288_, _05287_, _01279_);
  nor _28225_ (_05289_, \oc8051_symbolic_cxrom1.regarray[12] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28226_ (_05290_, _12416_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28227_ (_05291_, _05290_, _05289_);
  and _28228_ (_05292_, _05291_, _04585_);
  not _28229_ (_05293_, _05292_);
  nor _28230_ (_05294_, \oc8051_symbolic_cxrom1.regarray[10] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28231_ (_05295_, _11305_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28232_ (_05296_, _05295_, _05294_);
  and _28233_ (_05297_, _05296_, _04586_);
  nor _28234_ (_05298_, \oc8051_symbolic_cxrom1.regarray[14] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28235_ (_05299_, _12779_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28236_ (_05300_, _05299_, _05298_);
  and _28237_ (_05301_, _05300_, _04235_);
  nor _28238_ (_05302_, _05301_, _05297_);
  and _28239_ (_05303_, _05302_, _05293_);
  and _28240_ (_05304_, _05303_, _05288_);
  nor _28241_ (_05305_, _05304_, _05283_);
  and _28242_ (_05306_, _05305_, _05166_);
  nor _28243_ (_05307_, \oc8051_symbolic_cxrom1.regarray[2] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28244_ (_05308_, _10011_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28245_ (_05309_, _05308_, _05307_);
  and _28246_ (_05310_, _05309_, _04586_);
  nor _28247_ (_05311_, \oc8051_symbolic_cxrom1.regarray[4] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28248_ (_05312_, _10233_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28249_ (_05313_, _05312_, _05311_);
  and _28250_ (_05314_, _05313_, _04585_);
  nor _28251_ (_05315_, \oc8051_symbolic_cxrom1.regarray[6] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28252_ (_05316_, _10443_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28253_ (_05317_, _05316_, _05315_);
  and _28254_ (_05318_, _05317_, _04235_);
  nor _28255_ (_05319_, \oc8051_symbolic_cxrom1.regarray[0] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28256_ (_05320_, _09761_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28257_ (_05321_, _05320_, _05319_);
  and _28258_ (_05322_, _05321_, _05057_);
  or _28259_ (_05323_, _05322_, _05318_);
  or _28260_ (_05324_, _05323_, _05314_);
  or _28261_ (_05325_, _05324_, _05310_);
  and _28262_ (_05326_, _05325_, _01279_);
  nor _28263_ (_05327_, \oc8051_symbolic_cxrom1.regarray[10] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28264_ (_05328_, _11292_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28265_ (_05329_, _05328_, _05327_);
  and _28266_ (_05330_, _05329_, _04586_);
  nor _28267_ (_05331_, \oc8051_symbolic_cxrom1.regarray[12] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28268_ (_05332_, _12403_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28269_ (_05333_, _05332_, _05331_);
  and _28270_ (_05334_, _05333_, _04585_);
  nor _28271_ (_05335_, \oc8051_symbolic_cxrom1.regarray[14] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28272_ (_05336_, _12766_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28273_ (_05337_, _05336_, _05335_);
  and _28274_ (_05338_, _05337_, _04235_);
  nor _28275_ (_05339_, \oc8051_symbolic_cxrom1.regarray[8] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28276_ (_05340_, _10660_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28277_ (_05341_, _05340_, _05339_);
  and _28278_ (_05342_, _05341_, _05057_);
  or _28279_ (_05343_, _05342_, _05338_);
  or _28280_ (_05344_, _05343_, _05334_);
  or _28281_ (_05345_, _05344_, _05330_);
  and _28282_ (_05346_, _05345_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or _28283_ (_05347_, _05346_, _05326_);
  and _28284_ (_05348_, _05347_, _05166_);
  nor _28285_ (_05349_, _05348_, _05306_);
  and _28286_ (_05350_, _05349_, _05262_);
  nor _28287_ (_05351_, \oc8051_symbolic_cxrom1.regarray[2] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28288_ (_05352_, _09985_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28289_ (_05353_, _05352_, _05351_);
  and _28290_ (_05354_, _05353_, _04586_);
  nor _28291_ (_05355_, \oc8051_symbolic_cxrom1.regarray[4] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28292_ (_05356_, _10209_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28293_ (_05357_, _05356_, _05355_);
  and _28294_ (_05358_, _05357_, _04585_);
  nor _28295_ (_05359_, \oc8051_symbolic_cxrom1.regarray[0] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28296_ (_05360_, _09734_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28297_ (_05361_, _05360_, _05359_);
  and _28298_ (_05362_, _05361_, _05057_);
  nor _28299_ (_05363_, \oc8051_symbolic_cxrom1.regarray[6] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28300_ (_05364_, _10420_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28301_ (_05365_, _05364_, _05363_);
  and _28302_ (_05366_, _05365_, _04235_);
  or _28303_ (_05367_, _05366_, _05362_);
  or _28304_ (_05368_, _05367_, _05358_);
  or _28305_ (_05369_, _05368_, _05354_);
  and _28306_ (_05370_, _05369_, _01279_);
  nor _28307_ (_05371_, \oc8051_symbolic_cxrom1.regarray[10] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28308_ (_05372_, _11267_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28309_ (_05373_, _05372_, _05371_);
  and _28310_ (_05374_, _05373_, _04586_);
  nor _28311_ (_05375_, \oc8051_symbolic_cxrom1.regarray[12] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28312_ (_05376_, _12378_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28313_ (_05377_, _05376_, _05375_);
  and _28314_ (_05378_, _05377_, _04585_);
  nor _28315_ (_05379_, \oc8051_symbolic_cxrom1.regarray[8] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28316_ (_05380_, _10636_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28317_ (_05381_, _05380_, _05379_);
  and _28318_ (_05382_, _05381_, _05057_);
  nor _28319_ (_05383_, \oc8051_symbolic_cxrom1.regarray[14] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28320_ (_05384_, _12741_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28321_ (_05385_, _05384_, _05383_);
  and _28322_ (_05386_, _05385_, _04235_);
  or _28323_ (_05387_, _05386_, _05382_);
  or _28324_ (_05388_, _05387_, _05378_);
  or _28325_ (_05389_, _05388_, _05374_);
  and _28326_ (_05390_, _05389_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or _28327_ (_05391_, _05390_, _05370_);
  and _28328_ (_05392_, _05391_, _05166_);
  nor _28329_ (_05393_, \oc8051_symbolic_cxrom1.regarray[2] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28330_ (_05394_, _09998_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28331_ (_05395_, _05394_, _05393_);
  and _28332_ (_05396_, _05395_, _04586_);
  nor _28333_ (_05397_, \oc8051_symbolic_cxrom1.regarray[4] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28334_ (_05398_, _10221_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28335_ (_05399_, _05398_, _05397_);
  and _28336_ (_05400_, _05399_, _04585_);
  nor _28337_ (_05401_, \oc8051_symbolic_cxrom1.regarray[0] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28338_ (_05402_, _09749_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28339_ (_05403_, _05402_, _05401_);
  and _28340_ (_05404_, _05403_, _05057_);
  nor _28341_ (_05405_, \oc8051_symbolic_cxrom1.regarray[6] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28342_ (_05406_, _10431_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28343_ (_05407_, _05406_, _05405_);
  and _28344_ (_05408_, _05407_, _04235_);
  or _28345_ (_05409_, _05408_, _05404_);
  or _28346_ (_05410_, _05409_, _05400_);
  or _28347_ (_05411_, _05410_, _05396_);
  and _28348_ (_05412_, _05411_, _01279_);
  nor _28349_ (_05413_, \oc8051_symbolic_cxrom1.regarray[10] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28350_ (_05414_, _11279_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28351_ (_05415_, _05414_, _05413_);
  and _28352_ (_05416_, _05415_, _04586_);
  nor _28353_ (_05417_, \oc8051_symbolic_cxrom1.regarray[12] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28354_ (_05418_, _12391_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28355_ (_05419_, _05418_, _05417_);
  and _28356_ (_05420_, _05419_, _04585_);
  nor _28357_ (_05421_, \oc8051_symbolic_cxrom1.regarray[8] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28358_ (_05422_, _10649_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28359_ (_05423_, _05422_, _05421_);
  and _28360_ (_05424_, _05423_, _05057_);
  nor _28361_ (_05425_, \oc8051_symbolic_cxrom1.regarray[14] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28362_ (_05426_, _12754_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28363_ (_05427_, _05426_, _05425_);
  and _28364_ (_05428_, _05427_, _04235_);
  or _28365_ (_05429_, _05428_, _05424_);
  or _28366_ (_05430_, _05429_, _05420_);
  or _28367_ (_05431_, _05430_, _05416_);
  and _28368_ (_05432_, _05431_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or _28369_ (_05433_, _05432_, _05412_);
  and _28370_ (_05434_, _05433_, _05166_);
  nor _28371_ (_05435_, _05434_, _05392_);
  nor _28372_ (_05436_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_symbolic_cxrom1.regarray[0] [7]);
  and _28373_ (_05437_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _08600_);
  nor _28374_ (_05438_, _05437_, _05436_);
  and _28375_ (_05439_, _05438_, _05057_);
  nor _28376_ (_05440_, _05439_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _28377_ (_05441_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_symbolic_cxrom1.regarray[4] [7]);
  and _28378_ (_05442_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _08595_);
  nor _28379_ (_05443_, _05442_, _05441_);
  and _28380_ (_05444_, _05443_, _04585_);
  not _28381_ (_05445_, _05444_);
  nor _28382_ (_05446_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_symbolic_cxrom1.regarray[2] [7]);
  and _28383_ (_05447_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _08584_);
  nor _28384_ (_05448_, _05447_, _05446_);
  and _28385_ (_05449_, _05448_, _04586_);
  nor _28386_ (_05450_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_symbolic_cxrom1.regarray[6] [7]);
  and _28387_ (_05451_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _08590_);
  nor _28388_ (_05452_, _05451_, _05450_);
  and _28389_ (_05453_, _05452_, _04235_);
  nor _28390_ (_05454_, _05453_, _05449_);
  and _28391_ (_05455_, _05454_, _05445_);
  and _28392_ (_05456_, _05455_, _05440_);
  nor _28393_ (_05457_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_symbolic_cxrom1.regarray[8] [7]);
  and _28394_ (_05458_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _08576_);
  nor _28395_ (_05459_, _05458_, _05457_);
  and _28396_ (_05460_, _05459_, _05057_);
  nor _28397_ (_05461_, _05460_, _01279_);
  nor _28398_ (_05462_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_symbolic_cxrom1.regarray[12] [7]);
  and _28399_ (_05463_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _08571_);
  nor _28400_ (_05464_, _05463_, _05462_);
  and _28401_ (_05465_, _05464_, _04585_);
  not _28402_ (_05466_, _05465_);
  nor _28403_ (_05467_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_symbolic_cxrom1.regarray[10] [7]);
  and _28404_ (_05468_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _08565_);
  nor _28405_ (_05469_, _05468_, _05467_);
  and _28406_ (_05470_, _05469_, _04586_);
  nor _28407_ (_05471_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_symbolic_cxrom1.regarray[14] [7]);
  and _28408_ (_05472_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _08560_);
  nor _28409_ (_05473_, _05472_, _05471_);
  and _28410_ (_05474_, _05473_, _04235_);
  nor _28411_ (_05475_, _05474_, _05470_);
  and _28412_ (_05476_, _05475_, _05466_);
  and _28413_ (_05477_, _05476_, _05461_);
  nor _28414_ (_05478_, _05477_, _05456_);
  and _28415_ (_05479_, _05478_, _05166_);
  nor _28416_ (_05480_, \oc8051_symbolic_cxrom1.regarray[2] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28417_ (_05481_, _10042_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28418_ (_05482_, _05481_, _05480_);
  and _28419_ (_05483_, _05482_, _04586_);
  nor _28420_ (_05484_, \oc8051_symbolic_cxrom1.regarray[4] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28421_ (_05485_, _10258_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28422_ (_05486_, _05485_, _05484_);
  and _28423_ (_05487_, _05486_, _04585_);
  nor _28424_ (_05488_, \oc8051_symbolic_cxrom1.regarray[6] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28425_ (_05489_, _10469_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28426_ (_05490_, _05489_, _05488_);
  and _28427_ (_05491_, _05490_, _04235_);
  nor _28428_ (_05492_, \oc8051_symbolic_cxrom1.regarray[0] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28429_ (_05493_, _09792_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28430_ (_05494_, _05493_, _05492_);
  and _28431_ (_05495_, _05494_, _05057_);
  or _28432_ (_05496_, _05495_, _05491_);
  or _28433_ (_05497_, _05496_, _05487_);
  or _28434_ (_05498_, _05497_, _05483_);
  and _28435_ (_05499_, _05498_, _01279_);
  nor _28436_ (_05500_, \oc8051_symbolic_cxrom1.regarray[10] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28437_ (_05501_, _11318_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28438_ (_05502_, _05501_, _05500_);
  and _28439_ (_05503_, _05502_, _04586_);
  nor _28440_ (_05504_, \oc8051_symbolic_cxrom1.regarray[12] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28441_ (_05505_, _12429_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28442_ (_05506_, _05505_, _05504_);
  and _28443_ (_05507_, _05506_, _04585_);
  nor _28444_ (_05508_, \oc8051_symbolic_cxrom1.regarray[14] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28445_ (_05509_, _12794_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28446_ (_05510_, _05509_, _05508_);
  and _28447_ (_05511_, _05510_, _04235_);
  nor _28448_ (_05512_, \oc8051_symbolic_cxrom1.regarray[8] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28449_ (_05513_, _10685_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28450_ (_05514_, _05513_, _05512_);
  and _28451_ (_05515_, _05514_, _05057_);
  or _28452_ (_05516_, _05515_, _05511_);
  or _28453_ (_05517_, _05516_, _05507_);
  or _28454_ (_05518_, _05517_, _05503_);
  and _28455_ (_05519_, _05518_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or _28456_ (_05520_, _05519_, _05499_);
  and _28457_ (_05521_, _05520_, _05166_);
  not _28458_ (_05522_, _05521_);
  and _28459_ (_05523_, _05522_, _05479_);
  and _28460_ (_05524_, _05523_, _05435_);
  and _28461_ (_05525_, _05524_, _05350_);
  and _28462_ (_05526_, _05525_, _05173_);
  and _28463_ (_05527_, _05526_, _04881_);
  not _28464_ (_05528_, _05479_);
  nand _28465_ (_05529_, _05348_, _05305_);
  and _28466_ (_05530_, _05392_, _05217_);
  nor _28467_ (_05531_, _05530_, _05433_);
  nor _28468_ (_05532_, _05531_, _05529_);
  not _28469_ (_05533_, _05261_);
  and _28470_ (_05534_, _05435_, _05533_);
  and _28471_ (_05535_, _05534_, _05217_);
  not _28472_ (_05536_, _05260_);
  not _28473_ (_05537_, _05216_);
  not _28474_ (_05538_, _05433_);
  and _28475_ (_05539_, _05538_, _05392_);
  and _28476_ (_05540_, _05539_, _05537_);
  and _28477_ (_05541_, _05540_, _05536_);
  or _28478_ (_05542_, _05541_, _05535_);
  or _28479_ (_05543_, _05542_, _05532_);
  and _28480_ (_05544_, _05543_, _05521_);
  not _28481_ (_05545_, _05306_);
  nor _28482_ (_05546_, _05520_, _05545_);
  and _28483_ (_05547_, _05546_, _05540_);
  and _28484_ (_05548_, _05540_, _05261_);
  and _28485_ (_05549_, _05548_, _05545_);
  or _28486_ (_05550_, _05549_, _05547_);
  or _28487_ (_05551_, _05550_, _05544_);
  and _28488_ (_05552_, _05551_, _05528_);
  and _28489_ (_05553_, _05535_, _05545_);
  not _28490_ (_05554_, _05305_);
  and _28491_ (_05555_, _05521_, _05554_);
  and _28492_ (_05556_, _05555_, _05534_);
  and _28493_ (_05557_, _05521_, _05305_);
  and _28494_ (_05558_, _05557_, _05548_);
  or _28495_ (_05559_, _05558_, _05556_);
  or _28496_ (_05560_, _05559_, _05553_);
  and _28497_ (_05561_, _05560_, _05479_);
  and _28498_ (_05562_, _05348_, _05554_);
  and _28499_ (_05563_, _05562_, _05540_);
  not _28500_ (_05564_, _05348_);
  and _28501_ (_05565_, _05434_, _05564_);
  and _28502_ (_05566_, _05530_, _05564_);
  or _28503_ (_05567_, _05566_, _05565_);
  or _28504_ (_05568_, _05567_, _05563_);
  and _28505_ (_05569_, _05568_, _05523_);
  and _28506_ (_05570_, _05534_, _05306_);
  and _28507_ (_05571_, _05570_, _05523_);
  and _28508_ (_05572_, _05548_, _05564_);
  and _28509_ (_05573_, _05572_, _05521_);
  or _28510_ (_05574_, _05573_, _05571_);
  or _28511_ (_05575_, _05574_, _05569_);
  or _28512_ (_05576_, _05575_, _05561_);
  or _28513_ (_05577_, _05576_, _05552_);
  nor _28514_ (_05578_, _04359_, _00664_);
  and _28515_ (_05579_, _04359_, _00664_);
  or _28516_ (_05580_, _05579_, _05578_);
  or _28517_ (_05581_, _05580_, _04863_);
  and _28518_ (_05582_, _04249_, _01580_);
  nor _28519_ (_05583_, _04249_, _01580_);
  or _28520_ (_05584_, _05583_, _05582_);
  or _28521_ (_05585_, _05584_, _04757_);
  or _28522_ (_05586_, _05585_, _05581_);
  nor _28523_ (_05587_, _04363_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and _28524_ (_05588_, _04363_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nor _28525_ (_05589_, _05588_, _05587_);
  nor _28526_ (_05590_, _04368_, _01142_);
  and _28527_ (_05591_, _04368_, _01142_);
  or _28528_ (_05592_, _05591_, _05590_);
  nor _28529_ (_05593_, _04438_, _01128_);
  and _28530_ (_05594_, _04438_, _01128_);
  or _28531_ (_05595_, _05594_, _05593_);
  nor _28532_ (_05596_, _04393_, _01106_);
  and _28533_ (_05597_, _04393_, _01106_);
  or _28534_ (_05598_, _05597_, _05596_);
  or _28535_ (_05599_, _05598_, _05595_);
  and _28536_ (_05600_, _04525_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor _28537_ (_05601_, _04525_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or _28538_ (_05602_, _05601_, _05600_);
  and _28539_ (_05603_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nor _28540_ (_05604_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nor _28541_ (_05605_, _05604_, _05603_);
  nand _28542_ (_05606_, _05605_, _04819_);
  and _28543_ (_05607_, _04588_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor _28544_ (_05608_, _04588_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or _28545_ (_05609_, _05608_, _05607_);
  or _28546_ (_05610_, _05609_, _05606_);
  or _28547_ (_05611_, _05610_, _05602_);
  nor _28548_ (_05612_, _04482_, _01275_);
  and _28549_ (_05613_, _04482_, _01275_);
  or _28550_ (_05614_, _05613_, _05612_);
  or _28551_ (_05615_, _05614_, _05611_);
  nor _28552_ (_05616_, _04384_, _01872_);
  or _28553_ (_05617_, _05616_, _05615_);
  or _28554_ (_05618_, _05617_, _05599_);
  or _28555_ (_05619_, _05618_, _05592_);
  and _28556_ (_05620_, _04389_, _01076_);
  and _28557_ (_05621_, _04384_, _01872_);
  nor _28558_ (_05622_, _04389_, _01076_);
  or _28559_ (_05623_, _05622_, _05621_);
  or _28560_ (_05624_, _05623_, _05620_);
  or _28561_ (_05625_, _05624_, _04774_);
  or _28562_ (_05626_, _05625_, _05619_);
  or _28563_ (_05627_, _05626_, _05589_);
  or _28564_ (_05628_, _05627_, _05586_);
  and _28565_ (_05629_, _05628_, _05577_);
  and _28566_ (_05630_, _05261_, _05217_);
  and _28567_ (_05631_, _05630_, _05435_);
  and _28568_ (_05632_, _05541_, _05349_);
  or _28569_ (_05633_, _05632_, _05631_);
  nor _28570_ (_05634_, _05305_, _05260_);
  and _28571_ (_05635_, _05634_, _05392_);
  nor _28572_ (_05636_, _05635_, _05350_);
  nor _28573_ (_05637_, _05636_, _05479_);
  or _28574_ (_05638_, _05637_, _05633_);
  and _28575_ (_05639_, _05638_, _05522_);
  and _28576_ (_05640_, _05547_, _05564_);
  or _28577_ (_05641_, _05539_, _05306_);
  or _28578_ (_05642_, _05433_, _05536_);
  and _28579_ (_05643_, _05642_, _05521_);
  and _28580_ (_05644_, _05643_, _05641_);
  or _28581_ (_05645_, _05644_, _05640_);
  and _28582_ (_05646_, _05645_, _05479_);
  nand _28583_ (_05647_, _05478_, _05217_);
  nor _28584_ (_05648_, _05647_, _05642_);
  or _28585_ (_05649_, _05648_, _05566_);
  and _28586_ (_05650_, _05649_, _05521_);
  nor _28587_ (_05651_, _05521_, _05479_);
  nand _28588_ (_05652_, _05347_, _05545_);
  nor _28589_ (_05653_, _05652_, _05434_);
  or _28590_ (_05654_, _05653_, _05651_);
  and _28591_ (_05655_, _05654_, _05530_);
  and _28592_ (_05656_, _05522_, _05434_);
  not _28593_ (_05657_, _05478_);
  or _28594_ (_05658_, _05562_, _05657_);
  and _28595_ (_05659_, _05658_, _05656_);
  nor _28596_ (_05660_, _05478_, _05305_);
  and _28597_ (_05661_, _05660_, _05434_);
  and _28598_ (_05662_, _05565_, _05521_);
  or _28599_ (_05663_, _05662_, _05661_);
  or _28600_ (_05664_, _05663_, _05659_);
  or _28601_ (_05665_, _05664_, _05655_);
  or _28602_ (_05666_, _05665_, _05650_);
  or _28603_ (_05667_, _05666_, _05646_);
  or _28604_ (_05668_, _05667_, _05639_);
  nor _28605_ (_05669_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28606_ (_05670_, _04368_, _13796_);
  nor _28607_ (_05671_, _05670_, _05669_);
  and _28608_ (_05672_, _05671_, _01142_);
  and _28609_ (_05673_, _04247_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28610_ (_05674_, _05673_, _00601_);
  nor _28611_ (_05675_, _05673_, _00601_);
  or _28612_ (_05676_, _05675_, _05674_);
  nor _28613_ (_05677_, _05676_, _00584_);
  or _28614_ (_05678_, _05677_, _05672_);
  and _28615_ (_05679_, _04244_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28616_ (_05680_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  and _28617_ (_05681_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor _28618_ (_05682_, _05681_, _05680_);
  nand _28619_ (_05683_, _05682_, _05679_);
  or _28620_ (_05684_, _05682_, _05679_);
  and _28621_ (_05685_, _05684_, _05683_);
  and _28622_ (_05686_, _05676_, _00584_);
  or _28623_ (_05687_, _05686_, _05685_);
  or _28624_ (_05688_, _05687_, _05678_);
  nor _28625_ (_05689_, _05671_, _01142_);
  and _28626_ (_05690_, _04387_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28627_ (_05691_, _05690_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  and _28628_ (_05692_, _05690_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  nor _28629_ (_05693_, _05692_, _05691_);
  nor _28630_ (_05694_, _05693_, _01076_);
  and _28631_ (_05695_, _04259_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor _28632_ (_05696_, _04259_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or _28633_ (_05697_, _05696_, _05695_);
  or _28634_ (_05698_, _05697_, _05694_);
  and _28635_ (_05699_, _04236_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28636_ (_05700_, _05699_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nor _28637_ (_05701_, _05699_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nor _28638_ (_05702_, _05701_, _05700_);
  nor _28639_ (_05703_, _05702_, _01275_);
  and _28640_ (_05704_, _05702_, _01275_);
  or _28641_ (_05705_, _05704_, _05703_);
  and _28642_ (_05706_, _04386_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28643_ (_05707_, _05706_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nor _28644_ (_05708_, _05707_, _05690_);
  nor _28645_ (_05709_, _05708_, _01106_);
  and _28646_ (_05710_, _05700_, _01110_);
  nor _28647_ (_05711_, _05700_, _01110_);
  nor _28648_ (_05712_, _05711_, _05710_);
  nor _28649_ (_05713_, _05712_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  and _28650_ (_05714_, _05712_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nand _28651_ (_05715_, _05605_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  or _28652_ (_05716_, _05605_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28653_ (_05717_, _05716_, _05715_);
  or _28654_ (_05718_, _05717_, _04819_);
  nor _28655_ (_05719_, _04255_, _04811_);
  and _28656_ (_05720_, _04255_, _04811_);
  or _28657_ (_05721_, _05720_, _05719_);
  or _28658_ (_05722_, _05721_, _05718_);
  or _28659_ (_05723_, _05722_, _05714_);
  or _28660_ (_05724_, _05723_, _05713_);
  or _28661_ (_05725_, _05724_, _05709_);
  or _28662_ (_05726_, _05725_, _05705_);
  or _28663_ (_05727_, _05726_, _05698_);
  and _28664_ (_05728_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _13796_);
  and _28665_ (_05729_, _04378_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28666_ (_05730_, _05729_, _05728_);
  nor _28667_ (_05731_, _05730_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and _28668_ (_05732_, _05693_, _01076_);
  and _28669_ (_05733_, _05730_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  or _28670_ (_05734_, _05733_, _05732_);
  or _28671_ (_05735_, _05734_, _05731_);
  or _28672_ (_05736_, _05735_, _05727_);
  or _28673_ (_05737_, _05736_, _05689_);
  and _28674_ (_05738_, _05708_, _01106_);
  or _28675_ (_05739_, _04355_, _13796_);
  or _28676_ (_05740_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28677_ (_05741_, _05740_, _05739_);
  nor _28678_ (_05742_, _05741_, _01591_);
  or _28679_ (_05743_, _08066_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nand _28680_ (_05744_, _04363_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28681_ (_05745_, _05744_, _05743_);
  nor _28682_ (_05746_, _05745_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  or _28683_ (_05747_, _05746_, _05742_);
  or _28684_ (_05748_, _05747_, _05738_);
  or _28685_ (_05749_, _05748_, _05737_);
  nand _28686_ (_05750_, _04246_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28687_ (_05751_, _05750_, _00621_);
  nor _28688_ (_05752_, _05751_, _05673_);
  nor _28689_ (_05753_, _05752_, _01580_);
  and _28690_ (_05754_, _05752_, _01580_);
  or _28691_ (_05755_, _05754_, _05753_);
  and _28692_ (_05756_, _05741_, _01591_);
  or _28693_ (_05757_, _05756_, _05755_);
  and _28694_ (_05758_, _05699_, _04239_);
  and _28695_ (_05759_, _05758_, _01066_);
  nor _28696_ (_05760_, _05758_, _01066_);
  or _28697_ (_05761_, _05760_, _05759_);
  nor _28698_ (_05762_, _05761_, _01872_);
  and _28699_ (_05763_, _05761_, _01872_);
  or _28700_ (_05764_, _05763_, _05762_);
  and _28701_ (_05765_, _05745_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  or _28702_ (_05766_, _05765_, _05764_);
  or _28703_ (_05767_, _05766_, _05757_);
  or _28704_ (_05768_, _05767_, _05749_);
  or _28705_ (_05769_, _05768_, _05688_);
  and _28706_ (_05770_, _05769_, _05668_);
  and _28707_ (_05771_, _05558_, _05348_);
  and _28708_ (_05772_, _05529_, _05521_);
  and _28709_ (_05773_, _05772_, _05631_);
  or _28710_ (_05774_, _05773_, _05771_);
  and _28711_ (_05775_, _05774_, _05528_);
  and _28712_ (_05776_, _05435_, _05262_);
  and _28713_ (_05777_, _05776_, _05562_);
  and _28714_ (_05778_, _05572_, _05545_);
  or _28715_ (_05779_, _05778_, _05777_);
  and _28716_ (_05780_, _05779_, _05523_);
  or _28717_ (_05781_, _05780_, _05775_);
  and _28718_ (_05782_, _05053_, _04239_);
  and _28719_ (_05783_, _05782_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  and _28720_ (_05784_, _05783_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  and _28721_ (_05785_, _05784_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  and _28722_ (_05786_, _05785_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  nor _28723_ (_05787_, _05785_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  nor _28724_ (_05788_, _05787_, _05786_);
  nor _28725_ (_05789_, _05788_, _01602_);
  and _28726_ (_05790_, _05788_, _01602_);
  or _28727_ (_05791_, _05790_, _05789_);
  nor _28728_ (_05792_, _05784_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  nor _28729_ (_05793_, _05792_, _05785_);
  nor _28730_ (_05794_, _05793_, _01142_);
  not _28731_ (_05795_, _05786_);
  nor _28732_ (_05796_, _05795_, _05682_);
  or _28733_ (_05797_, _05796_, _05794_);
  and _28734_ (_05798_, _05793_, _01142_);
  and _28735_ (_05799_, _05795_, _05682_);
  or _28736_ (_05800_, _05799_, _05798_);
  or _28737_ (_05801_, _05800_, _05797_);
  nor _28738_ (_05802_, _05782_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor _28739_ (_05803_, _05802_, _05783_);
  nor _28740_ (_05804_, _05803_, _01872_);
  or _28741_ (_05805_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  nand _28742_ (_05806_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  and _28743_ (_05807_, _05806_, _05805_);
  nand _28744_ (_05808_, _05807_, _05783_);
  or _28745_ (_05809_, _05807_, _05783_);
  and _28746_ (_05810_, _05809_, _05808_);
  or _28747_ (_05811_, _05810_, _05804_);
  and _28748_ (_05812_, _05803_, _01872_);
  and _28749_ (_05813_, _05053_, _04237_);
  and _28750_ (_05814_, _05813_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nor _28751_ (_05815_, _05814_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  nor _28752_ (_05816_, _05815_, _05782_);
  and _28753_ (_05817_, _05816_, _01076_);
  or _28754_ (_05818_, _05817_, _05812_);
  or _28755_ (_05819_, _05818_, _05811_);
  nor _28756_ (_05820_, _05813_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nor _28757_ (_05821_, _05820_, _05814_);
  nor _28758_ (_05822_, _05821_, _01106_);
  and _28759_ (_05823_, _05821_, _01106_);
  nor _28760_ (_05824_, _05055_, _04802_);
  and _28761_ (_05825_, _05055_, _04802_);
  or _28762_ (_05826_, _05825_, _05824_);
  nand _28763_ (_05827_, _05717_, _04820_);
  and _28764_ (_05828_, _05059_, _04811_);
  nor _28765_ (_05829_, _05059_, _04811_);
  or _28766_ (_05830_, _05829_, _05828_);
  or _28767_ (_05831_, _05830_, _05827_);
  or _28768_ (_05832_, _05831_, _05826_);
  or _28769_ (_05833_, _05832_, _05823_);
  or _28770_ (_05834_, _05833_, _05822_);
  nor _28771_ (_05835_, _05816_, _01076_);
  or _28772_ (_05836_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nand _28773_ (_05837_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  and _28774_ (_05838_, _05837_, _05836_);
  and _28775_ (_05839_, _05053_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  or _28776_ (_05840_, _05839_, _05838_);
  nand _28777_ (_05841_, _05839_, _05838_);
  and _28778_ (_05842_, _05841_, _05840_);
  nor _28779_ (_05843_, _05053_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nor _28780_ (_05844_, _05843_, _05839_);
  and _28781_ (_05845_, _05844_, _01275_);
  nor _28782_ (_05846_, _05844_, _01275_);
  or _28783_ (_05847_, _05846_, _05845_);
  or _28784_ (_05848_, _05847_, _05842_);
  or _28785_ (_05849_, _05848_, _05835_);
  or _28786_ (_05850_, _05849_, _05834_);
  or _28787_ (_05851_, _05850_, _05819_);
  or _28788_ (_05852_, _05851_, _05801_);
  or _28789_ (_05853_, _05852_, _05791_);
  and _28790_ (_05854_, _05786_, _04245_);
  and _28791_ (_05855_, _05786_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor _28792_ (_05856_, _05855_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  nor _28793_ (_05857_, _05856_, _05854_);
  and _28794_ (_05858_, _05857_, _01591_);
  nor _28795_ (_05859_, _05857_, _01591_);
  or _28796_ (_05860_, _05859_, _05858_);
  or _28797_ (_05861_, _05860_, _05853_);
  and _28798_ (_05862_, _05854_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor _28799_ (_05863_, _05854_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor _28800_ (_05864_, _05863_, _05862_);
  nor _28801_ (_05865_, _05864_, _01580_);
  and _28802_ (_05866_, _05864_, _01580_);
  or _28803_ (_05867_, _05866_, _05865_);
  or _28804_ (_05868_, _05867_, _05861_);
  nor _28805_ (_05869_, _05862_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  and _28806_ (_05870_, _05862_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  nor _28807_ (_05871_, _05870_, _05869_);
  nor _28808_ (_05872_, _05871_, _00584_);
  and _28809_ (_05873_, _05871_, _00584_);
  or _28810_ (_05874_, _05873_, _05872_);
  or _28811_ (_05875_, _05874_, _05868_);
  and _28812_ (_05876_, _05875_, _05781_);
  or _28813_ (_05877_, _05876_, _05770_);
  or _28814_ (_05878_, _05877_, _05629_);
  and _28815_ (_05879_, _05878_, _05173_);
  or _28816_ (_05880_, _04670_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nand _28817_ (_05881_, _04670_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and _28818_ (_05882_, _05881_, _05880_);
  and _28819_ (_05883_, _04709_, _04977_);
  nor _28820_ (_05884_, _04709_, _04977_);
  or _28821_ (_05885_, _05884_, _05883_);
  or _28822_ (_05886_, _05885_, _05882_);
  or _28823_ (_05887_, _04578_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nand _28824_ (_05888_, _04578_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _28825_ (_05889_, _05888_, _05887_);
  and _28826_ (_05890_, _04631_, _04811_);
  nor _28827_ (_05891_, _04631_, _04811_);
  or _28828_ (_05892_, _05891_, _05890_);
  or _28829_ (_05893_, _05892_, _05889_);
  or _28830_ (_05894_, _05893_, _05886_);
  or _28831_ (_05895_, _04476_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nand _28832_ (_05896_, _04476_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  and _28833_ (_05897_, _05896_, _05895_);
  nor _28834_ (_05898_, _04521_, _01275_);
  and _28835_ (_05899_, _04521_, _01275_);
  or _28836_ (_05900_, _05899_, _05898_);
  or _28837_ (_05901_, _05900_, _05897_);
  and _28838_ (_05902_, _04349_, _01076_);
  nor _28839_ (_05903_, _04349_, _01076_);
  or _28840_ (_05904_, _05903_, _05902_);
  nor _28841_ (_05905_, _04431_, _01106_);
  and _28842_ (_05906_, _04431_, _01106_);
  or _28843_ (_05907_, _05906_, _05905_);
  or _28844_ (_05908_, _05907_, _05904_);
  or _28845_ (_05909_, _05908_, _05901_);
  or _28846_ (_05910_, _05909_, _05894_);
  or _28847_ (_05911_, _05479_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nand _28848_ (_05912_, _05479_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  and _28849_ (_05913_, _05912_, _05911_);
  or _28850_ (_05914_, _05913_, _05589_);
  or _28851_ (_05915_, _05306_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nand _28852_ (_05916_, _05306_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  and _28853_ (_05917_, _05916_, _05915_);
  nor _28854_ (_05918_, _05521_, _01150_);
  and _28855_ (_05919_, _05521_, _01150_);
  or _28856_ (_05920_, _05919_, _05918_);
  or _28857_ (_05921_, _05920_, _05917_);
  or _28858_ (_05922_, _05921_, _05914_);
  or _28859_ (_05923_, _05922_, _05586_);
  or _28860_ (_05924_, _05923_, _05910_);
  and _28861_ (_05925_, _05261_, _05537_);
  and _28862_ (_05926_, _05925_, _05435_);
  and _28863_ (_05927_, _05926_, _05173_);
  and _28864_ (_05928_, _05927_, _05924_);
  and _28865_ (_05929_, _05357_, _04586_);
  and _28866_ (_05930_, _05365_, _04585_);
  and _28867_ (_05931_, _05361_, _04235_);
  or _28868_ (_05932_, _05931_, _05930_);
  or _28869_ (_05933_, _05932_, _05929_);
  and _28870_ (_05934_, _05353_, _05057_);
  or _28871_ (_05935_, _05934_, _04526_);
  or _28872_ (_05936_, _05935_, _05933_);
  and _28873_ (_05937_, _05377_, _04586_);
  or _28874_ (_05938_, _05937_, _04525_);
  and _28875_ (_05939_, _05381_, _04235_);
  and _28876_ (_05940_, _05373_, _05057_);
  and _28877_ (_05941_, _05385_, _04585_);
  or _28878_ (_05942_, _05941_, _05940_);
  or _28879_ (_05943_, _05942_, _05939_);
  or _28880_ (_05944_, _05943_, _05938_);
  nand _28881_ (_05945_, _05944_, _05936_);
  nor _28882_ (_05946_, _05945_, _05147_);
  nand _28883_ (_05947_, _05946_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or _28884_ (_05948_, _05946_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and _28885_ (_05949_, _05948_, _05947_);
  and _28886_ (_05950_, _05399_, _04586_);
  or _28887_ (_05951_, _05950_, _04526_);
  and _28888_ (_05952_, _05403_, _04235_);
  and _28889_ (_05953_, _05395_, _05057_);
  and _28890_ (_05954_, _05407_, _04585_);
  or _28891_ (_05955_, _05954_, _05953_);
  or _28892_ (_05956_, _05955_, _05952_);
  or _28893_ (_05957_, _05956_, _05951_);
  and _28894_ (_05958_, _05419_, _04586_);
  or _28895_ (_05959_, _05958_, _04525_);
  and _28896_ (_05960_, _05423_, _04235_);
  and _28897_ (_05961_, _05415_, _05057_);
  and _28898_ (_05962_, _05427_, _04585_);
  or _28899_ (_05963_, _05962_, _05961_);
  or _28900_ (_05964_, _05963_, _05960_);
  or _28901_ (_05965_, _05964_, _05959_);
  nand _28902_ (_05966_, _05965_, _05957_);
  nor _28903_ (_05967_, _05966_, _05147_);
  nor _28904_ (_05968_, _05967_, _04802_);
  and _28905_ (_05969_, _05967_, _04802_);
  or _28906_ (_05970_, _05969_, _05968_);
  or _28907_ (_05971_, _05970_, _05949_);
  and _28908_ (_05972_, _05181_, _04586_);
  or _28909_ (_05973_, _05972_, _04526_);
  and _28910_ (_05974_, _05176_, _04235_);
  and _28911_ (_05975_, _05186_, _05057_);
  and _28912_ (_05976_, _05190_, _04585_);
  or _28913_ (_05977_, _05976_, _05975_);
  or _28914_ (_05978_, _05977_, _05974_);
  or _28915_ (_05979_, _05978_, _05973_);
  and _28916_ (_05980_, _05202_, _04586_);
  or _28917_ (_05981_, _05980_, _04525_);
  and _28918_ (_05982_, _05197_, _04235_);
  and _28919_ (_05983_, _05207_, _05057_);
  and _28920_ (_05984_, _05211_, _04585_);
  or _28921_ (_05985_, _05984_, _05983_);
  or _28922_ (_05986_, _05985_, _05982_);
  or _28923_ (_05987_, _05986_, _05981_);
  nand _28924_ (_05988_, _05987_, _05979_);
  nor _28925_ (_05989_, _05988_, _05147_);
  and _28926_ (_05990_, _05989_, _04827_);
  nor _28927_ (_05991_, _05989_, _04827_);
  or _28928_ (_05992_, _05991_, _05990_);
  and _28929_ (_05993_, _05225_, _04586_);
  or _28930_ (_05994_, _05993_, _04526_);
  and _28931_ (_05995_, _05220_, _04235_);
  and _28932_ (_05996_, _05230_, _05057_);
  and _28933_ (_05997_, _05234_, _04585_);
  or _28934_ (_05998_, _05997_, _05996_);
  or _28935_ (_05999_, _05998_, _05995_);
  or _28936_ (_06000_, _05999_, _05994_);
  and _28937_ (_06001_, _05246_, _04586_);
  or _28938_ (_06002_, _06001_, _04525_);
  and _28939_ (_06003_, _05241_, _04235_);
  and _28940_ (_06004_, _05251_, _05057_);
  and _28941_ (_06005_, _05255_, _04585_);
  or _28942_ (_06006_, _06005_, _06004_);
  or _28943_ (_06007_, _06006_, _06003_);
  or _28944_ (_06008_, _06007_, _06002_);
  nand _28945_ (_06009_, _06008_, _06000_);
  nor _28946_ (_06010_, _06009_, _05147_);
  nor _28947_ (_06011_, _06010_, _04977_);
  and _28948_ (_06012_, _06010_, _04977_);
  or _28949_ (_06013_, _06012_, _06011_);
  or _28950_ (_06014_, _06013_, _05992_);
  or _28951_ (_06015_, _06014_, _05971_);
  not _28952_ (_06016_, _05147_);
  and _28953_ (_06017_, _05313_, _04586_);
  nor _28954_ (_06018_, _06017_, _04526_);
  and _28955_ (_06019_, _05321_, _04235_);
  not _28956_ (_06020_, _06019_);
  and _28957_ (_06021_, _05309_, _05057_);
  and _28958_ (_06022_, _05317_, _04585_);
  nor _28959_ (_06023_, _06022_, _06021_);
  and _28960_ (_06024_, _06023_, _06020_);
  and _28961_ (_06025_, _06024_, _06018_);
  and _28962_ (_06026_, _05337_, _04585_);
  and _28963_ (_06027_, _05333_, _04586_);
  and _28964_ (_06028_, _05341_, _04235_);
  or _28965_ (_06029_, _06028_, _06027_);
  nor _28966_ (_06030_, _06029_, _06026_);
  and _28967_ (_06031_, _05329_, _05057_);
  nor _28968_ (_06032_, _06031_, _04525_);
  and _28969_ (_06033_, _06032_, _06030_);
  nor _28970_ (_06034_, _06033_, _06025_);
  and _28971_ (_06035_, _06034_, _06016_);
  nand _28972_ (_06036_, _06035_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  or _28973_ (_06037_, _06035_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  and _28974_ (_06038_, _06037_, _06036_);
  and _28975_ (_06039_, _05296_, _05057_);
  and _28976_ (_06040_, _05300_, _04585_);
  and _28977_ (_06041_, _05286_, _04235_);
  and _28978_ (_06042_, _05291_, _04586_);
  or _28979_ (_06043_, _06042_, _06041_);
  or _28980_ (_06044_, _06043_, _06040_);
  or _28981_ (_06045_, _06044_, _06039_);
  and _28982_ (_06046_, _06045_, _04526_);
  and _28983_ (_06047_, _05275_, _05057_);
  and _28984_ (_06048_, _05279_, _04585_);
  and _28985_ (_06049_, _05265_, _04235_);
  and _28986_ (_06050_, _05270_, _04586_);
  or _28987_ (_06051_, _06050_, _06049_);
  or _28988_ (_06052_, _06051_, _06048_);
  or _28989_ (_06053_, _06052_, _06047_);
  and _28990_ (_06054_, _06053_, _04525_);
  or _28991_ (_06055_, _06054_, _06046_);
  and _28992_ (_06056_, _06055_, _06016_);
  and _28993_ (_06057_, _06056_, _01128_);
  nor _28994_ (_06058_, _06056_, _01128_);
  or _28995_ (_06059_, _06058_, _06057_);
  or _28996_ (_06060_, _06059_, _06038_);
  and _28997_ (_06061_, _05510_, _04585_);
  and _28998_ (_06062_, _05506_, _04586_);
  nor _28999_ (_06063_, _06062_, _06061_);
  and _29000_ (_06064_, _05502_, _05057_);
  and _29001_ (_06065_, _05514_, _01279_);
  nor _29002_ (_06066_, _06065_, _06064_);
  and _29003_ (_06067_, _06066_, _06063_);
  nor _29004_ (_06068_, _06067_, _04525_);
  and _29005_ (_06069_, _05490_, _04585_);
  and _29006_ (_06070_, _05486_, _04586_);
  nor _29007_ (_06071_, _06070_, _06069_);
  and _29008_ (_06072_, _05482_, _05057_);
  and _29009_ (_06073_, _05494_, _04235_);
  nor _29010_ (_06074_, _06073_, _06072_);
  and _29011_ (_06075_, _06074_, _06071_);
  nor _29012_ (_06076_, _06075_, _04526_);
  nor _29013_ (_06077_, _06076_, _06068_);
  nor _29014_ (_06078_, _06077_, _05147_);
  and _29015_ (_06079_, _06078_, _01106_);
  nor _29016_ (_06080_, _06078_, _01106_);
  or _29017_ (_06081_, _06080_, _06079_);
  and _29018_ (_06082_, _05459_, _01279_);
  and _29019_ (_06083_, _05469_, _05057_);
  and _29020_ (_06084_, _05464_, _04586_);
  and _29021_ (_06085_, _05473_, _04585_);
  or _29022_ (_06086_, _06085_, _06084_);
  or _29023_ (_06087_, _06086_, _06083_);
  or _29024_ (_06088_, _06087_, _06082_);
  and _29025_ (_06089_, _06088_, _04526_);
  and _29026_ (_06090_, _05438_, _04235_);
  and _29027_ (_06091_, _05443_, _04586_);
  and _29028_ (_06092_, _05448_, _05057_);
  and _29029_ (_06093_, _05452_, _04585_);
  or _29030_ (_06094_, _06093_, _06092_);
  or _29031_ (_06095_, _06094_, _06091_);
  or _29032_ (_06096_, _06095_, _06090_);
  and _29033_ (_06097_, _06096_, _04525_);
  or _29034_ (_06098_, _06097_, _06089_);
  and _29035_ (_06099_, _06098_, _06016_);
  nand _29036_ (_06100_, _06099_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  or _29037_ (_06101_, _06099_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  and _29038_ (_06102_, _06101_, _06100_);
  or _29039_ (_06103_, _06102_, _06081_);
  or _29040_ (_06104_, _06103_, _06060_);
  or _29041_ (_06105_, _06104_, _06015_);
  or _29042_ (_06106_, _04670_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nand _29043_ (_06107_, _04670_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and _29044_ (_06108_, _06107_, _06106_);
  nor _29045_ (_06109_, _04709_, _01872_);
  and _29046_ (_06110_, _04709_, _01872_);
  or _29047_ (_06111_, _06110_, _06109_);
  or _29048_ (_06112_, _06111_, _06108_);
  or _29049_ (_06113_, _04578_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nand _29050_ (_06114_, _04578_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and _29051_ (_06115_, _06114_, _06113_);
  and _29052_ (_06116_, _04631_, _01142_);
  nor _29053_ (_06117_, _04631_, _01142_);
  or _29054_ (_06118_, _06117_, _06116_);
  or _29055_ (_06119_, _06118_, _06115_);
  or _29056_ (_06120_, _06119_, _06112_);
  or _29057_ (_06121_, _04476_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nand _29058_ (_06122_, _04476_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and _29059_ (_06123_, _06122_, _06121_);
  nor _29060_ (_06124_, _04521_, _00664_);
  and _29061_ (_06125_, _04521_, _00664_);
  or _29062_ (_06126_, _06125_, _06124_);
  or _29063_ (_06127_, _06126_, _06123_);
  and _29064_ (_06128_, _04349_, _00584_);
  nor _29065_ (_06129_, _04349_, _00584_);
  or _29066_ (_06130_, _06129_, _06128_);
  and _29067_ (_06131_, _04431_, _01580_);
  nor _29068_ (_06132_, _04431_, _01580_);
  or _29069_ (_06133_, _06132_, _06131_);
  or _29070_ (_06134_, _06133_, _06130_);
  or _29071_ (_06135_, _06134_, _06127_);
  or _29072_ (_06136_, _06135_, _06120_);
  or _29073_ (_06137_, _06136_, _06105_);
  and _29074_ (_06138_, _05651_, _05553_);
  and _29075_ (_06139_, _06138_, _05173_);
  and _29076_ (_06140_, _06139_, _06137_);
  or _29077_ (_06141_, _06140_, _05928_);
  or _29078_ (_06142_, _06141_, _05879_);
  or _29079_ (property_invalid, _06142_, _05527_);
  and _29080_ (_06143_, _05167_, first_instr);
  or _29081_ (_00000_, _06143_, rst);
  and _29082_ (_06144_, _07046_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  nor _29083_ (_06145_, _10494_, _07046_);
  or _29084_ (_06146_, _06145_, _06144_);
  and _29085_ (_04894_, _06146_, _06444_);
  and _29086_ (_06147_, _07029_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and _29087_ (_06148_, _06147_, _07026_);
  and _29088_ (_06149_, _07011_, _06996_);
  nor _29089_ (_06150_, _06149_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  nor _29090_ (_06151_, _06150_, _09507_);
  or _29091_ (_06152_, _06151_, _07017_);
  or _29092_ (_06153_, _06152_, _06148_);
  nor _29093_ (_06154_, _07035_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  nor _29094_ (_06155_, _06154_, _06985_);
  and _29095_ (_06156_, _06155_, _06153_);
  nor _29096_ (_06157_, _10494_, _02538_);
  or _29097_ (_06158_, _06157_, _06156_);
  or _29098_ (_06159_, _06158_, _06989_);
  or _29099_ (_06160_, _09503_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and _29100_ (_06161_, _06160_, _06444_);
  and _29101_ (_04910_, _06161_, _06159_);
  and _29102_ (_06162_, _07029_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and _29103_ (_06163_, _06162_, _07026_);
  and _29104_ (_06164_, _02515_, _03116_);
  nor _29105_ (_06165_, _06164_, _06149_);
  or _29106_ (_06166_, _06165_, _07017_);
  or _29107_ (_06167_, _06166_, _06163_);
  or _29108_ (_06168_, _07035_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and _29109_ (_06169_, _06168_, _02538_);
  and _29110_ (_06170_, _06169_, _06167_);
  nor _29111_ (_06171_, _02538_, _06666_);
  or _29112_ (_06172_, _06171_, _06989_);
  or _29113_ (_06173_, _06172_, _06170_);
  nand _29114_ (_06174_, _06989_, _03116_);
  and _29115_ (_06175_, _06174_, _06444_);
  and _29116_ (_04916_, _06175_, _06173_);
  and _29117_ (_06176_, _07011_, _07002_);
  or _29118_ (_06177_, _06176_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and _29119_ (_06178_, _06177_, _04189_);
  and _29120_ (_06179_, _07029_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and _29121_ (_06180_, _06179_, _07026_);
  or _29122_ (_06181_, _06180_, _06178_);
  and _29123_ (_06182_, _06181_, _07035_);
  and _29124_ (_06183_, _07017_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  or _29125_ (_06184_, _06183_, _06985_);
  or _29126_ (_06185_, _06184_, _06182_);
  or _29127_ (_06186_, _02538_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and _29128_ (_06187_, _06186_, _09503_);
  and _29129_ (_06188_, _06187_, _06185_);
  nor _29130_ (_06189_, _07188_, _09503_);
  or _29131_ (_06190_, _06189_, _06188_);
  and _29132_ (_04926_, _06190_, _06444_);
  not _29133_ (_06191_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  nand _29134_ (_06192_, _07011_, _07001_);
  and _29135_ (_06193_, _06192_, _06191_);
  or _29136_ (_06194_, _06193_, _06176_);
  nor _29137_ (_06195_, _07028_, _02903_);
  nand _29138_ (_06196_, _06195_, _07026_);
  and _29139_ (_06197_, _06196_, _06194_);
  nor _29140_ (_06198_, _06197_, _07017_);
  and _29141_ (_06199_, _07017_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  or _29142_ (_06200_, _06199_, _06985_);
  or _29143_ (_06201_, _06200_, _06198_);
  nand _29144_ (_06202_, _06985_, _06191_);
  and _29145_ (_06203_, _06202_, _09503_);
  and _29146_ (_06204_, _06203_, _06201_);
  nor _29147_ (_06205_, _07300_, _09503_);
  or _29148_ (_06206_, _06205_, _06204_);
  and _29149_ (_04935_, _06206_, _06444_);
  and _29150_ (_06207_, _07029_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and _29151_ (_06208_, _06207_, _07026_);
  and _29152_ (_06209_, _07011_, _07000_);
  or _29153_ (_06210_, _06209_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and _29154_ (_06211_, _06210_, _06192_);
  or _29155_ (_06212_, _06211_, _07017_);
  or _29156_ (_06213_, _06212_, _06208_);
  nor _29157_ (_06214_, _07035_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  nor _29158_ (_06215_, _06214_, _06985_);
  and _29159_ (_06216_, _06215_, _06213_);
  and _29160_ (_06217_, _06985_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or _29161_ (_06218_, _06217_, _06989_);
  or _29162_ (_06219_, _06218_, _06216_);
  nand _29163_ (_06220_, _11589_, _06989_);
  and _29164_ (_06221_, _06220_, _06444_);
  and _29165_ (_04937_, _06221_, _06219_);
  and _29166_ (_06222_, _08064_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nor _29167_ (_06223_, _08064_, _01275_);
  or _29168_ (_06224_, _06223_, _06222_);
  and _29169_ (_04943_, _06224_, _06444_);
  and _29170_ (_06225_, _07029_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  and _29171_ (_06226_, _06225_, _07026_);
  and _29172_ (_06227_, _07011_, _06999_);
  nor _29173_ (_06228_, _06227_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  nor _29174_ (_06229_, _06228_, _06209_);
  or _29175_ (_06230_, _06229_, _07017_);
  or _29176_ (_06231_, _06230_, _06226_);
  nor _29177_ (_06232_, _07035_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  nor _29178_ (_06233_, _06232_, _06985_);
  and _29179_ (_06234_, _06233_, _06231_);
  and _29180_ (_06235_, _06985_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  or _29181_ (_06236_, _06235_, _06989_);
  or _29182_ (_06237_, _06236_, _06234_);
  nand _29183_ (_06238_, _07069_, _06989_);
  and _29184_ (_06239_, _06238_, _06444_);
  and _29185_ (_04945_, _06239_, _06237_);
  and _29186_ (_06240_, _08064_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nor _29187_ (_06241_, _08064_, _04802_);
  or _29188_ (_06242_, _06241_, _06240_);
  and _29189_ (_04950_, _06242_, _06444_);
  or _29190_ (_06243_, _00936_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  or _29191_ (_06244_, _03404_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  nand _29192_ (_06245_, _06244_, _06243_);
  nor _29193_ (_06246_, _06245_, _06442_);
  and _29194_ (_06247_, _03410_, _07070_);
  or _29195_ (_06248_, _06247_, _06246_);
  and _29196_ (_06249_, _04154_, _11882_);
  or _29197_ (_06250_, _06249_, _06248_);
  and _29198_ (_04960_, _06250_, _06444_);
  and _29199_ (_06251_, _07029_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  and _29200_ (_06252_, _06251_, _07026_);
  and _29201_ (_06253_, _07011_, _06998_);
  nor _29202_ (_06254_, _06253_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nor _29203_ (_06255_, _06254_, _06227_);
  or _29204_ (_06256_, _06255_, _07017_);
  or _29205_ (_06257_, _06256_, _06252_);
  nor _29206_ (_06258_, _07035_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  nor _29207_ (_06259_, _06258_, _06985_);
  and _29208_ (_06260_, _06259_, _06257_);
  and _29209_ (_06261_, _06985_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  or _29210_ (_06262_, _06261_, _06989_);
  or _29211_ (_06263_, _06262_, _06260_);
  nand _29212_ (_06264_, _09526_, _06989_);
  and _29213_ (_06265_, _06264_, _06444_);
  and _29214_ (_04966_, _06265_, _06263_);
  or _29215_ (_06266_, _00936_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  not _29216_ (_06267_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  nand _29217_ (_06268_, _00936_, _06267_);
  nand _29218_ (_06269_, _06268_, _06266_);
  nor _29219_ (_06270_, _06269_, _06442_);
  and _29220_ (_06271_, _03410_, _09527_);
  or _29221_ (_06272_, _06271_, _06270_);
  and _29222_ (_06273_, _04154_, _07070_);
  or _29223_ (_06274_, _06273_, _06272_);
  and _29224_ (_04984_, _06274_, _06444_);
  or _29225_ (_06275_, _00935_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  nand _29226_ (_06276_, _00935_, _06267_);
  and _29227_ (_06277_, _06276_, _06275_);
  and _29228_ (_06278_, _06277_, _13849_);
  and _29229_ (_06279_, _13847_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  or _29230_ (_06280_, _06279_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  and _29231_ (_06281_, _06280_, _13836_);
  nor _29232_ (_06282_, _06281_, _06278_);
  nor _29233_ (_06283_, _06282_, _06442_);
  and _29234_ (_06284_, _03977_, _09527_);
  or _29235_ (_06285_, _06284_, _06283_);
  and _29236_ (_04986_, _06285_, _06444_);
  and _29237_ (_06286_, _08064_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nor _29238_ (_06287_, _08064_, _04811_);
  or _29239_ (_06288_, _06287_, _06286_);
  and _29240_ (_04990_, _06288_, _06444_);
  and _29241_ (_06289_, _08064_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nor _29242_ (_06290_, _08064_, _04827_);
  or _29243_ (_06291_, _06290_, _06289_);
  and _29244_ (_05020_, _06291_, _06444_);
  and _29245_ (_06292_, _08064_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor _29246_ (_06293_, _08064_, _04977_);
  or _29247_ (_06294_, _06293_, _06292_);
  and _29248_ (_05031_, _06294_, _06444_);
  dff _29249_ (first_instr, _00000_, clk);
  dff _29250_ (\oc8051_symbolic_cxrom1.regarray[10] [0], _14555_, clk);
  dff _29251_ (\oc8051_symbolic_cxrom1.regarray[10] [1], _14556_, clk);
  dff _29252_ (\oc8051_symbolic_cxrom1.regarray[10] [2], _14557_, clk);
  dff _29253_ (\oc8051_symbolic_cxrom1.regarray[10] [3], _14558_, clk);
  dff _29254_ (\oc8051_symbolic_cxrom1.regarray[10] [4], _14559_, clk);
  dff _29255_ (\oc8051_symbolic_cxrom1.regarray[10] [5], _14560_, clk);
  dff _29256_ (\oc8051_symbolic_cxrom1.regarray[10] [6], _14561_, clk);
  dff _29257_ (\oc8051_symbolic_cxrom1.regarray[10] [7], _14562_, clk);
  dff _29258_ (\oc8051_symbolic_cxrom1.regarray[9] [0], _14600_, clk);
  dff _29259_ (\oc8051_symbolic_cxrom1.regarray[9] [1], _14601_, clk);
  dff _29260_ (\oc8051_symbolic_cxrom1.regarray[9] [2], _14602_, clk);
  dff _29261_ (\oc8051_symbolic_cxrom1.regarray[9] [3], _14603_, clk);
  dff _29262_ (\oc8051_symbolic_cxrom1.regarray[9] [4], _14604_, clk);
  dff _29263_ (\oc8051_symbolic_cxrom1.regarray[9] [5], _14605_, clk);
  dff _29264_ (\oc8051_symbolic_cxrom1.regarray[9] [6], _14606_, clk);
  dff _29265_ (\oc8051_symbolic_cxrom1.regarray[9] [7], _14607_, clk);
  dff _29266_ (\oc8051_symbolic_cxrom1.regarray[8] [0], _09446_, clk);
  dff _29267_ (\oc8051_symbolic_cxrom1.regarray[8] [1], _09449_, clk);
  dff _29268_ (\oc8051_symbolic_cxrom1.regarray[8] [2], _14594_, clk);
  dff _29269_ (\oc8051_symbolic_cxrom1.regarray[8] [3], _14595_, clk);
  dff _29270_ (\oc8051_symbolic_cxrom1.regarray[8] [4], _14596_, clk);
  dff _29271_ (\oc8051_symbolic_cxrom1.regarray[8] [5], _14597_, clk);
  dff _29272_ (\oc8051_symbolic_cxrom1.regarray[8] [6], _14598_, clk);
  dff _29273_ (\oc8051_symbolic_cxrom1.regarray[8] [7], _14599_, clk);
  dff _29274_ (\oc8051_symbolic_cxrom1.regarray[7] [0], _14586_, clk);
  dff _29275_ (\oc8051_symbolic_cxrom1.regarray[7] [1], _14587_, clk);
  dff _29276_ (\oc8051_symbolic_cxrom1.regarray[7] [2], _14588_, clk);
  dff _29277_ (\oc8051_symbolic_cxrom1.regarray[7] [3], _14589_, clk);
  dff _29278_ (\oc8051_symbolic_cxrom1.regarray[7] [4], _14590_, clk);
  dff _29279_ (\oc8051_symbolic_cxrom1.regarray[7] [5], _14591_, clk);
  dff _29280_ (\oc8051_symbolic_cxrom1.regarray[7] [6], _14592_, clk);
  dff _29281_ (\oc8051_symbolic_cxrom1.regarray[7] [7], _14593_, clk);
  dff _29282_ (\oc8051_symbolic_cxrom1.regarray[11] [0], _14563_, clk);
  dff _29283_ (\oc8051_symbolic_cxrom1.regarray[11] [1], _14564_, clk);
  dff _29284_ (\oc8051_symbolic_cxrom1.regarray[11] [2], _14565_, clk);
  dff _29285_ (\oc8051_symbolic_cxrom1.regarray[11] [3], _14566_, clk);
  dff _29286_ (\oc8051_symbolic_cxrom1.regarray[11] [4], _14567_, clk);
  dff _29287_ (\oc8051_symbolic_cxrom1.regarray[11] [5], _14568_, clk);
  dff _29288_ (\oc8051_symbolic_cxrom1.regarray[11] [6], _14569_, clk);
  dff _29289_ (\oc8051_symbolic_cxrom1.regarray[11] [7], _14570_, clk);
  dff _29290_ (\oc8051_symbolic_cxrom1.regarray[6] [0], _09240_, clk);
  dff _29291_ (\oc8051_symbolic_cxrom1.regarray[6] [1], _09245_, clk);
  dff _29292_ (\oc8051_symbolic_cxrom1.regarray[6] [2], _09248_, clk);
  dff _29293_ (\oc8051_symbolic_cxrom1.regarray[6] [3], _09253_, clk);
  dff _29294_ (\oc8051_symbolic_cxrom1.regarray[6] [4], _09258_, clk);
  dff _29295_ (\oc8051_symbolic_cxrom1.regarray[6] [5], _09261_, clk);
  dff _29296_ (\oc8051_symbolic_cxrom1.regarray[6] [6], _09265_, clk);
  dff _29297_ (\oc8051_symbolic_cxrom1.regarray[6] [7], _09270_, clk);
  dff _29298_ (\oc8051_symbolic_cxrom1.regarray[5] [0], _09148_, clk);
  dff _29299_ (\oc8051_symbolic_cxrom1.regarray[5] [1], _09150_, clk);
  dff _29300_ (\oc8051_symbolic_cxrom1.regarray[5] [2], _09153_, clk);
  dff _29301_ (\oc8051_symbolic_cxrom1.regarray[5] [3], _09156_, clk);
  dff _29302_ (\oc8051_symbolic_cxrom1.regarray[5] [4], _09159_, clk);
  dff _29303_ (\oc8051_symbolic_cxrom1.regarray[5] [5], _09162_, clk);
  dff _29304_ (\oc8051_symbolic_cxrom1.regarray[5] [6], _09166_, clk);
  dff _29305_ (\oc8051_symbolic_cxrom1.regarray[5] [7], _09170_, clk);
  dff _29306_ (\oc8051_symbolic_cxrom1.regarray[1] [0], _08741_, clk);
  dff _29307_ (\oc8051_symbolic_cxrom1.regarray[1] [1], _08743_, clk);
  dff _29308_ (\oc8051_symbolic_cxrom1.regarray[1] [2], _08745_, clk);
  dff _29309_ (\oc8051_symbolic_cxrom1.regarray[1] [3], _08750_, clk);
  dff _29310_ (\oc8051_symbolic_cxrom1.regarray[1] [4], _08755_, clk);
  dff _29311_ (\oc8051_symbolic_cxrom1.regarray[1] [5], _08757_, clk);
  dff _29312_ (\oc8051_symbolic_cxrom1.regarray[1] [6], _08762_, clk);
  dff _29313_ (\oc8051_symbolic_cxrom1.regarray[1] [7], _08767_, clk);
  dff _29314_ (\oc8051_symbolic_cxrom1.regarray[0] [0], _08621_, clk);
  dff _29315_ (\oc8051_symbolic_cxrom1.regarray[0] [1], _08625_, clk);
  dff _29316_ (\oc8051_symbolic_cxrom1.regarray[0] [2], _08629_, clk);
  dff _29317_ (\oc8051_symbolic_cxrom1.regarray[0] [3], _08633_, clk);
  dff _29318_ (\oc8051_symbolic_cxrom1.regarray[0] [4], _08637_, clk);
  dff _29319_ (\oc8051_symbolic_cxrom1.regarray[0] [5], _08641_, clk);
  dff _29320_ (\oc8051_symbolic_cxrom1.regarray[0] [6], _08647_, clk);
  dff _29321_ (\oc8051_symbolic_cxrom1.regarray[0] [7], _08650_, clk);
  dff _29322_ (\oc8051_symbolic_cxrom1.regarray[3] [0], _14581_, clk);
  dff _29323_ (\oc8051_symbolic_cxrom1.regarray[3] [1], _08943_, clk);
  dff _29324_ (\oc8051_symbolic_cxrom1.regarray[3] [2], _08945_, clk);
  dff _29325_ (\oc8051_symbolic_cxrom1.regarray[3] [3], _08948_, clk);
  dff _29326_ (\oc8051_symbolic_cxrom1.regarray[3] [4], _08951_, clk);
  dff _29327_ (\oc8051_symbolic_cxrom1.regarray[3] [5], _08954_, clk);
  dff _29328_ (\oc8051_symbolic_cxrom1.regarray[3] [6], _08957_, clk);
  dff _29329_ (\oc8051_symbolic_cxrom1.regarray[3] [7], _08960_, clk);
  dff _29330_ (\oc8051_symbolic_cxrom1.regarray[2] [0], _08851_, clk);
  dff _29331_ (\oc8051_symbolic_cxrom1.regarray[2] [1], _08854_, clk);
  dff _29332_ (\oc8051_symbolic_cxrom1.regarray[2] [2], _08858_, clk);
  dff _29333_ (\oc8051_symbolic_cxrom1.regarray[2] [3], _08861_, clk);
  dff _29334_ (\oc8051_symbolic_cxrom1.regarray[2] [4], _08864_, clk);
  dff _29335_ (\oc8051_symbolic_cxrom1.regarray[2] [5], _14580_, clk);
  dff _29336_ (\oc8051_symbolic_cxrom1.regarray[2] [6], _08873_, clk);
  dff _29337_ (\oc8051_symbolic_cxrom1.regarray[2] [7], _08876_, clk);
  dff _29338_ (\oc8051_symbolic_cxrom1.regarray[4] [0], _09044_, clk);
  dff _29339_ (\oc8051_symbolic_cxrom1.regarray[4] [1], _09047_, clk);
  dff _29340_ (\oc8051_symbolic_cxrom1.regarray[4] [2], _14582_, clk);
  dff _29341_ (\oc8051_symbolic_cxrom1.regarray[4] [3], _14583_, clk);
  dff _29342_ (\oc8051_symbolic_cxrom1.regarray[4] [4], _14584_, clk);
  dff _29343_ (\oc8051_symbolic_cxrom1.regarray[4] [5], _14585_, clk);
  dff _29344_ (\oc8051_symbolic_cxrom1.regarray[4] [6], _09058_, clk);
  dff _29345_ (\oc8051_symbolic_cxrom1.regarray[4] [7], _09061_, clk);
  dff _29346_ (\oc8051_symbolic_cxrom1.regvalid [0], _07097_, clk);
  dff _29347_ (\oc8051_symbolic_cxrom1.regvalid [1], _07129_, clk);
  dff _29348_ (\oc8051_symbolic_cxrom1.regvalid [2], _07165_, clk);
  dff _29349_ (\oc8051_symbolic_cxrom1.regvalid [3], _07212_, clk);
  dff _29350_ (\oc8051_symbolic_cxrom1.regvalid [4], _07279_, clk);
  dff _29351_ (\oc8051_symbolic_cxrom1.regvalid [5], _07337_, clk);
  dff _29352_ (\oc8051_symbolic_cxrom1.regvalid [6], _07395_, clk);
  dff _29353_ (\oc8051_symbolic_cxrom1.regvalid [7], _07485_, clk);
  dff _29354_ (\oc8051_symbolic_cxrom1.regvalid [8], _07563_, clk);
  dff _29355_ (\oc8051_symbolic_cxrom1.regvalid [9], _07663_, clk);
  dff _29356_ (\oc8051_symbolic_cxrom1.regvalid [10], _07759_, clk);
  dff _29357_ (\oc8051_symbolic_cxrom1.regvalid [11], _07867_, clk);
  dff _29358_ (\oc8051_symbolic_cxrom1.regvalid [12], _07977_, clk);
  dff _29359_ (\oc8051_symbolic_cxrom1.regvalid [13], _08118_, clk);
  dff _29360_ (\oc8051_symbolic_cxrom1.regvalid [14], _08240_, clk);
  dff _29361_ (\oc8051_symbolic_cxrom1.regvalid [15], _07051_, clk);
  dff _29362_ (\oc8051_symbolic_cxrom1.regarray[15] [0], _14572_, clk);
  dff _29363_ (\oc8051_symbolic_cxrom1.regarray[15] [1], _14573_, clk);
  dff _29364_ (\oc8051_symbolic_cxrom1.regarray[15] [2], _14574_, clk);
  dff _29365_ (\oc8051_symbolic_cxrom1.regarray[15] [3], _14575_, clk);
  dff _29366_ (\oc8051_symbolic_cxrom1.regarray[15] [4], _14576_, clk);
  dff _29367_ (\oc8051_symbolic_cxrom1.regarray[15] [5], _14577_, clk);
  dff _29368_ (\oc8051_symbolic_cxrom1.regarray[15] [6], _14578_, clk);
  dff _29369_ (\oc8051_symbolic_cxrom1.regarray[15] [7], _14579_, clk);
  dff _29370_ (\oc8051_symbolic_cxrom1.regarray[14] [0], _09955_, clk);
  dff _29371_ (\oc8051_symbolic_cxrom1.regarray[14] [1], _09960_, clk);
  dff _29372_ (\oc8051_symbolic_cxrom1.regarray[14] [2], _09964_, clk);
  dff _29373_ (\oc8051_symbolic_cxrom1.regarray[14] [3], _09969_, clk);
  dff _29374_ (\oc8051_symbolic_cxrom1.regarray[14] [4], _09974_, clk);
  dff _29375_ (\oc8051_symbolic_cxrom1.regarray[14] [5], _09976_, clk);
  dff _29376_ (\oc8051_symbolic_cxrom1.regarray[14] [6], _09981_, clk);
  dff _29377_ (\oc8051_symbolic_cxrom1.regarray[14] [7], _09983_, clk);
  dff _29378_ (\oc8051_symbolic_cxrom1.regarray[13] [0], _14571_, clk);
  dff _29379_ (\oc8051_symbolic_cxrom1.regarray[13] [1], _09872_, clk);
  dff _29380_ (\oc8051_symbolic_cxrom1.regarray[13] [2], _09877_, clk);
  dff _29381_ (\oc8051_symbolic_cxrom1.regarray[13] [3], _09880_, clk);
  dff _29382_ (\oc8051_symbolic_cxrom1.regarray[13] [4], _09884_, clk);
  dff _29383_ (\oc8051_symbolic_cxrom1.regarray[13] [5], _09887_, clk);
  dff _29384_ (\oc8051_symbolic_cxrom1.regarray[13] [6], _09890_, clk);
  dff _29385_ (\oc8051_symbolic_cxrom1.regarray[13] [7], _09894_, clk);
  dff _29386_ (\oc8051_symbolic_cxrom1.regarray[12] [0], _09784_, clk);
  dff _29387_ (\oc8051_symbolic_cxrom1.regarray[12] [1], _09786_, clk);
  dff _29388_ (\oc8051_symbolic_cxrom1.regarray[12] [2], _09789_, clk);
  dff _29389_ (\oc8051_symbolic_cxrom1.regarray[12] [3], _09791_, clk);
  dff _29390_ (\oc8051_symbolic_cxrom1.regarray[12] [4], _09793_, clk);
  dff _29391_ (\oc8051_symbolic_cxrom1.regarray[12] [5], _09796_, clk);
  dff _29392_ (\oc8051_symbolic_cxrom1.regarray[12] [6], _09799_, clk);
  dff _29393_ (\oc8051_symbolic_cxrom1.regarray[12] [7], _09801_, clk);
  dff _29394_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _13422_, clk);
  dff _29395_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _13050_, clk);
  dff _29396_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _13046_, clk);
  dff _29397_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _12889_, clk);
  dff _29398_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4], _04074_, clk);
  dff _29399_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5], _04203_, clk);
  dff _29400_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], _04088_, clk);
  dff _29401_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1], _04192_, clk);
  dff _29402_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0], _03293_, clk);
  dff _29403_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1], _11898_, clk);
  dff _29404_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2], _11916_, clk);
  dff _29405_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3], _11913_, clk);
  dff _29406_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4], _04094_, clk);
  dff _29407_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5], _12057_, clk);
  dff _29408_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6], _12317_, clk);
  dff _29409_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7], _04195_, clk);
  dff _29410_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], _11176_, clk);
  dff _29411_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _12304_, clk);
  dff _29412_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0], _11252_, clk);
  dff _29413_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1], _11248_, clk);
  dff _29414_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2], _11222_, clk);
  dff _29415_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3], _11308_, clk);
  dff _29416_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4], _11304_, clk);
  dff _29417_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5], _11298_, clk);
  dff _29418_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6], _11219_, clk);
  dff _29419_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7], _07878_, clk);
  dff _29420_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8], _11141_, clk);
  dff _29421_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9], _11159_, clk);
  dff _29422_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10], _11154_, clk);
  dff _29423_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11], _11239_, clk);
  dff _29424_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12], _11214_, clk);
  dff _29425_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13], _11198_, clk);
  dff _29426_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [0], _06713_, clk);
  dff _29427_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [1], _06715_, clk);
  dff _29428_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [2], _06717_, clk);
  dff _29429_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [3], _06719_, clk);
  dff _29430_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [4], _06721_, clk);
  dff _29431_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [5], _06724_, clk);
  dff _29432_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [6], _06726_, clk);
  dff _29433_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [7], _06566_, clk);
  dff _29434_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [2], _04491_, clk);
  dff _29435_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [7], _06569_, clk);
  dff _29436_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [0], _08694_, clk);
  dff _29437_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [6], _03747_, clk);
  dff _29438_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [7], _00282_, clk);
  dff _29439_ (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], _03794_, clk);
  dff _29440_ (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], _03758_, clk);
  dff _29441_ (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], _03623_, clk);
  dff _29442_ (\oc8051_top_1.oc8051_decoder1.mem_act [0], _03688_, clk);
  dff _29443_ (\oc8051_top_1.oc8051_decoder1.mem_act [1], _03715_, clk);
  dff _29444_ (\oc8051_top_1.oc8051_decoder1.mem_act [2], _03625_, clk);
  dff _29445_ (\oc8051_top_1.oc8051_decoder1.state [0], _03718_, clk);
  dff _29446_ (\oc8051_top_1.oc8051_decoder1.state [1], _03627_, clk);
  dff _29447_ (\oc8051_top_1.oc8051_decoder1.op [0], _03831_, clk);
  dff _29448_ (\oc8051_top_1.oc8051_decoder1.op [1], _03833_, clk);
  dff _29449_ (\oc8051_top_1.oc8051_decoder1.op [2], _03835_, clk);
  dff _29450_ (\oc8051_top_1.oc8051_decoder1.op [3], _03837_, clk);
  dff _29451_ (\oc8051_top_1.oc8051_decoder1.op [4], _03839_, clk);
  dff _29452_ (\oc8051_top_1.oc8051_decoder1.op [5], _03840_, clk);
  dff _29453_ (\oc8051_top_1.oc8051_decoder1.op [6], _03851_, clk);
  dff _29454_ (\oc8051_top_1.oc8051_decoder1.op [7], _03630_, clk);
  dff _29455_ (\oc8051_top_1.oc8051_decoder1.src_sel3 , _03632_, clk);
  dff _29456_ (\oc8051_top_1.oc8051_decoder1.wr_sfr [0], _03537_, clk);
  dff _29457_ (\oc8051_top_1.oc8051_decoder1.wr_sfr [1], _03634_, clk);
  dff _29458_ (\oc8051_top_1.oc8051_decoder1.src_sel2 [0], _03545_, clk);
  dff _29459_ (\oc8051_top_1.oc8051_decoder1.src_sel2 [1], _03637_, clk);
  dff _29460_ (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _03554_, clk);
  dff _29461_ (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _03573_, clk);
  dff _29462_ (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], _03646_, clk);
  dff _29463_ (\oc8051_top_1.oc8051_decoder1.src_sel1 [0], _03710_, clk);
  dff _29464_ (\oc8051_top_1.oc8051_decoder1.src_sel1 [1], _03743_, clk);
  dff _29465_ (\oc8051_top_1.oc8051_decoder1.src_sel1 [2], _03648_, clk);
  dff _29466_ (\oc8051_top_1.oc8051_decoder1.cy_sel [0], _03816_, clk);
  dff _29467_ (\oc8051_top_1.oc8051_decoder1.cy_sel [1], _03653_, clk);
  dff _29468_ (\oc8051_top_1.oc8051_decoder1.alu_op [0], _03981_, clk);
  dff _29469_ (\oc8051_top_1.oc8051_decoder1.alu_op [1], _03989_, clk);
  dff _29470_ (\oc8051_top_1.oc8051_decoder1.alu_op [2], _03994_, clk);
  dff _29471_ (\oc8051_top_1.oc8051_decoder1.alu_op [3], _03656_, clk);
  dff _29472_ (\oc8051_top_1.oc8051_decoder1.psw_set [0], _04011_, clk);
  dff _29473_ (\oc8051_top_1.oc8051_decoder1.psw_set [1], _03658_, clk);
  dff _29474_ (\oc8051_top_1.oc8051_decoder1.wr , _03660_, clk);
  dff _29475_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [0], _03765_, clk);
  dff _29476_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [1], _14515_, clk);
  dff _29477_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [2], _11806_, clk);
  dff _29478_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [3], _09234_, clk);
  dff _29479_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [4], _13300_, clk);
  dff _29480_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [5], _09050_, clk);
  dff _29481_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [6], _04105_, clk);
  dff _29482_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [7], _14356_, clk);
  dff _29483_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [0], _01247_, clk);
  dff _29484_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [1], _04204_, clk);
  dff _29485_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [2], _13148_, clk);
  dff _29486_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [3], _04208_, clk);
  dff _29487_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [4], _02269_, clk);
  dff _29488_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [5], _07623_, clk);
  dff _29489_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [6], _04210_, clk);
  dff _29490_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [7], _04025_, clk);
  dff _29491_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [0], _03036_, clk);
  dff _29492_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [1], _00471_, clk);
  dff _29493_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [2], _10727_, clk);
  dff _29494_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [3], _00509_, clk);
  dff _29495_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [4], _03325_, clk);
  dff _29496_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [5], _12642_, clk);
  dff _29497_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [6], _12351_, clk);
  dff _29498_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [7], _02763_, clk);
  dff _29499_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [0], _03321_, clk);
  dff _29500_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [1], _03357_, clk);
  dff _29501_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [2], _13161_, clk);
  dff _29502_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [3], _01641_, clk);
  dff _29503_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [4], _00504_, clk);
  dff _29504_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [5], _03429_, clk);
  dff _29505_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [6], _01734_, clk);
  dff _29506_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [7], _03986_, clk);
  dff _29507_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [0], _08409_, clk);
  dff _29508_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [1], _07824_, clk);
  dff _29509_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [2], _04095_, clk);
  dff _29510_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [3], _01560_, clk);
  dff _29511_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [4], _12259_, clk);
  dff _29512_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [5], _12465_, clk);
  dff _29513_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [6], _03425_, clk);
  dff _29514_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [7], _02146_, clk);
  dff _29515_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [0], _10802_, clk);
  dff _29516_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [1], _11722_, clk);
  dff _29517_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [2], _03944_, clk);
  dff _29518_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [3], _12752_, clk);
  dff _29519_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [4], _03344_, clk);
  dff _29520_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [5], _03996_, clk);
  dff _29521_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [6], _04894_, clk);
  dff _29522_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [7], _04587_, clk);
  dff _29523_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [0], _02645_, clk);
  dff _29524_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [1], _13387_, clk);
  dff _29525_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [2], _01183_, clk);
  dff _29526_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [3], _08690_, clk);
  dff _29527_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [4], _13150_, clk);
  dff _29528_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [5], _11956_, clk);
  dff _29529_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [6], _09410_, clk);
  dff _29530_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [7], _12599_, clk);
  dff _29531_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [0], _01218_, clk);
  dff _29532_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [1], _12864_, clk);
  dff _29533_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [2], _10905_, clk);
  dff _29534_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [3], _13551_, clk);
  dff _29535_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [4], _07954_, clk);
  dff _29536_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [5], _06471_, clk);
  dff _29537_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [6], _02266_, clk);
  dff _29538_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [7], _01157_, clk);
  dff _29539_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [0], _08075_, clk);
  dff _29540_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [1], _07992_, clk);
  dff _29541_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [2], _07809_, clk);
  dff _29542_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [3], _07964_, clk);
  dff _29543_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [4], _03532_, clk);
  dff _29544_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [0], _05031_, clk);
  dff _29545_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [1], _05020_, clk);
  dff _29546_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [2], _04990_, clk);
  dff _29547_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [3], _04950_, clk);
  dff _29548_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [4], _04943_, clk);
  dff _29549_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [5], _00650_, clk);
  dff _29550_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [6], _04566_, clk);
  dff _29551_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [7], _02945_, clk);
  dff _29552_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [8], _02908_, clk);
  dff _29553_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [9], _02898_, clk);
  dff _29554_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [10], _00676_, clk);
  dff _29555_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [11], _02090_, clk);
  dff _29556_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [12], _01790_, clk);
  dff _29557_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [13], _02042_, clk);
  dff _29558_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [14], _01974_, clk);
  dff _29559_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [15], _14073_, clk);
  dff _29560_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _11397_, clk);
  dff _29561_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _10809_, clk);
  dff _29562_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _00691_, clk);
  dff _29563_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _01394_, clk);
  dff _29564_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _01378_, clk);
  dff _29565_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _00572_, clk);
  dff _29566_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _00569_, clk);
  dff _29567_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _00475_, clk);
  dff _29568_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _00447_, clk);
  dff _29569_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _00688_, clk);
  dff _29570_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _00671_, clk);
  dff _29571_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _06473_, clk);
  dff _29572_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _14524_, clk);
  dff _29573_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _14522_, clk);
  dff _29574_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _14348_, clk);
  dff _29575_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _14207_, clk);
  dff _29576_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [0], _04313_, clk);
  dff _29577_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [1], _04533_, clk);
  dff _29578_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [2], _04362_, clk);
  dff _29579_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [3], _09949_, clk);
  dff _29580_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [4], _09624_, clk);
  dff _29581_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [5], _09742_, clk);
  dff _29582_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [6], _03700_, clk);
  dff _29583_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [7], _03692_, clk);
  dff _29584_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [8], _09962_, clk);
  dff _29585_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [9], _04057_, clk);
  dff _29586_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [10], _04052_, clk);
  dff _29587_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [11], _04050_, clk);
  dff _29588_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [12], _09958_, clk);
  dff _29589_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [13], _03147_, clk);
  dff _29590_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [14], _00724_, clk);
  dff _29591_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [15], _02566_, clk);
  dff _29592_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [16], _01803_, clk);
  dff _29593_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [17], _01708_, clk);
  dff _29594_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [18], _09972_, clk);
  dff _29595_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [19], _03460_, clk);
  dff _29596_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [20], _03502_, clk);
  dff _29597_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [21], _03495_, clk);
  dff _29598_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [22], _09967_, clk);
  dff _29599_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [23], _09619_, clk);
  dff _29600_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [24], _13974_, clk);
  dff _29601_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [25], _13783_, clk);
  dff _29602_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [26], _13897_, clk);
  dff _29603_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [27], _13805_, clk);
  dff _29604_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [28], _09979_, clk);
  dff _29605_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [29], _00434_, clk);
  dff _29606_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [30], _00088_, clk);
  dff _29607_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [31], _13965_, clk);
  dff _29608_ (\oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _14177_, clk);
  dff _29609_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [0], _09996_, clk);
  dff _29610_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [1], _09610_, clk);
  dff _29611_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [2], _09730_, clk);
  dff _29612_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [3], _14055_, clk);
  dff _29613_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [4], _14295_, clk);
  dff _29614_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [5], _01145_, clk);
  dff _29615_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [6], _09849_, clk);
  dff _29616_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [7], _03523_, clk);
  dff _29617_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [0], _09852_, clk);
  dff _29618_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [1], _09673_, clk);
  dff _29619_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [3], _00608_, clk);
  dff _29620_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [4], _09859_, clk);
  dff _29621_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [5], _10040_, clk);
  dff _29622_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [6], _09590_, clk);
  dff _29623_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [1], _09863_, clk);
  dff _29624_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [2], _09668_, clk);
  dff _29625_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [3], _04000_, clk);
  dff _29626_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [4], _03812_, clk);
  dff _29627_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [5], _03802_, clk);
  dff _29628_ (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _00272_, clk);
  dff _29629_ (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _03752_, clk);
  dff _29630_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [0], _10012_, clk);
  dff _29631_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [1], _04582_, clk);
  dff _29632_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _04576_, clk);
  dff _29633_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [3], _04564_, clk);
  dff _29634_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [4], _04562_, clk);
  dff _29635_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [5], _10009_, clk);
  dff _29636_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [6], _09725_, clk);
  dff _29637_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [7], _04131_, clk);
  dff _29638_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [8], _04126_, clk);
  dff _29639_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [9], _04123_, clk);
  dff _29640_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [10], _04113_, clk);
  dff _29641_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [11], _04109_, clk);
  dff _29642_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [12], _10017_, clk);
  dff _29643_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [13], _04226_, clk);
  dff _29644_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [14], _04222_, clk);
  dff _29645_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [15], _03733_, clk);
  dff _29646_ (\oc8051_top_1.oc8051_memory_interface1.pc [0], _03385_, clk);
  dff _29647_ (\oc8051_top_1.oc8051_memory_interface1.pc [1], _03360_, clk);
  dff _29648_ (\oc8051_top_1.oc8051_memory_interface1.pc [2], _03355_, clk);
  dff _29649_ (\oc8051_top_1.oc8051_memory_interface1.pc [3], _10029_, clk);
  dff _29650_ (\oc8051_top_1.oc8051_memory_interface1.pc [4], _03842_, clk);
  dff _29651_ (\oc8051_top_1.oc8051_memory_interface1.pc [5], _03712_, clk);
  dff _29652_ (\oc8051_top_1.oc8051_memory_interface1.pc [6], _03669_, clk);
  dff _29653_ (\oc8051_top_1.oc8051_memory_interface1.pc [7], _03621_, clk);
  dff _29654_ (\oc8051_top_1.oc8051_memory_interface1.pc [8], _10025_, clk);
  dff _29655_ (\oc8051_top_1.oc8051_memory_interface1.pc [9], _09598_, clk);
  dff _29656_ (\oc8051_top_1.oc8051_memory_interface1.pc [10], _02046_, clk);
  dff _29657_ (\oc8051_top_1.oc8051_memory_interface1.pc [11], _01846_, clk);
  dff _29658_ (\oc8051_top_1.oc8051_memory_interface1.pc [12], _02013_, clk);
  dff _29659_ (\oc8051_top_1.oc8051_memory_interface1.pc [13], _01854_, clk);
  dff _29660_ (\oc8051_top_1.oc8051_memory_interface1.pc [14], _01849_, clk);
  dff _29661_ (\oc8051_top_1.oc8051_memory_interface1.pc [15], _03720_, clk);
  dff _29662_ (\oc8051_top_1.oc8051_memory_interface1.int_ack , _13966_, clk);
  dff _29663_ (\oc8051_top_1.oc8051_memory_interface1.int_ack_t , _03309_, clk);
  dff _29664_ (\oc8051_top_1.oc8051_memory_interface1.int_ack_buff , _03331_, clk);
  dff _29665_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], _00999_, clk);
  dff _29666_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], _00976_, clk);
  dff _29667_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _10037_, clk);
  dff _29668_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], _01716_, clk);
  dff _29669_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _01684_, clk);
  dff _29670_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], _01679_, clk);
  dff _29671_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _01676_, clk);
  dff _29672_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _03304_, clk);
  dff _29673_ (\oc8051_top_1.oc8051_memory_interface1.op_pos [0], _09594_, clk);
  dff _29674_ (\oc8051_top_1.oc8051_memory_interface1.op_pos [1], _00655_, clk);
  dff _29675_ (\oc8051_top_1.oc8051_memory_interface1.op_pos [2], _03295_, clk);
  dff _29676_ (\oc8051_top_1.oc8051_memory_interface1.reti , _03428_, clk);
  dff _29677_ (\oc8051_top_1.oc8051_memory_interface1.cdata [0], _10053_, clk);
  dff _29678_ (\oc8051_top_1.oc8051_memory_interface1.cdata [1], _00189_, clk);
  dff _29679_ (\oc8051_top_1.oc8051_memory_interface1.cdata [2], _00151_, clk);
  dff _29680_ (\oc8051_top_1.oc8051_memory_interface1.cdata [3], _00177_, clk);
  dff _29681_ (\oc8051_top_1.oc8051_memory_interface1.cdata [4], _00166_, clk);
  dff _29682_ (\oc8051_top_1.oc8051_memory_interface1.cdata [5], _00164_, clk);
  dff _29683_ (\oc8051_top_1.oc8051_memory_interface1.cdata [6], _00162_, clk);
  dff _29684_ (\oc8051_top_1.oc8051_memory_interface1.cdata [7], _03414_, clk);
  dff _29685_ (\oc8051_top_1.oc8051_memory_interface1.cdone , _03406_, clk);
  dff _29686_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst , _03398_, clk);
  dff _29687_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], _14197_, clk);
  dff _29688_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], _14182_, clk);
  dff _29689_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], _14180_, clk);
  dff _29690_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], _00278_, clk);
  dff _29691_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [0], _13138_, clk);
  dff _29692_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [1], _13108_, clk);
  dff _29693_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [2], _13078_, clk);
  dff _29694_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [3], _13038_, clk);
  dff _29695_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [4], _10345_, clk);
  dff _29696_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [5], _09571_, clk);
  dff _29697_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [6], _12049_, clk);
  dff _29698_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [7], _12027_, clk);
  dff _29699_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [8], _11988_, clk);
  dff _29700_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [9], _10357_, clk);
  dff _29701_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [10], _12409_, clk);
  dff _29702_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [11], _12334_, clk);
  dff _29703_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [12], _12407_, clk);
  dff _29704_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [13], _12380_, clk);
  dff _29705_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [14], _12375_, clk);
  dff _29706_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [15], _12356_, clk);
  dff _29707_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [16], _12341_, clk);
  dff _29708_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [17], _10354_, clk);
  dff _29709_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [18], _09566_, clk);
  dff _29710_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [19], _09708_, clk);
  dff _29711_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [20], _11506_, clk);
  dff _29712_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [21], _11462_, clk);
  dff _29713_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [22], _10364_, clk);
  dff _29714_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [23], _11748_, clk);
  dff _29715_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [24], _11783_, clk);
  dff _29716_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [25], _11768_, clk);
  dff _29717_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [26], _11752_, clk);
  dff _29718_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [27], _10362_, clk);
  dff _29719_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [28], _09561_, clk);
  dff _29720_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [29], _10922_, clk);
  dff _29721_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [30], _01936_, clk);
  dff _29722_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [31], _02583_, clk);
  dff _29723_ (\oc8051_top_1.oc8051_memory_interface1.dmem_wait , _03150_, clk);
  dff _29724_ (\oc8051_top_1.oc8051_memory_interface1.istb_t , _03144_, clk);
  dff _29725_ (\oc8051_top_1.oc8051_memory_interface1.imem_wait , _03132_, clk);
  dff _29726_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _01786_, clk);
  dff _29727_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _01752_, clk);
  dff _29728_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _01697_, clk);
  dff _29729_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _01650_, clk);
  dff _29730_ (\oc8051_top_1.oc8051_memory_interface1.rd_ind , _00287_, clk);
  dff _29731_ (\oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0], clk);
  dff _29732_ (\oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1], clk);
  dff _29733_ (\oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2], clk);
  dff _29734_ (\oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3], clk);
  dff _29735_ (\oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4], clk);
  dff _29736_ (\oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5], clk);
  dff _29737_ (\oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6], clk);
  dff _29738_ (\oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7], clk);
  dff _29739_ (\oc8051_top_1.oc8051_rom1.data_o [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8], clk);
  dff _29740_ (\oc8051_top_1.oc8051_rom1.data_o [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9], clk);
  dff _29741_ (\oc8051_top_1.oc8051_rom1.data_o [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10], clk);
  dff _29742_ (\oc8051_top_1.oc8051_rom1.data_o [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11], clk);
  dff _29743_ (\oc8051_top_1.oc8051_rom1.data_o [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12], clk);
  dff _29744_ (\oc8051_top_1.oc8051_rom1.data_o [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13], clk);
  dff _29745_ (\oc8051_top_1.oc8051_rom1.data_o [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14], clk);
  dff _29746_ (\oc8051_top_1.oc8051_rom1.data_o [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15], clk);
  dff _29747_ (\oc8051_top_1.oc8051_rom1.data_o [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16], clk);
  dff _29748_ (\oc8051_top_1.oc8051_rom1.data_o [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17], clk);
  dff _29749_ (\oc8051_top_1.oc8051_rom1.data_o [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18], clk);
  dff _29750_ (\oc8051_top_1.oc8051_rom1.data_o [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19], clk);
  dff _29751_ (\oc8051_top_1.oc8051_rom1.data_o [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20], clk);
  dff _29752_ (\oc8051_top_1.oc8051_rom1.data_o [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21], clk);
  dff _29753_ (\oc8051_top_1.oc8051_rom1.data_o [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22], clk);
  dff _29754_ (\oc8051_top_1.oc8051_rom1.data_o [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23], clk);
  dff _29755_ (\oc8051_top_1.oc8051_rom1.data_o [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24], clk);
  dff _29756_ (\oc8051_top_1.oc8051_rom1.data_o [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25], clk);
  dff _29757_ (\oc8051_top_1.oc8051_rom1.data_o [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26], clk);
  dff _29758_ (\oc8051_top_1.oc8051_rom1.data_o [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27], clk);
  dff _29759_ (\oc8051_top_1.oc8051_rom1.data_o [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28], clk);
  dff _29760_ (\oc8051_top_1.oc8051_rom1.data_o [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29], clk);
  dff _29761_ (\oc8051_top_1.oc8051_rom1.data_o [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30], clk);
  dff _29762_ (\oc8051_top_1.oc8051_rom1.data_o [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31], clk);
  dff _29763_ (\oc8051_top_1.oc8051_sfr1.pres_ow , _04220_, clk);
  dff _29764_ (\oc8051_top_1.oc8051_sfr1.prescaler [0], _01806_, clk);
  dff _29765_ (\oc8051_top_1.oc8051_sfr1.prescaler [1], _14012_, clk);
  dff _29766_ (\oc8051_top_1.oc8051_sfr1.prescaler [2], _14009_, clk);
  dff _29767_ (\oc8051_top_1.oc8051_sfr1.prescaler [3], _04218_, clk);
  dff _29768_ (\oc8051_top_1.oc8051_sfr1.bit_out , _04214_, clk);
  dff _29769_ (\oc8051_top_1.oc8051_sfr1.wait_data , _04557_, clk);
  dff _29770_ (\oc8051_top_1.oc8051_sfr1.dat0 [0], _01810_, clk);
  dff _29771_ (\oc8051_top_1.oc8051_sfr1.dat0 [1], _13548_, clk);
  dff _29772_ (\oc8051_top_1.oc8051_sfr1.dat0 [2], _13525_, clk);
  dff _29773_ (\oc8051_top_1.oc8051_sfr1.dat0 [3], _13519_, clk);
  dff _29774_ (\oc8051_top_1.oc8051_sfr1.dat0 [4], _01808_, clk);
  dff _29775_ (\oc8051_top_1.oc8051_sfr1.dat0 [5], _01164_, clk);
  dff _29776_ (\oc8051_top_1.oc8051_sfr1.dat0 [6], _13364_, clk);
  dff _29777_ (\oc8051_top_1.oc8051_sfr1.dat0 [7], _04366_, clk);
  dff _29778_ (\oc8051_top_1.oc8051_sfr1.wr_bit_r , _04364_, clk);
  dff _29779_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], _06433_, clk);
  dff _29780_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], _06429_, clk);
  dff _29781_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], _03350_, clk);
  dff _29782_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3], _06536_, clk);
  dff _29783_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4], _06533_, clk);
  dff _29784_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], _06517_, clk);
  dff _29785_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], _03307_, clk);
  dff _29786_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], _09630_, clk);
  dff _29787_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0], _03705_, clk);
  dff _29788_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1], _03804_, clk);
  dff _29789_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2], _03824_, clk);
  dff _29790_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3], _03807_, clk);
  dff _29791_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4], _03678_, clk);
  dff _29792_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5], _03708_, clk);
  dff _29793_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6], _03737_, clk);
  dff _29794_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7], _04377_, clk);
  dff _29795_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], _07710_, clk);
  dff _29796_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], _07705_, clk);
  dff _29797_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], _07702_, clk);
  dff _29798_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], _07678_, clk);
  dff _29799_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], _07658_, clk);
  dff _29800_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], _07648_, clk);
  dff _29801_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], _07645_, clk);
  dff _29802_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7], _13596_, clk);
  dff _29803_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0], _07449_, clk);
  dff _29804_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1], _07514_, clk);
  dff _29805_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2], _07498_, clk);
  dff _29806_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3], _07494_, clk);
  dff _29807_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4], _07469_, clk);
  dff _29808_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5], _07455_, clk);
  dff _29809_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6], _07452_, clk);
  dff _29810_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7], _13589_, clk);
  dff _29811_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff , _02560_, clk);
  dff _29812_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], _00371_, clk);
  dff _29813_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], _00368_, clk);
  dff _29814_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _00350_, clk);
  dff _29815_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3], _00345_, clk);
  dff _29816_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4], _00342_, clk);
  dff _29817_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], _00339_, clk);
  dff _29818_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _00331_, clk);
  dff _29819_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _12487_, clk);
  dff _29820_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], _00326_, clk);
  dff _29821_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _12749_, clk);
  dff _29822_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc , _12769_, clk);
  dff _29823_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _00299_, clk);
  dff _29824_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _00295_, clk);
  dff _29825_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], _03515_, clk);
  dff _29826_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _00276_, clk);
  dff _29827_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _00274_, clk);
  dff _29828_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], _13339_, clk);
  dff _29829_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], _00256_, clk);
  dff _29830_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _00252_, clk);
  dff _29831_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , _04592_, clk);
  dff _29832_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , _04803_, clk);
  dff _29833_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , _04826_, clk);
  dff _29834_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , _01342_, clk);
  dff _29835_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0], _00211_, clk);
  dff _29836_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1], _00205_, clk);
  dff _29837_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2], _00191_, clk);
  dff _29838_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], _04530_, clk);
  dff _29839_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0], _00172_, clk);
  dff _29840_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], _00169_, clk);
  dff _29841_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], _00153_, clk);
  dff _29842_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3], _00143_, clk);
  dff _29843_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4], _00149_, clk);
  dff _29844_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5], _00147_, clk);
  dff _29845_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6], _00145_, clk);
  dff _29846_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _04535_, clk);
  dff _29847_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0], _00085_, clk);
  dff _29848_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1], _00082_, clk);
  dff _29849_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2], _00066_, clk);
  dff _29850_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3], _00064_, clk);
  dff _29851_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4], _00061_, clk);
  dff _29852_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5], _00056_, clk);
  dff _29853_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6], _00038_, clk);
  dff _29854_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7], _04538_, clk);
  dff _29855_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0], _02924_, clk);
  dff _29856_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1], _02893_, clk);
  dff _29857_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2], _03074_, clk);
  dff _29858_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3], _02926_, clk);
  dff _29859_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4], _03072_, clk);
  dff _29860_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5], _02890_, clk);
  dff _29861_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6], _03070_, clk);
  dff _29862_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7], _14416_, clk);
  dff _29863_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0], _02921_, clk);
  dff _29864_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1], _03080_, clk);
  dff _29865_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2], _02888_, clk);
  dff _29866_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3], _03076_, clk);
  dff _29867_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4], _03042_, clk);
  dff _29868_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5], _03040_, clk);
  dff _29869_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6], _02919_, clk);
  dff _29870_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7], _14346_, clk);
  dff _29871_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0], _03084_, clk);
  dff _29872_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1], _02883_, clk);
  dff _29873_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2], _03081_, clk);
  dff _29874_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3], _03046_, clk);
  dff _29875_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4], _03044_, clk);
  dff _29876_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5], _02886_, clk);
  dff _29877_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6], _03078_, clk);
  dff _29878_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7], _07328_, clk);
  dff _29879_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0], _02914_, clk);
  dff _29880_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1], _02879_, clk);
  dff _29881_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2], _03091_, clk);
  dff _29882_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3], _02916_, clk);
  dff _29883_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4], _03088_, clk);
  dff _29884_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5], _02881_, clk);
  dff _29885_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6], _03086_, clk);
  dff _29886_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7], _00501_, clk);
  dff _29887_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1], _03869_, clk);
  dff _29888_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], _03860_, clk);
  dff _29889_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3], _03828_, clk);
  dff _29890_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4], _03784_, clk);
  dff _29891_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5], _03640_, clk);
  dff _29892_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6], _03547_, clk);
  dff _29893_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], _02905_, clk);
  dff _29894_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop , _03196_, clk);
  dff _29895_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], _04806_, clk);
  dff _29896_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], _04808_, clk);
  dff _29897_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2], _04810_, clk);
  dff _29898_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3], _04812_, clk);
  dff _29899_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4], _04814_, clk);
  dff _29900_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5], _04822_, clk);
  dff _29901_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6], _04824_, clk);
  dff _29902_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7], _03300_, clk);
  dff _29903_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , _02670_, clk);
  dff _29904_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff , _02679_, clk);
  dff _29905_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0], _14392_, clk);
  dff _29906_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1], _14040_, clk);
  dff _29907_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2], _14032_, clk);
  dff _29908_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3], _14037_, clk);
  dff _29909_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4], _14026_, clk);
  dff _29910_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], _14021_, clk);
  dff _29911_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6], _14023_, clk);
  dff _29912_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7], _02676_, clk);
  dff _29913_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0], _14047_, clk);
  dff _29914_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1], _13996_, clk);
  dff _29915_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2], _14000_, clk);
  dff _29916_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3], _13988_, clk);
  dff _29917_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4], _13991_, clk);
  dff _29918_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5], _13981_, clk);
  dff _29919_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6], _13978_, clk);
  dff _29920_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7], _02673_, clk);
  dff _29921_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , _02666_, clk);
  dff _29922_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _02664_, clk);
  dff _29923_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0], _13925_, clk);
  dff _29924_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1], _13928_, clk);
  dff _29925_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2], _13834_, clk);
  dff _29926_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3], _13829_, clk);
  dff _29927_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4], _13831_, clk);
  dff _29928_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], _13727_, clk);
  dff _29929_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6], _13721_, clk);
  dff _29930_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7], _02661_, clk);
  dff _29931_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0], _13714_, clk);
  dff _29932_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1], _13747_, clk);
  dff _29933_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2], _13739_, clk);
  dff _29934_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3], _13745_, clk);
  dff _29935_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4], _13742_, clk);
  dff _29936_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5], _13690_, clk);
  dff _29937_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6], _13693_, clk);
  dff _29938_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7], _02652_, clk);
  dff _29939_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 , _02658_, clk);
  dff _29940_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _13675_, clk);
  dff _29941_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], _13637_, clk);
  dff _29942_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2], _13634_, clk);
  dff _29943_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3], _13661_, clk);
  dff _29944_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _13665_, clk);
  dff _29945_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], _13844_, clk);
  dff _29946_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6], _13839_, clk);
  dff _29947_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7], _02649_, clk);
  dff _29948_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r , _10560_, clk);
  dff _29949_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _08140_, clk);
  dff _29950_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , _08189_, clk);
  dff _29951_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r , _08204_, clk);
  dff _29952_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0], _03962_, clk);
  dff _29953_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1], _03958_, clk);
  dff _29954_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2], _03935_, clk);
  dff _29955_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3], _03911_, clk);
  dff _29956_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4], _03923_, clk);
  dff _29957_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5], _03917_, clk);
  dff _29958_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6], _03914_, clk);
  dff _29959_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7], _08719_, clk);
  dff _29960_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0], _03864_, clk);
  dff _29961_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1], _03787_, clk);
  dff _29962_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2], _03821_, clk);
  dff _29963_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3], _03800_, clk);
  dff _29964_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4], _03797_, clk);
  dff _29965_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5], _03791_, clk);
  dff _29966_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6], _03756_, clk);
  dff _29967_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7], _08068_, clk);
  dff _29968_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 , _08149_, clk);
  dff _29969_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0], _03685_, clk);
  dff _29970_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1], _03667_, clk);
  dff _29971_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2], _03663_, clk);
  dff _29972_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3], _03651_, clk);
  dff _29973_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4], _03644_, clk);
  dff _29974_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5], _04916_, clk);
  dff _29975_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6], _04910_, clk);
  dff _29976_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7], _08219_, clk);
  dff _29977_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0], _04966_, clk);
  dff _29978_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1], _04945_, clk);
  dff _29979_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2], _04937_, clk);
  dff _29980_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3], _04935_, clk);
  dff _29981_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4], _04926_, clk);
  dff _29982_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5], _04597_, clk);
  dff _29983_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6], _04595_, clk);
  dff _29984_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7], _11388_, clk);
  dff _29985_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set , _09435_, clk);
  dff _29986_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0], _04555_, clk);
  dff _29987_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1], _04551_, clk);
  dff _29988_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2], _04548_, clk);
  dff _29989_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3], _04545_, clk);
  dff _29990_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], _03606_, clk);
  dff _29991_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], _03599_, clk);
  dff _29992_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6], _03597_, clk);
  dff _29993_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], _09333_, clk);
  dff _29994_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0], _07970_, clk);
  dff _29995_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1], _07876_, clk);
  dff _29996_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2], _07849_, clk);
  dff _29997_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _07863_, clk);
  dff _29998_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _07860_, clk);
  dff _29999_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _07855_, clk);
  dff _30000_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _07852_, clk);
  dff _30001_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _07909_, clk);
  dff _30002_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8], _07934_, clk);
  dff _30003_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9], _07983_, clk);
  dff _30004_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], _07973_, clk);
  dff _30005_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _13023_, clk);
  dff _30006_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf , _12089_, clk);
  dff _30007_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , _12083_, clk);
  dff _30008_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , _00247_, clk);
  dff _30009_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive , _12133_, clk);
  dff _30010_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _12159_, clk);
  dff _30011_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r , _12153_, clk);
  dff _30012_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], _02250_, clk);
  dff _30013_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1], _12143_, clk);
  dff _30014_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], _02236_, clk);
  dff _30015_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], _08701_, clk);
  dff _30016_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _03483_, clk);
  dff _30017_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3], _12140_, clk);
  dff _30018_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0], _00550_, clk);
  dff _30019_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1], _00544_, clk);
  dff _30020_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2], _14544_, clk);
  dff _30021_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3], _14365_, clk);
  dff _30022_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4], _13011_, clk);
  dff _30023_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5], _12870_, clk);
  dff _30024_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6], _11894_, clk);
  dff _30025_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7], _00239_, clk);
  dff _30026_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr , _12010_, clk);
  dff _30027_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr , _12007_, clk);
  dff _30028_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans , _12000_, clk);
  dff _30029_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , _11992_, clk);
  dff _30030_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0], _14257_, clk);
  dff _30031_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1], _10468_, clk);
  dff _30032_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2], _06950_, clk);
  dff _30033_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3], _11985_, clk);
  dff _30034_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0], _04986_, clk);
  dff _30035_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1], _04984_, clk);
  dff _30036_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], _04960_, clk);
  dff _30037_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3], _04590_, clk);
  dff _30038_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4], _04580_, clk);
  dff _30039_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5], _04573_, clk);
  dff _30040_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6], _04383_, clk);
  dff _30041_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7], _04379_, clk);
  dff _30042_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8], _04369_, clk);
  dff _30043_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], _04206_, clk);
  dff _30044_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10], _00280_, clk);
  dff _30045_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0], _03118_, clk);
  dff _30046_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1], _03061_, clk);
  dff _30047_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2], _03049_, clk);
  dff _30048_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3], _02632_, clk);
  dff _30049_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4], _02313_, clk);
  dff _30050_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5], _02191_, clk);
  dff _30051_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6], _02204_, clk);
  dff _30052_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], _12036_, clk);
  dff _30053_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0], _01702_, clk);
  dff _30054_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], _01700_, clk);
  dff _30055_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2], _00629_, clk);
  dff _30056_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3], _01159_, clk);
  dff _30057_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], _00701_, clk);
  dff _30058_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5], _00695_, clk);
  dff _30059_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6], _13754_, clk);
  dff _30060_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], _12053_, clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_for_ajmp [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_out [0], \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_out [1], \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [0], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [1], \oc8051_top_1.oc8051_memory_interface1.imm2_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [2], \oc8051_top_1.oc8051_memory_interface1.imm2_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [3], \oc8051_top_1.oc8051_memory_interface1.imm2_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [4], \oc8051_top_1.oc8051_memory_interface1.imm2_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [5], \oc8051_top_1.oc8051_memory_interface1.imm2_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [6], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [7], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [0], \oc8051_top_1.oc8051_memory_interface1.imm_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [1], \oc8051_top_1.oc8051_memory_interface1.imm_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [2], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [3], \oc8051_top_1.oc8051_memory_interface1.imm_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [4], \oc8051_top_1.oc8051_memory_interface1.imm_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [5], \oc8051_top_1.oc8051_memory_interface1.imm_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [6], \oc8051_top_1.oc8051_memory_interface1.imm_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [7], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [0], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [6], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [7], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [2], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [7], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [0], ABINPUT[1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [1], ABINPUT[2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [2], ABINPUT[3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [3], ABINPUT[4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [4], ABINPUT[5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [5], ABINPUT[6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [6], ABINPUT[7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [7], ABINPUT[8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.oc8051_memory_interface1.bit_in , ABINPUT[0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.rst , rst);
  buf(\oc8051_top_1.oc8051_memory_interface1.clk , clk);
  buf(\oc8051_top_1.oc8051_indi_addr1.wr_bit_r , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_indi_addr1.rst , rst);
  buf(\oc8051_top_1.oc8051_indi_addr1.clk , clk);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.oc8051_rom1.clk , clk);
  buf(\oc8051_top_1.oc8051_rom1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk , clk);
  buf(\oc8051_top_1.oc8051_decoder1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.oc8051_decoder1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.oc8051_decoder1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.ip [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_sfr1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [0], \oc8051_top_1.oc8051_memory_interface1.imm_r [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [1], \oc8051_top_1.oc8051_memory_interface1.imm_r [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [3], \oc8051_top_1.oc8051_memory_interface1.imm_r [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [4], \oc8051_top_1.oc8051_memory_interface1.imm_r [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [5], \oc8051_top_1.oc8051_memory_interface1.imm_r [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [6], \oc8051_top_1.oc8051_memory_interface1.imm_r [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3_r [1], \oc8051_top_1.oc8051_memory_interface1.imm2_r [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3_r [2], \oc8051_top_1.oc8051_memory_interface1.imm2_r [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3_r [3], \oc8051_top_1.oc8051_memory_interface1.imm2_r [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3_r [4], \oc8051_top_1.oc8051_memory_interface1.imm2_r [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3_r [5], \oc8051_top_1.oc8051_memory_interface1.imm2_r [5]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_in , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_symbolic_cxrom1.clk , clk);
  buf(\oc8051_symbolic_cxrom1.rst , rst);
  buf(\oc8051_symbolic_cxrom1.word_in [0], word_in[0]);
  buf(\oc8051_symbolic_cxrom1.word_in [1], word_in[1]);
  buf(\oc8051_symbolic_cxrom1.word_in [2], word_in[2]);
  buf(\oc8051_symbolic_cxrom1.word_in [3], word_in[3]);
  buf(\oc8051_symbolic_cxrom1.word_in [4], word_in[4]);
  buf(\oc8051_symbolic_cxrom1.word_in [5], word_in[5]);
  buf(\oc8051_symbolic_cxrom1.word_in [6], word_in[6]);
  buf(\oc8051_symbolic_cxrom1.word_in [7], word_in[7]);
  buf(\oc8051_symbolic_cxrom1.word_in [8], word_in[8]);
  buf(\oc8051_symbolic_cxrom1.word_in [9], word_in[9]);
  buf(\oc8051_symbolic_cxrom1.word_in [10], word_in[10]);
  buf(\oc8051_symbolic_cxrom1.word_in [11], word_in[11]);
  buf(\oc8051_symbolic_cxrom1.word_in [12], word_in[12]);
  buf(\oc8051_symbolic_cxrom1.word_in [13], word_in[13]);
  buf(\oc8051_symbolic_cxrom1.word_in [14], word_in[14]);
  buf(\oc8051_symbolic_cxrom1.word_in [15], word_in[15]);
  buf(\oc8051_symbolic_cxrom1.word_in [16], word_in[16]);
  buf(\oc8051_symbolic_cxrom1.word_in [17], word_in[17]);
  buf(\oc8051_symbolic_cxrom1.word_in [18], word_in[18]);
  buf(\oc8051_symbolic_cxrom1.word_in [19], word_in[19]);
  buf(\oc8051_symbolic_cxrom1.word_in [20], word_in[20]);
  buf(\oc8051_symbolic_cxrom1.word_in [21], word_in[21]);
  buf(\oc8051_symbolic_cxrom1.word_in [22], word_in[22]);
  buf(\oc8051_symbolic_cxrom1.word_in [23], word_in[23]);
  buf(\oc8051_symbolic_cxrom1.word_in [24], word_in[24]);
  buf(\oc8051_symbolic_cxrom1.word_in [25], word_in[25]);
  buf(\oc8051_symbolic_cxrom1.word_in [26], word_in[26]);
  buf(\oc8051_symbolic_cxrom1.word_in [27], word_in[27]);
  buf(\oc8051_symbolic_cxrom1.word_in [28], word_in[28]);
  buf(\oc8051_symbolic_cxrom1.word_in [29], word_in[29]);
  buf(\oc8051_symbolic_cxrom1.word_in [30], word_in[30]);
  buf(\oc8051_symbolic_cxrom1.word_in [31], word_in[31]);
  buf(\oc8051_symbolic_cxrom1.pc1 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc1 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_symbolic_cxrom1.pc1 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_symbolic_cxrom1.pc1 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_symbolic_cxrom1.pc1 [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_symbolic_cxrom1.pc1 [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_symbolic_cxrom1.pc1 [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_symbolic_cxrom1.pc1 [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_symbolic_cxrom1.pc1 [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_symbolic_cxrom1.pc1 [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_symbolic_cxrom1.pc1 [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_symbolic_cxrom1.pc1 [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_symbolic_cxrom1.pc1 [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_symbolic_cxrom1.pc1 [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_symbolic_cxrom1.pc1 [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_symbolic_cxrom1.pc1 [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_symbolic_cxrom1.pc2 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_symbolic_cxrom1.pc2 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_symbolic_cxrom1.pc2 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_symbolic_cxrom1.pc2 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_symbolic_cxrom1.pc2 [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_symbolic_cxrom1.pc2 [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_symbolic_cxrom1.pc2 [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_symbolic_cxrom1.pc2 [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_symbolic_cxrom1.pc2 [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_symbolic_cxrom1.pc2 [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_symbolic_cxrom1.pc2 [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_symbolic_cxrom1.pc2 [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_symbolic_cxrom1.pc2 [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_symbolic_cxrom1.pc2 [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_symbolic_cxrom1.pc2 [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_symbolic_cxrom1.pc2 [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [0], word_in[0]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [1], word_in[1]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [2], word_in[2]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [3], word_in[3]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [4], word_in[4]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [5], word_in[5]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [6], word_in[6]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [7], word_in[7]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [0], word_in[8]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [1], word_in[9]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [2], word_in[10]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [3], word_in[11]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [4], word_in[12]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [5], word_in[13]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [6], word_in[14]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [7], word_in[15]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [0], word_in[16]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [1], word_in[17]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [2], word_in[18]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [3], word_in[19]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [4], word_in[20]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [5], word_in[21]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [6], word_in[22]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [7], word_in[23]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [0], word_in[24]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [1], word_in[25]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [2], word_in[26]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [3], word_in[27]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [4], word_in[28]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [5], word_in[29]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [6], word_in[30]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [7], word_in[31]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_symbolic_cxrom1.pc10 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc10 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_symbolic_cxrom1.pc10 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_symbolic_cxrom1.pc10 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_symbolic_cxrom1.pc12 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc12 [1], pc1_plus_2[1]);
  buf(\oc8051_symbolic_cxrom1.pc12 [2], pc1_plus_2[2]);
  buf(\oc8051_symbolic_cxrom1.pc12 [3], pc1_plus_2[3]);
  buf(\oc8051_symbolic_cxrom1.pc20 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_symbolic_cxrom1.pc20 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_symbolic_cxrom1.pc20 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_symbolic_cxrom1.pc20 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_symbolic_cxrom1.pc22 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.oc8051_comp1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_comp1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_comp1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_comp1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_comp1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_comp1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_comp1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_comp1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_comp1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_alu1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div1 , \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div0 , \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [4], \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [5], \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.uart_int , \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.t2_int , \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [0], \oc8051_top_1.oc8051_sfr1.psw [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.p , \oc8051_top_1.oc8051_sfr1.psw [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk , clk);
  buf(\oc8051_top_1.ABINPUT [0], ABINPUT[0]);
  buf(\oc8051_top_1.ABINPUT [1], ABINPUT[1]);
  buf(\oc8051_top_1.ABINPUT [2], ABINPUT[2]);
  buf(\oc8051_top_1.ABINPUT [3], ABINPUT[3]);
  buf(\oc8051_top_1.ABINPUT [4], ABINPUT[4]);
  buf(\oc8051_top_1.ABINPUT [5], ABINPUT[5]);
  buf(\oc8051_top_1.ABINPUT [6], ABINPUT[6]);
  buf(\oc8051_top_1.ABINPUT [7], ABINPUT[7]);
  buf(\oc8051_top_1.ABINPUT [8], ABINPUT[8]);
  buf(\oc8051_top_1.wb_rst_i , rst);
  buf(\oc8051_top_1.wb_clk_i , clk);
  buf(\oc8051_top_1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.bit_data , ABINPUT[0]);
  buf(\oc8051_top_1.rd_ind , \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  buf(\oc8051_top_1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.sfr_out [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.sfr_out [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.sfr_out [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.sfr_out [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.sfr_out [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.sfr_out [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.sfr_out [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.sfr_out [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.ram_data [0], ABINPUT[1]);
  buf(\oc8051_top_1.ram_data [1], ABINPUT[2]);
  buf(\oc8051_top_1.ram_data [2], ABINPUT[3]);
  buf(\oc8051_top_1.ram_data [3], ABINPUT[4]);
  buf(\oc8051_top_1.ram_data [4], ABINPUT[5]);
  buf(\oc8051_top_1.ram_data [5], ABINPUT[6]);
  buf(\oc8051_top_1.ram_data [6], ABINPUT[7]);
  buf(\oc8051_top_1.ram_data [7], ABINPUT[8]);
  buf(\oc8051_top_1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.src_sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.src_sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_top_1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_top_1.pc_log [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_top_1.pc_log [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_top_1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_top_1.pc_log [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_top_1.pc_log [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_top_1.pc_log [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_top_1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_top_1.pc_log [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_top_1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_top_1.pc_log [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_top_1.pc_log [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_top_1.pc_log [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_top_1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_top_1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_top_1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_top_1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_top_1.pc_log_prev [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_top_1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_top_1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_top_1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_top_1.pc_log_prev [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_top_1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_top_1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_top_1.pc_log_prev [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_top_1.pc_log_prev [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_top_1.pc_log_prev [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_top_1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_top_1.pc_log_prev [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_top_1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_top_1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.t2ex_i , t2ex_i);
  buf(\oc8051_top_1.t2_i , t2_i);
  buf(\oc8051_top_1.t1_i , t1_i);
  buf(\oc8051_top_1.t0_i , t0_i);
  buf(\oc8051_top_1.rxd_i , rxd_i);
  buf(\oc8051_top_1.p3_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.p3_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.p3_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.p3_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.p3_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.p3_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.p3_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.p3_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.p3_i [0], p3_in[0]);
  buf(\oc8051_top_1.p3_i [1], p3_in[1]);
  buf(\oc8051_top_1.p3_i [2], p3_in[2]);
  buf(\oc8051_top_1.p3_i [3], p3_in[3]);
  buf(\oc8051_top_1.p3_i [4], p3_in[4]);
  buf(\oc8051_top_1.p3_i [5], p3_in[5]);
  buf(\oc8051_top_1.p3_i [6], p3_in[6]);
  buf(\oc8051_top_1.p3_i [7], p3_in[7]);
  buf(\oc8051_top_1.p2_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.p2_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.p2_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.p2_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.p2_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.p2_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.p2_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.p2_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.p2_i [0], p2_in[0]);
  buf(\oc8051_top_1.p2_i [1], p2_in[1]);
  buf(\oc8051_top_1.p2_i [2], p2_in[2]);
  buf(\oc8051_top_1.p2_i [3], p2_in[3]);
  buf(\oc8051_top_1.p2_i [4], p2_in[4]);
  buf(\oc8051_top_1.p2_i [5], p2_in[5]);
  buf(\oc8051_top_1.p2_i [6], p2_in[6]);
  buf(\oc8051_top_1.p2_i [7], p2_in[7]);
  buf(\oc8051_top_1.p1_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.p1_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.p1_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.p1_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.p1_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.p1_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.p1_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.p1_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.p1_i [0], p1_in[0]);
  buf(\oc8051_top_1.p1_i [1], p1_in[1]);
  buf(\oc8051_top_1.p1_i [2], p1_in[2]);
  buf(\oc8051_top_1.p1_i [3], p1_in[3]);
  buf(\oc8051_top_1.p1_i [4], p1_in[4]);
  buf(\oc8051_top_1.p1_i [5], p1_in[5]);
  buf(\oc8051_top_1.p1_i [6], p1_in[6]);
  buf(\oc8051_top_1.p1_i [7], p1_in[7]);
  buf(\oc8051_top_1.p0_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.p0_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.p0_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.p0_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.p0_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.p0_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.p0_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.p0_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.p0_i [0], p0_in[0]);
  buf(\oc8051_top_1.p0_i [1], p0_in[1]);
  buf(\oc8051_top_1.p0_i [2], p0_in[2]);
  buf(\oc8051_top_1.p0_i [3], p0_in[3]);
  buf(\oc8051_top_1.p0_i [4], p0_in[4]);
  buf(\oc8051_top_1.p0_i [5], p0_in[5]);
  buf(\oc8051_top_1.p0_i [6], p0_in[6]);
  buf(\oc8051_top_1.p0_i [7], p0_in[7]);
  buf(\oc8051_top_1.cxrom_data_out [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.cxrom_data_out [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.cxrom_data_out [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.cxrom_data_out [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.cxrom_data_out [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.cxrom_data_out [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.cxrom_data_out [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.cxrom_data_out [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.cxrom_data_out [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.cxrom_data_out [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.cxrom_data_out [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.cxrom_data_out [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.cxrom_data_out [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.cxrom_data_out [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.cxrom_data_out [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.cxrom_data_out [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.cxrom_data_out [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.cxrom_data_out [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.cxrom_data_out [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.cxrom_data_out [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.cxrom_data_out [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.cxrom_data_out [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.cxrom_data_out [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.cxrom_data_out [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.cxrom_data_out [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.cxrom_data_out [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.cxrom_data_out [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.cxrom_data_out [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.cxrom_data_out [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.cxrom_data_out [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.cxrom_data_out [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.cxrom_data_out [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk , clk);
  buf(pc1_plus_2[0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(pc1[0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(pc1[1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(pc1[2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(pc1[3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(pc1[4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(pc1[5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(pc1[6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(pc1[7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(pc1[8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(pc1[9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(pc1[10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(pc1[11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(pc1[12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(pc1[13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(pc1[14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(pc1[15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(pc2[0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(pc2[1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(pc2[2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(pc2[3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(pc2[4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(pc2[5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(pc2[6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(pc2[7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(pc2[8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(pc2[9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(pc2[10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(pc2[11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(pc2[12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(pc2[13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(pc2[14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(pc2[15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(cxrom_data_out[0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(cxrom_data_out[1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(cxrom_data_out[2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(cxrom_data_out[3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(cxrom_data_out[4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(cxrom_data_out[5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(cxrom_data_out[6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(cxrom_data_out[7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(cxrom_data_out[8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(cxrom_data_out[9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(cxrom_data_out[10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(cxrom_data_out[11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(cxrom_data_out[12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(cxrom_data_out[13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(cxrom_data_out[14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(cxrom_data_out[15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(cxrom_data_out[16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(cxrom_data_out[17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(cxrom_data_out[18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(cxrom_data_out[19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(cxrom_data_out[20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(cxrom_data_out[21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(cxrom_data_out[22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(cxrom_data_out[23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(cxrom_data_out[24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(cxrom_data_out[25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(cxrom_data_out[26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(cxrom_data_out[27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(cxrom_data_out[28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(cxrom_data_out[29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(cxrom_data_out[30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(cxrom_data_out[31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk , clk);
  buf(p3_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(p3_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(p3_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(p3_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(p3_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(p3_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(p3_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(p3_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(p2_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(p2_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(p2_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(p2_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(p2_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(p2_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(p2_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(p2_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(p1_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(p1_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(p1_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(p1_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(p1_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(p1_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(p1_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(p1_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(p0_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(p0_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(p0_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(p0_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(p0_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(p0_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(p0_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(p0_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
endmodule
