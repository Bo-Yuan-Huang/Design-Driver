
module oc8051_gm_top(clk, rst, word_in, p0_in, p1_in, p2_in, p3_in, rxd_i, t0_i, t1_i, t2_i, t2ex_i, property_invalid_pc);
  wire _00000_;
  wire _00001_;
  wire _00002_;
  wire _00003_;
  wire _00004_;
  wire _00005_;
  wire _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  wire _08001_;
  wire _08002_;
  wire _08003_;
  wire _08004_;
  wire _08005_;
  wire _08006_;
  wire _08007_;
  wire _08008_;
  wire _08009_;
  wire _08010_;
  wire _08011_;
  wire _08012_;
  wire _08013_;
  wire _08014_;
  wire _08015_;
  wire _08016_;
  wire _08017_;
  wire _08018_;
  wire _08019_;
  wire _08020_;
  wire _08021_;
  wire _08022_;
  wire _08023_;
  wire _08024_;
  wire _08025_;
  wire _08026_;
  wire _08027_;
  wire _08028_;
  wire _08029_;
  wire _08030_;
  wire _08031_;
  wire _08032_;
  wire _08033_;
  wire _08034_;
  wire _08035_;
  wire _08036_;
  wire _08037_;
  wire _08038_;
  wire _08039_;
  wire _08040_;
  wire _08041_;
  wire _08042_;
  wire _08043_;
  wire _08044_;
  wire _08045_;
  wire _08046_;
  wire _08047_;
  wire _08048_;
  wire _08049_;
  wire _08050_;
  wire _08051_;
  wire _08052_;
  wire _08053_;
  wire _08054_;
  wire _08055_;
  wire _08056_;
  wire _08057_;
  wire _08058_;
  wire _08059_;
  wire _08060_;
  wire _08061_;
  wire _08062_;
  wire _08063_;
  wire _08064_;
  wire _08065_;
  wire _08066_;
  wire _08067_;
  wire _08068_;
  wire _08069_;
  wire _08070_;
  wire _08071_;
  wire _08072_;
  wire _08073_;
  wire _08074_;
  wire _08075_;
  wire _08076_;
  wire _08077_;
  wire _08078_;
  wire _08079_;
  wire _08080_;
  wire _08081_;
  wire _08082_;
  wire _08083_;
  wire _08084_;
  wire _08085_;
  wire _08086_;
  wire _08087_;
  wire _08088_;
  wire _08089_;
  wire _08090_;
  wire _08091_;
  wire _08092_;
  wire _08093_;
  wire _08094_;
  wire _08095_;
  wire _08096_;
  wire _08097_;
  wire _08098_;
  wire _08099_;
  wire _08100_;
  wire _08101_;
  wire _08102_;
  wire _08103_;
  wire _08104_;
  wire _08105_;
  wire _08106_;
  wire _08107_;
  wire _08108_;
  wire _08109_;
  wire _08110_;
  wire _08111_;
  wire _08112_;
  wire _08113_;
  wire _08114_;
  wire _08115_;
  wire _08116_;
  wire _08117_;
  wire _08118_;
  wire _08119_;
  wire _08120_;
  wire _08121_;
  wire _08122_;
  wire _08123_;
  wire _08124_;
  wire _08125_;
  wire _08126_;
  wire _08127_;
  wire _08128_;
  wire _08129_;
  wire _08130_;
  wire _08131_;
  wire _08132_;
  wire _08133_;
  wire _08134_;
  wire _08135_;
  wire _08136_;
  wire _08137_;
  wire _08138_;
  wire _08139_;
  wire _08140_;
  wire _08141_;
  wire _08142_;
  wire _08143_;
  wire _08144_;
  wire _08145_;
  wire _08146_;
  wire _08147_;
  wire _08148_;
  wire _08149_;
  wire _08150_;
  wire _08151_;
  wire _08152_;
  wire _08153_;
  wire _08154_;
  wire _08155_;
  wire _08156_;
  wire _08157_;
  wire _08158_;
  wire _08159_;
  wire _08160_;
  wire _08161_;
  wire _08162_;
  wire _08163_;
  wire _08164_;
  wire _08165_;
  wire _08166_;
  wire _08167_;
  wire _08168_;
  wire _08169_;
  wire _08170_;
  wire _08171_;
  wire _08172_;
  wire _08173_;
  wire _08174_;
  wire _08175_;
  wire _08176_;
  wire _08177_;
  wire _08178_;
  wire _08179_;
  wire _08180_;
  wire _08181_;
  wire _08182_;
  wire _08183_;
  wire _08184_;
  wire _08185_;
  wire _08186_;
  wire _08187_;
  wire _08188_;
  wire _08189_;
  wire _08190_;
  wire _08191_;
  wire _08192_;
  wire _08193_;
  wire _08194_;
  wire _08195_;
  wire _08196_;
  wire _08197_;
  wire _08198_;
  wire _08199_;
  wire _08200_;
  wire _08201_;
  wire _08202_;
  wire _08203_;
  wire _08204_;
  wire _08205_;
  wire _08206_;
  wire _08207_;
  wire _08208_;
  wire _08209_;
  wire _08210_;
  wire _08211_;
  wire _08212_;
  wire _08213_;
  wire _08214_;
  wire _08215_;
  wire _08216_;
  wire _08217_;
  wire _08218_;
  wire _08219_;
  wire _08220_;
  wire _08221_;
  wire _08222_;
  wire _08223_;
  wire _08224_;
  wire _08225_;
  wire _08226_;
  wire _08227_;
  wire _08228_;
  wire _08229_;
  wire _08230_;
  wire _08231_;
  wire _08232_;
  wire _08233_;
  wire _08234_;
  wire _08235_;
  wire _08236_;
  wire _08237_;
  wire _08238_;
  wire _08239_;
  wire _08240_;
  wire _08241_;
  wire _08242_;
  wire _08243_;
  wire _08244_;
  wire _08245_;
  wire _08246_;
  wire _08247_;
  wire _08248_;
  wire _08249_;
  wire _08250_;
  wire _08251_;
  wire _08252_;
  wire _08253_;
  wire _08254_;
  wire _08255_;
  wire _08256_;
  wire _08257_;
  wire _08258_;
  wire _08259_;
  wire _08260_;
  wire _08261_;
  wire _08262_;
  wire _08263_;
  wire _08264_;
  wire _08265_;
  wire _08266_;
  wire _08267_;
  wire _08268_;
  wire _08269_;
  wire _08270_;
  wire _08271_;
  wire _08272_;
  wire _08273_;
  wire _08274_;
  wire _08275_;
  wire _08276_;
  wire _08277_;
  wire _08278_;
  wire _08279_;
  wire _08280_;
  wire _08281_;
  wire _08282_;
  wire _08283_;
  wire _08284_;
  wire _08285_;
  wire _08286_;
  wire _08287_;
  wire _08288_;
  wire _08289_;
  wire _08290_;
  wire _08291_;
  wire _08292_;
  wire _08293_;
  wire _08294_;
  wire _08295_;
  wire _08296_;
  wire _08297_;
  wire _08298_;
  wire _08299_;
  wire _08300_;
  wire _08301_;
  wire _08302_;
  wire _08303_;
  wire _08304_;
  wire _08305_;
  wire _08306_;
  wire _08307_;
  wire _08308_;
  wire _08309_;
  wire _08310_;
  wire _08311_;
  wire _08312_;
  wire _08313_;
  wire _08314_;
  wire _08315_;
  wire _08316_;
  wire _08317_;
  wire _08318_;
  wire _08319_;
  wire _08320_;
  wire _08321_;
  wire _08322_;
  wire _08323_;
  wire _08324_;
  wire _08325_;
  wire _08326_;
  wire _08327_;
  wire _08328_;
  wire _08329_;
  wire _08330_;
  wire _08331_;
  wire _08332_;
  wire _08333_;
  wire _08334_;
  wire _08335_;
  wire _08336_;
  wire _08337_;
  wire _08338_;
  wire _08339_;
  wire _08340_;
  wire _08341_;
  wire _08342_;
  wire _08343_;
  wire _08344_;
  wire _08345_;
  wire _08346_;
  wire _08347_;
  wire _08348_;
  wire _08349_;
  wire _08350_;
  wire _08351_;
  wire _08352_;
  wire _08353_;
  wire _08354_;
  wire _08355_;
  wire _08356_;
  wire _08357_;
  wire _08358_;
  wire _08359_;
  wire _08360_;
  wire _08361_;
  wire _08362_;
  wire _08363_;
  wire _08364_;
  wire _08365_;
  wire _08366_;
  wire _08367_;
  wire _08368_;
  wire _08369_;
  wire _08370_;
  wire _08371_;
  wire _08372_;
  wire _08373_;
  wire _08374_;
  wire _08375_;
  wire _08376_;
  wire _08377_;
  wire _08378_;
  wire _08379_;
  wire _08380_;
  wire _08381_;
  wire _08382_;
  wire _08383_;
  wire _08384_;
  wire _08385_;
  wire _08386_;
  wire _08387_;
  wire _08388_;
  wire _08389_;
  wire _08390_;
  wire _08391_;
  wire _08392_;
  wire _08393_;
  wire _08394_;
  wire _08395_;
  wire _08396_;
  wire _08397_;
  wire _08398_;
  wire _08399_;
  wire _08400_;
  wire _08401_;
  wire _08402_;
  wire _08403_;
  wire _08404_;
  wire _08405_;
  wire _08406_;
  wire _08407_;
  wire _08408_;
  wire _08409_;
  wire _08410_;
  wire _08411_;
  wire _08412_;
  wire _08413_;
  wire _08414_;
  wire _08415_;
  wire _08416_;
  wire _08417_;
  wire _08418_;
  wire _08419_;
  wire _08420_;
  wire _08421_;
  wire _08422_;
  wire _08423_;
  wire _08424_;
  wire _08425_;
  wire _08426_;
  wire _08427_;
  wire _08428_;
  wire _08429_;
  wire _08430_;
  wire _08431_;
  wire _08432_;
  wire _08433_;
  wire _08434_;
  wire _08435_;
  wire _08436_;
  wire _08437_;
  wire _08438_;
  wire _08439_;
  wire _08440_;
  wire _08441_;
  wire _08442_;
  wire _08443_;
  wire _08444_;
  wire _08445_;
  wire _08446_;
  wire _08447_;
  wire _08448_;
  wire _08449_;
  wire _08450_;
  wire _08451_;
  wire _08452_;
  wire _08453_;
  wire _08454_;
  wire _08455_;
  wire _08456_;
  wire _08457_;
  wire _08458_;
  wire _08459_;
  wire _08460_;
  wire _08461_;
  wire _08462_;
  wire _08463_;
  wire _08464_;
  wire _08465_;
  wire _08466_;
  wire _08467_;
  wire _08468_;
  wire _08469_;
  wire _08470_;
  wire _08471_;
  wire _08472_;
  wire _08473_;
  wire _08474_;
  wire _08475_;
  wire _08476_;
  wire _08477_;
  wire _08478_;
  wire _08479_;
  wire _08480_;
  wire _08481_;
  wire _08482_;
  wire _08483_;
  wire _08484_;
  wire _08485_;
  wire _08486_;
  wire _08487_;
  wire _08488_;
  wire _08489_;
  wire _08490_;
  wire _08491_;
  wire _08492_;
  wire _08493_;
  wire _08494_;
  wire _08495_;
  wire _08496_;
  wire _08497_;
  wire _08498_;
  wire _08499_;
  wire _08500_;
  wire _08501_;
  wire _08502_;
  wire _08503_;
  wire _08504_;
  wire _08505_;
  wire _08506_;
  wire _08507_;
  wire _08508_;
  wire _08509_;
  wire _08510_;
  wire _08511_;
  wire _08512_;
  wire _08513_;
  wire _08514_;
  wire _08515_;
  wire _08516_;
  wire _08517_;
  wire _08518_;
  wire _08519_;
  wire _08520_;
  wire _08521_;
  wire _08522_;
  wire _08523_;
  wire _08524_;
  wire _08525_;
  wire _08526_;
  wire _08527_;
  wire _08528_;
  wire _08529_;
  wire _08530_;
  wire _08531_;
  wire _08532_;
  wire _08533_;
  wire _08534_;
  wire _08535_;
  wire _08536_;
  wire _08537_;
  wire _08538_;
  wire _08539_;
  wire _08540_;
  wire _08541_;
  wire _08542_;
  wire _08543_;
  wire _08544_;
  wire _08545_;
  wire _08546_;
  wire _08547_;
  wire _08548_;
  wire _08549_;
  wire _08550_;
  wire _08551_;
  wire _08552_;
  wire _08553_;
  wire _08554_;
  wire _08555_;
  wire _08556_;
  wire _08557_;
  wire _08558_;
  wire _08559_;
  wire _08560_;
  wire _08561_;
  wire _08562_;
  wire _08563_;
  wire _08564_;
  wire _08565_;
  wire _08566_;
  wire _08567_;
  wire _08568_;
  wire _08569_;
  wire _08570_;
  wire _08571_;
  wire _08572_;
  wire _08573_;
  wire _08574_;
  wire _08575_;
  wire _08576_;
  wire _08577_;
  wire _08578_;
  wire _08579_;
  wire _08580_;
  wire _08581_;
  wire _08582_;
  wire _08583_;
  wire _08584_;
  wire _08585_;
  wire _08586_;
  wire _08587_;
  wire _08588_;
  wire _08589_;
  wire _08590_;
  wire _08591_;
  wire _08592_;
  wire _08593_;
  wire _08594_;
  wire _08595_;
  wire _08596_;
  wire _08597_;
  wire _08598_;
  wire _08599_;
  wire _08600_;
  wire _08601_;
  wire _08602_;
  wire _08603_;
  wire _08604_;
  wire _08605_;
  wire _08606_;
  wire _08607_;
  wire _08608_;
  wire _08609_;
  wire _08610_;
  wire _08611_;
  wire _08612_;
  wire _08613_;
  wire _08614_;
  wire _08615_;
  wire _08616_;
  wire _08617_;
  wire _08618_;
  wire _08619_;
  wire _08620_;
  wire _08621_;
  wire _08622_;
  wire _08623_;
  wire _08624_;
  wire _08625_;
  wire _08626_;
  wire _08627_;
  wire _08628_;
  wire _08629_;
  wire _08630_;
  wire _08631_;
  wire _08632_;
  wire _08633_;
  wire _08634_;
  wire _08635_;
  wire _08636_;
  wire _08637_;
  wire _08638_;
  wire _08639_;
  wire _08640_;
  wire _08641_;
  wire _08642_;
  wire _08643_;
  wire _08644_;
  wire _08645_;
  wire _08646_;
  wire _08647_;
  wire _08648_;
  wire _08649_;
  wire _08650_;
  wire _08651_;
  wire _08652_;
  wire _08653_;
  wire _08654_;
  wire _08655_;
  wire _08656_;
  wire _08657_;
  wire _08658_;
  wire _08659_;
  wire _08660_;
  wire _08661_;
  wire _08662_;
  wire _08663_;
  wire _08664_;
  wire _08665_;
  wire _08666_;
  wire _08667_;
  wire _08668_;
  wire _08669_;
  wire _08670_;
  wire _08671_;
  wire _08672_;
  wire _08673_;
  wire _08674_;
  wire _08675_;
  wire _08676_;
  wire _08677_;
  wire _08678_;
  wire _08679_;
  wire _08680_;
  wire _08681_;
  wire _08682_;
  wire _08683_;
  wire _08684_;
  wire _08685_;
  wire _08686_;
  wire _08687_;
  wire _08688_;
  wire _08689_;
  wire _08690_;
  wire _08691_;
  wire _08692_;
  wire _08693_;
  wire _08694_;
  wire _08695_;
  wire _08696_;
  wire _08697_;
  wire _08698_;
  wire _08699_;
  wire _08700_;
  wire _08701_;
  wire _08702_;
  wire _08703_;
  wire _08704_;
  wire _08705_;
  wire _08706_;
  wire _08707_;
  wire _08708_;
  wire _08709_;
  wire _08710_;
  wire _08711_;
  wire _08712_;
  wire _08713_;
  wire _08714_;
  wire _08715_;
  wire _08716_;
  wire _08717_;
  wire _08718_;
  wire _08719_;
  wire _08720_;
  wire _08721_;
  wire _08722_;
  wire _08723_;
  wire _08724_;
  wire _08725_;
  wire _08726_;
  wire _08727_;
  wire _08728_;
  wire _08729_;
  wire _08730_;
  wire _08731_;
  wire _08732_;
  wire _08733_;
  wire _08734_;
  wire _08735_;
  wire _08736_;
  wire _08737_;
  wire _08738_;
  wire _08739_;
  wire _08740_;
  wire _08741_;
  wire _08742_;
  wire _08743_;
  wire _08744_;
  wire _08745_;
  wire _08746_;
  wire _08747_;
  wire _08748_;
  wire _08749_;
  wire _08750_;
  wire _08751_;
  wire _08752_;
  wire _08753_;
  wire _08754_;
  wire _08755_;
  wire _08756_;
  wire _08757_;
  wire _08758_;
  wire _08759_;
  wire _08760_;
  wire _08761_;
  wire _08762_;
  wire _08763_;
  wire _08764_;
  wire _08765_;
  wire _08766_;
  wire _08767_;
  wire _08768_;
  wire _08769_;
  wire _08770_;
  wire _08771_;
  wire _08772_;
  wire _08773_;
  wire _08774_;
  wire _08775_;
  wire _08776_;
  wire _08777_;
  wire _08778_;
  wire _08779_;
  wire _08780_;
  wire _08781_;
  wire _08782_;
  wire _08783_;
  wire _08784_;
  wire _08785_;
  wire _08786_;
  wire _08787_;
  wire _08788_;
  wire _08789_;
  wire _08790_;
  wire _08791_;
  wire _08792_;
  wire _08793_;
  wire _08794_;
  wire _08795_;
  wire _08796_;
  wire _08797_;
  wire _08798_;
  wire _08799_;
  wire _08800_;
  wire _08801_;
  wire _08802_;
  wire _08803_;
  wire _08804_;
  wire _08805_;
  wire _08806_;
  wire _08807_;
  wire _08808_;
  wire _08809_;
  wire _08810_;
  wire _08811_;
  wire _08812_;
  wire _08813_;
  wire _08814_;
  wire _08815_;
  wire _08816_;
  wire _08817_;
  wire _08818_;
  wire _08819_;
  wire _08820_;
  wire _08821_;
  wire _08822_;
  wire _08823_;
  wire _08824_;
  wire _08825_;
  wire _08826_;
  wire _08827_;
  wire _08828_;
  wire _08829_;
  wire _08830_;
  wire _08831_;
  wire _08832_;
  wire _08833_;
  wire _08834_;
  wire _08835_;
  wire _08836_;
  wire _08837_;
  wire _08838_;
  wire _08839_;
  wire _08840_;
  wire _08841_;
  wire _08842_;
  wire _08843_;
  wire _08844_;
  wire _08845_;
  wire _08846_;
  wire _08847_;
  wire _08848_;
  wire _08849_;
  wire _08850_;
  wire _08851_;
  wire _08852_;
  wire _08853_;
  wire _08854_;
  wire _08855_;
  wire _08856_;
  wire _08857_;
  wire _08858_;
  wire _08859_;
  wire _08860_;
  wire _08861_;
  wire _08862_;
  wire _08863_;
  wire _08864_;
  wire _08865_;
  wire _08866_;
  wire _08867_;
  wire _08868_;
  wire _08869_;
  wire _08870_;
  wire _08871_;
  wire _08872_;
  wire _08873_;
  wire _08874_;
  wire _08875_;
  wire _08876_;
  wire _08877_;
  wire _08878_;
  wire _08879_;
  wire _08880_;
  wire _08881_;
  wire _08882_;
  wire _08883_;
  wire _08884_;
  wire _08885_;
  wire _08886_;
  wire _08887_;
  wire _08888_;
  wire _08889_;
  wire _08890_;
  wire _08891_;
  wire _08892_;
  wire _08893_;
  wire _08894_;
  wire _08895_;
  wire _08896_;
  wire _08897_;
  wire _08898_;
  wire _08899_;
  wire _08900_;
  wire _08901_;
  wire _08902_;
  wire _08903_;
  wire _08904_;
  wire _08905_;
  wire _08906_;
  wire _08907_;
  wire _08908_;
  wire _08909_;
  wire _08910_;
  wire _08911_;
  wire _08912_;
  wire _08913_;
  wire _08914_;
  wire _08915_;
  wire _08916_;
  wire _08917_;
  wire _08918_;
  wire _08919_;
  wire _08920_;
  wire _08921_;
  wire _08922_;
  wire _08923_;
  wire _08924_;
  wire _08925_;
  wire _08926_;
  wire _08927_;
  wire _08928_;
  wire _08929_;
  wire _08930_;
  wire _08931_;
  wire _08932_;
  wire _08933_;
  wire _08934_;
  wire _08935_;
  wire _08936_;
  wire _08937_;
  wire _08938_;
  wire _08939_;
  wire _08940_;
  wire _08941_;
  wire _08942_;
  wire _08943_;
  wire _08944_;
  wire _08945_;
  wire _08946_;
  wire _08947_;
  wire _08948_;
  wire _08949_;
  wire _08950_;
  wire _08951_;
  wire _08952_;
  wire _08953_;
  wire _08954_;
  wire _08955_;
  wire _08956_;
  wire _08957_;
  wire _08958_;
  wire _08959_;
  wire _08960_;
  wire _08961_;
  wire _08962_;
  wire _08963_;
  wire _08964_;
  wire _08965_;
  wire _08966_;
  wire _08967_;
  wire _08968_;
  wire _08969_;
  wire _08970_;
  wire _08971_;
  wire _08972_;
  wire _08973_;
  wire _08974_;
  wire _08975_;
  wire _08976_;
  wire _08977_;
  wire _08978_;
  wire _08979_;
  wire _08980_;
  wire _08981_;
  wire _08982_;
  wire _08983_;
  wire _08984_;
  wire _08985_;
  wire _08986_;
  wire _08987_;
  wire _08988_;
  wire _08989_;
  wire _08990_;
  wire _08991_;
  wire _08992_;
  wire _08993_;
  wire _08994_;
  wire _08995_;
  wire _08996_;
  wire _08997_;
  wire _08998_;
  wire _08999_;
  wire _09000_;
  wire _09001_;
  wire _09002_;
  wire _09003_;
  wire _09004_;
  wire _09005_;
  wire _09006_;
  wire _09007_;
  wire _09008_;
  wire _09009_;
  wire _09010_;
  wire _09011_;
  wire _09012_;
  wire _09013_;
  wire _09014_;
  wire _09015_;
  wire _09016_;
  wire _09017_;
  wire _09018_;
  wire _09019_;
  wire _09020_;
  wire _09021_;
  wire _09022_;
  wire _09023_;
  wire _09024_;
  wire _09025_;
  wire _09026_;
  wire _09027_;
  wire _09028_;
  wire _09029_;
  wire _09030_;
  wire _09031_;
  wire _09032_;
  wire _09033_;
  wire _09034_;
  wire _09035_;
  wire _09036_;
  wire _09037_;
  wire _09038_;
  wire _09039_;
  wire _09040_;
  wire _09041_;
  wire _09042_;
  wire _09043_;
  wire _09044_;
  wire _09045_;
  wire _09046_;
  wire _09047_;
  wire _09048_;
  wire _09049_;
  wire _09050_;
  wire _09051_;
  wire _09052_;
  wire _09053_;
  wire _09054_;
  wire _09055_;
  wire _09056_;
  wire _09057_;
  wire _09058_;
  wire _09059_;
  wire _09060_;
  wire _09061_;
  wire _09062_;
  wire _09063_;
  wire _09064_;
  wire _09065_;
  wire _09066_;
  wire _09067_;
  wire _09068_;
  wire _09069_;
  wire _09070_;
  wire _09071_;
  wire _09072_;
  wire _09073_;
  wire _09074_;
  wire _09075_;
  wire _09076_;
  wire _09077_;
  wire _09078_;
  wire _09079_;
  wire _09080_;
  wire _09081_;
  wire _09082_;
  wire _09083_;
  wire _09084_;
  wire _09085_;
  wire _09086_;
  wire _09087_;
  wire _09088_;
  wire _09089_;
  wire _09090_;
  wire _09091_;
  wire _09092_;
  wire _09093_;
  wire _09094_;
  wire _09095_;
  wire _09096_;
  wire _09097_;
  wire _09098_;
  wire _09099_;
  wire _09100_;
  wire _09101_;
  wire _09102_;
  wire _09103_;
  wire _09104_;
  wire _09105_;
  wire _09106_;
  wire _09107_;
  wire _09108_;
  wire _09109_;
  wire _09110_;
  wire _09111_;
  wire _09112_;
  wire _09113_;
  wire _09114_;
  wire _09115_;
  wire _09116_;
  wire _09117_;
  wire _09118_;
  wire _09119_;
  wire _09120_;
  wire _09121_;
  wire _09122_;
  wire _09123_;
  wire _09124_;
  wire _09125_;
  wire _09126_;
  wire _09127_;
  wire _09128_;
  wire _09129_;
  wire _09130_;
  wire _09131_;
  wire _09132_;
  wire _09133_;
  wire _09134_;
  wire _09135_;
  wire _09136_;
  wire _09137_;
  wire _09138_;
  wire _09139_;
  wire _09140_;
  wire _09141_;
  wire _09142_;
  wire _09143_;
  wire _09144_;
  wire _09145_;
  wire _09146_;
  wire _09147_;
  wire _09148_;
  wire _09149_;
  wire _09150_;
  wire _09151_;
  wire _09152_;
  wire _09153_;
  wire _09154_;
  wire _09155_;
  wire _09156_;
  wire _09157_;
  wire _09158_;
  wire _09159_;
  wire _09160_;
  wire _09161_;
  wire _09162_;
  wire _09163_;
  wire _09164_;
  wire _09165_;
  wire _09166_;
  wire _09167_;
  wire _09168_;
  wire _09169_;
  wire _09170_;
  wire _09171_;
  wire _09172_;
  wire _09173_;
  wire _09174_;
  wire _09175_;
  wire _09176_;
  wire _09177_;
  wire _09178_;
  wire _09179_;
  wire _09180_;
  wire _09181_;
  wire _09182_;
  wire _09183_;
  wire _09184_;
  wire _09185_;
  wire _09186_;
  wire _09187_;
  wire _09188_;
  wire _09189_;
  wire _09190_;
  wire _09191_;
  wire _09192_;
  wire _09193_;
  wire _09194_;
  wire _09195_;
  wire _09196_;
  wire _09197_;
  wire _09198_;
  wire _09199_;
  wire _09200_;
  wire _09201_;
  wire _09202_;
  wire _09203_;
  wire _09204_;
  wire _09205_;
  wire _09206_;
  wire _09207_;
  wire _09208_;
  wire _09209_;
  wire _09210_;
  wire _09211_;
  wire _09212_;
  wire _09213_;
  wire _09214_;
  wire _09215_;
  wire _09216_;
  wire _09217_;
  wire _09218_;
  wire _09219_;
  wire _09220_;
  wire _09221_;
  wire _09222_;
  wire _09223_;
  wire _09224_;
  wire _09225_;
  wire _09226_;
  wire _09227_;
  wire _09228_;
  wire _09229_;
  wire _09230_;
  wire _09231_;
  wire _09232_;
  wire _09233_;
  wire _09234_;
  wire _09235_;
  wire _09236_;
  wire _09237_;
  wire _09238_;
  wire _09239_;
  wire _09240_;
  wire _09241_;
  wire _09242_;
  wire _09243_;
  wire _09244_;
  wire _09245_;
  wire _09246_;
  wire _09247_;
  wire _09248_;
  wire _09249_;
  wire _09250_;
  wire _09251_;
  wire _09252_;
  wire _09253_;
  wire _09254_;
  wire _09255_;
  wire _09256_;
  wire _09257_;
  wire _09258_;
  wire _09259_;
  wire _09260_;
  wire _09261_;
  wire _09262_;
  wire _09263_;
  wire _09264_;
  wire _09265_;
  wire _09266_;
  wire _09267_;
  wire _09268_;
  wire _09269_;
  wire _09270_;
  wire _09271_;
  wire _09272_;
  wire _09273_;
  wire _09274_;
  wire _09275_;
  wire _09276_;
  wire _09277_;
  wire _09278_;
  wire _09279_;
  wire _09280_;
  wire _09281_;
  wire _09282_;
  wire _09283_;
  wire _09284_;
  wire _09285_;
  wire _09286_;
  wire _09287_;
  wire _09288_;
  wire _09289_;
  wire _09290_;
  wire _09291_;
  wire _09292_;
  wire _09293_;
  wire _09294_;
  wire _09295_;
  wire _09296_;
  wire _09297_;
  wire _09298_;
  wire _09299_;
  wire _09300_;
  wire _09301_;
  wire _09302_;
  wire _09303_;
  wire _09304_;
  wire _09305_;
  wire _09306_;
  wire _09307_;
  wire _09308_;
  wire _09309_;
  wire _09310_;
  wire _09311_;
  wire _09312_;
  wire _09313_;
  wire _09314_;
  wire _09315_;
  wire _09316_;
  wire _09317_;
  wire _09318_;
  wire _09319_;
  wire _09320_;
  wire _09321_;
  wire _09322_;
  wire _09323_;
  wire _09324_;
  wire _09325_;
  wire _09326_;
  wire _09327_;
  wire _09328_;
  wire _09329_;
  wire _09330_;
  wire _09331_;
  wire _09332_;
  wire _09333_;
  wire _09334_;
  wire _09335_;
  wire _09336_;
  wire _09337_;
  wire _09338_;
  wire _09339_;
  wire _09340_;
  wire _09341_;
  wire _09342_;
  wire _09343_;
  wire _09344_;
  wire _09345_;
  wire _09346_;
  wire _09347_;
  wire _09348_;
  wire _09349_;
  wire _09350_;
  wire _09351_;
  wire _09352_;
  wire _09353_;
  wire _09354_;
  wire _09355_;
  wire _09356_;
  wire _09357_;
  wire _09358_;
  wire _09359_;
  wire _09360_;
  wire _09361_;
  wire _09362_;
  wire _09363_;
  wire _09364_;
  wire _09365_;
  wire _09366_;
  wire _09367_;
  wire _09368_;
  wire _09369_;
  wire _09370_;
  wire _09371_;
  wire _09372_;
  wire _09373_;
  wire _09374_;
  wire _09375_;
  wire _09376_;
  wire _09377_;
  wire _09378_;
  wire _09379_;
  wire _09380_;
  wire _09381_;
  wire _09382_;
  wire _09383_;
  wire _09384_;
  wire _09385_;
  wire _09386_;
  wire _09387_;
  wire _09388_;
  wire _09389_;
  wire _09390_;
  wire _09391_;
  wire _09392_;
  wire _09393_;
  wire _09394_;
  wire _09395_;
  wire _09396_;
  wire _09397_;
  wire _09398_;
  wire _09399_;
  wire _09400_;
  wire _09401_;
  wire _09402_;
  wire _09403_;
  wire _09404_;
  wire _09405_;
  wire _09406_;
  wire _09407_;
  wire _09408_;
  wire _09409_;
  wire _09410_;
  wire _09411_;
  wire _09412_;
  wire _09413_;
  wire _09414_;
  wire _09415_;
  wire _09416_;
  wire _09417_;
  wire _09418_;
  wire _09419_;
  wire _09420_;
  wire _09421_;
  wire _09422_;
  wire _09423_;
  wire _09424_;
  wire _09425_;
  wire _09426_;
  wire _09427_;
  wire _09428_;
  wire _09429_;
  wire _09430_;
  wire _09431_;
  wire _09432_;
  wire _09433_;
  wire _09434_;
  wire _09435_;
  wire _09436_;
  wire _09437_;
  wire _09438_;
  wire _09439_;
  wire _09440_;
  wire _09441_;
  wire _09442_;
  wire _09443_;
  wire _09444_;
  wire _09445_;
  wire _09446_;
  wire _09447_;
  wire _09448_;
  wire _09449_;
  wire _09450_;
  wire _09451_;
  wire _09452_;
  wire _09453_;
  wire _09454_;
  wire _09455_;
  wire _09456_;
  wire _09457_;
  wire _09458_;
  wire _09459_;
  wire _09460_;
  wire _09461_;
  wire _09462_;
  wire _09463_;
  wire _09464_;
  wire _09465_;
  wire _09466_;
  wire _09467_;
  wire _09468_;
  wire _09469_;
  wire _09470_;
  wire _09471_;
  wire _09472_;
  wire _09473_;
  wire _09474_;
  wire _09475_;
  wire _09476_;
  wire _09477_;
  wire _09478_;
  wire _09479_;
  wire _09480_;
  wire _09481_;
  wire _09482_;
  wire _09483_;
  wire _09484_;
  wire _09485_;
  wire _09486_;
  wire _09487_;
  wire _09488_;
  wire _09489_;
  wire _09490_;
  wire _09491_;
  wire _09492_;
  wire _09493_;
  wire _09494_;
  wire _09495_;
  wire _09496_;
  wire _09497_;
  wire _09498_;
  wire _09499_;
  wire _09500_;
  wire _09501_;
  wire _09502_;
  wire _09503_;
  wire _09504_;
  wire _09505_;
  wire _09506_;
  wire _09507_;
  wire _09508_;
  wire _09509_;
  wire _09510_;
  wire _09511_;
  wire _09512_;
  wire _09513_;
  wire _09514_;
  wire _09515_;
  wire _09516_;
  wire _09517_;
  wire _09518_;
  wire _09519_;
  wire _09520_;
  wire _09521_;
  wire _09522_;
  wire _09523_;
  wire _09524_;
  wire _09525_;
  wire _09526_;
  wire _09527_;
  wire _09528_;
  wire _09529_;
  wire _09530_;
  wire _09531_;
  wire _09532_;
  wire _09533_;
  wire _09534_;
  wire _09535_;
  wire _09536_;
  wire _09537_;
  wire _09538_;
  wire _09539_;
  wire _09540_;
  wire _09541_;
  wire _09542_;
  wire _09543_;
  wire _09544_;
  wire _09545_;
  wire _09546_;
  wire _09547_;
  wire _09548_;
  wire _09549_;
  wire _09550_;
  wire _09551_;
  wire _09552_;
  wire _09553_;
  wire _09554_;
  wire _09555_;
  wire _09556_;
  wire _09557_;
  wire _09558_;
  wire _09559_;
  wire _09560_;
  wire _09561_;
  wire _09562_;
  wire _09563_;
  wire _09564_;
  wire _09565_;
  wire _09566_;
  wire _09567_;
  wire _09568_;
  wire _09569_;
  wire _09570_;
  wire _09571_;
  wire _09572_;
  wire _09573_;
  wire _09574_;
  wire _09575_;
  wire _09576_;
  wire _09577_;
  wire _09578_;
  wire _09579_;
  wire _09580_;
  wire _09581_;
  wire _09582_;
  wire _09583_;
  wire _09584_;
  wire _09585_;
  wire _09586_;
  wire _09587_;
  wire _09588_;
  wire _09589_;
  wire _09590_;
  wire _09591_;
  wire _09592_;
  wire _09593_;
  wire _09594_;
  wire _09595_;
  wire _09596_;
  wire _09597_;
  wire _09598_;
  wire _09599_;
  wire _09600_;
  wire _09601_;
  wire _09602_;
  wire _09603_;
  wire _09604_;
  wire _09605_;
  wire _09606_;
  wire _09607_;
  wire _09608_;
  wire _09609_;
  wire _09610_;
  wire _09611_;
  wire _09612_;
  wire _09613_;
  wire _09614_;
  wire _09615_;
  wire _09616_;
  wire _09617_;
  wire _09618_;
  wire _09619_;
  wire _09620_;
  wire _09621_;
  wire _09622_;
  wire _09623_;
  wire _09624_;
  wire _09625_;
  wire _09626_;
  wire _09627_;
  wire _09628_;
  wire _09629_;
  wire _09630_;
  wire _09631_;
  wire _09632_;
  wire _09633_;
  wire _09634_;
  wire _09635_;
  wire _09636_;
  wire _09637_;
  wire _09638_;
  wire _09639_;
  wire _09640_;
  wire _09641_;
  wire _09642_;
  wire _09643_;
  wire _09644_;
  wire _09645_;
  wire _09646_;
  wire _09647_;
  wire _09648_;
  wire _09649_;
  wire _09650_;
  wire _09651_;
  wire _09652_;
  wire _09653_;
  wire _09654_;
  wire _09655_;
  wire _09656_;
  wire _09657_;
  wire _09658_;
  wire _09659_;
  wire _09660_;
  wire _09661_;
  wire _09662_;
  wire _09663_;
  wire _09664_;
  wire _09665_;
  wire _09666_;
  wire _09667_;
  wire _09668_;
  wire _09669_;
  wire _09670_;
  wire _09671_;
  wire _09672_;
  wire _09673_;
  wire _09674_;
  wire _09675_;
  wire _09676_;
  wire _09677_;
  wire _09678_;
  wire _09679_;
  wire _09680_;
  wire _09681_;
  wire _09682_;
  wire _09683_;
  wire _09684_;
  wire _09685_;
  wire _09686_;
  wire _09687_;
  wire _09688_;
  wire _09689_;
  wire _09690_;
  wire _09691_;
  wire _09692_;
  wire _09693_;
  wire _09694_;
  wire _09695_;
  wire _09696_;
  wire _09697_;
  wire _09698_;
  wire _09699_;
  wire _09700_;
  wire _09701_;
  wire _09702_;
  wire _09703_;
  wire _09704_;
  wire _09705_;
  wire _09706_;
  wire _09707_;
  wire _09708_;
  wire _09709_;
  wire _09710_;
  wire _09711_;
  wire _09712_;
  wire _09713_;
  wire _09714_;
  wire _09715_;
  wire _09716_;
  wire _09717_;
  wire _09718_;
  wire _09719_;
  wire _09720_;
  wire _09721_;
  wire _09722_;
  wire _09723_;
  wire _09724_;
  wire _09725_;
  wire _09726_;
  wire _09727_;
  wire _09728_;
  wire _09729_;
  wire _09730_;
  wire _09731_;
  wire _09732_;
  wire _09733_;
  wire _09734_;
  wire _09735_;
  wire _09736_;
  wire _09737_;
  wire _09738_;
  wire _09739_;
  wire _09740_;
  wire _09741_;
  wire _09742_;
  wire _09743_;
  wire _09744_;
  wire _09745_;
  wire _09746_;
  wire _09747_;
  wire _09748_;
  wire _09749_;
  wire _09750_;
  wire _09751_;
  wire _09752_;
  wire _09753_;
  wire _09754_;
  wire _09755_;
  wire _09756_;
  wire _09757_;
  wire _09758_;
  wire _09759_;
  wire _09760_;
  wire _09761_;
  wire _09762_;
  wire _09763_;
  wire _09764_;
  wire _09765_;
  wire _09766_;
  wire _09767_;
  wire _09768_;
  wire _09769_;
  wire _09770_;
  wire _09771_;
  wire _09772_;
  wire _09773_;
  wire _09774_;
  wire _09775_;
  wire _09776_;
  wire _09777_;
  wire _09778_;
  wire _09779_;
  wire _09780_;
  wire _09781_;
  wire _09782_;
  wire _09783_;
  wire _09784_;
  wire _09785_;
  wire _09786_;
  wire _09787_;
  wire _09788_;
  wire _09789_;
  wire _09790_;
  wire _09791_;
  wire _09792_;
  wire _09793_;
  wire _09794_;
  wire _09795_;
  wire _09796_;
  wire _09797_;
  wire _09798_;
  wire _09799_;
  wire _09800_;
  wire _09801_;
  wire _09802_;
  wire _09803_;
  wire _09804_;
  wire _09805_;
  wire _09806_;
  wire _09807_;
  wire _09808_;
  wire _09809_;
  wire _09810_;
  wire _09811_;
  wire _09812_;
  wire _09813_;
  wire _09814_;
  wire _09815_;
  wire _09816_;
  wire _09817_;
  wire _09818_;
  wire _09819_;
  wire _09820_;
  wire _09821_;
  wire _09822_;
  wire _09823_;
  wire _09824_;
  wire _09825_;
  wire _09826_;
  wire _09827_;
  wire _09828_;
  wire _09829_;
  wire _09830_;
  wire _09831_;
  wire _09832_;
  wire _09833_;
  wire _09834_;
  wire _09835_;
  wire _09836_;
  wire _09837_;
  wire _09838_;
  wire _09839_;
  wire _09840_;
  wire _09841_;
  wire _09842_;
  wire _09843_;
  wire _09844_;
  wire _09845_;
  wire _09846_;
  wire _09847_;
  wire _09848_;
  wire _09849_;
  wire _09850_;
  wire _09851_;
  wire _09852_;
  wire _09853_;
  wire _09854_;
  wire _09855_;
  wire _09856_;
  wire _09857_;
  wire _09858_;
  wire _09859_;
  wire _09860_;
  wire _09861_;
  wire _09862_;
  wire _09863_;
  wire _09864_;
  wire _09865_;
  wire _09866_;
  wire _09867_;
  wire _09868_;
  wire _09869_;
  wire _09870_;
  wire _09871_;
  wire _09872_;
  wire _09873_;
  wire _09874_;
  wire _09875_;
  wire _09876_;
  wire _09877_;
  wire _09878_;
  wire _09879_;
  wire _09880_;
  wire _09881_;
  wire _09882_;
  wire _09883_;
  wire _09884_;
  wire _09885_;
  wire _09886_;
  wire _09887_;
  wire _09888_;
  wire _09889_;
  wire _09890_;
  wire _09891_;
  wire _09892_;
  wire _09893_;
  wire _09894_;
  wire _09895_;
  wire _09896_;
  wire _09897_;
  wire _09898_;
  wire _09899_;
  wire _09900_;
  wire _09901_;
  wire _09902_;
  wire _09903_;
  wire _09904_;
  wire _09905_;
  wire _09906_;
  wire _09907_;
  wire _09908_;
  wire _09909_;
  wire _09910_;
  wire _09911_;
  wire _09912_;
  wire _09913_;
  wire _09914_;
  wire _09915_;
  wire _09916_;
  wire _09917_;
  wire _09918_;
  wire _09919_;
  wire _09920_;
  wire _09921_;
  wire _09922_;
  wire _09923_;
  wire _09924_;
  wire _09925_;
  wire _09926_;
  wire _09927_;
  wire _09928_;
  wire _09929_;
  wire _09930_;
  wire _09931_;
  wire _09932_;
  wire _09933_;
  wire _09934_;
  wire _09935_;
  wire _09936_;
  wire _09937_;
  wire _09938_;
  wire _09939_;
  wire _09940_;
  wire _09941_;
  wire _09942_;
  wire _09943_;
  wire _09944_;
  wire _09945_;
  wire _09946_;
  wire _09947_;
  wire _09948_;
  wire _09949_;
  wire _09950_;
  wire _09951_;
  wire _09952_;
  wire _09953_;
  wire _09954_;
  wire _09955_;
  wire _09956_;
  wire _09957_;
  wire _09958_;
  wire _09959_;
  wire _09960_;
  wire _09961_;
  wire _09962_;
  wire _09963_;
  wire _09964_;
  wire _09965_;
  wire _09966_;
  wire _09967_;
  wire _09968_;
  wire _09969_;
  wire _09970_;
  wire _09971_;
  wire _09972_;
  wire _09973_;
  wire _09974_;
  wire _09975_;
  wire _09976_;
  wire _09977_;
  wire _09978_;
  wire _09979_;
  wire _09980_;
  wire _09981_;
  wire _09982_;
  wire _09983_;
  wire _09984_;
  wire _09985_;
  wire _09986_;
  wire _09987_;
  wire _09988_;
  wire _09989_;
  wire _09990_;
  wire _09991_;
  wire _09992_;
  wire _09993_;
  wire _09994_;
  wire _09995_;
  wire _09996_;
  wire _09997_;
  wire _09998_;
  wire _09999_;
  wire _10000_;
  wire _10001_;
  wire _10002_;
  wire _10003_;
  wire _10004_;
  wire _10005_;
  wire _10006_;
  wire _10007_;
  wire _10008_;
  wire _10009_;
  wire _10010_;
  wire _10011_;
  wire _10012_;
  wire _10013_;
  wire _10014_;
  wire _10015_;
  wire _10016_;
  wire _10017_;
  wire _10018_;
  wire _10019_;
  wire _10020_;
  wire _10021_;
  wire _10022_;
  wire _10023_;
  wire _10024_;
  wire _10025_;
  wire _10026_;
  wire _10027_;
  wire _10028_;
  wire _10029_;
  wire _10030_;
  wire _10031_;
  wire _10032_;
  wire _10033_;
  wire _10034_;
  wire _10035_;
  wire _10036_;
  wire _10037_;
  wire _10038_;
  wire _10039_;
  wire _10040_;
  wire _10041_;
  wire _10042_;
  wire _10043_;
  wire _10044_;
  wire _10045_;
  wire _10046_;
  wire _10047_;
  wire _10048_;
  wire _10049_;
  wire _10050_;
  wire _10051_;
  wire _10052_;
  wire _10053_;
  wire _10054_;
  wire _10055_;
  wire _10056_;
  wire _10057_;
  wire _10058_;
  wire _10059_;
  wire _10060_;
  wire _10061_;
  wire _10062_;
  wire _10063_;
  wire _10064_;
  wire _10065_;
  wire _10066_;
  wire _10067_;
  wire _10068_;
  wire _10069_;
  wire _10070_;
  wire _10071_;
  wire _10072_;
  wire _10073_;
  wire _10074_;
  wire _10075_;
  wire _10076_;
  wire _10077_;
  wire _10078_;
  wire _10079_;
  wire _10080_;
  wire _10081_;
  wire _10082_;
  wire _10083_;
  wire _10084_;
  wire _10085_;
  wire _10086_;
  wire _10087_;
  wire _10088_;
  wire _10089_;
  wire _10090_;
  wire _10091_;
  wire _10092_;
  wire _10093_;
  wire _10094_;
  wire _10095_;
  wire _10096_;
  wire _10097_;
  wire _10098_;
  wire _10099_;
  wire _10100_;
  wire _10101_;
  wire _10102_;
  wire _10103_;
  wire _10104_;
  wire _10105_;
  wire _10106_;
  wire _10107_;
  wire _10108_;
  wire _10109_;
  wire _10110_;
  wire _10111_;
  wire _10112_;
  wire _10113_;
  wire _10114_;
  wire _10115_;
  wire _10116_;
  wire _10117_;
  wire _10118_;
  wire _10119_;
  wire _10120_;
  wire _10121_;
  wire _10122_;
  wire _10123_;
  wire _10124_;
  wire _10125_;
  wire _10126_;
  wire _10127_;
  wire _10128_;
  wire _10129_;
  wire _10130_;
  wire _10131_;
  wire _10132_;
  wire _10133_;
  wire _10134_;
  wire _10135_;
  wire _10136_;
  wire _10137_;
  wire _10138_;
  wire _10139_;
  wire _10140_;
  wire _10141_;
  wire _10142_;
  wire _10143_;
  wire _10144_;
  wire _10145_;
  wire _10146_;
  wire _10147_;
  wire _10148_;
  wire _10149_;
  wire _10150_;
  wire _10151_;
  wire _10152_;
  wire _10153_;
  wire _10154_;
  wire _10155_;
  wire _10156_;
  wire _10157_;
  wire _10158_;
  wire _10159_;
  wire _10160_;
  wire _10161_;
  wire _10162_;
  wire _10163_;
  wire _10164_;
  wire _10165_;
  wire _10166_;
  wire _10167_;
  wire _10168_;
  wire _10169_;
  wire _10170_;
  wire _10171_;
  wire _10172_;
  wire _10173_;
  wire _10174_;
  wire _10175_;
  wire _10176_;
  wire _10177_;
  wire _10178_;
  wire _10179_;
  wire _10180_;
  wire _10181_;
  wire _10182_;
  wire _10183_;
  wire _10184_;
  wire _10185_;
  wire _10186_;
  wire _10187_;
  wire _10188_;
  wire _10189_;
  wire _10190_;
  wire _10191_;
  wire _10192_;
  wire _10193_;
  wire _10194_;
  wire _10195_;
  wire _10196_;
  wire _10197_;
  wire _10198_;
  wire _10199_;
  wire _10200_;
  wire _10201_;
  wire _10202_;
  wire _10203_;
  wire _10204_;
  wire _10205_;
  wire _10206_;
  wire _10207_;
  wire _10208_;
  wire _10209_;
  wire _10210_;
  wire _10211_;
  wire _10212_;
  wire _10213_;
  wire _10214_;
  wire _10215_;
  wire _10216_;
  wire _10217_;
  wire _10218_;
  wire _10219_;
  wire _10220_;
  wire _10221_;
  wire _10222_;
  wire _10223_;
  wire _10224_;
  wire _10225_;
  wire _10226_;
  wire _10227_;
  wire _10228_;
  wire _10229_;
  wire _10230_;
  wire _10231_;
  wire _10232_;
  wire _10233_;
  wire _10234_;
  wire _10235_;
  wire _10236_;
  wire _10237_;
  wire _10238_;
  wire _10239_;
  wire _10240_;
  wire _10241_;
  wire _10242_;
  wire _10243_;
  wire _10244_;
  wire _10245_;
  wire _10246_;
  wire _10247_;
  wire _10248_;
  wire _10249_;
  wire _10250_;
  wire _10251_;
  wire _10252_;
  wire _10253_;
  wire _10254_;
  wire _10255_;
  wire _10256_;
  wire _10257_;
  wire _10258_;
  wire _10259_;
  wire _10260_;
  wire _10261_;
  wire _10262_;
  wire _10263_;
  wire _10264_;
  wire _10265_;
  wire _10266_;
  wire _10267_;
  wire _10268_;
  wire _10269_;
  wire _10270_;
  wire _10271_;
  wire _10272_;
  wire _10273_;
  wire _10274_;
  wire _10275_;
  wire _10276_;
  wire _10277_;
  wire _10278_;
  wire _10279_;
  wire _10280_;
  wire _10281_;
  wire _10282_;
  wire _10283_;
  wire _10284_;
  wire _10285_;
  wire _10286_;
  wire _10287_;
  wire _10288_;
  wire _10289_;
  wire _10290_;
  wire _10291_;
  wire _10292_;
  wire _10293_;
  wire _10294_;
  wire _10295_;
  wire _10296_;
  wire _10297_;
  wire _10298_;
  wire _10299_;
  wire _10300_;
  wire _10301_;
  wire _10302_;
  wire _10303_;
  wire _10304_;
  wire _10305_;
  wire _10306_;
  wire _10307_;
  wire _10308_;
  wire _10309_;
  wire _10310_;
  wire _10311_;
  wire _10312_;
  wire _10313_;
  wire _10314_;
  wire _10315_;
  wire _10316_;
  wire _10317_;
  wire _10318_;
  wire _10319_;
  wire _10320_;
  wire _10321_;
  wire _10322_;
  wire _10323_;
  wire _10324_;
  wire _10325_;
  wire _10326_;
  wire _10327_;
  wire _10328_;
  wire _10329_;
  wire _10330_;
  wire _10331_;
  wire _10332_;
  wire _10333_;
  wire _10334_;
  wire _10335_;
  wire _10336_;
  wire _10337_;
  wire _10338_;
  wire _10339_;
  wire _10340_;
  wire _10341_;
  wire _10342_;
  wire _10343_;
  wire _10344_;
  wire _10345_;
  wire _10346_;
  wire _10347_;
  wire _10348_;
  wire _10349_;
  wire _10350_;
  wire _10351_;
  wire _10352_;
  wire _10353_;
  wire _10354_;
  wire _10355_;
  wire _10356_;
  wire _10357_;
  wire _10358_;
  wire _10359_;
  wire _10360_;
  wire _10361_;
  wire _10362_;
  wire _10363_;
  wire _10364_;
  wire _10365_;
  wire _10366_;
  wire _10367_;
  wire _10368_;
  wire _10369_;
  wire _10370_;
  wire _10371_;
  wire _10372_;
  wire _10373_;
  wire _10374_;
  wire _10375_;
  wire _10376_;
  wire _10377_;
  wire _10378_;
  wire _10379_;
  wire _10380_;
  wire _10381_;
  wire _10382_;
  wire _10383_;
  wire _10384_;
  wire _10385_;
  wire _10386_;
  wire _10387_;
  wire _10388_;
  wire _10389_;
  wire _10390_;
  wire _10391_;
  wire _10392_;
  wire _10393_;
  wire _10394_;
  wire _10395_;
  wire _10396_;
  wire _10397_;
  wire _10398_;
  wire _10399_;
  wire _10400_;
  wire _10401_;
  wire _10402_;
  wire _10403_;
  wire _10404_;
  wire _10405_;
  wire _10406_;
  wire _10407_;
  wire _10408_;
  wire _10409_;
  wire _10410_;
  wire _10411_;
  wire _10412_;
  wire _10413_;
  wire _10414_;
  wire _10415_;
  wire _10416_;
  wire _10417_;
  wire _10418_;
  wire _10419_;
  wire _10420_;
  wire _10421_;
  wire _10422_;
  wire _10423_;
  wire _10424_;
  wire _10425_;
  wire _10426_;
  wire _10427_;
  wire _10428_;
  wire _10429_;
  wire _10430_;
  wire _10431_;
  wire _10432_;
  wire _10433_;
  wire _10434_;
  wire _10435_;
  wire _10436_;
  wire _10437_;
  wire _10438_;
  wire _10439_;
  wire _10440_;
  wire _10441_;
  wire _10442_;
  wire _10443_;
  wire _10444_;
  wire _10445_;
  wire _10446_;
  wire _10447_;
  wire _10448_;
  wire _10449_;
  wire _10450_;
  wire _10451_;
  wire _10452_;
  wire _10453_;
  wire _10454_;
  wire _10455_;
  wire _10456_;
  wire _10457_;
  wire _10458_;
  wire _10459_;
  wire _10460_;
  wire _10461_;
  wire _10462_;
  wire _10463_;
  wire _10464_;
  wire _10465_;
  wire _10466_;
  wire _10467_;
  wire _10468_;
  wire _10469_;
  wire _10470_;
  wire _10471_;
  wire _10472_;
  wire _10473_;
  wire _10474_;
  wire _10475_;
  wire _10476_;
  wire _10477_;
  wire _10478_;
  wire _10479_;
  wire _10480_;
  wire _10481_;
  wire _10482_;
  wire _10483_;
  wire _10484_;
  wire _10485_;
  wire _10486_;
  wire _10487_;
  wire _10488_;
  wire _10489_;
  wire _10490_;
  wire _10491_;
  wire _10492_;
  wire _10493_;
  wire _10494_;
  wire _10495_;
  wire _10496_;
  wire _10497_;
  wire _10498_;
  wire _10499_;
  wire _10500_;
  wire _10501_;
  wire _10502_;
  wire _10503_;
  wire _10504_;
  wire _10505_;
  wire _10506_;
  wire _10507_;
  wire _10508_;
  wire _10509_;
  wire _10510_;
  wire _10511_;
  wire _10512_;
  wire _10513_;
  wire _10514_;
  wire _10515_;
  wire _10516_;
  wire _10517_;
  wire _10518_;
  wire _10519_;
  wire _10520_;
  wire _10521_;
  wire _10522_;
  wire _10523_;
  wire _10524_;
  wire _10525_;
  wire _10526_;
  wire _10527_;
  wire _10528_;
  wire _10529_;
  wire _10530_;
  wire _10531_;
  wire _10532_;
  wire _10533_;
  wire _10534_;
  wire _10535_;
  wire _10536_;
  wire _10537_;
  wire _10538_;
  wire _10539_;
  wire _10540_;
  wire _10541_;
  wire _10542_;
  wire _10543_;
  wire _10544_;
  wire _10545_;
  wire _10546_;
  wire _10547_;
  wire _10548_;
  wire _10549_;
  wire _10550_;
  wire _10551_;
  wire _10552_;
  wire _10553_;
  wire _10554_;
  wire _10555_;
  wire _10556_;
  wire _10557_;
  wire _10558_;
  wire _10559_;
  wire _10560_;
  wire _10561_;
  wire _10562_;
  wire _10563_;
  wire _10564_;
  wire _10565_;
  wire _10566_;
  wire _10567_;
  wire _10568_;
  wire _10569_;
  wire _10570_;
  wire _10571_;
  wire _10572_;
  wire _10573_;
  wire _10574_;
  wire _10575_;
  wire _10576_;
  wire _10577_;
  wire _10578_;
  wire _10579_;
  wire _10580_;
  wire _10581_;
  wire _10582_;
  wire _10583_;
  wire _10584_;
  wire _10585_;
  wire _10586_;
  wire _10587_;
  wire _10588_;
  wire _10589_;
  wire _10590_;
  wire _10591_;
  wire _10592_;
  wire _10593_;
  wire _10594_;
  wire _10595_;
  wire _10596_;
  wire _10597_;
  wire _10598_;
  wire _10599_;
  wire _10600_;
  wire _10601_;
  wire _10602_;
  wire _10603_;
  wire _10604_;
  wire _10605_;
  wire _10606_;
  wire _10607_;
  wire _10608_;
  wire _10609_;
  wire _10610_;
  wire _10611_;
  wire _10612_;
  wire _10613_;
  wire _10614_;
  wire _10615_;
  wire _10616_;
  wire _10617_;
  wire _10618_;
  wire _10619_;
  wire _10620_;
  wire _10621_;
  wire _10622_;
  wire _10623_;
  wire _10624_;
  wire _10625_;
  wire _10626_;
  wire _10627_;
  wire _10628_;
  wire _10629_;
  wire _10630_;
  wire _10631_;
  wire _10632_;
  wire _10633_;
  wire _10634_;
  wire _10635_;
  wire _10636_;
  wire _10637_;
  wire _10638_;
  wire _10639_;
  wire _10640_;
  wire _10641_;
  wire _10642_;
  wire _10643_;
  wire _10644_;
  wire _10645_;
  wire _10646_;
  wire _10647_;
  wire _10648_;
  wire _10649_;
  wire _10650_;
  wire _10651_;
  wire _10652_;
  wire _10653_;
  wire _10654_;
  wire _10655_;
  wire _10656_;
  wire _10657_;
  wire _10658_;
  wire _10659_;
  wire _10660_;
  wire _10661_;
  wire _10662_;
  wire _10663_;
  wire _10664_;
  wire _10665_;
  wire _10666_;
  wire _10667_;
  wire _10668_;
  wire _10669_;
  wire _10670_;
  wire _10671_;
  wire _10672_;
  wire _10673_;
  wire _10674_;
  wire _10675_;
  wire _10676_;
  wire _10677_;
  wire _10678_;
  wire _10679_;
  wire _10680_;
  wire _10681_;
  wire _10682_;
  wire _10683_;
  wire _10684_;
  wire _10685_;
  wire _10686_;
  wire _10687_;
  wire _10688_;
  wire _10689_;
  wire _10690_;
  wire _10691_;
  wire _10692_;
  wire _10693_;
  wire _10694_;
  wire _10695_;
  wire _10696_;
  wire _10697_;
  wire _10698_;
  wire _10699_;
  wire _10700_;
  wire _10701_;
  wire _10702_;
  wire _10703_;
  wire _10704_;
  wire _10705_;
  wire _10706_;
  wire _10707_;
  wire _10708_;
  wire _10709_;
  wire _10710_;
  wire _10711_;
  wire _10712_;
  wire _10713_;
  wire _10714_;
  wire _10715_;
  wire _10716_;
  wire _10717_;
  wire _10718_;
  wire _10719_;
  wire _10720_;
  wire _10721_;
  wire _10722_;
  wire _10723_;
  wire _10724_;
  wire _10725_;
  wire _10726_;
  wire _10727_;
  wire _10728_;
  wire _10729_;
  wire _10730_;
  wire _10731_;
  wire _10732_;
  wire _10733_;
  wire _10734_;
  wire _10735_;
  wire _10736_;
  wire _10737_;
  wire _10738_;
  wire _10739_;
  wire _10740_;
  wire _10741_;
  wire _10742_;
  wire _10743_;
  wire _10744_;
  wire _10745_;
  wire _10746_;
  wire _10747_;
  wire _10748_;
  wire _10749_;
  wire _10750_;
  wire _10751_;
  wire _10752_;
  wire _10753_;
  wire _10754_;
  wire _10755_;
  wire _10756_;
  wire _10757_;
  wire _10758_;
  wire _10759_;
  wire _10760_;
  wire _10761_;
  wire _10762_;
  wire _10763_;
  wire _10764_;
  wire _10765_;
  wire _10766_;
  wire _10767_;
  wire _10768_;
  wire _10769_;
  wire _10770_;
  wire _10771_;
  wire _10772_;
  wire _10773_;
  wire _10774_;
  wire _10775_;
  wire _10776_;
  wire _10777_;
  wire _10778_;
  wire _10779_;
  wire _10780_;
  wire _10781_;
  wire _10782_;
  wire _10783_;
  wire _10784_;
  wire _10785_;
  wire _10786_;
  wire _10787_;
  wire _10788_;
  wire _10789_;
  wire _10790_;
  wire _10791_;
  wire _10792_;
  wire _10793_;
  wire _10794_;
  wire _10795_;
  wire _10796_;
  wire _10797_;
  wire _10798_;
  wire _10799_;
  wire _10800_;
  wire _10801_;
  wire _10802_;
  wire _10803_;
  wire _10804_;
  wire _10805_;
  wire _10806_;
  wire _10807_;
  wire _10808_;
  wire _10809_;
  wire _10810_;
  wire _10811_;
  wire _10812_;
  wire _10813_;
  wire _10814_;
  wire _10815_;
  wire _10816_;
  wire _10817_;
  wire _10818_;
  wire _10819_;
  wire _10820_;
  wire _10821_;
  wire _10822_;
  wire _10823_;
  wire _10824_;
  wire _10825_;
  wire _10826_;
  wire _10827_;
  wire _10828_;
  wire _10829_;
  wire _10830_;
  wire _10831_;
  wire _10832_;
  wire _10833_;
  wire _10834_;
  wire _10835_;
  wire _10836_;
  wire _10837_;
  wire _10838_;
  wire _10839_;
  wire _10840_;
  wire _10841_;
  wire _10842_;
  wire _10843_;
  wire _10844_;
  wire _10845_;
  wire _10846_;
  wire _10847_;
  wire _10848_;
  wire _10849_;
  wire _10850_;
  wire _10851_;
  wire _10852_;
  wire _10853_;
  wire _10854_;
  wire _10855_;
  wire _10856_;
  wire _10857_;
  wire _10858_;
  wire _10859_;
  wire _10860_;
  wire _10861_;
  wire _10862_;
  wire _10863_;
  wire _10864_;
  wire _10865_;
  wire _10866_;
  wire _10867_;
  wire _10868_;
  wire _10869_;
  wire _10870_;
  wire _10871_;
  wire _10872_;
  wire _10873_;
  wire _10874_;
  wire _10875_;
  wire _10876_;
  wire _10877_;
  wire _10878_;
  wire _10879_;
  wire _10880_;
  wire _10881_;
  wire _10882_;
  wire _10883_;
  wire _10884_;
  wire _10885_;
  wire _10886_;
  wire _10887_;
  wire _10888_;
  wire _10889_;
  wire _10890_;
  wire _10891_;
  wire _10892_;
  wire _10893_;
  wire _10894_;
  wire _10895_;
  wire _10896_;
  wire _10897_;
  wire _10898_;
  wire _10899_;
  wire _10900_;
  wire _10901_;
  wire _10902_;
  wire _10903_;
  wire _10904_;
  wire _10905_;
  wire _10906_;
  wire _10907_;
  wire _10908_;
  wire _10909_;
  wire _10910_;
  wire _10911_;
  wire _10912_;
  wire _10913_;
  wire _10914_;
  wire _10915_;
  wire _10916_;
  wire _10917_;
  wire _10918_;
  wire _10919_;
  wire _10920_;
  wire _10921_;
  wire _10922_;
  wire _10923_;
  wire _10924_;
  wire _10925_;
  wire _10926_;
  wire _10927_;
  wire _10928_;
  wire _10929_;
  wire _10930_;
  wire _10931_;
  wire _10932_;
  wire _10933_;
  wire _10934_;
  wire _10935_;
  wire _10936_;
  wire _10937_;
  wire _10938_;
  wire _10939_;
  wire _10940_;
  wire _10941_;
  wire _10942_;
  wire _10943_;
  wire _10944_;
  wire _10945_;
  wire _10946_;
  wire _10947_;
  wire _10948_;
  wire _10949_;
  wire _10950_;
  wire _10951_;
  wire _10952_;
  wire _10953_;
  wire _10954_;
  wire _10955_;
  wire _10956_;
  wire _10957_;
  wire _10958_;
  wire _10959_;
  wire _10960_;
  wire _10961_;
  wire _10962_;
  wire _10963_;
  wire _10964_;
  wire _10965_;
  wire _10966_;
  wire _10967_;
  wire _10968_;
  wire _10969_;
  wire _10970_;
  wire _10971_;
  wire _10972_;
  wire _10973_;
  wire _10974_;
  wire _10975_;
  wire _10976_;
  wire _10977_;
  wire _10978_;
  wire _10979_;
  wire _10980_;
  wire _10981_;
  wire _10982_;
  wire _10983_;
  wire _10984_;
  wire _10985_;
  wire _10986_;
  wire _10987_;
  wire _10988_;
  wire _10989_;
  wire _10990_;
  wire _10991_;
  wire _10992_;
  wire _10993_;
  wire _10994_;
  wire _10995_;
  wire _10996_;
  wire _10997_;
  wire _10998_;
  wire _10999_;
  wire _11000_;
  wire _11001_;
  wire _11002_;
  wire _11003_;
  wire _11004_;
  wire _11005_;
  wire _11006_;
  wire _11007_;
  wire _11008_;
  wire _11009_;
  wire _11010_;
  wire _11011_;
  wire _11012_;
  wire _11013_;
  wire _11014_;
  wire _11015_;
  wire _11016_;
  wire _11017_;
  wire _11018_;
  wire _11019_;
  wire _11020_;
  wire _11021_;
  wire _11022_;
  wire _11023_;
  wire _11024_;
  wire _11025_;
  wire _11026_;
  wire _11027_;
  wire _11028_;
  wire _11029_;
  wire _11030_;
  wire _11031_;
  wire _11032_;
  wire _11033_;
  wire _11034_;
  wire _11035_;
  wire _11036_;
  wire _11037_;
  wire _11038_;
  wire _11039_;
  wire _11040_;
  wire _11041_;
  wire _11042_;
  wire _11043_;
  wire _11044_;
  wire _11045_;
  wire _11046_;
  wire _11047_;
  wire _11048_;
  wire _11049_;
  wire _11050_;
  wire _11051_;
  wire _11052_;
  wire _11053_;
  wire _11054_;
  wire _11055_;
  wire _11056_;
  wire _11057_;
  wire _11058_;
  wire _11059_;
  wire _11060_;
  wire _11061_;
  wire _11062_;
  wire _11063_;
  wire _11064_;
  wire _11065_;
  wire _11066_;
  wire _11067_;
  wire _11068_;
  wire _11069_;
  wire _11070_;
  wire _11071_;
  wire _11072_;
  wire _11073_;
  wire _11074_;
  wire _11075_;
  wire _11076_;
  wire _11077_;
  wire _11078_;
  wire _11079_;
  wire _11080_;
  wire _11081_;
  wire _11082_;
  wire _11083_;
  wire _11084_;
  wire _11085_;
  wire _11086_;
  wire _11087_;
  wire _11088_;
  wire _11089_;
  wire _11090_;
  wire _11091_;
  wire _11092_;
  wire _11093_;
  wire _11094_;
  wire _11095_;
  wire _11096_;
  wire _11097_;
  wire _11098_;
  wire _11099_;
  wire _11100_;
  wire _11101_;
  wire _11102_;
  wire _11103_;
  wire _11104_;
  wire _11105_;
  wire _11106_;
  wire _11107_;
  wire _11108_;
  wire _11109_;
  wire _11110_;
  wire _11111_;
  wire _11112_;
  wire _11113_;
  wire _11114_;
  wire _11115_;
  wire _11116_;
  wire _11117_;
  wire _11118_;
  wire _11119_;
  wire _11120_;
  wire _11121_;
  wire _11122_;
  wire _11123_;
  wire _11124_;
  wire _11125_;
  wire _11126_;
  wire _11127_;
  wire _11128_;
  wire _11129_;
  wire _11130_;
  wire _11131_;
  wire _11132_;
  wire _11133_;
  wire _11134_;
  wire _11135_;
  wire _11136_;
  wire _11137_;
  wire _11138_;
  wire _11139_;
  wire _11140_;
  wire _11141_;
  wire _11142_;
  wire _11143_;
  wire _11144_;
  wire _11145_;
  wire _11146_;
  wire _11147_;
  wire _11148_;
  wire _11149_;
  wire _11150_;
  wire _11151_;
  wire _11152_;
  wire _11153_;
  wire _11154_;
  wire _11155_;
  wire _11156_;
  wire _11157_;
  wire _11158_;
  wire _11159_;
  wire _11160_;
  wire _11161_;
  wire _11162_;
  wire _11163_;
  wire _11164_;
  wire _11165_;
  wire _11166_;
  wire _11167_;
  wire _11168_;
  wire _11169_;
  wire _11170_;
  wire _11171_;
  wire _11172_;
  wire _11173_;
  wire _11174_;
  wire _11175_;
  wire _11176_;
  wire _11177_;
  wire _11178_;
  wire _11179_;
  wire _11180_;
  wire _11181_;
  wire _11182_;
  wire _11183_;
  wire _11184_;
  wire _11185_;
  wire _11186_;
  wire _11187_;
  wire _11188_;
  wire _11189_;
  wire _11190_;
  wire _11191_;
  wire _11192_;
  wire _11193_;
  wire _11194_;
  wire _11195_;
  wire _11196_;
  wire _11197_;
  wire _11198_;
  wire _11199_;
  wire _11200_;
  wire _11201_;
  wire _11202_;
  wire _11203_;
  wire _11204_;
  wire _11205_;
  wire _11206_;
  wire _11207_;
  wire _11208_;
  wire _11209_;
  wire _11210_;
  wire _11211_;
  wire _11212_;
  wire _11213_;
  wire _11214_;
  wire _11215_;
  wire _11216_;
  wire _11217_;
  wire _11218_;
  wire _11219_;
  wire _11220_;
  wire _11221_;
  wire _11222_;
  wire _11223_;
  wire _11224_;
  wire _11225_;
  wire _11226_;
  wire _11227_;
  wire _11228_;
  wire _11229_;
  wire _11230_;
  wire _11231_;
  wire _11232_;
  wire _11233_;
  wire _11234_;
  wire _11235_;
  wire _11236_;
  wire _11237_;
  wire _11238_;
  wire _11239_;
  wire _11240_;
  wire _11241_;
  wire _11242_;
  wire _11243_;
  wire _11244_;
  wire _11245_;
  wire _11246_;
  wire _11247_;
  wire _11248_;
  wire _11249_;
  wire _11250_;
  wire _11251_;
  wire _11252_;
  wire _11253_;
  wire _11254_;
  wire _11255_;
  wire _11256_;
  wire _11257_;
  wire _11258_;
  wire _11259_;
  wire _11260_;
  wire _11261_;
  wire _11262_;
  wire _11263_;
  wire _11264_;
  wire _11265_;
  wire _11266_;
  wire _11267_;
  wire _11268_;
  wire _11269_;
  wire _11270_;
  wire _11271_;
  wire _11272_;
  wire _11273_;
  wire _11274_;
  wire _11275_;
  wire _11276_;
  wire _11277_;
  wire _11278_;
  wire _11279_;
  wire _11280_;
  wire _11281_;
  wire _11282_;
  wire _11283_;
  wire _11284_;
  wire _11285_;
  wire _11286_;
  wire _11287_;
  wire _11288_;
  wire _11289_;
  wire _11290_;
  wire _11291_;
  wire _11292_;
  wire _11293_;
  wire _11294_;
  wire _11295_;
  wire _11296_;
  wire _11297_;
  wire _11298_;
  wire _11299_;
  wire _11300_;
  wire _11301_;
  wire _11302_;
  wire _11303_;
  wire _11304_;
  wire _11305_;
  wire _11306_;
  wire _11307_;
  wire _11308_;
  wire _11309_;
  wire _11310_;
  wire _11311_;
  wire _11312_;
  wire _11313_;
  wire _11314_;
  wire _11315_;
  wire _11316_;
  wire _11317_;
  wire _11318_;
  wire _11319_;
  wire _11320_;
  wire _11321_;
  wire _11322_;
  wire _11323_;
  wire _11324_;
  wire _11325_;
  wire _11326_;
  wire _11327_;
  wire _11328_;
  wire _11329_;
  wire _11330_;
  wire _11331_;
  wire _11332_;
  wire _11333_;
  wire _11334_;
  wire _11335_;
  wire _11336_;
  wire _11337_;
  wire _11338_;
  wire _11339_;
  wire _11340_;
  wire _11341_;
  wire _11342_;
  wire _11343_;
  wire _11344_;
  wire _11345_;
  wire _11346_;
  wire _11347_;
  wire _11348_;
  wire _11349_;
  wire _11350_;
  wire _11351_;
  wire _11352_;
  wire _11353_;
  wire _11354_;
  wire _11355_;
  wire _11356_;
  wire _11357_;
  wire _11358_;
  wire _11359_;
  wire _11360_;
  wire _11361_;
  wire _11362_;
  wire _11363_;
  wire _11364_;
  wire _11365_;
  wire _11366_;
  wire _11367_;
  wire _11368_;
  wire _11369_;
  wire _11370_;
  wire _11371_;
  wire _11372_;
  wire _11373_;
  wire _11374_;
  wire _11375_;
  wire _11376_;
  wire _11377_;
  wire _11378_;
  wire _11379_;
  wire _11380_;
  wire _11381_;
  wire _11382_;
  wire _11383_;
  wire _11384_;
  wire _11385_;
  wire _11386_;
  wire _11387_;
  wire _11388_;
  wire _11389_;
  wire _11390_;
  wire _11391_;
  wire _11392_;
  wire _11393_;
  wire _11394_;
  wire _11395_;
  wire _11396_;
  wire _11397_;
  wire _11398_;
  wire _11399_;
  wire _11400_;
  wire _11401_;
  wire _11402_;
  wire _11403_;
  wire _11404_;
  wire _11405_;
  wire _11406_;
  wire _11407_;
  wire _11408_;
  wire _11409_;
  wire _11410_;
  wire _11411_;
  wire _11412_;
  wire _11413_;
  wire _11414_;
  wire _11415_;
  wire _11416_;
  wire _11417_;
  wire _11418_;
  wire _11419_;
  wire _11420_;
  wire _11421_;
  wire _11422_;
  wire _11423_;
  wire _11424_;
  wire _11425_;
  wire _11426_;
  wire _11427_;
  wire _11428_;
  wire _11429_;
  wire _11430_;
  wire _11431_;
  wire _11432_;
  wire _11433_;
  wire _11434_;
  wire _11435_;
  wire _11436_;
  wire _11437_;
  wire _11438_;
  wire _11439_;
  wire _11440_;
  wire _11441_;
  wire _11442_;
  wire _11443_;
  wire _11444_;
  wire _11445_;
  wire _11446_;
  wire _11447_;
  wire _11448_;
  wire _11449_;
  wire _11450_;
  wire _11451_;
  wire _11452_;
  wire _11453_;
  wire _11454_;
  wire _11455_;
  wire _11456_;
  wire _11457_;
  wire _11458_;
  wire _11459_;
  wire _11460_;
  wire _11461_;
  wire _11462_;
  wire _11463_;
  wire _11464_;
  wire _11465_;
  wire _11466_;
  wire _11467_;
  wire _11468_;
  wire _11469_;
  wire _11470_;
  wire _11471_;
  wire _11472_;
  wire _11473_;
  wire _11474_;
  wire _11475_;
  wire _11476_;
  wire _11477_;
  wire _11478_;
  wire _11479_;
  wire _11480_;
  wire _11481_;
  wire _11482_;
  wire _11483_;
  wire _11484_;
  wire _11485_;
  wire _11486_;
  wire _11487_;
  wire _11488_;
  wire _11489_;
  wire _11490_;
  wire _11491_;
  wire _11492_;
  wire _11493_;
  wire _11494_;
  wire _11495_;
  wire _11496_;
  wire _11497_;
  wire _11498_;
  wire _11499_;
  wire _11500_;
  wire _11501_;
  wire _11502_;
  wire _11503_;
  wire _11504_;
  wire _11505_;
  wire _11506_;
  wire _11507_;
  wire _11508_;
  wire _11509_;
  wire _11510_;
  wire _11511_;
  wire _11512_;
  wire _11513_;
  wire _11514_;
  wire _11515_;
  wire _11516_;
  wire _11517_;
  wire _11518_;
  wire _11519_;
  wire _11520_;
  wire _11521_;
  wire _11522_;
  wire _11523_;
  wire _11524_;
  wire _11525_;
  wire _11526_;
  wire _11527_;
  wire _11528_;
  wire _11529_;
  wire _11530_;
  wire _11531_;
  wire _11532_;
  wire _11533_;
  wire _11534_;
  wire _11535_;
  wire _11536_;
  wire _11537_;
  wire _11538_;
  wire _11539_;
  wire _11540_;
  wire _11541_;
  wire _11542_;
  wire _11543_;
  wire _11544_;
  wire _11545_;
  wire _11546_;
  wire _11547_;
  wire _11548_;
  wire _11549_;
  wire _11550_;
  wire _11551_;
  wire _11552_;
  wire _11553_;
  wire _11554_;
  wire _11555_;
  wire _11556_;
  wire _11557_;
  wire _11558_;
  wire _11559_;
  wire _11560_;
  wire _11561_;
  wire _11562_;
  wire _11563_;
  wire _11564_;
  wire _11565_;
  wire _11566_;
  wire _11567_;
  wire _11568_;
  wire _11569_;
  wire _11570_;
  wire _11571_;
  wire _11572_;
  wire _11573_;
  wire _11574_;
  wire _11575_;
  wire _11576_;
  wire _11577_;
  wire _11578_;
  wire _11579_;
  wire _11580_;
  wire _11581_;
  wire _11582_;
  wire _11583_;
  wire _11584_;
  wire _11585_;
  wire _11586_;
  wire _11587_;
  wire _11588_;
  wire _11589_;
  wire _11590_;
  wire _11591_;
  wire _11592_;
  wire _11593_;
  wire _11594_;
  wire _11595_;
  wire _11596_;
  wire _11597_;
  wire _11598_;
  wire _11599_;
  wire _11600_;
  wire _11601_;
  wire _11602_;
  wire _11603_;
  wire _11604_;
  wire _11605_;
  wire _11606_;
  wire _11607_;
  wire _11608_;
  wire _11609_;
  wire _11610_;
  wire _11611_;
  wire _11612_;
  wire _11613_;
  wire _11614_;
  wire _11615_;
  wire _11616_;
  wire _11617_;
  wire _11618_;
  wire _11619_;
  wire _11620_;
  wire _11621_;
  wire _11622_;
  wire _11623_;
  wire _11624_;
  wire _11625_;
  wire _11626_;
  wire _11627_;
  wire _11628_;
  wire _11629_;
  wire _11630_;
  wire _11631_;
  wire _11632_;
  wire _11633_;
  wire _11634_;
  wire _11635_;
  wire _11636_;
  wire _11637_;
  wire _11638_;
  wire _11639_;
  wire _11640_;
  wire _11641_;
  wire _11642_;
  wire _11643_;
  wire _11644_;
  wire _11645_;
  wire _11646_;
  wire _11647_;
  wire _11648_;
  wire _11649_;
  wire _11650_;
  wire _11651_;
  wire _11652_;
  wire _11653_;
  wire _11654_;
  wire _11655_;
  wire _11656_;
  wire _11657_;
  wire _11658_;
  wire _11659_;
  wire _11660_;
  wire _11661_;
  wire _11662_;
  wire _11663_;
  wire _11664_;
  wire _11665_;
  wire _11666_;
  wire _11667_;
  wire _11668_;
  wire _11669_;
  wire _11670_;
  wire _11671_;
  wire _11672_;
  wire _11673_;
  wire _11674_;
  wire _11675_;
  wire _11676_;
  wire _11677_;
  wire _11678_;
  wire _11679_;
  wire _11680_;
  wire _11681_;
  wire _11682_;
  wire _11683_;
  wire _11684_;
  wire _11685_;
  wire _11686_;
  wire _11687_;
  wire _11688_;
  wire _11689_;
  wire _11690_;
  wire _11691_;
  wire _11692_;
  wire _11693_;
  wire _11694_;
  wire _11695_;
  wire _11696_;
  wire _11697_;
  wire _11698_;
  wire _11699_;
  wire _11700_;
  wire _11701_;
  wire _11702_;
  wire _11703_;
  wire _11704_;
  wire _11705_;
  wire _11706_;
  wire _11707_;
  wire _11708_;
  wire _11709_;
  wire _11710_;
  wire _11711_;
  wire _11712_;
  wire _11713_;
  wire _11714_;
  wire _11715_;
  wire _11716_;
  wire _11717_;
  wire _11718_;
  wire _11719_;
  wire _11720_;
  wire _11721_;
  wire _11722_;
  wire _11723_;
  wire _11724_;
  wire _11725_;
  wire _11726_;
  wire _11727_;
  wire _11728_;
  wire _11729_;
  wire _11730_;
  wire _11731_;
  wire _11732_;
  wire _11733_;
  wire _11734_;
  wire _11735_;
  wire _11736_;
  wire _11737_;
  wire _11738_;
  wire _11739_;
  wire _11740_;
  wire _11741_;
  wire _11742_;
  wire _11743_;
  wire _11744_;
  wire _11745_;
  wire _11746_;
  wire _11747_;
  wire _11748_;
  wire _11749_;
  wire _11750_;
  wire _11751_;
  wire _11752_;
  wire _11753_;
  wire _11754_;
  wire _11755_;
  wire _11756_;
  wire _11757_;
  wire _11758_;
  wire _11759_;
  wire _11760_;
  wire _11761_;
  wire _11762_;
  wire _11763_;
  wire _11764_;
  wire _11765_;
  wire _11766_;
  wire _11767_;
  wire _11768_;
  wire _11769_;
  wire _11770_;
  wire _11771_;
  wire _11772_;
  wire _11773_;
  wire _11774_;
  wire _11775_;
  wire _11776_;
  wire _11777_;
  wire _11778_;
  wire _11779_;
  wire _11780_;
  wire _11781_;
  wire _11782_;
  wire _11783_;
  wire _11784_;
  wire _11785_;
  wire _11786_;
  wire _11787_;
  wire _11788_;
  wire _11789_;
  wire _11790_;
  wire _11791_;
  wire _11792_;
  wire _11793_;
  wire _11794_;
  wire _11795_;
  wire _11796_;
  wire _11797_;
  wire _11798_;
  wire _11799_;
  wire _11800_;
  wire _11801_;
  wire _11802_;
  wire _11803_;
  wire _11804_;
  wire _11805_;
  wire _11806_;
  wire _11807_;
  wire _11808_;
  wire _11809_;
  wire _11810_;
  wire _11811_;
  wire _11812_;
  wire _11813_;
  wire _11814_;
  wire _11815_;
  wire _11816_;
  wire _11817_;
  wire _11818_;
  wire _11819_;
  wire _11820_;
  wire _11821_;
  wire _11822_;
  wire _11823_;
  wire _11824_;
  wire _11825_;
  wire _11826_;
  wire _11827_;
  wire _11828_;
  wire _11829_;
  wire _11830_;
  wire _11831_;
  wire _11832_;
  wire _11833_;
  wire _11834_;
  wire _11835_;
  wire _11836_;
  wire _11837_;
  wire _11838_;
  wire _11839_;
  wire _11840_;
  wire _11841_;
  wire _11842_;
  wire _11843_;
  wire _11844_;
  wire _11845_;
  wire _11846_;
  wire _11847_;
  wire _11848_;
  wire _11849_;
  wire _11850_;
  wire _11851_;
  wire _11852_;
  wire _11853_;
  wire _11854_;
  wire _11855_;
  wire _11856_;
  wire _11857_;
  wire _11858_;
  wire _11859_;
  wire _11860_;
  wire _11861_;
  wire _11862_;
  wire _11863_;
  wire _11864_;
  wire _11865_;
  wire _11866_;
  wire _11867_;
  wire _11868_;
  wire _11869_;
  wire _11870_;
  wire _11871_;
  wire _11872_;
  wire _11873_;
  wire _11874_;
  wire _11875_;
  wire _11876_;
  wire _11877_;
  wire _11878_;
  wire _11879_;
  wire _11880_;
  wire _11881_;
  wire _11882_;
  wire _11883_;
  wire _11884_;
  wire _11885_;
  wire _11886_;
  wire _11887_;
  wire _11888_;
  wire _11889_;
  wire _11890_;
  wire _11891_;
  wire _11892_;
  wire _11893_;
  wire _11894_;
  wire _11895_;
  wire _11896_;
  wire _11897_;
  wire _11898_;
  wire _11899_;
  wire _11900_;
  wire _11901_;
  wire _11902_;
  wire _11903_;
  wire _11904_;
  wire _11905_;
  wire _11906_;
  wire _11907_;
  wire _11908_;
  wire _11909_;
  wire _11910_;
  wire _11911_;
  wire _11912_;
  wire _11913_;
  wire _11914_;
  wire _11915_;
  wire _11916_;
  wire _11917_;
  wire _11918_;
  wire _11919_;
  wire _11920_;
  wire _11921_;
  wire _11922_;
  wire _11923_;
  wire _11924_;
  wire _11925_;
  wire _11926_;
  wire _11927_;
  wire _11928_;
  wire _11929_;
  wire _11930_;
  wire _11931_;
  wire _11932_;
  wire _11933_;
  wire _11934_;
  wire _11935_;
  wire _11936_;
  wire _11937_;
  wire _11938_;
  wire _11939_;
  wire _11940_;
  wire _11941_;
  wire _11942_;
  wire _11943_;
  wire _11944_;
  wire _11945_;
  wire _11946_;
  wire _11947_;
  wire _11948_;
  wire _11949_;
  wire _11950_;
  wire _11951_;
  wire _11952_;
  wire _11953_;
  wire _11954_;
  wire _11955_;
  wire _11956_;
  wire _11957_;
  wire _11958_;
  wire _11959_;
  wire _11960_;
  wire _11961_;
  wire _11962_;
  wire _11963_;
  wire _11964_;
  wire _11965_;
  wire _11966_;
  wire _11967_;
  wire _11968_;
  wire _11969_;
  wire _11970_;
  wire _11971_;
  wire _11972_;
  wire _11973_;
  wire _11974_;
  wire _11975_;
  wire _11976_;
  wire _11977_;
  wire _11978_;
  wire _11979_;
  wire _11980_;
  wire _11981_;
  wire _11982_;
  wire _11983_;
  wire _11984_;
  wire _11985_;
  wire _11986_;
  wire _11987_;
  wire _11988_;
  wire _11989_;
  wire _11990_;
  wire _11991_;
  wire _11992_;
  wire _11993_;
  wire _11994_;
  wire _11995_;
  wire _11996_;
  wire _11997_;
  wire _11998_;
  wire _11999_;
  wire _12000_;
  wire _12001_;
  wire _12002_;
  wire _12003_;
  wire _12004_;
  wire _12005_;
  wire _12006_;
  wire _12007_;
  wire _12008_;
  wire _12009_;
  wire _12010_;
  wire _12011_;
  wire _12012_;
  wire _12013_;
  wire _12014_;
  wire _12015_;
  wire _12016_;
  wire _12017_;
  wire _12018_;
  wire _12019_;
  wire _12020_;
  wire _12021_;
  wire _12022_;
  wire _12023_;
  wire _12024_;
  wire _12025_;
  wire _12026_;
  wire _12027_;
  wire _12028_;
  wire _12029_;
  wire _12030_;
  wire _12031_;
  wire _12032_;
  wire _12033_;
  wire _12034_;
  wire _12035_;
  wire _12036_;
  wire _12037_;
  wire _12038_;
  wire _12039_;
  wire _12040_;
  wire _12041_;
  wire _12042_;
  wire _12043_;
  wire _12044_;
  wire _12045_;
  wire _12046_;
  wire _12047_;
  wire _12048_;
  wire _12049_;
  wire _12050_;
  wire _12051_;
  wire _12052_;
  wire _12053_;
  wire _12054_;
  wire _12055_;
  wire _12056_;
  wire _12057_;
  wire _12058_;
  wire _12059_;
  wire _12060_;
  wire _12061_;
  wire _12062_;
  wire _12063_;
  wire _12064_;
  wire _12065_;
  wire _12066_;
  wire _12067_;
  wire _12068_;
  wire _12069_;
  wire _12070_;
  wire _12071_;
  wire _12072_;
  wire _12073_;
  wire _12074_;
  wire _12075_;
  wire _12076_;
  wire _12077_;
  wire _12078_;
  wire _12079_;
  wire _12080_;
  wire _12081_;
  wire _12082_;
  wire _12083_;
  wire _12084_;
  wire _12085_;
  wire _12086_;
  wire _12087_;
  wire _12088_;
  wire _12089_;
  wire _12090_;
  wire _12091_;
  wire _12092_;
  wire _12093_;
  wire _12094_;
  wire _12095_;
  wire _12096_;
  wire _12097_;
  wire _12098_;
  wire _12099_;
  wire _12100_;
  wire _12101_;
  wire _12102_;
  wire _12103_;
  wire _12104_;
  wire _12105_;
  wire _12106_;
  wire _12107_;
  wire _12108_;
  wire _12109_;
  wire _12110_;
  wire _12111_;
  wire _12112_;
  wire _12113_;
  wire _12114_;
  wire _12115_;
  wire _12116_;
  wire _12117_;
  wire _12118_;
  wire _12119_;
  wire _12120_;
  wire _12121_;
  wire _12122_;
  wire _12123_;
  wire _12124_;
  wire _12125_;
  wire _12126_;
  wire _12127_;
  wire _12128_;
  wire _12129_;
  wire _12130_;
  wire _12131_;
  wire _12132_;
  wire _12133_;
  wire _12134_;
  wire _12135_;
  wire _12136_;
  wire _12137_;
  wire _12138_;
  wire _12139_;
  wire _12140_;
  wire _12141_;
  wire _12142_;
  wire _12143_;
  wire _12144_;
  wire _12145_;
  wire _12146_;
  wire _12147_;
  wire _12148_;
  wire _12149_;
  wire _12150_;
  wire _12151_;
  wire _12152_;
  wire _12153_;
  wire _12154_;
  wire _12155_;
  wire _12156_;
  wire _12157_;
  wire _12158_;
  wire _12159_;
  wire _12160_;
  wire _12161_;
  wire _12162_;
  wire _12163_;
  wire _12164_;
  wire _12165_;
  wire _12166_;
  wire _12167_;
  wire _12168_;
  wire _12169_;
  wire _12170_;
  wire _12171_;
  wire _12172_;
  wire _12173_;
  wire _12174_;
  wire _12175_;
  wire _12176_;
  wire _12177_;
  wire _12178_;
  wire _12179_;
  wire _12180_;
  wire _12181_;
  wire _12182_;
  wire _12183_;
  wire _12184_;
  wire _12185_;
  wire _12186_;
  wire _12187_;
  wire _12188_;
  wire _12189_;
  wire _12190_;
  wire _12191_;
  wire _12192_;
  wire _12193_;
  wire _12194_;
  wire _12195_;
  wire _12196_;
  wire _12197_;
  wire _12198_;
  wire _12199_;
  wire _12200_;
  wire _12201_;
  wire _12202_;
  wire _12203_;
  wire _12204_;
  wire _12205_;
  wire _12206_;
  wire _12207_;
  wire _12208_;
  wire _12209_;
  wire _12210_;
  wire _12211_;
  wire _12212_;
  wire _12213_;
  wire _12214_;
  wire _12215_;
  wire _12216_;
  wire _12217_;
  wire _12218_;
  wire _12219_;
  wire _12220_;
  wire _12221_;
  wire _12222_;
  wire _12223_;
  wire _12224_;
  wire _12225_;
  wire _12226_;
  wire _12227_;
  wire _12228_;
  wire _12229_;
  wire _12230_;
  wire _12231_;
  wire _12232_;
  wire _12233_;
  wire _12234_;
  wire _12235_;
  wire _12236_;
  wire _12237_;
  wire _12238_;
  wire _12239_;
  wire _12240_;
  wire _12241_;
  wire _12242_;
  wire _12243_;
  wire _12244_;
  wire _12245_;
  wire _12246_;
  wire _12247_;
  wire _12248_;
  wire _12249_;
  wire _12250_;
  wire _12251_;
  wire _12252_;
  wire _12253_;
  wire _12254_;
  wire _12255_;
  wire _12256_;
  wire _12257_;
  wire _12258_;
  wire _12259_;
  wire _12260_;
  wire _12261_;
  wire _12262_;
  wire _12263_;
  wire _12264_;
  wire _12265_;
  wire _12266_;
  wire _12267_;
  wire _12268_;
  wire _12269_;
  wire _12270_;
  wire _12271_;
  wire _12272_;
  wire _12273_;
  wire _12274_;
  wire _12275_;
  wire _12276_;
  wire _12277_;
  wire _12278_;
  wire _12279_;
  wire _12280_;
  wire _12281_;
  wire _12282_;
  wire _12283_;
  wire _12284_;
  wire _12285_;
  wire _12286_;
  wire _12287_;
  wire _12288_;
  wire _12289_;
  wire _12290_;
  wire _12291_;
  wire _12292_;
  wire _12293_;
  wire _12294_;
  wire _12295_;
  wire _12296_;
  wire _12297_;
  wire _12298_;
  wire _12299_;
  wire _12300_;
  wire _12301_;
  wire _12302_;
  wire _12303_;
  wire _12304_;
  wire _12305_;
  wire _12306_;
  wire _12307_;
  wire _12308_;
  wire _12309_;
  wire _12310_;
  wire _12311_;
  wire _12312_;
  wire _12313_;
  wire _12314_;
  wire _12315_;
  wire _12316_;
  wire _12317_;
  wire _12318_;
  wire _12319_;
  wire _12320_;
  wire _12321_;
  wire _12322_;
  wire _12323_;
  wire _12324_;
  wire _12325_;
  wire _12326_;
  wire _12327_;
  wire _12328_;
  wire _12329_;
  wire _12330_;
  wire _12331_;
  wire _12332_;
  wire _12333_;
  wire _12334_;
  wire _12335_;
  wire _12336_;
  wire _12337_;
  wire _12338_;
  wire _12339_;
  wire _12340_;
  wire _12341_;
  wire _12342_;
  wire _12343_;
  wire _12344_;
  wire _12345_;
  wire _12346_;
  wire _12347_;
  wire _12348_;
  wire _12349_;
  wire _12350_;
  wire _12351_;
  wire _12352_;
  wire _12353_;
  wire _12354_;
  wire _12355_;
  wire _12356_;
  wire _12357_;
  wire _12358_;
  wire _12359_;
  wire _12360_;
  wire _12361_;
  wire _12362_;
  wire _12363_;
  wire _12364_;
  wire _12365_;
  wire _12366_;
  wire _12367_;
  wire _12368_;
  wire _12369_;
  wire _12370_;
  wire _12371_;
  wire _12372_;
  wire _12373_;
  wire _12374_;
  wire _12375_;
  wire _12376_;
  wire _12377_;
  wire _12378_;
  wire _12379_;
  wire _12380_;
  wire _12381_;
  wire _12382_;
  wire _12383_;
  wire _12384_;
  wire _12385_;
  wire _12386_;
  wire _12387_;
  wire _12388_;
  wire _12389_;
  wire _12390_;
  wire _12391_;
  wire _12392_;
  wire _12393_;
  wire _12394_;
  wire _12395_;
  wire _12396_;
  wire _12397_;
  wire _12398_;
  wire _12399_;
  wire _12400_;
  wire _12401_;
  wire _12402_;
  wire _12403_;
  wire _12404_;
  wire _12405_;
  wire _12406_;
  wire _12407_;
  wire _12408_;
  wire _12409_;
  wire _12410_;
  wire _12411_;
  wire _12412_;
  wire _12413_;
  wire _12414_;
  wire _12415_;
  wire _12416_;
  wire _12417_;
  wire _12418_;
  wire _12419_;
  wire _12420_;
  wire _12421_;
  wire _12422_;
  wire _12423_;
  wire _12424_;
  wire _12425_;
  wire _12426_;
  wire _12427_;
  wire _12428_;
  wire _12429_;
  wire _12430_;
  wire _12431_;
  wire _12432_;
  wire _12433_;
  wire _12434_;
  wire _12435_;
  wire _12436_;
  wire _12437_;
  wire _12438_;
  wire _12439_;
  wire _12440_;
  wire _12441_;
  wire _12442_;
  wire _12443_;
  wire _12444_;
  wire _12445_;
  wire _12446_;
  wire _12447_;
  wire _12448_;
  wire _12449_;
  wire _12450_;
  wire _12451_;
  wire _12452_;
  wire _12453_;
  wire _12454_;
  wire _12455_;
  wire _12456_;
  wire _12457_;
  wire _12458_;
  wire _12459_;
  wire _12460_;
  wire _12461_;
  wire _12462_;
  wire _12463_;
  wire _12464_;
  wire _12465_;
  wire _12466_;
  wire _12467_;
  wire _12468_;
  wire _12469_;
  wire _12470_;
  wire _12471_;
  wire _12472_;
  wire _12473_;
  wire _12474_;
  wire _12475_;
  wire _12476_;
  wire _12477_;
  wire _12478_;
  wire _12479_;
  wire _12480_;
  wire _12481_;
  wire _12482_;
  wire _12483_;
  wire _12484_;
  wire _12485_;
  wire _12486_;
  wire _12487_;
  wire _12488_;
  wire _12489_;
  wire _12490_;
  wire _12491_;
  wire _12492_;
  wire _12493_;
  wire _12494_;
  wire _12495_;
  wire _12496_;
  wire _12497_;
  wire _12498_;
  wire _12499_;
  wire _12500_;
  wire _12501_;
  wire _12502_;
  wire _12503_;
  wire _12504_;
  wire _12505_;
  wire _12506_;
  wire _12507_;
  wire _12508_;
  wire _12509_;
  wire _12510_;
  wire _12511_;
  wire _12512_;
  wire _12513_;
  wire _12514_;
  wire _12515_;
  wire _12516_;
  wire _12517_;
  wire _12518_;
  wire _12519_;
  wire _12520_;
  wire _12521_;
  wire _12522_;
  wire _12523_;
  wire _12524_;
  wire _12525_;
  wire _12526_;
  wire _12527_;
  wire _12528_;
  wire _12529_;
  wire _12530_;
  wire _12531_;
  wire _12532_;
  wire _12533_;
  wire _12534_;
  wire _12535_;
  wire _12536_;
  wire _12537_;
  wire _12538_;
  wire _12539_;
  wire _12540_;
  wire _12541_;
  wire _12542_;
  wire _12543_;
  wire _12544_;
  wire _12545_;
  wire _12546_;
  wire _12547_;
  wire _12548_;
  wire _12549_;
  wire _12550_;
  wire _12551_;
  wire _12552_;
  wire _12553_;
  wire _12554_;
  wire _12555_;
  wire _12556_;
  wire _12557_;
  wire _12558_;
  wire _12559_;
  wire _12560_;
  wire _12561_;
  wire _12562_;
  wire _12563_;
  wire _12564_;
  wire _12565_;
  wire _12566_;
  wire _12567_;
  wire _12568_;
  wire _12569_;
  wire _12570_;
  wire _12571_;
  wire _12572_;
  wire _12573_;
  wire _12574_;
  wire _12575_;
  wire _12576_;
  wire _12577_;
  wire _12578_;
  wire _12579_;
  wire _12580_;
  wire _12581_;
  wire _12582_;
  wire _12583_;
  wire _12584_;
  wire _12585_;
  wire _12586_;
  wire _12587_;
  wire _12588_;
  wire _12589_;
  wire _12590_;
  wire _12591_;
  wire _12592_;
  wire _12593_;
  wire _12594_;
  wire _12595_;
  wire _12596_;
  wire _12597_;
  wire _12598_;
  wire _12599_;
  wire _12600_;
  wire _12601_;
  wire _12602_;
  wire _12603_;
  wire _12604_;
  wire _12605_;
  wire _12606_;
  wire _12607_;
  wire _12608_;
  wire _12609_;
  wire _12610_;
  wire _12611_;
  wire _12612_;
  wire _12613_;
  wire _12614_;
  wire _12615_;
  wire _12616_;
  wire _12617_;
  wire _12618_;
  wire _12619_;
  wire _12620_;
  wire _12621_;
  wire _12622_;
  wire _12623_;
  wire _12624_;
  wire _12625_;
  wire _12626_;
  wire _12627_;
  wire _12628_;
  wire _12629_;
  wire _12630_;
  wire _12631_;
  wire _12632_;
  wire _12633_;
  wire _12634_;
  wire _12635_;
  wire _12636_;
  wire _12637_;
  wire _12638_;
  wire _12639_;
  wire _12640_;
  wire _12641_;
  wire _12642_;
  wire _12643_;
  wire _12644_;
  wire _12645_;
  wire _12646_;
  wire _12647_;
  wire _12648_;
  wire _12649_;
  wire _12650_;
  wire _12651_;
  wire _12652_;
  wire _12653_;
  wire _12654_;
  wire _12655_;
  wire _12656_;
  wire _12657_;
  wire _12658_;
  wire _12659_;
  wire _12660_;
  wire _12661_;
  wire _12662_;
  wire _12663_;
  wire _12664_;
  wire _12665_;
  wire _12666_;
  wire _12667_;
  wire _12668_;
  wire _12669_;
  wire _12670_;
  wire _12671_;
  wire _12672_;
  wire _12673_;
  wire _12674_;
  wire _12675_;
  wire _12676_;
  wire _12677_;
  wire _12678_;
  wire _12679_;
  wire _12680_;
  wire _12681_;
  wire _12682_;
  wire _12683_;
  wire _12684_;
  wire _12685_;
  wire _12686_;
  wire _12687_;
  wire _12688_;
  wire _12689_;
  wire _12690_;
  wire _12691_;
  wire _12692_;
  wire _12693_;
  wire _12694_;
  wire _12695_;
  wire _12696_;
  wire _12697_;
  wire _12698_;
  wire _12699_;
  wire _12700_;
  wire _12701_;
  wire _12702_;
  wire _12703_;
  wire _12704_;
  wire _12705_;
  wire _12706_;
  wire _12707_;
  wire _12708_;
  wire _12709_;
  wire _12710_;
  wire _12711_;
  wire _12712_;
  wire _12713_;
  wire _12714_;
  wire _12715_;
  wire _12716_;
  wire _12717_;
  wire _12718_;
  wire _12719_;
  wire _12720_;
  wire _12721_;
  wire _12722_;
  wire _12723_;
  wire _12724_;
  wire _12725_;
  wire _12726_;
  wire _12727_;
  wire _12728_;
  wire _12729_;
  wire _12730_;
  wire _12731_;
  wire _12732_;
  wire _12733_;
  wire _12734_;
  wire _12735_;
  wire _12736_;
  wire _12737_;
  wire _12738_;
  wire _12739_;
  wire _12740_;
  wire _12741_;
  wire _12742_;
  wire _12743_;
  wire _12744_;
  wire _12745_;
  wire _12746_;
  wire _12747_;
  wire _12748_;
  wire _12749_;
  wire _12750_;
  wire _12751_;
  wire _12752_;
  wire _12753_;
  wire _12754_;
  wire _12755_;
  wire _12756_;
  wire _12757_;
  wire _12758_;
  wire _12759_;
  wire _12760_;
  wire _12761_;
  wire _12762_;
  wire _12763_;
  wire _12764_;
  wire _12765_;
  wire _12766_;
  wire _12767_;
  wire _12768_;
  wire _12769_;
  wire _12770_;
  wire _12771_;
  wire _12772_;
  wire _12773_;
  wire _12774_;
  wire _12775_;
  wire _12776_;
  wire _12777_;
  wire _12778_;
  wire _12779_;
  wire _12780_;
  wire _12781_;
  wire _12782_;
  wire _12783_;
  wire _12784_;
  wire _12785_;
  wire _12786_;
  wire _12787_;
  wire _12788_;
  wire _12789_;
  wire _12790_;
  wire _12791_;
  wire _12792_;
  wire _12793_;
  wire _12794_;
  wire _12795_;
  wire _12796_;
  wire _12797_;
  wire _12798_;
  wire _12799_;
  wire _12800_;
  wire _12801_;
  wire _12802_;
  wire _12803_;
  wire _12804_;
  wire _12805_;
  wire _12806_;
  wire _12807_;
  wire _12808_;
  wire _12809_;
  wire _12810_;
  wire _12811_;
  wire _12812_;
  wire _12813_;
  wire _12814_;
  wire _12815_;
  wire _12816_;
  wire _12817_;
  wire _12818_;
  wire _12819_;
  wire _12820_;
  wire _12821_;
  wire _12822_;
  wire _12823_;
  wire _12824_;
  wire _12825_;
  wire _12826_;
  wire _12827_;
  wire _12828_;
  wire _12829_;
  wire _12830_;
  wire _12831_;
  wire _12832_;
  wire _12833_;
  wire _12834_;
  wire _12835_;
  wire _12836_;
  wire _12837_;
  wire _12838_;
  wire _12839_;
  wire _12840_;
  wire _12841_;
  wire _12842_;
  wire _12843_;
  wire _12844_;
  wire _12845_;
  wire _12846_;
  wire _12847_;
  wire _12848_;
  wire _12849_;
  wire _12850_;
  wire _12851_;
  wire _12852_;
  wire _12853_;
  wire _12854_;
  wire _12855_;
  wire _12856_;
  wire _12857_;
  wire _12858_;
  wire _12859_;
  wire _12860_;
  wire _12861_;
  wire _12862_;
  wire _12863_;
  wire _12864_;
  wire _12865_;
  wire _12866_;
  wire _12867_;
  wire _12868_;
  wire _12869_;
  wire _12870_;
  wire _12871_;
  wire _12872_;
  wire _12873_;
  wire _12874_;
  wire _12875_;
  wire _12876_;
  wire _12877_;
  wire _12878_;
  wire _12879_;
  wire _12880_;
  wire _12881_;
  wire _12882_;
  wire _12883_;
  wire _12884_;
  wire _12885_;
  wire _12886_;
  wire _12887_;
  wire _12888_;
  wire _12889_;
  wire _12890_;
  wire _12891_;
  wire _12892_;
  wire _12893_;
  wire _12894_;
  wire _12895_;
  wire _12896_;
  wire _12897_;
  wire _12898_;
  wire _12899_;
  wire _12900_;
  wire _12901_;
  wire _12902_;
  wire _12903_;
  wire _12904_;
  wire _12905_;
  wire _12906_;
  wire _12907_;
  wire _12908_;
  wire _12909_;
  wire _12910_;
  wire _12911_;
  wire _12912_;
  wire _12913_;
  wire _12914_;
  wire _12915_;
  wire _12916_;
  wire _12917_;
  wire _12918_;
  wire _12919_;
  wire _12920_;
  wire _12921_;
  wire _12922_;
  wire _12923_;
  wire _12924_;
  wire _12925_;
  wire _12926_;
  wire _12927_;
  wire _12928_;
  wire _12929_;
  wire _12930_;
  wire _12931_;
  wire _12932_;
  wire _12933_;
  wire _12934_;
  wire _12935_;
  wire _12936_;
  wire _12937_;
  wire _12938_;
  wire _12939_;
  wire _12940_;
  wire _12941_;
  wire _12942_;
  wire _12943_;
  wire _12944_;
  wire _12945_;
  wire _12946_;
  wire _12947_;
  wire _12948_;
  wire _12949_;
  wire _12950_;
  wire _12951_;
  wire _12952_;
  wire _12953_;
  wire _12954_;
  wire _12955_;
  wire _12956_;
  wire _12957_;
  wire _12958_;
  wire _12959_;
  wire _12960_;
  wire _12961_;
  wire _12962_;
  wire _12963_;
  wire _12964_;
  wire _12965_;
  wire _12966_;
  wire _12967_;
  wire _12968_;
  wire _12969_;
  wire _12970_;
  wire _12971_;
  wire _12972_;
  wire _12973_;
  wire _12974_;
  wire _12975_;
  wire _12976_;
  wire _12977_;
  wire _12978_;
  wire _12979_;
  wire _12980_;
  wire _12981_;
  wire _12982_;
  wire _12983_;
  wire _12984_;
  wire _12985_;
  wire _12986_;
  wire _12987_;
  wire _12988_;
  wire _12989_;
  wire _12990_;
  wire _12991_;
  wire _12992_;
  wire _12993_;
  wire _12994_;
  wire _12995_;
  wire _12996_;
  wire _12997_;
  wire _12998_;
  wire _12999_;
  wire _13000_;
  wire _13001_;
  wire _13002_;
  wire _13003_;
  wire _13004_;
  wire _13005_;
  wire _13006_;
  wire _13007_;
  wire _13008_;
  wire _13009_;
  wire _13010_;
  wire _13011_;
  wire _13012_;
  wire _13013_;
  wire _13014_;
  wire _13015_;
  wire _13016_;
  wire _13017_;
  wire _13018_;
  wire _13019_;
  wire _13020_;
  wire _13021_;
  wire _13022_;
  wire _13023_;
  wire _13024_;
  wire _13025_;
  wire _13026_;
  wire _13027_;
  wire _13028_;
  wire _13029_;
  wire _13030_;
  wire _13031_;
  wire _13032_;
  wire _13033_;
  wire _13034_;
  wire _13035_;
  wire _13036_;
  wire _13037_;
  wire _13038_;
  wire _13039_;
  wire _13040_;
  wire _13041_;
  wire _13042_;
  wire _13043_;
  wire _13044_;
  wire _13045_;
  wire _13046_;
  wire _13047_;
  wire _13048_;
  wire _13049_;
  wire _13050_;
  wire _13051_;
  wire _13052_;
  wire _13053_;
  wire _13054_;
  wire _13055_;
  wire _13056_;
  wire _13057_;
  wire _13058_;
  wire _13059_;
  wire _13060_;
  wire _13061_;
  wire _13062_;
  wire _13063_;
  wire _13064_;
  wire _13065_;
  wire _13066_;
  wire _13067_;
  wire _13068_;
  wire _13069_;
  wire _13070_;
  wire _13071_;
  wire _13072_;
  wire _13073_;
  wire _13074_;
  wire _13075_;
  wire _13076_;
  wire _13077_;
  wire _13078_;
  wire _13079_;
  wire _13080_;
  wire _13081_;
  wire _13082_;
  wire _13083_;
  wire _13084_;
  wire _13085_;
  wire _13086_;
  wire _13087_;
  wire _13088_;
  wire _13089_;
  wire _13090_;
  wire _13091_;
  wire _13092_;
  wire _13093_;
  wire _13094_;
  wire _13095_;
  wire _13096_;
  wire _13097_;
  wire _13098_;
  wire _13099_;
  wire _13100_;
  wire _13101_;
  wire _13102_;
  wire _13103_;
  wire _13104_;
  wire _13105_;
  wire _13106_;
  wire _13107_;
  wire _13108_;
  wire _13109_;
  wire _13110_;
  wire _13111_;
  wire _13112_;
  wire _13113_;
  wire _13114_;
  wire _13115_;
  wire _13116_;
  wire _13117_;
  wire _13118_;
  wire _13119_;
  wire _13120_;
  wire _13121_;
  wire _13122_;
  wire _13123_;
  wire _13124_;
  wire _13125_;
  wire _13126_;
  wire _13127_;
  wire _13128_;
  wire _13129_;
  wire _13130_;
  wire _13131_;
  wire _13132_;
  wire _13133_;
  wire _13134_;
  wire _13135_;
  wire _13136_;
  wire _13137_;
  wire _13138_;
  wire _13139_;
  wire _13140_;
  wire _13141_;
  wire _13142_;
  wire _13143_;
  wire _13144_;
  wire _13145_;
  wire _13146_;
  wire _13147_;
  wire _13148_;
  wire _13149_;
  wire _13150_;
  wire _13151_;
  wire _13152_;
  wire _13153_;
  wire _13154_;
  wire _13155_;
  wire _13156_;
  wire _13157_;
  wire _13158_;
  wire _13159_;
  wire _13160_;
  wire _13161_;
  wire _13162_;
  wire _13163_;
  wire _13164_;
  wire _13165_;
  wire _13166_;
  wire _13167_;
  wire _13168_;
  wire _13169_;
  wire _13170_;
  wire _13171_;
  wire _13172_;
  wire _13173_;
  wire _13174_;
  wire _13175_;
  wire _13176_;
  wire _13177_;
  wire _13178_;
  wire _13179_;
  wire _13180_;
  wire _13181_;
  wire _13182_;
  wire _13183_;
  wire _13184_;
  wire _13185_;
  wire _13186_;
  wire _13187_;
  wire _13188_;
  wire _13189_;
  wire _13190_;
  wire _13191_;
  wire _13192_;
  wire _13193_;
  wire _13194_;
  wire _13195_;
  wire _13196_;
  wire _13197_;
  wire _13198_;
  wire _13199_;
  wire _13200_;
  wire _13201_;
  wire _13202_;
  wire _13203_;
  wire _13204_;
  wire _13205_;
  wire _13206_;
  wire _13207_;
  wire _13208_;
  wire _13209_;
  wire _13210_;
  wire _13211_;
  wire _13212_;
  wire _13213_;
  wire _13214_;
  wire _13215_;
  wire _13216_;
  wire _13217_;
  wire _13218_;
  wire _13219_;
  wire _13220_;
  wire _13221_;
  wire _13222_;
  wire _13223_;
  wire _13224_;
  wire _13225_;
  wire _13226_;
  wire _13227_;
  wire _13228_;
  wire _13229_;
  wire _13230_;
  wire _13231_;
  wire _13232_;
  wire _13233_;
  wire _13234_;
  wire _13235_;
  wire _13236_;
  wire _13237_;
  wire _13238_;
  wire _13239_;
  wire _13240_;
  wire _13241_;
  wire _13242_;
  wire _13243_;
  wire _13244_;
  wire _13245_;
  wire _13246_;
  wire _13247_;
  wire _13248_;
  wire _13249_;
  wire _13250_;
  wire _13251_;
  wire _13252_;
  wire _13253_;
  wire _13254_;
  wire _13255_;
  wire _13256_;
  wire _13257_;
  wire _13258_;
  wire _13259_;
  wire _13260_;
  wire _13261_;
  wire _13262_;
  wire _13263_;
  wire _13264_;
  wire _13265_;
  wire _13266_;
  wire _13267_;
  wire _13268_;
  wire _13269_;
  wire _13270_;
  wire _13271_;
  wire _13272_;
  wire _13273_;
  wire _13274_;
  wire _13275_;
  wire _13276_;
  wire _13277_;
  wire _13278_;
  wire _13279_;
  wire _13280_;
  wire _13281_;
  wire _13282_;
  wire _13283_;
  wire _13284_;
  wire _13285_;
  wire _13286_;
  wire _13287_;
  wire _13288_;
  wire _13289_;
  wire _13290_;
  wire _13291_;
  wire _13292_;
  wire _13293_;
  wire _13294_;
  wire _13295_;
  wire _13296_;
  wire _13297_;
  wire _13298_;
  wire _13299_;
  wire _13300_;
  wire _13301_;
  wire _13302_;
  wire _13303_;
  wire _13304_;
  wire _13305_;
  wire _13306_;
  wire _13307_;
  wire _13308_;
  wire _13309_;
  wire _13310_;
  wire _13311_;
  wire _13312_;
  wire _13313_;
  wire _13314_;
  wire _13315_;
  wire _13316_;
  wire _13317_;
  wire _13318_;
  wire _13319_;
  wire _13320_;
  wire _13321_;
  wire _13322_;
  wire _13323_;
  wire _13324_;
  wire _13325_;
  wire _13326_;
  wire _13327_;
  wire _13328_;
  wire _13329_;
  wire _13330_;
  wire _13331_;
  wire _13332_;
  wire _13333_;
  wire _13334_;
  wire _13335_;
  wire _13336_;
  wire _13337_;
  wire _13338_;
  wire _13339_;
  wire _13340_;
  wire _13341_;
  wire _13342_;
  wire _13343_;
  wire _13344_;
  wire _13345_;
  wire _13346_;
  wire _13347_;
  wire _13348_;
  wire _13349_;
  wire _13350_;
  wire _13351_;
  wire _13352_;
  wire _13353_;
  wire _13354_;
  wire _13355_;
  wire _13356_;
  wire _13357_;
  wire _13358_;
  wire _13359_;
  wire _13360_;
  wire _13361_;
  wire _13362_;
  wire _13363_;
  wire _13364_;
  wire _13365_;
  wire _13366_;
  wire _13367_;
  wire _13368_;
  wire _13369_;
  wire _13370_;
  wire _13371_;
  wire _13372_;
  wire _13373_;
  wire _13374_;
  wire _13375_;
  wire _13376_;
  wire _13377_;
  wire _13378_;
  wire _13379_;
  wire _13380_;
  wire _13381_;
  wire _13382_;
  wire _13383_;
  wire _13384_;
  wire _13385_;
  wire _13386_;
  wire _13387_;
  wire _13388_;
  wire _13389_;
  wire _13390_;
  wire _13391_;
  wire _13392_;
  wire _13393_;
  wire _13394_;
  wire _13395_;
  wire _13396_;
  wire _13397_;
  wire _13398_;
  wire _13399_;
  wire _13400_;
  wire _13401_;
  wire _13402_;
  wire _13403_;
  wire _13404_;
  wire _13405_;
  wire _13406_;
  wire _13407_;
  wire _13408_;
  wire _13409_;
  wire _13410_;
  wire _13411_;
  wire _13412_;
  wire _13413_;
  wire _13414_;
  wire _13415_;
  wire _13416_;
  wire _13417_;
  wire _13418_;
  wire _13419_;
  wire _13420_;
  wire _13421_;
  wire _13422_;
  wire _13423_;
  wire _13424_;
  wire _13425_;
  wire _13426_;
  wire _13427_;
  wire _13428_;
  wire _13429_;
  wire _13430_;
  wire _13431_;
  wire _13432_;
  wire _13433_;
  wire _13434_;
  wire _13435_;
  wire _13436_;
  wire _13437_;
  wire _13438_;
  wire _13439_;
  wire _13440_;
  wire _13441_;
  wire _13442_;
  wire _13443_;
  wire _13444_;
  wire _13445_;
  wire _13446_;
  wire _13447_;
  wire _13448_;
  wire _13449_;
  wire _13450_;
  wire _13451_;
  wire _13452_;
  wire _13453_;
  wire _13454_;
  wire _13455_;
  wire _13456_;
  wire _13457_;
  wire _13458_;
  wire _13459_;
  wire _13460_;
  wire _13461_;
  wire _13462_;
  wire _13463_;
  wire _13464_;
  wire _13465_;
  wire _13466_;
  wire _13467_;
  wire _13468_;
  wire _13469_;
  wire _13470_;
  wire _13471_;
  wire _13472_;
  wire _13473_;
  wire _13474_;
  wire _13475_;
  wire _13476_;
  wire _13477_;
  wire _13478_;
  wire _13479_;
  wire _13480_;
  wire _13481_;
  wire _13482_;
  wire _13483_;
  wire _13484_;
  wire _13485_;
  wire _13486_;
  wire _13487_;
  wire _13488_;
  wire _13489_;
  wire _13490_;
  wire _13491_;
  wire _13492_;
  wire _13493_;
  wire _13494_;
  wire _13495_;
  wire _13496_;
  wire _13497_;
  wire _13498_;
  wire _13499_;
  wire _13500_;
  wire _13501_;
  wire _13502_;
  wire _13503_;
  wire _13504_;
  wire _13505_;
  wire _13506_;
  wire _13507_;
  wire _13508_;
  wire _13509_;
  wire _13510_;
  wire _13511_;
  wire _13512_;
  wire _13513_;
  wire _13514_;
  wire _13515_;
  wire _13516_;
  wire _13517_;
  wire _13518_;
  wire _13519_;
  wire _13520_;
  wire _13521_;
  wire _13522_;
  wire _13523_;
  wire _13524_;
  wire _13525_;
  wire _13526_;
  wire _13527_;
  wire _13528_;
  wire _13529_;
  wire _13530_;
  wire _13531_;
  wire _13532_;
  wire _13533_;
  wire _13534_;
  wire _13535_;
  wire _13536_;
  wire _13537_;
  wire _13538_;
  wire _13539_;
  wire _13540_;
  wire _13541_;
  wire _13542_;
  wire _13543_;
  wire _13544_;
  wire _13545_;
  wire _13546_;
  wire _13547_;
  wire _13548_;
  wire _13549_;
  wire _13550_;
  wire _13551_;
  wire _13552_;
  wire _13553_;
  wire _13554_;
  wire _13555_;
  wire _13556_;
  wire _13557_;
  wire _13558_;
  wire _13559_;
  wire _13560_;
  wire _13561_;
  wire _13562_;
  wire _13563_;
  wire _13564_;
  wire _13565_;
  wire _13566_;
  wire _13567_;
  wire _13568_;
  wire _13569_;
  wire _13570_;
  wire _13571_;
  wire _13572_;
  wire _13573_;
  wire _13574_;
  wire _13575_;
  wire _13576_;
  wire _13577_;
  wire _13578_;
  wire _13579_;
  wire _13580_;
  wire _13581_;
  wire _13582_;
  wire _13583_;
  wire _13584_;
  wire _13585_;
  wire _13586_;
  wire _13587_;
  wire _13588_;
  wire _13589_;
  wire _13590_;
  wire _13591_;
  wire _13592_;
  wire _13593_;
  wire _13594_;
  wire _13595_;
  wire _13596_;
  wire _13597_;
  wire _13598_;
  wire _13599_;
  wire _13600_;
  wire _13601_;
  wire _13602_;
  wire _13603_;
  wire _13604_;
  wire _13605_;
  wire _13606_;
  wire _13607_;
  wire _13608_;
  wire _13609_;
  wire _13610_;
  wire _13611_;
  wire _13612_;
  wire _13613_;
  wire _13614_;
  wire _13615_;
  wire _13616_;
  wire _13617_;
  wire _13618_;
  wire _13619_;
  wire _13620_;
  wire _13621_;
  wire _13622_;
  wire _13623_;
  wire _13624_;
  wire _13625_;
  wire _13626_;
  wire _13627_;
  wire _13628_;
  wire _13629_;
  wire _13630_;
  wire _13631_;
  wire _13632_;
  wire _13633_;
  wire _13634_;
  wire _13635_;
  wire _13636_;
  wire _13637_;
  wire _13638_;
  wire _13639_;
  wire _13640_;
  wire _13641_;
  wire _13642_;
  wire _13643_;
  wire _13644_;
  wire _13645_;
  wire _13646_;
  wire _13647_;
  wire _13648_;
  wire _13649_;
  wire _13650_;
  wire _13651_;
  wire _13652_;
  wire _13653_;
  wire _13654_;
  wire _13655_;
  wire _13656_;
  wire _13657_;
  wire _13658_;
  wire _13659_;
  wire _13660_;
  wire _13661_;
  wire _13662_;
  wire _13663_;
  wire _13664_;
  wire _13665_;
  wire _13666_;
  wire _13667_;
  wire _13668_;
  wire _13669_;
  wire _13670_;
  wire _13671_;
  wire _13672_;
  wire _13673_;
  wire _13674_;
  wire _13675_;
  wire _13676_;
  wire _13677_;
  wire _13678_;
  wire _13679_;
  wire _13680_;
  wire _13681_;
  wire _13682_;
  wire _13683_;
  wire _13684_;
  wire _13685_;
  wire _13686_;
  wire _13687_;
  wire _13688_;
  wire _13689_;
  wire _13690_;
  wire _13691_;
  wire _13692_;
  wire _13693_;
  wire _13694_;
  wire _13695_;
  wire _13696_;
  wire _13697_;
  wire _13698_;
  wire _13699_;
  wire _13700_;
  wire _13701_;
  wire _13702_;
  wire _13703_;
  wire _13704_;
  wire _13705_;
  wire _13706_;
  wire _13707_;
  wire _13708_;
  wire _13709_;
  wire _13710_;
  wire _13711_;
  wire _13712_;
  wire _13713_;
  wire _13714_;
  wire _13715_;
  wire _13716_;
  wire _13717_;
  wire _13718_;
  wire _13719_;
  wire _13720_;
  wire _13721_;
  wire _13722_;
  wire _13723_;
  wire _13724_;
  wire _13725_;
  wire _13726_;
  wire _13727_;
  wire _13728_;
  wire _13729_;
  wire _13730_;
  wire _13731_;
  wire _13732_;
  wire _13733_;
  wire _13734_;
  wire _13735_;
  wire _13736_;
  wire _13737_;
  wire _13738_;
  wire _13739_;
  wire _13740_;
  wire _13741_;
  wire _13742_;
  wire _13743_;
  wire _13744_;
  wire _13745_;
  wire _13746_;
  wire _13747_;
  wire _13748_;
  wire _13749_;
  wire _13750_;
  wire _13751_;
  wire _13752_;
  wire _13753_;
  wire _13754_;
  wire _13755_;
  wire _13756_;
  wire _13757_;
  wire _13758_;
  wire _13759_;
  wire _13760_;
  wire _13761_;
  wire _13762_;
  wire _13763_;
  wire _13764_;
  wire _13765_;
  wire _13766_;
  wire _13767_;
  wire _13768_;
  wire _13769_;
  wire _13770_;
  wire _13771_;
  wire _13772_;
  wire _13773_;
  wire _13774_;
  wire _13775_;
  wire _13776_;
  wire _13777_;
  wire _13778_;
  wire _13779_;
  wire _13780_;
  wire _13781_;
  wire _13782_;
  wire _13783_;
  wire _13784_;
  wire _13785_;
  wire _13786_;
  wire _13787_;
  wire _13788_;
  wire _13789_;
  wire _13790_;
  wire _13791_;
  wire _13792_;
  wire _13793_;
  wire _13794_;
  wire _13795_;
  wire _13796_;
  wire _13797_;
  wire _13798_;
  wire _13799_;
  wire _13800_;
  wire _13801_;
  wire _13802_;
  wire _13803_;
  wire _13804_;
  wire _13805_;
  wire _13806_;
  wire _13807_;
  wire _13808_;
  wire _13809_;
  wire _13810_;
  wire _13811_;
  wire _13812_;
  wire _13813_;
  wire _13814_;
  wire _13815_;
  wire _13816_;
  wire _13817_;
  wire _13818_;
  wire _13819_;
  wire _13820_;
  wire _13821_;
  wire _13822_;
  wire _13823_;
  wire _13824_;
  wire _13825_;
  wire _13826_;
  wire _13827_;
  wire _13828_;
  wire _13829_;
  wire _13830_;
  wire _13831_;
  wire _13832_;
  wire _13833_;
  wire _13834_;
  wire _13835_;
  wire _13836_;
  wire _13837_;
  wire _13838_;
  wire _13839_;
  wire _13840_;
  wire _13841_;
  wire _13842_;
  wire _13843_;
  wire _13844_;
  wire _13845_;
  wire _13846_;
  wire _13847_;
  wire _13848_;
  wire _13849_;
  wire _13850_;
  wire _13851_;
  wire _13852_;
  wire _13853_;
  wire _13854_;
  wire _13855_;
  wire _13856_;
  wire _13857_;
  wire _13858_;
  wire _13859_;
  wire _13860_;
  wire _13861_;
  wire _13862_;
  wire _13863_;
  wire _13864_;
  wire _13865_;
  wire _13866_;
  wire _13867_;
  wire _13868_;
  wire _13869_;
  wire _13870_;
  wire _13871_;
  wire _13872_;
  wire _13873_;
  wire _13874_;
  wire _13875_;
  wire _13876_;
  wire _13877_;
  wire _13878_;
  wire _13879_;
  wire _13880_;
  wire _13881_;
  wire _13882_;
  wire _13883_;
  wire _13884_;
  wire _13885_;
  wire _13886_;
  wire _13887_;
  wire _13888_;
  wire _13889_;
  wire _13890_;
  wire _13891_;
  wire _13892_;
  wire _13893_;
  wire _13894_;
  wire _13895_;
  wire _13896_;
  wire _13897_;
  wire _13898_;
  wire _13899_;
  wire _13900_;
  wire _13901_;
  wire _13902_;
  wire _13903_;
  wire _13904_;
  wire _13905_;
  wire _13906_;
  wire _13907_;
  wire _13908_;
  wire _13909_;
  wire _13910_;
  wire _13911_;
  wire _13912_;
  wire _13913_;
  wire _13914_;
  wire _13915_;
  wire _13916_;
  wire _13917_;
  wire _13918_;
  wire _13919_;
  wire _13920_;
  wire _13921_;
  wire _13922_;
  wire _13923_;
  wire _13924_;
  wire _13925_;
  wire _13926_;
  wire _13927_;
  wire _13928_;
  wire _13929_;
  wire _13930_;
  wire _13931_;
  wire _13932_;
  wire _13933_;
  wire _13934_;
  wire _13935_;
  wire _13936_;
  wire _13937_;
  wire _13938_;
  wire _13939_;
  wire _13940_;
  wire _13941_;
  wire _13942_;
  wire _13943_;
  wire _13944_;
  wire _13945_;
  wire _13946_;
  wire _13947_;
  wire _13948_;
  wire _13949_;
  wire _13950_;
  wire _13951_;
  wire _13952_;
  wire _13953_;
  wire _13954_;
  wire _13955_;
  wire _13956_;
  wire _13957_;
  wire _13958_;
  wire _13959_;
  wire _13960_;
  wire _13961_;
  wire _13962_;
  wire _13963_;
  wire _13964_;
  wire _13965_;
  wire _13966_;
  wire _13967_;
  wire _13968_;
  wire _13969_;
  wire _13970_;
  wire _13971_;
  wire _13972_;
  wire _13973_;
  wire _13974_;
  wire _13975_;
  wire _13976_;
  wire _13977_;
  wire _13978_;
  wire _13979_;
  wire _13980_;
  wire _13981_;
  wire _13982_;
  wire _13983_;
  wire _13984_;
  wire _13985_;
  wire _13986_;
  wire _13987_;
  wire _13988_;
  wire _13989_;
  wire _13990_;
  wire _13991_;
  wire _13992_;
  wire _13993_;
  wire _13994_;
  wire _13995_;
  wire _13996_;
  wire _13997_;
  wire _13998_;
  wire _13999_;
  wire _14000_;
  wire _14001_;
  wire _14002_;
  wire _14003_;
  wire _14004_;
  wire _14005_;
  wire _14006_;
  wire _14007_;
  wire _14008_;
  wire _14009_;
  wire _14010_;
  wire _14011_;
  wire _14012_;
  wire _14013_;
  wire _14014_;
  wire _14015_;
  wire _14016_;
  wire _14017_;
  wire _14018_;
  wire _14019_;
  wire _14020_;
  wire _14021_;
  wire _14022_;
  wire _14023_;
  wire _14024_;
  wire _14025_;
  wire _14026_;
  wire _14027_;
  wire _14028_;
  wire _14029_;
  wire _14030_;
  wire _14031_;
  wire _14032_;
  wire _14033_;
  wire _14034_;
  wire _14035_;
  wire _14036_;
  wire _14037_;
  wire _14038_;
  wire _14039_;
  wire _14040_;
  wire _14041_;
  wire _14042_;
  wire _14043_;
  wire _14044_;
  wire _14045_;
  wire _14046_;
  wire _14047_;
  wire _14048_;
  wire _14049_;
  wire _14050_;
  wire _14051_;
  wire _14052_;
  wire _14053_;
  wire _14054_;
  wire _14055_;
  wire _14056_;
  wire _14057_;
  wire _14058_;
  wire _14059_;
  wire _14060_;
  wire _14061_;
  wire _14062_;
  wire _14063_;
  wire _14064_;
  wire _14065_;
  wire _14066_;
  wire _14067_;
  wire _14068_;
  wire _14069_;
  wire _14070_;
  wire _14071_;
  wire _14072_;
  wire _14073_;
  wire _14074_;
  wire _14075_;
  wire _14076_;
  wire _14077_;
  wire _14078_;
  wire _14079_;
  wire _14080_;
  wire _14081_;
  wire _14082_;
  wire _14083_;
  wire _14084_;
  wire _14085_;
  wire _14086_;
  wire _14087_;
  wire _14088_;
  wire _14089_;
  wire _14090_;
  wire _14091_;
  wire _14092_;
  wire _14093_;
  wire _14094_;
  wire _14095_;
  wire _14096_;
  wire _14097_;
  wire _14098_;
  wire _14099_;
  wire _14100_;
  wire _14101_;
  wire _14102_;
  wire _14103_;
  wire _14104_;
  wire _14105_;
  wire _14106_;
  wire _14107_;
  wire _14108_;
  wire _14109_;
  wire _14110_;
  wire _14111_;
  wire _14112_;
  wire _14113_;
  wire _14114_;
  wire _14115_;
  wire _14116_;
  wire _14117_;
  wire _14118_;
  wire _14119_;
  wire _14120_;
  wire _14121_;
  wire _14122_;
  wire _14123_;
  wire _14124_;
  wire _14125_;
  wire _14126_;
  wire _14127_;
  wire _14128_;
  wire _14129_;
  wire _14130_;
  wire _14131_;
  wire _14132_;
  wire _14133_;
  wire _14134_;
  wire _14135_;
  wire _14136_;
  wire _14137_;
  wire _14138_;
  wire _14139_;
  wire _14140_;
  wire _14141_;
  wire _14142_;
  wire _14143_;
  wire _14144_;
  wire _14145_;
  wire _14146_;
  wire _14147_;
  wire _14148_;
  wire _14149_;
  wire _14150_;
  wire _14151_;
  wire _14152_;
  wire _14153_;
  wire _14154_;
  wire _14155_;
  wire _14156_;
  wire _14157_;
  wire _14158_;
  wire _14159_;
  wire _14160_;
  wire _14161_;
  wire _14162_;
  wire _14163_;
  wire _14164_;
  wire _14165_;
  wire _14166_;
  wire _14167_;
  wire _14168_;
  wire _14169_;
  wire _14170_;
  wire _14171_;
  wire _14172_;
  wire _14173_;
  wire _14174_;
  wire _14175_;
  wire _14176_;
  wire _14177_;
  wire _14178_;
  wire _14179_;
  wire _14180_;
  wire _14181_;
  wire _14182_;
  wire _14183_;
  wire _14184_;
  wire _14185_;
  wire _14186_;
  wire _14187_;
  wire _14188_;
  wire _14189_;
  wire _14190_;
  wire _14191_;
  wire _14192_;
  wire _14193_;
  wire _14194_;
  wire _14195_;
  wire _14196_;
  wire _14197_;
  wire _14198_;
  wire _14199_;
  wire _14200_;
  wire _14201_;
  wire _14202_;
  wire _14203_;
  wire _14204_;
  wire _14205_;
  wire _14206_;
  wire _14207_;
  wire _14208_;
  wire _14209_;
  wire _14210_;
  wire _14211_;
  wire _14212_;
  wire _14213_;
  wire _14214_;
  wire _14215_;
  wire _14216_;
  wire _14217_;
  wire _14218_;
  wire _14219_;
  wire _14220_;
  wire _14221_;
  wire _14222_;
  wire _14223_;
  wire _14224_;
  wire _14225_;
  wire _14226_;
  wire _14227_;
  wire _14228_;
  wire _14229_;
  wire _14230_;
  wire _14231_;
  wire _14232_;
  wire _14233_;
  wire _14234_;
  wire _14235_;
  wire _14236_;
  wire _14237_;
  wire _14238_;
  wire _14239_;
  wire _14240_;
  wire _14241_;
  wire _14242_;
  wire _14243_;
  wire _14244_;
  wire _14245_;
  wire _14246_;
  wire _14247_;
  wire _14248_;
  wire _14249_;
  wire _14250_;
  wire _14251_;
  wire _14252_;
  wire _14253_;
  wire _14254_;
  wire _14255_;
  wire _14256_;
  wire _14257_;
  wire _14258_;
  wire _14259_;
  wire _14260_;
  wire _14261_;
  wire _14262_;
  wire _14263_;
  wire _14264_;
  wire _14265_;
  wire _14266_;
  wire _14267_;
  wire _14268_;
  wire _14269_;
  wire _14270_;
  wire _14271_;
  wire _14272_;
  wire _14273_;
  wire _14274_;
  wire _14275_;
  wire _14276_;
  wire _14277_;
  wire _14278_;
  wire _14279_;
  wire _14280_;
  wire _14281_;
  wire _14282_;
  wire _14283_;
  wire _14284_;
  wire _14285_;
  wire _14286_;
  wire _14287_;
  wire _14288_;
  wire _14289_;
  wire _14290_;
  wire _14291_;
  wire _14292_;
  wire _14293_;
  wire _14294_;
  wire _14295_;
  wire _14296_;
  wire _14297_;
  wire _14298_;
  wire _14299_;
  wire _14300_;
  wire _14301_;
  wire _14302_;
  wire _14303_;
  wire _14304_;
  wire _14305_;
  wire _14306_;
  wire _14307_;
  wire _14308_;
  wire _14309_;
  wire _14310_;
  wire _14311_;
  wire _14312_;
  wire _14313_;
  wire _14314_;
  wire _14315_;
  wire _14316_;
  wire _14317_;
  wire _14318_;
  wire _14319_;
  wire _14320_;
  wire _14321_;
  wire _14322_;
  wire _14323_;
  wire _14324_;
  wire _14325_;
  wire _14326_;
  wire _14327_;
  wire _14328_;
  wire _14329_;
  wire _14330_;
  wire _14331_;
  wire _14332_;
  wire _14333_;
  wire _14334_;
  wire _14335_;
  wire _14336_;
  wire _14337_;
  wire _14338_;
  wire _14339_;
  wire _14340_;
  wire _14341_;
  wire _14342_;
  wire _14343_;
  wire _14344_;
  wire _14345_;
  wire _14346_;
  wire _14347_;
  wire _14348_;
  wire _14349_;
  wire _14350_;
  wire _14351_;
  wire _14352_;
  wire _14353_;
  wire _14354_;
  wire _14355_;
  wire _14356_;
  wire _14357_;
  wire _14358_;
  wire _14359_;
  wire _14360_;
  wire _14361_;
  wire _14362_;
  wire _14363_;
  wire _14364_;
  wire _14365_;
  wire _14366_;
  wire _14367_;
  wire _14368_;
  wire _14369_;
  wire _14370_;
  wire _14371_;
  wire _14372_;
  wire _14373_;
  wire _14374_;
  wire _14375_;
  wire _14376_;
  wire _14377_;
  wire _14378_;
  wire _14379_;
  wire _14380_;
  wire _14381_;
  wire _14382_;
  wire _14383_;
  wire _14384_;
  wire _14385_;
  wire _14386_;
  wire _14387_;
  wire _14388_;
  wire _14389_;
  wire _14390_;
  wire _14391_;
  wire _14392_;
  wire _14393_;
  wire _14394_;
  wire _14395_;
  wire _14396_;
  wire _14397_;
  wire _14398_;
  wire _14399_;
  wire _14400_;
  wire _14401_;
  wire _14402_;
  wire _14403_;
  wire _14404_;
  wire _14405_;
  wire _14406_;
  wire _14407_;
  wire _14408_;
  wire _14409_;
  wire _14410_;
  wire _14411_;
  wire _14412_;
  wire _14413_;
  wire _14414_;
  wire _14415_;
  wire _14416_;
  wire _14417_;
  wire _14418_;
  wire _14419_;
  wire _14420_;
  wire _14421_;
  wire _14422_;
  wire _14423_;
  wire _14424_;
  wire _14425_;
  wire _14426_;
  wire _14427_;
  wire _14428_;
  wire _14429_;
  wire _14430_;
  wire _14431_;
  wire _14432_;
  wire _14433_;
  wire _14434_;
  wire _14435_;
  wire _14436_;
  wire _14437_;
  wire _14438_;
  wire _14439_;
  wire _14440_;
  wire _14441_;
  wire _14442_;
  wire _14443_;
  wire _14444_;
  wire _14445_;
  wire _14446_;
  wire _14447_;
  wire _14448_;
  wire _14449_;
  wire _14450_;
  wire _14451_;
  wire _14452_;
  wire _14453_;
  wire _14454_;
  wire _14455_;
  wire _14456_;
  wire _14457_;
  wire _14458_;
  wire _14459_;
  wire _14460_;
  wire _14461_;
  wire _14462_;
  wire _14463_;
  wire _14464_;
  wire _14465_;
  wire _14466_;
  wire _14467_;
  wire _14468_;
  wire _14469_;
  wire _14470_;
  wire _14471_;
  wire _14472_;
  wire _14473_;
  wire _14474_;
  wire _14475_;
  wire _14476_;
  wire _14477_;
  wire _14478_;
  wire _14479_;
  wire _14480_;
  wire _14481_;
  wire _14482_;
  wire _14483_;
  wire _14484_;
  wire _14485_;
  wire _14486_;
  wire _14487_;
  wire _14488_;
  wire _14489_;
  wire _14490_;
  wire _14491_;
  wire _14492_;
  wire _14493_;
  wire _14494_;
  wire _14495_;
  wire _14496_;
  wire _14497_;
  wire _14498_;
  wire _14499_;
  wire _14500_;
  wire _14501_;
  wire _14502_;
  wire _14503_;
  wire _14504_;
  wire _14505_;
  wire _14506_;
  wire _14507_;
  wire _14508_;
  wire _14509_;
  wire _14510_;
  wire _14511_;
  wire _14512_;
  wire _14513_;
  wire _14514_;
  wire _14515_;
  wire _14516_;
  wire _14517_;
  wire _14518_;
  wire _14519_;
  wire _14520_;
  wire _14521_;
  wire _14522_;
  wire _14523_;
  wire _14524_;
  wire _14525_;
  wire _14526_;
  wire _14527_;
  wire _14528_;
  wire _14529_;
  wire _14530_;
  wire _14531_;
  wire _14532_;
  wire _14533_;
  wire _14534_;
  wire _14535_;
  wire _14536_;
  wire _14537_;
  wire _14538_;
  wire _14539_;
  wire _14540_;
  wire _14541_;
  wire _14542_;
  wire _14543_;
  wire _14544_;
  wire _14545_;
  wire _14546_;
  wire _14547_;
  wire _14548_;
  wire _14549_;
  wire _14550_;
  wire _14551_;
  wire _14552_;
  wire _14553_;
  wire _14554_;
  wire _14555_;
  wire _14556_;
  wire _14557_;
  wire _14558_;
  wire _14559_;
  wire _14560_;
  wire _14561_;
  wire _14562_;
  wire _14563_;
  wire _14564_;
  wire _14565_;
  wire _14566_;
  wire _14567_;
  wire _14568_;
  wire _14569_;
  wire _14570_;
  wire _14571_;
  wire _14572_;
  wire _14573_;
  wire _14574_;
  wire _14575_;
  wire _14576_;
  wire _14577_;
  wire _14578_;
  wire _14579_;
  wire _14580_;
  wire _14581_;
  wire _14582_;
  wire _14583_;
  wire _14584_;
  wire _14585_;
  wire _14586_;
  wire _14587_;
  wire _14588_;
  wire _14589_;
  wire _14590_;
  wire _14591_;
  wire _14592_;
  wire _14593_;
  wire _14594_;
  wire _14595_;
  wire _14596_;
  wire _14597_;
  wire _14598_;
  wire _14599_;
  wire _14600_;
  wire _14601_;
  wire _14602_;
  wire _14603_;
  wire _14604_;
  wire _14605_;
  wire _14606_;
  wire _14607_;
  wire _14608_;
  wire _14609_;
  wire _14610_;
  wire _14611_;
  wire _14612_;
  wire _14613_;
  wire _14614_;
  wire _14615_;
  wire _14616_;
  wire _14617_;
  wire _14618_;
  wire _14619_;
  wire _14620_;
  wire _14621_;
  wire _14622_;
  wire _14623_;
  wire _14624_;
  wire _14625_;
  wire _14626_;
  wire _14627_;
  wire _14628_;
  wire _14629_;
  wire _14630_;
  wire _14631_;
  wire _14632_;
  wire _14633_;
  wire _14634_;
  wire _14635_;
  wire _14636_;
  wire _14637_;
  wire _14638_;
  wire _14639_;
  wire _14640_;
  wire _14641_;
  wire _14642_;
  wire _14643_;
  wire _14644_;
  wire _14645_;
  wire _14646_;
  wire _14647_;
  wire _14648_;
  wire _14649_;
  wire _14650_;
  wire _14651_;
  wire _14652_;
  wire _14653_;
  wire _14654_;
  wire _14655_;
  wire _14656_;
  wire _14657_;
  wire _14658_;
  wire _14659_;
  wire _14660_;
  wire _14661_;
  wire _14662_;
  wire _14663_;
  wire _14664_;
  wire _14665_;
  wire _14666_;
  wire _14667_;
  wire _14668_;
  wire _14669_;
  wire _14670_;
  wire _14671_;
  wire _14672_;
  wire _14673_;
  wire _14674_;
  wire _14675_;
  wire _14676_;
  wire _14677_;
  wire _14678_;
  wire _14679_;
  wire _14680_;
  wire _14681_;
  wire _14682_;
  wire _14683_;
  wire _14684_;
  wire _14685_;
  wire _14686_;
  wire _14687_;
  wire _14688_;
  wire _14689_;
  wire _14690_;
  wire _14691_;
  wire _14692_;
  wire _14693_;
  wire _14694_;
  wire _14695_;
  wire _14696_;
  wire _14697_;
  wire _14698_;
  wire _14699_;
  wire _14700_;
  wire _14701_;
  wire _14702_;
  wire _14703_;
  wire _14704_;
  wire _14705_;
  wire _14706_;
  wire _14707_;
  wire _14708_;
  wire _14709_;
  wire _14710_;
  wire _14711_;
  wire _14712_;
  wire _14713_;
  wire _14714_;
  wire _14715_;
  wire _14716_;
  wire _14717_;
  wire _14718_;
  wire _14719_;
  wire _14720_;
  wire _14721_;
  wire _14722_;
  wire _14723_;
  wire _14724_;
  wire _14725_;
  wire _14726_;
  wire _14727_;
  wire _14728_;
  wire _14729_;
  wire _14730_;
  wire _14731_;
  wire _14732_;
  wire _14733_;
  wire _14734_;
  wire _14735_;
  wire _14736_;
  wire _14737_;
  wire _14738_;
  wire _14739_;
  wire _14740_;
  wire _14741_;
  wire _14742_;
  wire _14743_;
  wire _14744_;
  wire _14745_;
  wire _14746_;
  wire _14747_;
  wire _14748_;
  wire _14749_;
  wire _14750_;
  wire _14751_;
  wire _14752_;
  wire _14753_;
  wire _14754_;
  wire _14755_;
  wire _14756_;
  wire _14757_;
  wire _14758_;
  wire _14759_;
  wire _14760_;
  wire _14761_;
  wire _14762_;
  wire _14763_;
  wire _14764_;
  wire _14765_;
  wire _14766_;
  wire _14767_;
  wire _14768_;
  wire _14769_;
  wire _14770_;
  wire _14771_;
  wire _14772_;
  wire _14773_;
  wire _14774_;
  wire _14775_;
  wire _14776_;
  wire _14777_;
  wire _14778_;
  wire _14779_;
  wire _14780_;
  wire _14781_;
  wire _14782_;
  wire _14783_;
  wire _14784_;
  wire _14785_;
  wire _14786_;
  wire _14787_;
  wire _14788_;
  wire _14789_;
  wire _14790_;
  wire _14791_;
  wire _14792_;
  wire _14793_;
  wire _14794_;
  wire _14795_;
  wire _14796_;
  wire _14797_;
  wire _14798_;
  wire _14799_;
  wire _14800_;
  wire _14801_;
  wire _14802_;
  wire _14803_;
  wire _14804_;
  wire _14805_;
  wire _14806_;
  wire _14807_;
  wire _14808_;
  wire _14809_;
  wire _14810_;
  wire _14811_;
  wire _14812_;
  wire _14813_;
  wire _14814_;
  wire _14815_;
  wire _14816_;
  wire _14817_;
  wire _14818_;
  wire _14819_;
  wire _14820_;
  wire _14821_;
  wire _14822_;
  wire _14823_;
  wire _14824_;
  wire _14825_;
  wire _14826_;
  wire _14827_;
  wire _14828_;
  wire _14829_;
  wire _14830_;
  wire _14831_;
  wire _14832_;
  wire _14833_;
  wire _14834_;
  wire _14835_;
  wire _14836_;
  wire _14837_;
  wire _14838_;
  wire _14839_;
  wire _14840_;
  wire _14841_;
  wire _14842_;
  wire _14843_;
  wire _14844_;
  wire _14845_;
  wire _14846_;
  wire _14847_;
  wire _14848_;
  wire _14849_;
  wire _14850_;
  wire _14851_;
  wire _14852_;
  wire _14853_;
  wire _14854_;
  wire _14855_;
  wire _14856_;
  wire _14857_;
  wire _14858_;
  wire _14859_;
  wire _14860_;
  wire _14861_;
  wire _14862_;
  wire _14863_;
  wire _14864_;
  wire _14865_;
  wire _14866_;
  wire _14867_;
  wire _14868_;
  wire _14869_;
  wire _14870_;
  wire _14871_;
  wire _14872_;
  wire _14873_;
  wire _14874_;
  wire _14875_;
  wire _14876_;
  wire _14877_;
  wire _14878_;
  wire _14879_;
  wire _14880_;
  wire _14881_;
  wire _14882_;
  wire _14883_;
  wire _14884_;
  wire _14885_;
  wire _14886_;
  wire _14887_;
  wire _14888_;
  wire _14889_;
  wire _14890_;
  wire _14891_;
  wire _14892_;
  wire _14893_;
  wire _14894_;
  wire _14895_;
  wire _14896_;
  wire _14897_;
  wire _14898_;
  wire _14899_;
  wire _14900_;
  wire _14901_;
  wire _14902_;
  wire _14903_;
  wire _14904_;
  wire _14905_;
  wire _14906_;
  wire _14907_;
  wire _14908_;
  wire _14909_;
  wire _14910_;
  wire _14911_;
  wire _14912_;
  wire _14913_;
  wire _14914_;
  wire _14915_;
  wire _14916_;
  wire _14917_;
  wire _14918_;
  wire _14919_;
  wire _14920_;
  wire _14921_;
  wire _14922_;
  wire _14923_;
  wire _14924_;
  wire _14925_;
  wire _14926_;
  wire _14927_;
  wire _14928_;
  wire _14929_;
  wire _14930_;
  wire _14931_;
  wire _14932_;
  wire _14933_;
  wire _14934_;
  wire _14935_;
  wire _14936_;
  wire _14937_;
  wire _14938_;
  wire _14939_;
  wire _14940_;
  wire _14941_;
  wire _14942_;
  wire _14943_;
  wire _14944_;
  wire _14945_;
  wire _14946_;
  wire _14947_;
  wire _14948_;
  wire _14949_;
  wire _14950_;
  wire _14951_;
  wire _14952_;
  wire _14953_;
  wire _14954_;
  wire _14955_;
  wire _14956_;
  wire _14957_;
  wire _14958_;
  wire _14959_;
  wire _14960_;
  wire _14961_;
  wire _14962_;
  wire _14963_;
  wire _14964_;
  wire _14965_;
  wire _14966_;
  wire _14967_;
  wire _14968_;
  wire _14969_;
  wire _14970_;
  wire _14971_;
  wire _14972_;
  wire _14973_;
  wire _14974_;
  wire _14975_;
  wire _14976_;
  wire _14977_;
  wire _14978_;
  wire _14979_;
  wire _14980_;
  wire _14981_;
  wire _14982_;
  wire _14983_;
  wire _14984_;
  wire _14985_;
  wire _14986_;
  wire _14987_;
  wire _14988_;
  wire _14989_;
  wire _14990_;
  wire _14991_;
  wire _14992_;
  wire _14993_;
  wire _14994_;
  wire _14995_;
  wire _14996_;
  wire _14997_;
  wire _14998_;
  wire _14999_;
  wire _15000_;
  wire _15001_;
  wire _15002_;
  wire _15003_;
  wire _15004_;
  wire _15005_;
  wire _15006_;
  wire _15007_;
  wire _15008_;
  wire _15009_;
  wire _15010_;
  wire _15011_;
  wire _15012_;
  wire _15013_;
  wire _15014_;
  wire _15015_;
  wire _15016_;
  wire _15017_;
  wire _15018_;
  wire _15019_;
  wire _15020_;
  wire _15021_;
  wire _15022_;
  wire _15023_;
  wire _15024_;
  wire _15025_;
  wire _15026_;
  wire _15027_;
  wire _15028_;
  wire _15029_;
  wire _15030_;
  wire _15031_;
  wire _15032_;
  wire _15033_;
  wire _15034_;
  wire _15035_;
  wire _15036_;
  wire _15037_;
  wire _15038_;
  wire _15039_;
  wire _15040_;
  wire _15041_;
  wire _15042_;
  wire _15043_;
  wire _15044_;
  wire _15045_;
  wire _15046_;
  wire _15047_;
  wire _15048_;
  wire _15049_;
  wire _15050_;
  wire _15051_;
  wire _15052_;
  wire _15053_;
  wire _15054_;
  wire _15055_;
  wire _15056_;
  wire _15057_;
  wire _15058_;
  wire _15059_;
  wire _15060_;
  wire _15061_;
  wire _15062_;
  wire _15063_;
  wire _15064_;
  wire _15065_;
  wire _15066_;
  wire _15067_;
  wire _15068_;
  wire _15069_;
  wire _15070_;
  wire _15071_;
  wire _15072_;
  wire _15073_;
  wire _15074_;
  wire _15075_;
  wire _15076_;
  wire _15077_;
  wire _15078_;
  wire _15079_;
  wire _15080_;
  wire _15081_;
  wire _15082_;
  wire _15083_;
  wire _15084_;
  wire _15085_;
  wire _15086_;
  wire _15087_;
  wire _15088_;
  wire _15089_;
  wire _15090_;
  wire _15091_;
  wire _15092_;
  wire _15093_;
  wire _15094_;
  wire _15095_;
  wire _15096_;
  wire _15097_;
  wire _15098_;
  wire _15099_;
  wire _15100_;
  wire _15101_;
  wire _15102_;
  wire _15103_;
  wire _15104_;
  wire _15105_;
  wire _15106_;
  wire _15107_;
  wire _15108_;
  wire _15109_;
  wire _15110_;
  wire _15111_;
  wire _15112_;
  wire _15113_;
  wire _15114_;
  wire _15115_;
  wire _15116_;
  wire _15117_;
  wire _15118_;
  wire _15119_;
  wire _15120_;
  wire _15121_;
  wire _15122_;
  wire _15123_;
  wire _15124_;
  wire _15125_;
  wire _15126_;
  wire _15127_;
  wire _15128_;
  wire _15129_;
  wire _15130_;
  wire _15131_;
  wire _15132_;
  wire _15133_;
  wire _15134_;
  wire _15135_;
  wire _15136_;
  wire _15137_;
  wire _15138_;
  wire _15139_;
  wire _15140_;
  wire _15141_;
  wire _15142_;
  wire _15143_;
  wire _15144_;
  wire _15145_;
  wire _15146_;
  wire _15147_;
  wire _15148_;
  wire _15149_;
  wire _15150_;
  wire _15151_;
  wire _15152_;
  wire _15153_;
  wire _15154_;
  wire _15155_;
  wire _15156_;
  wire _15157_;
  wire _15158_;
  wire _15159_;
  wire _15160_;
  wire _15161_;
  wire _15162_;
  wire _15163_;
  wire _15164_;
  wire _15165_;
  wire _15166_;
  wire _15167_;
  wire _15168_;
  wire _15169_;
  wire _15170_;
  wire _15171_;
  wire _15172_;
  wire _15173_;
  wire _15174_;
  wire _15175_;
  wire _15176_;
  wire _15177_;
  wire _15178_;
  wire _15179_;
  wire _15180_;
  wire _15181_;
  wire _15182_;
  wire _15183_;
  wire _15184_;
  wire _15185_;
  wire _15186_;
  wire _15187_;
  wire _15188_;
  wire _15189_;
  wire _15190_;
  wire _15191_;
  wire _15192_;
  wire _15193_;
  wire _15194_;
  wire _15195_;
  wire _15196_;
  wire _15197_;
  wire _15198_;
  wire _15199_;
  wire _15200_;
  wire _15201_;
  wire _15202_;
  wire _15203_;
  wire _15204_;
  wire _15205_;
  wire _15206_;
  wire _15207_;
  wire _15208_;
  wire _15209_;
  wire _15210_;
  wire _15211_;
  wire _15212_;
  wire _15213_;
  wire _15214_;
  wire _15215_;
  wire _15216_;
  wire _15217_;
  wire _15218_;
  wire _15219_;
  wire _15220_;
  wire _15221_;
  wire _15222_;
  wire _15223_;
  wire _15224_;
  wire _15225_;
  wire _15226_;
  wire _15227_;
  wire _15228_;
  wire _15229_;
  wire _15230_;
  wire _15231_;
  wire _15232_;
  wire _15233_;
  wire _15234_;
  wire _15235_;
  wire _15236_;
  wire _15237_;
  wire _15238_;
  wire _15239_;
  wire _15240_;
  wire _15241_;
  wire _15242_;
  wire _15243_;
  wire _15244_;
  wire _15245_;
  wire _15246_;
  wire _15247_;
  wire _15248_;
  wire _15249_;
  wire _15250_;
  wire _15251_;
  wire _15252_;
  wire _15253_;
  wire _15254_;
  wire _15255_;
  wire _15256_;
  wire _15257_;
  wire _15258_;
  wire _15259_;
  wire _15260_;
  wire _15261_;
  wire _15262_;
  wire _15263_;
  wire _15264_;
  wire _15265_;
  wire _15266_;
  wire _15267_;
  wire _15268_;
  wire _15269_;
  wire _15270_;
  wire _15271_;
  wire _15272_;
  wire _15273_;
  wire _15274_;
  wire _15275_;
  wire _15276_;
  wire _15277_;
  wire _15278_;
  wire _15279_;
  wire _15280_;
  wire _15281_;
  wire _15282_;
  wire _15283_;
  wire _15284_;
  wire _15285_;
  wire _15286_;
  wire _15287_;
  wire _15288_;
  wire _15289_;
  wire _15290_;
  wire _15291_;
  wire _15292_;
  wire _15293_;
  wire _15294_;
  wire _15295_;
  wire _15296_;
  wire _15297_;
  wire _15298_;
  wire _15299_;
  wire _15300_;
  wire _15301_;
  wire _15302_;
  wire _15303_;
  wire _15304_;
  wire _15305_;
  wire _15306_;
  wire _15307_;
  wire _15308_;
  wire _15309_;
  wire _15310_;
  wire _15311_;
  wire _15312_;
  wire _15313_;
  wire _15314_;
  wire _15315_;
  wire _15316_;
  wire _15317_;
  wire _15318_;
  wire _15319_;
  wire _15320_;
  wire _15321_;
  wire _15322_;
  wire _15323_;
  wire _15324_;
  wire _15325_;
  wire _15326_;
  wire _15327_;
  wire _15328_;
  wire _15329_;
  wire _15330_;
  wire _15331_;
  wire _15332_;
  wire _15333_;
  wire _15334_;
  wire _15335_;
  wire _15336_;
  wire _15337_;
  wire _15338_;
  wire _15339_;
  wire _15340_;
  wire _15341_;
  wire _15342_;
  wire _15343_;
  wire _15344_;
  wire _15345_;
  wire _15346_;
  wire _15347_;
  wire _15348_;
  wire _15349_;
  wire _15350_;
  wire _15351_;
  wire _15352_;
  wire _15353_;
  wire _15354_;
  wire _15355_;
  wire _15356_;
  wire _15357_;
  wire _15358_;
  wire _15359_;
  wire _15360_;
  wire _15361_;
  wire _15362_;
  wire _15363_;
  wire _15364_;
  wire _15365_;
  wire _15366_;
  wire _15367_;
  wire _15368_;
  wire _15369_;
  wire _15370_;
  wire _15371_;
  wire _15372_;
  wire _15373_;
  wire _15374_;
  wire _15375_;
  wire _15376_;
  wire _15377_;
  wire _15378_;
  wire _15379_;
  wire _15380_;
  wire _15381_;
  wire _15382_;
  wire _15383_;
  wire _15384_;
  wire _15385_;
  wire _15386_;
  wire _15387_;
  wire _15388_;
  wire _15389_;
  wire _15390_;
  wire _15391_;
  wire _15392_;
  wire _15393_;
  wire _15394_;
  wire _15395_;
  wire _15396_;
  wire _15397_;
  wire _15398_;
  wire _15399_;
  wire _15400_;
  wire _15401_;
  wire _15402_;
  wire _15403_;
  wire _15404_;
  wire _15405_;
  wire _15406_;
  wire _15407_;
  wire _15408_;
  wire _15409_;
  wire _15410_;
  wire _15411_;
  wire _15412_;
  wire _15413_;
  wire _15414_;
  wire _15415_;
  wire _15416_;
  wire _15417_;
  wire _15418_;
  wire _15419_;
  wire _15420_;
  wire _15421_;
  wire _15422_;
  wire _15423_;
  wire _15424_;
  wire _15425_;
  wire _15426_;
  wire _15427_;
  wire _15428_;
  wire _15429_;
  wire _15430_;
  wire _15431_;
  wire _15432_;
  wire _15433_;
  wire _15434_;
  wire _15435_;
  wire _15436_;
  wire _15437_;
  wire _15438_;
  wire _15439_;
  wire _15440_;
  wire _15441_;
  wire _15442_;
  wire _15443_;
  wire _15444_;
  wire _15445_;
  wire _15446_;
  wire _15447_;
  wire _15448_;
  wire _15449_;
  wire _15450_;
  wire _15451_;
  wire _15452_;
  wire _15453_;
  wire _15454_;
  wire _15455_;
  wire _15456_;
  wire _15457_;
  wire _15458_;
  wire _15459_;
  wire _15460_;
  wire _15461_;
  wire _15462_;
  wire _15463_;
  wire _15464_;
  wire _15465_;
  wire _15466_;
  wire _15467_;
  wire _15468_;
  wire _15469_;
  wire _15470_;
  wire _15471_;
  wire _15472_;
  wire _15473_;
  wire _15474_;
  wire _15475_;
  wire _15476_;
  wire _15477_;
  wire _15478_;
  wire _15479_;
  wire _15480_;
  wire _15481_;
  wire _15482_;
  wire _15483_;
  wire _15484_;
  wire _15485_;
  wire _15486_;
  wire _15487_;
  wire _15488_;
  wire _15489_;
  wire _15490_;
  wire _15491_;
  wire _15492_;
  wire _15493_;
  wire _15494_;
  wire _15495_;
  wire _15496_;
  wire _15497_;
  wire _15498_;
  wire _15499_;
  wire _15500_;
  wire _15501_;
  wire _15502_;
  wire _15503_;
  wire _15504_;
  wire _15505_;
  wire _15506_;
  wire _15507_;
  wire _15508_;
  wire _15509_;
  wire _15510_;
  wire _15511_;
  wire _15512_;
  wire _15513_;
  wire _15514_;
  wire _15515_;
  wire _15516_;
  wire _15517_;
  wire _15518_;
  wire _15519_;
  wire _15520_;
  wire _15521_;
  wire _15522_;
  wire _15523_;
  wire _15524_;
  wire _15525_;
  wire _15526_;
  wire _15527_;
  wire _15528_;
  wire _15529_;
  wire _15530_;
  wire _15531_;
  wire _15532_;
  wire _15533_;
  wire _15534_;
  wire _15535_;
  wire _15536_;
  wire _15537_;
  wire _15538_;
  wire _15539_;
  wire _15540_;
  wire _15541_;
  wire _15542_;
  wire _15543_;
  wire _15544_;
  wire _15545_;
  wire _15546_;
  wire _15547_;
  wire _15548_;
  wire _15549_;
  wire _15550_;
  wire _15551_;
  wire _15552_;
  wire _15553_;
  wire _15554_;
  wire _15555_;
  wire _15556_;
  wire _15557_;
  wire _15558_;
  wire _15559_;
  wire _15560_;
  wire _15561_;
  wire _15562_;
  wire _15563_;
  wire _15564_;
  wire _15565_;
  wire _15566_;
  wire _15567_;
  wire _15568_;
  wire _15569_;
  wire _15570_;
  wire _15571_;
  wire _15572_;
  wire _15573_;
  wire _15574_;
  wire _15575_;
  wire _15576_;
  wire _15577_;
  wire _15578_;
  wire _15579_;
  wire _15580_;
  wire _15581_;
  wire _15582_;
  wire _15583_;
  wire _15584_;
  wire _15585_;
  wire _15586_;
  wire _15587_;
  wire _15588_;
  wire _15589_;
  wire _15590_;
  wire _15591_;
  wire _15592_;
  wire _15593_;
  wire _15594_;
  wire _15595_;
  wire _15596_;
  wire _15597_;
  wire _15598_;
  wire _15599_;
  wire _15600_;
  wire _15601_;
  wire _15602_;
  wire _15603_;
  wire _15604_;
  wire _15605_;
  wire _15606_;
  wire _15607_;
  wire _15608_;
  wire _15609_;
  wire _15610_;
  wire _15611_;
  wire _15612_;
  wire _15613_;
  wire _15614_;
  wire _15615_;
  wire _15616_;
  wire _15617_;
  wire _15618_;
  wire _15619_;
  wire _15620_;
  wire _15621_;
  wire _15622_;
  wire _15623_;
  wire _15624_;
  wire _15625_;
  wire _15626_;
  wire _15627_;
  wire _15628_;
  wire _15629_;
  wire _15630_;
  wire _15631_;
  wire _15632_;
  wire _15633_;
  wire _15634_;
  wire _15635_;
  wire _15636_;
  wire _15637_;
  wire _15638_;
  wire _15639_;
  wire _15640_;
  wire _15641_;
  wire _15642_;
  wire _15643_;
  wire _15644_;
  wire _15645_;
  wire _15646_;
  wire _15647_;
  wire _15648_;
  wire _15649_;
  wire _15650_;
  wire _15651_;
  wire _15652_;
  wire _15653_;
  wire _15654_;
  wire _15655_;
  wire _15656_;
  wire _15657_;
  wire _15658_;
  wire _15659_;
  wire _15660_;
  wire _15661_;
  wire _15662_;
  wire _15663_;
  wire _15664_;
  wire _15665_;
  wire _15666_;
  wire _15667_;
  wire _15668_;
  wire _15669_;
  wire _15670_;
  wire _15671_;
  wire _15672_;
  wire _15673_;
  wire _15674_;
  wire _15675_;
  wire _15676_;
  wire _15677_;
  wire _15678_;
  wire _15679_;
  wire _15680_;
  wire _15681_;
  wire _15682_;
  wire _15683_;
  wire _15684_;
  wire _15685_;
  wire _15686_;
  wire _15687_;
  wire _15688_;
  wire _15689_;
  wire _15690_;
  wire _15691_;
  wire _15692_;
  wire _15693_;
  wire _15694_;
  wire _15695_;
  wire _15696_;
  wire _15697_;
  wire _15698_;
  wire _15699_;
  wire _15700_;
  wire _15701_;
  wire _15702_;
  wire _15703_;
  wire _15704_;
  wire _15705_;
  wire _15706_;
  wire _15707_;
  wire _15708_;
  wire _15709_;
  wire _15710_;
  wire _15711_;
  wire _15712_;
  wire _15713_;
  wire _15714_;
  wire _15715_;
  wire _15716_;
  wire _15717_;
  wire _15718_;
  wire _15719_;
  wire _15720_;
  wire _15721_;
  wire _15722_;
  wire _15723_;
  wire _15724_;
  wire _15725_;
  wire _15726_;
  wire _15727_;
  wire _15728_;
  wire _15729_;
  wire _15730_;
  wire _15731_;
  wire _15732_;
  wire _15733_;
  wire _15734_;
  wire _15735_;
  wire _15736_;
  wire _15737_;
  wire _15738_;
  wire _15739_;
  wire _15740_;
  wire _15741_;
  wire _15742_;
  wire _15743_;
  wire _15744_;
  wire _15745_;
  wire _15746_;
  wire _15747_;
  wire _15748_;
  wire _15749_;
  wire _15750_;
  wire _15751_;
  wire _15752_;
  wire _15753_;
  wire _15754_;
  wire _15755_;
  wire _15756_;
  wire _15757_;
  wire _15758_;
  wire _15759_;
  wire _15760_;
  wire _15761_;
  wire _15762_;
  wire _15763_;
  wire _15764_;
  wire _15765_;
  wire _15766_;
  wire _15767_;
  wire _15768_;
  wire _15769_;
  wire _15770_;
  wire _15771_;
  wire _15772_;
  wire _15773_;
  wire _15774_;
  wire _15775_;
  wire _15776_;
  wire _15777_;
  wire _15778_;
  wire _15779_;
  wire _15780_;
  wire _15781_;
  wire _15782_;
  wire _15783_;
  wire _15784_;
  wire _15785_;
  wire _15786_;
  wire _15787_;
  wire _15788_;
  wire _15789_;
  wire _15790_;
  wire _15791_;
  wire _15792_;
  wire _15793_;
  wire _15794_;
  wire _15795_;
  wire _15796_;
  wire _15797_;
  wire _15798_;
  wire _15799_;
  wire _15800_;
  wire _15801_;
  wire _15802_;
  wire _15803_;
  wire _15804_;
  wire _15805_;
  wire _15806_;
  wire _15807_;
  wire _15808_;
  wire _15809_;
  wire _15810_;
  wire _15811_;
  wire _15812_;
  wire _15813_;
  wire _15814_;
  wire _15815_;
  wire _15816_;
  wire _15817_;
  wire _15818_;
  wire _15819_;
  wire _15820_;
  wire _15821_;
  wire _15822_;
  wire _15823_;
  wire _15824_;
  wire _15825_;
  wire _15826_;
  wire _15827_;
  wire _15828_;
  wire _15829_;
  wire _15830_;
  wire _15831_;
  wire _15832_;
  wire _15833_;
  wire _15834_;
  wire _15835_;
  wire _15836_;
  wire _15837_;
  wire _15838_;
  wire _15839_;
  wire _15840_;
  wire _15841_;
  wire _15842_;
  wire _15843_;
  wire _15844_;
  wire _15845_;
  wire _15846_;
  wire _15847_;
  wire _15848_;
  wire _15849_;
  wire _15850_;
  wire _15851_;
  wire _15852_;
  wire _15853_;
  wire _15854_;
  wire _15855_;
  wire _15856_;
  wire _15857_;
  wire _15858_;
  wire _15859_;
  wire _15860_;
  wire _15861_;
  wire _15862_;
  wire _15863_;
  wire _15864_;
  wire _15865_;
  wire _15866_;
  wire _15867_;
  wire _15868_;
  wire _15869_;
  wire _15870_;
  wire _15871_;
  wire _15872_;
  wire _15873_;
  wire _15874_;
  wire _15875_;
  wire _15876_;
  wire _15877_;
  wire _15878_;
  wire _15879_;
  wire _15880_;
  wire _15881_;
  wire _15882_;
  wire _15883_;
  wire _15884_;
  wire _15885_;
  wire _15886_;
  wire _15887_;
  wire _15888_;
  wire _15889_;
  wire _15890_;
  wire _15891_;
  wire _15892_;
  wire _15893_;
  wire _15894_;
  wire _15895_;
  wire _15896_;
  wire _15897_;
  wire _15898_;
  wire _15899_;
  wire _15900_;
  wire _15901_;
  wire _15902_;
  wire _15903_;
  wire _15904_;
  wire _15905_;
  wire _15906_;
  wire _15907_;
  wire _15908_;
  wire _15909_;
  wire _15910_;
  wire _15911_;
  wire _15912_;
  wire _15913_;
  wire _15914_;
  wire _15915_;
  wire _15916_;
  wire _15917_;
  wire _15918_;
  wire _15919_;
  wire _15920_;
  wire _15921_;
  wire _15922_;
  wire _15923_;
  wire _15924_;
  wire _15925_;
  wire _15926_;
  wire _15927_;
  wire _15928_;
  wire _15929_;
  wire _15930_;
  wire _15931_;
  wire _15932_;
  wire _15933_;
  wire _15934_;
  wire _15935_;
  wire _15936_;
  wire _15937_;
  wire _15938_;
  wire _15939_;
  wire _15940_;
  wire _15941_;
  wire _15942_;
  wire _15943_;
  wire _15944_;
  wire _15945_;
  wire _15946_;
  wire _15947_;
  wire _15948_;
  wire _15949_;
  wire _15950_;
  wire _15951_;
  wire _15952_;
  wire _15953_;
  wire _15954_;
  wire _15955_;
  wire _15956_;
  wire _15957_;
  wire _15958_;
  wire _15959_;
  wire _15960_;
  wire _15961_;
  wire _15962_;
  wire _15963_;
  wire _15964_;
  wire _15965_;
  wire _15966_;
  wire _15967_;
  wire _15968_;
  wire _15969_;
  wire _15970_;
  wire _15971_;
  wire _15972_;
  wire _15973_;
  wire _15974_;
  wire _15975_;
  wire _15976_;
  wire _15977_;
  wire _15978_;
  wire _15979_;
  wire _15980_;
  wire _15981_;
  wire _15982_;
  wire _15983_;
  wire _15984_;
  wire _15985_;
  wire _15986_;
  wire _15987_;
  wire _15988_;
  wire _15989_;
  wire _15990_;
  wire _15991_;
  wire _15992_;
  wire _15993_;
  wire _15994_;
  wire _15995_;
  wire _15996_;
  wire _15997_;
  wire _15998_;
  wire _15999_;
  wire _16000_;
  wire _16001_;
  wire _16002_;
  wire _16003_;
  wire _16004_;
  wire _16005_;
  wire _16006_;
  wire _16007_;
  wire _16008_;
  wire _16009_;
  wire _16010_;
  wire _16011_;
  wire _16012_;
  wire _16013_;
  wire _16014_;
  wire _16015_;
  wire _16016_;
  wire _16017_;
  wire _16018_;
  wire _16019_;
  wire _16020_;
  wire _16021_;
  wire _16022_;
  wire _16023_;
  wire _16024_;
  wire _16025_;
  wire _16026_;
  wire _16027_;
  wire _16028_;
  wire _16029_;
  wire _16030_;
  wire _16031_;
  wire _16032_;
  wire _16033_;
  wire _16034_;
  wire _16035_;
  wire _16036_;
  wire _16037_;
  wire _16038_;
  wire _16039_;
  wire _16040_;
  wire _16041_;
  wire _16042_;
  wire _16043_;
  wire _16044_;
  wire _16045_;
  wire _16046_;
  wire _16047_;
  wire _16048_;
  wire _16049_;
  wire _16050_;
  wire _16051_;
  wire _16052_;
  wire _16053_;
  wire _16054_;
  wire _16055_;
  wire _16056_;
  wire _16057_;
  wire _16058_;
  wire _16059_;
  wire _16060_;
  wire _16061_;
  wire _16062_;
  wire _16063_;
  wire _16064_;
  wire _16065_;
  wire _16066_;
  wire _16067_;
  wire _16068_;
  wire _16069_;
  wire _16070_;
  wire _16071_;
  wire _16072_;
  wire _16073_;
  wire _16074_;
  wire _16075_;
  wire _16076_;
  wire _16077_;
  wire _16078_;
  wire _16079_;
  wire _16080_;
  wire _16081_;
  wire _16082_;
  wire _16083_;
  wire _16084_;
  wire _16085_;
  wire _16086_;
  wire _16087_;
  wire _16088_;
  wire _16089_;
  wire _16090_;
  wire _16091_;
  wire _16092_;
  wire _16093_;
  wire _16094_;
  wire _16095_;
  wire _16096_;
  wire _16097_;
  wire _16098_;
  wire _16099_;
  wire _16100_;
  wire _16101_;
  wire _16102_;
  wire _16103_;
  wire _16104_;
  wire _16105_;
  wire _16106_;
  wire _16107_;
  wire _16108_;
  wire _16109_;
  wire _16110_;
  wire _16111_;
  wire _16112_;
  wire _16113_;
  wire _16114_;
  wire _16115_;
  wire _16116_;
  wire _16117_;
  wire _16118_;
  wire _16119_;
  wire _16120_;
  wire _16121_;
  wire _16122_;
  wire _16123_;
  wire _16124_;
  wire _16125_;
  wire _16126_;
  wire _16127_;
  wire _16128_;
  wire _16129_;
  wire _16130_;
  wire _16131_;
  wire _16132_;
  wire _16133_;
  wire _16134_;
  wire _16135_;
  wire _16136_;
  wire _16137_;
  wire _16138_;
  wire _16139_;
  wire _16140_;
  wire _16141_;
  wire _16142_;
  wire _16143_;
  wire _16144_;
  wire _16145_;
  wire _16146_;
  wire _16147_;
  wire _16148_;
  wire _16149_;
  wire _16150_;
  wire _16151_;
  wire _16152_;
  wire _16153_;
  wire _16154_;
  wire _16155_;
  wire _16156_;
  wire _16157_;
  wire _16158_;
  wire _16159_;
  wire _16160_;
  wire _16161_;
  wire _16162_;
  wire _16163_;
  wire _16164_;
  wire _16165_;
  wire _16166_;
  wire _16167_;
  wire _16168_;
  wire _16169_;
  wire _16170_;
  wire _16171_;
  wire _16172_;
  wire _16173_;
  wire _16174_;
  wire _16175_;
  wire _16176_;
  wire _16177_;
  wire _16178_;
  wire _16179_;
  wire _16180_;
  wire _16181_;
  wire _16182_;
  wire _16183_;
  wire _16184_;
  wire _16185_;
  wire _16186_;
  wire _16187_;
  wire _16188_;
  wire _16189_;
  wire _16190_;
  wire _16191_;
  wire _16192_;
  wire _16193_;
  wire _16194_;
  wire _16195_;
  wire _16196_;
  wire _16197_;
  wire _16198_;
  wire _16199_;
  wire _16200_;
  wire _16201_;
  wire _16202_;
  wire _16203_;
  wire _16204_;
  wire _16205_;
  wire _16206_;
  wire _16207_;
  wire _16208_;
  wire _16209_;
  wire _16210_;
  wire _16211_;
  wire _16212_;
  wire _16213_;
  wire _16214_;
  wire _16215_;
  wire _16216_;
  wire _16217_;
  wire _16218_;
  wire _16219_;
  wire _16220_;
  wire _16221_;
  wire _16222_;
  wire _16223_;
  wire _16224_;
  wire _16225_;
  wire _16226_;
  wire _16227_;
  wire _16228_;
  wire _16229_;
  wire _16230_;
  wire _16231_;
  wire _16232_;
  wire _16233_;
  wire _16234_;
  wire _16235_;
  wire _16236_;
  wire _16237_;
  wire _16238_;
  wire _16239_;
  wire _16240_;
  wire _16241_;
  wire _16242_;
  wire _16243_;
  wire _16244_;
  wire _16245_;
  wire _16246_;
  wire _16247_;
  wire _16248_;
  wire _16249_;
  wire _16250_;
  wire _16251_;
  wire _16252_;
  wire _16253_;
  wire _16254_;
  wire _16255_;
  wire _16256_;
  wire _16257_;
  wire _16258_;
  wire _16259_;
  wire _16260_;
  wire _16261_;
  wire _16262_;
  wire _16263_;
  wire _16264_;
  wire _16265_;
  wire _16266_;
  wire _16267_;
  wire _16268_;
  wire _16269_;
  wire _16270_;
  wire _16271_;
  wire _16272_;
  wire _16273_;
  wire _16274_;
  wire _16275_;
  wire _16276_;
  wire _16277_;
  wire _16278_;
  wire _16279_;
  wire _16280_;
  wire _16281_;
  wire _16282_;
  wire _16283_;
  wire _16284_;
  wire _16285_;
  wire _16286_;
  wire _16287_;
  wire _16288_;
  wire _16289_;
  wire _16290_;
  wire _16291_;
  wire _16292_;
  wire _16293_;
  wire _16294_;
  wire _16295_;
  wire _16296_;
  wire _16297_;
  wire _16298_;
  wire _16299_;
  wire _16300_;
  wire _16301_;
  wire _16302_;
  wire _16303_;
  wire _16304_;
  wire _16305_;
  wire _16306_;
  wire _16307_;
  wire _16308_;
  wire _16309_;
  wire _16310_;
  wire _16311_;
  wire _16312_;
  wire _16313_;
  wire _16314_;
  wire _16315_;
  wire _16316_;
  wire _16317_;
  wire _16318_;
  wire _16319_;
  wire _16320_;
  wire _16321_;
  wire _16322_;
  wire _16323_;
  wire _16324_;
  wire _16325_;
  wire _16326_;
  wire _16327_;
  wire _16328_;
  wire _16329_;
  wire _16330_;
  wire _16331_;
  wire _16332_;
  wire _16333_;
  wire _16334_;
  wire _16335_;
  wire _16336_;
  wire _16337_;
  wire _16338_;
  wire _16339_;
  wire _16340_;
  wire _16341_;
  wire _16342_;
  wire _16343_;
  wire _16344_;
  wire _16345_;
  wire _16346_;
  wire _16347_;
  wire _16348_;
  wire _16349_;
  wire _16350_;
  wire _16351_;
  wire _16352_;
  wire _16353_;
  wire _16354_;
  wire _16355_;
  wire _16356_;
  wire _16357_;
  wire _16358_;
  wire _16359_;
  wire _16360_;
  wire _16361_;
  wire _16362_;
  wire _16363_;
  wire _16364_;
  wire _16365_;
  wire _16366_;
  wire _16367_;
  wire _16368_;
  wire _16369_;
  wire _16370_;
  wire _16371_;
  wire _16372_;
  wire _16373_;
  wire _16374_;
  wire _16375_;
  wire _16376_;
  wire _16377_;
  wire _16378_;
  wire _16379_;
  wire _16380_;
  wire _16381_;
  wire _16382_;
  wire _16383_;
  wire _16384_;
  wire _16385_;
  wire _16386_;
  wire _16387_;
  wire _16388_;
  wire _16389_;
  wire _16390_;
  wire _16391_;
  wire _16392_;
  wire _16393_;
  wire _16394_;
  wire _16395_;
  wire _16396_;
  wire _16397_;
  wire _16398_;
  wire _16399_;
  wire _16400_;
  wire _16401_;
  wire _16402_;
  wire _16403_;
  wire _16404_;
  wire _16405_;
  wire _16406_;
  wire _16407_;
  wire _16408_;
  wire _16409_;
  wire _16410_;
  wire _16411_;
  wire _16412_;
  wire _16413_;
  wire _16414_;
  wire _16415_;
  wire _16416_;
  wire _16417_;
  wire _16418_;
  wire _16419_;
  wire _16420_;
  wire _16421_;
  wire _16422_;
  wire _16423_;
  wire _16424_;
  wire _16425_;
  wire _16426_;
  wire _16427_;
  wire _16428_;
  wire _16429_;
  wire _16430_;
  wire _16431_;
  wire _16432_;
  wire _16433_;
  wire _16434_;
  wire _16435_;
  wire _16436_;
  wire _16437_;
  wire _16438_;
  wire _16439_;
  wire _16440_;
  wire _16441_;
  wire _16442_;
  wire _16443_;
  wire _16444_;
  wire _16445_;
  wire _16446_;
  wire _16447_;
  wire _16448_;
  wire _16449_;
  wire _16450_;
  wire _16451_;
  wire _16452_;
  wire _16453_;
  wire _16454_;
  wire _16455_;
  wire _16456_;
  wire _16457_;
  wire _16458_;
  wire _16459_;
  wire _16460_;
  wire _16461_;
  wire _16462_;
  wire _16463_;
  wire _16464_;
  wire _16465_;
  wire _16466_;
  wire _16467_;
  wire _16468_;
  wire _16469_;
  wire _16470_;
  wire _16471_;
  wire _16472_;
  wire _16473_;
  wire _16474_;
  wire _16475_;
  wire _16476_;
  wire _16477_;
  wire _16478_;
  wire _16479_;
  wire _16480_;
  wire _16481_;
  wire _16482_;
  wire _16483_;
  wire _16484_;
  wire _16485_;
  wire _16486_;
  wire _16487_;
  wire _16488_;
  wire _16489_;
  wire _16490_;
  wire _16491_;
  wire _16492_;
  wire _16493_;
  wire _16494_;
  wire _16495_;
  wire _16496_;
  wire _16497_;
  wire _16498_;
  wire _16499_;
  wire _16500_;
  wire _16501_;
  wire _16502_;
  wire _16503_;
  wire _16504_;
  wire _16505_;
  wire _16506_;
  wire _16507_;
  wire _16508_;
  wire _16509_;
  wire _16510_;
  wire _16511_;
  wire _16512_;
  wire _16513_;
  wire _16514_;
  wire _16515_;
  wire _16516_;
  wire _16517_;
  wire _16518_;
  wire _16519_;
  wire _16520_;
  wire _16521_;
  wire _16522_;
  wire _16523_;
  wire _16524_;
  wire _16525_;
  wire _16526_;
  wire _16527_;
  wire _16528_;
  wire _16529_;
  wire _16530_;
  wire _16531_;
  wire _16532_;
  wire _16533_;
  wire _16534_;
  wire _16535_;
  wire _16536_;
  wire _16537_;
  wire _16538_;
  wire _16539_;
  wire _16540_;
  wire _16541_;
  wire _16542_;
  wire _16543_;
  wire _16544_;
  wire _16545_;
  wire _16546_;
  wire _16547_;
  wire _16548_;
  wire _16549_;
  wire _16550_;
  wire _16551_;
  wire _16552_;
  wire _16553_;
  wire _16554_;
  wire _16555_;
  wire _16556_;
  wire _16557_;
  wire _16558_;
  wire _16559_;
  wire _16560_;
  wire _16561_;
  wire _16562_;
  wire _16563_;
  wire _16564_;
  wire _16565_;
  wire _16566_;
  wire _16567_;
  wire _16568_;
  wire _16569_;
  wire _16570_;
  wire _16571_;
  wire _16572_;
  wire _16573_;
  wire _16574_;
  wire _16575_;
  wire _16576_;
  wire _16577_;
  wire _16578_;
  wire _16579_;
  wire _16580_;
  wire _16581_;
  wire _16582_;
  wire _16583_;
  wire _16584_;
  wire _16585_;
  wire _16586_;
  wire _16587_;
  wire _16588_;
  wire _16589_;
  wire _16590_;
  wire _16591_;
  wire _16592_;
  wire _16593_;
  wire _16594_;
  wire _16595_;
  wire _16596_;
  wire _16597_;
  wire _16598_;
  wire _16599_;
  wire _16600_;
  wire _16601_;
  wire _16602_;
  wire _16603_;
  wire _16604_;
  wire _16605_;
  wire _16606_;
  wire _16607_;
  wire _16608_;
  wire _16609_;
  wire _16610_;
  wire _16611_;
  wire _16612_;
  wire _16613_;
  wire _16614_;
  wire _16615_;
  wire _16616_;
  wire _16617_;
  wire _16618_;
  wire _16619_;
  wire _16620_;
  wire _16621_;
  wire _16622_;
  wire _16623_;
  wire _16624_;
  wire _16625_;
  wire _16626_;
  wire _16627_;
  wire _16628_;
  wire _16629_;
  wire _16630_;
  wire _16631_;
  wire _16632_;
  wire _16633_;
  wire _16634_;
  wire _16635_;
  wire _16636_;
  wire _16637_;
  wire _16638_;
  wire _16639_;
  wire _16640_;
  wire _16641_;
  wire _16642_;
  wire _16643_;
  wire _16644_;
  wire _16645_;
  wire _16646_;
  wire _16647_;
  wire _16648_;
  wire _16649_;
  wire _16650_;
  wire _16651_;
  wire _16652_;
  wire _16653_;
  wire _16654_;
  wire _16655_;
  wire _16656_;
  wire _16657_;
  wire _16658_;
  wire _16659_;
  wire _16660_;
  wire _16661_;
  wire _16662_;
  wire _16663_;
  wire _16664_;
  wire _16665_;
  wire _16666_;
  wire _16667_;
  wire _16668_;
  wire _16669_;
  wire _16670_;
  wire _16671_;
  wire _16672_;
  wire _16673_;
  wire _16674_;
  wire _16675_;
  wire _16676_;
  wire _16677_;
  wire _16678_;
  wire _16679_;
  wire _16680_;
  wire _16681_;
  wire _16682_;
  wire _16683_;
  wire _16684_;
  wire _16685_;
  wire _16686_;
  wire _16687_;
  wire _16688_;
  wire _16689_;
  wire _16690_;
  wire _16691_;
  wire _16692_;
  wire _16693_;
  wire _16694_;
  wire _16695_;
  wire _16696_;
  wire _16697_;
  wire _16698_;
  wire _16699_;
  wire _16700_;
  wire _16701_;
  wire _16702_;
  wire _16703_;
  wire _16704_;
  wire _16705_;
  wire _16706_;
  wire _16707_;
  wire _16708_;
  wire _16709_;
  wire _16710_;
  wire _16711_;
  wire _16712_;
  wire _16713_;
  wire _16714_;
  wire _16715_;
  wire _16716_;
  wire _16717_;
  wire _16718_;
  wire _16719_;
  wire _16720_;
  wire _16721_;
  wire _16722_;
  wire _16723_;
  wire _16724_;
  wire _16725_;
  wire _16726_;
  wire _16727_;
  wire _16728_;
  wire _16729_;
  wire _16730_;
  wire _16731_;
  wire _16732_;
  wire _16733_;
  wire _16734_;
  wire _16735_;
  wire _16736_;
  wire _16737_;
  wire _16738_;
  wire _16739_;
  wire _16740_;
  wire _16741_;
  wire _16742_;
  wire _16743_;
  wire _16744_;
  wire _16745_;
  wire _16746_;
  wire _16747_;
  wire _16748_;
  wire _16749_;
  wire _16750_;
  wire _16751_;
  wire _16752_;
  wire _16753_;
  wire _16754_;
  wire _16755_;
  wire _16756_;
  wire _16757_;
  wire _16758_;
  wire _16759_;
  wire _16760_;
  wire _16761_;
  wire _16762_;
  wire _16763_;
  wire _16764_;
  wire _16765_;
  wire _16766_;
  wire _16767_;
  wire _16768_;
  wire _16769_;
  wire _16770_;
  wire _16771_;
  wire _16772_;
  wire _16773_;
  wire _16774_;
  wire _16775_;
  wire _16776_;
  wire _16777_;
  wire _16778_;
  wire _16779_;
  wire _16780_;
  wire _16781_;
  wire _16782_;
  wire _16783_;
  wire _16784_;
  wire _16785_;
  wire _16786_;
  wire _16787_;
  wire _16788_;
  wire _16789_;
  wire _16790_;
  wire _16791_;
  wire _16792_;
  wire _16793_;
  wire _16794_;
  wire _16795_;
  wire _16796_;
  wire _16797_;
  wire _16798_;
  wire _16799_;
  wire _16800_;
  wire _16801_;
  wire _16802_;
  wire _16803_;
  wire _16804_;
  wire _16805_;
  wire _16806_;
  wire _16807_;
  wire _16808_;
  wire _16809_;
  wire _16810_;
  wire _16811_;
  wire _16812_;
  wire _16813_;
  wire _16814_;
  wire _16815_;
  wire _16816_;
  wire _16817_;
  wire _16818_;
  wire _16819_;
  wire _16820_;
  wire _16821_;
  wire _16822_;
  wire _16823_;
  wire _16824_;
  wire _16825_;
  wire _16826_;
  wire _16827_;
  wire _16828_;
  wire _16829_;
  wire _16830_;
  wire _16831_;
  wire _16832_;
  wire _16833_;
  wire _16834_;
  wire _16835_;
  wire _16836_;
  wire _16837_;
  wire _16838_;
  wire _16839_;
  wire _16840_;
  wire _16841_;
  wire _16842_;
  wire _16843_;
  wire _16844_;
  wire _16845_;
  wire _16846_;
  wire _16847_;
  wire _16848_;
  wire _16849_;
  wire _16850_;
  wire _16851_;
  wire _16852_;
  wire _16853_;
  wire _16854_;
  wire _16855_;
  wire _16856_;
  wire _16857_;
  wire _16858_;
  wire _16859_;
  wire _16860_;
  wire _16861_;
  wire _16862_;
  wire _16863_;
  wire _16864_;
  wire _16865_;
  wire _16866_;
  wire _16867_;
  wire _16868_;
  wire _16869_;
  wire _16870_;
  wire _16871_;
  wire _16872_;
  wire _16873_;
  wire _16874_;
  wire _16875_;
  wire _16876_;
  wire _16877_;
  wire _16878_;
  wire _16879_;
  wire _16880_;
  wire _16881_;
  wire _16882_;
  wire _16883_;
  wire _16884_;
  wire _16885_;
  wire _16886_;
  wire _16887_;
  wire _16888_;
  wire _16889_;
  wire _16890_;
  wire _16891_;
  wire _16892_;
  wire _16893_;
  wire _16894_;
  wire _16895_;
  wire _16896_;
  wire _16897_;
  wire _16898_;
  wire _16899_;
  wire _16900_;
  wire _16901_;
  wire _16902_;
  wire _16903_;
  wire _16904_;
  wire _16905_;
  wire _16906_;
  wire _16907_;
  wire _16908_;
  wire _16909_;
  wire _16910_;
  wire _16911_;
  wire _16912_;
  wire _16913_;
  wire _16914_;
  wire _16915_;
  wire _16916_;
  wire _16917_;
  wire _16918_;
  wire _16919_;
  wire _16920_;
  wire _16921_;
  wire _16922_;
  wire _16923_;
  wire _16924_;
  wire _16925_;
  wire _16926_;
  wire _16927_;
  wire _16928_;
  wire _16929_;
  wire _16930_;
  wire _16931_;
  wire _16932_;
  wire _16933_;
  wire _16934_;
  wire _16935_;
  wire _16936_;
  wire _16937_;
  wire _16938_;
  wire _16939_;
  wire _16940_;
  wire _16941_;
  wire _16942_;
  wire _16943_;
  wire _16944_;
  wire _16945_;
  wire _16946_;
  wire _16947_;
  wire _16948_;
  wire _16949_;
  wire _16950_;
  wire _16951_;
  wire _16952_;
  wire _16953_;
  wire _16954_;
  wire _16955_;
  wire _16956_;
  wire _16957_;
  wire _16958_;
  wire _16959_;
  wire _16960_;
  wire _16961_;
  wire _16962_;
  wire _16963_;
  wire _16964_;
  wire _16965_;
  wire _16966_;
  wire _16967_;
  wire _16968_;
  wire _16969_;
  wire _16970_;
  wire _16971_;
  wire _16972_;
  wire _16973_;
  wire _16974_;
  wire _16975_;
  wire _16976_;
  wire _16977_;
  wire _16978_;
  wire _16979_;
  wire _16980_;
  wire _16981_;
  wire _16982_;
  wire _16983_;
  wire _16984_;
  wire _16985_;
  wire _16986_;
  wire _16987_;
  wire _16988_;
  wire _16989_;
  wire _16990_;
  wire _16991_;
  wire _16992_;
  wire _16993_;
  wire _16994_;
  wire _16995_;
  wire _16996_;
  wire _16997_;
  wire _16998_;
  wire _16999_;
  wire _17000_;
  wire _17001_;
  wire _17002_;
  wire _17003_;
  wire _17004_;
  wire _17005_;
  wire _17006_;
  wire _17007_;
  wire _17008_;
  wire _17009_;
  wire _17010_;
  wire _17011_;
  wire _17012_;
  wire _17013_;
  wire _17014_;
  wire _17015_;
  wire _17016_;
  wire _17017_;
  wire _17018_;
  wire _17019_;
  wire _17020_;
  wire _17021_;
  wire _17022_;
  wire _17023_;
  wire _17024_;
  wire _17025_;
  wire _17026_;
  wire _17027_;
  wire _17028_;
  wire _17029_;
  wire _17030_;
  wire _17031_;
  wire _17032_;
  wire _17033_;
  wire _17034_;
  wire _17035_;
  wire _17036_;
  wire _17037_;
  wire _17038_;
  wire _17039_;
  wire _17040_;
  wire _17041_;
  wire _17042_;
  wire _17043_;
  wire _17044_;
  wire _17045_;
  wire _17046_;
  wire _17047_;
  wire _17048_;
  wire _17049_;
  wire _17050_;
  wire _17051_;
  wire _17052_;
  wire _17053_;
  wire _17054_;
  wire _17055_;
  wire _17056_;
  wire _17057_;
  wire _17058_;
  wire _17059_;
  wire _17060_;
  wire _17061_;
  wire _17062_;
  wire _17063_;
  wire _17064_;
  wire _17065_;
  wire _17066_;
  wire _17067_;
  wire _17068_;
  wire _17069_;
  wire _17070_;
  wire _17071_;
  wire _17072_;
  wire _17073_;
  wire _17074_;
  wire _17075_;
  wire _17076_;
  wire _17077_;
  wire _17078_;
  wire _17079_;
  wire _17080_;
  wire _17081_;
  wire _17082_;
  wire _17083_;
  wire _17084_;
  wire _17085_;
  wire _17086_;
  wire _17087_;
  wire _17088_;
  wire _17089_;
  wire _17090_;
  wire _17091_;
  wire _17092_;
  wire _17093_;
  wire _17094_;
  wire _17095_;
  wire _17096_;
  wire _17097_;
  wire _17098_;
  wire _17099_;
  wire _17100_;
  wire _17101_;
  wire _17102_;
  wire _17103_;
  wire _17104_;
  wire _17105_;
  wire _17106_;
  wire _17107_;
  wire _17108_;
  wire _17109_;
  wire _17110_;
  wire _17111_;
  wire _17112_;
  wire _17113_;
  wire _17114_;
  wire _17115_;
  wire _17116_;
  wire _17117_;
  wire _17118_;
  wire _17119_;
  wire _17120_;
  wire _17121_;
  wire _17122_;
  wire _17123_;
  wire _17124_;
  wire _17125_;
  wire _17126_;
  wire _17127_;
  wire _17128_;
  wire _17129_;
  wire _17130_;
  wire _17131_;
  wire _17132_;
  wire _17133_;
  wire _17134_;
  wire _17135_;
  wire _17136_;
  wire _17137_;
  wire _17138_;
  wire _17139_;
  wire _17140_;
  wire _17141_;
  wire _17142_;
  wire _17143_;
  wire _17144_;
  wire _17145_;
  wire _17146_;
  wire _17147_;
  wire _17148_;
  wire _17149_;
  wire _17150_;
  wire _17151_;
  wire _17152_;
  wire _17153_;
  wire _17154_;
  wire _17155_;
  wire _17156_;
  wire _17157_;
  wire _17158_;
  wire _17159_;
  wire _17160_;
  wire _17161_;
  wire _17162_;
  wire _17163_;
  wire _17164_;
  wire _17165_;
  wire _17166_;
  wire _17167_;
  wire _17168_;
  wire _17169_;
  wire _17170_;
  wire _17171_;
  wire _17172_;
  wire _17173_;
  wire _17174_;
  wire _17175_;
  wire _17176_;
  wire _17177_;
  wire _17178_;
  wire _17179_;
  wire _17180_;
  wire _17181_;
  wire _17182_;
  wire _17183_;
  wire _17184_;
  wire _17185_;
  wire _17186_;
  wire _17187_;
  wire _17188_;
  wire _17189_;
  wire _17190_;
  wire _17191_;
  wire _17192_;
  wire _17193_;
  wire _17194_;
  wire _17195_;
  wire _17196_;
  wire _17197_;
  wire _17198_;
  wire _17199_;
  wire _17200_;
  wire _17201_;
  wire _17202_;
  wire _17203_;
  wire _17204_;
  wire _17205_;
  wire _17206_;
  wire _17207_;
  wire _17208_;
  wire _17209_;
  wire _17210_;
  wire _17211_;
  wire _17212_;
  wire _17213_;
  wire _17214_;
  wire _17215_;
  wire _17216_;
  wire _17217_;
  wire _17218_;
  wire _17219_;
  wire _17220_;
  wire _17221_;
  wire _17222_;
  wire _17223_;
  wire _17224_;
  wire _17225_;
  wire _17226_;
  wire _17227_;
  wire _17228_;
  wire _17229_;
  wire _17230_;
  wire _17231_;
  wire _17232_;
  wire _17233_;
  wire _17234_;
  wire _17235_;
  wire _17236_;
  wire _17237_;
  wire _17238_;
  wire _17239_;
  wire _17240_;
  wire _17241_;
  wire _17242_;
  wire _17243_;
  wire _17244_;
  wire _17245_;
  wire _17246_;
  wire _17247_;
  wire _17248_;
  wire _17249_;
  wire _17250_;
  wire _17251_;
  wire _17252_;
  wire _17253_;
  wire _17254_;
  wire _17255_;
  wire _17256_;
  wire _17257_;
  wire _17258_;
  wire _17259_;
  wire _17260_;
  wire _17261_;
  wire _17262_;
  wire _17263_;
  wire _17264_;
  wire _17265_;
  wire _17266_;
  wire _17267_;
  wire _17268_;
  wire _17269_;
  wire _17270_;
  wire _17271_;
  wire _17272_;
  wire _17273_;
  wire _17274_;
  wire _17275_;
  wire _17276_;
  wire _17277_;
  wire _17278_;
  wire _17279_;
  wire _17280_;
  wire _17281_;
  wire _17282_;
  wire _17283_;
  wire _17284_;
  wire _17285_;
  wire _17286_;
  wire _17287_;
  wire _17288_;
  wire _17289_;
  wire _17290_;
  wire _17291_;
  wire _17292_;
  wire _17293_;
  wire _17294_;
  wire _17295_;
  wire _17296_;
  wire _17297_;
  wire _17298_;
  wire _17299_;
  wire _17300_;
  wire _17301_;
  wire _17302_;
  wire _17303_;
  wire _17304_;
  wire _17305_;
  wire _17306_;
  wire _17307_;
  wire _17308_;
  wire _17309_;
  wire _17310_;
  wire _17311_;
  wire _17312_;
  wire _17313_;
  wire _17314_;
  wire _17315_;
  wire _17316_;
  wire _17317_;
  wire _17318_;
  wire _17319_;
  wire _17320_;
  wire _17321_;
  wire _17322_;
  wire _17323_;
  wire _17324_;
  wire _17325_;
  wire _17326_;
  wire _17327_;
  wire _17328_;
  wire _17329_;
  wire _17330_;
  wire _17331_;
  wire _17332_;
  wire _17333_;
  wire _17334_;
  wire _17335_;
  wire _17336_;
  wire _17337_;
  wire _17338_;
  wire _17339_;
  wire _17340_;
  wire _17341_;
  wire _17342_;
  wire _17343_;
  wire _17344_;
  wire _17345_;
  wire _17346_;
  wire _17347_;
  wire _17348_;
  wire _17349_;
  wire _17350_;
  wire _17351_;
  wire _17352_;
  wire _17353_;
  wire _17354_;
  wire _17355_;
  wire _17356_;
  wire _17357_;
  wire _17358_;
  wire _17359_;
  wire _17360_;
  wire _17361_;
  wire _17362_;
  wire _17363_;
  wire _17364_;
  wire _17365_;
  wire _17366_;
  wire _17367_;
  wire _17368_;
  wire _17369_;
  wire _17370_;
  wire _17371_;
  wire _17372_;
  wire _17373_;
  wire _17374_;
  wire _17375_;
  wire _17376_;
  wire _17377_;
  wire _17378_;
  wire _17379_;
  wire _17380_;
  wire _17381_;
  wire _17382_;
  wire _17383_;
  wire _17384_;
  wire _17385_;
  wire _17386_;
  wire _17387_;
  wire _17388_;
  wire _17389_;
  wire _17390_;
  wire _17391_;
  wire _17392_;
  wire _17393_;
  wire _17394_;
  wire _17395_;
  wire _17396_;
  wire _17397_;
  wire _17398_;
  wire _17399_;
  wire _17400_;
  wire _17401_;
  wire _17402_;
  wire _17403_;
  wire _17404_;
  wire _17405_;
  wire _17406_;
  wire _17407_;
  wire _17408_;
  wire _17409_;
  wire _17410_;
  wire _17411_;
  wire _17412_;
  wire _17413_;
  wire _17414_;
  wire _17415_;
  wire _17416_;
  wire _17417_;
  wire _17418_;
  wire _17419_;
  wire _17420_;
  wire _17421_;
  wire _17422_;
  wire _17423_;
  wire _17424_;
  wire _17425_;
  wire _17426_;
  wire _17427_;
  wire _17428_;
  wire _17429_;
  wire _17430_;
  wire _17431_;
  wire _17432_;
  wire _17433_;
  wire _17434_;
  wire _17435_;
  wire _17436_;
  wire _17437_;
  wire _17438_;
  wire _17439_;
  wire _17440_;
  wire _17441_;
  wire _17442_;
  wire _17443_;
  wire _17444_;
  wire _17445_;
  wire _17446_;
  wire _17447_;
  wire _17448_;
  wire _17449_;
  wire _17450_;
  wire _17451_;
  wire _17452_;
  wire _17453_;
  wire _17454_;
  wire _17455_;
  wire _17456_;
  wire _17457_;
  wire _17458_;
  wire _17459_;
  wire _17460_;
  wire _17461_;
  wire _17462_;
  wire _17463_;
  wire _17464_;
  wire _17465_;
  wire _17466_;
  wire _17467_;
  wire _17468_;
  wire _17469_;
  wire _17470_;
  wire _17471_;
  wire _17472_;
  wire _17473_;
  wire _17474_;
  wire _17475_;
  wire _17476_;
  wire _17477_;
  wire _17478_;
  wire _17479_;
  wire _17480_;
  wire _17481_;
  wire _17482_;
  wire _17483_;
  wire _17484_;
  wire _17485_;
  wire _17486_;
  wire _17487_;
  wire _17488_;
  wire _17489_;
  wire _17490_;
  wire _17491_;
  wire _17492_;
  wire _17493_;
  wire _17494_;
  wire _17495_;
  wire _17496_;
  wire _17497_;
  wire _17498_;
  wire _17499_;
  wire _17500_;
  wire _17501_;
  wire _17502_;
  wire _17503_;
  wire _17504_;
  wire _17505_;
  wire _17506_;
  wire _17507_;
  wire _17508_;
  wire _17509_;
  wire _17510_;
  wire _17511_;
  wire _17512_;
  wire _17513_;
  wire _17514_;
  wire _17515_;
  wire _17516_;
  wire _17517_;
  wire _17518_;
  wire _17519_;
  wire _17520_;
  wire _17521_;
  wire _17522_;
  wire _17523_;
  wire _17524_;
  wire _17525_;
  wire _17526_;
  wire _17527_;
  wire _17528_;
  wire _17529_;
  wire _17530_;
  wire _17531_;
  wire _17532_;
  wire _17533_;
  wire _17534_;
  wire _17535_;
  wire _17536_;
  wire _17537_;
  wire _17538_;
  wire _17539_;
  wire _17540_;
  wire _17541_;
  wire _17542_;
  wire _17543_;
  wire _17544_;
  wire _17545_;
  wire _17546_;
  wire _17547_;
  wire _17548_;
  wire _17549_;
  wire _17550_;
  wire _17551_;
  wire _17552_;
  wire _17553_;
  wire _17554_;
  wire _17555_;
  wire _17556_;
  wire _17557_;
  wire _17558_;
  wire _17559_;
  wire _17560_;
  wire _17561_;
  wire _17562_;
  wire _17563_;
  wire _17564_;
  wire _17565_;
  wire _17566_;
  wire _17567_;
  wire _17568_;
  wire _17569_;
  wire _17570_;
  wire _17571_;
  wire _17572_;
  wire _17573_;
  wire _17574_;
  wire _17575_;
  wire _17576_;
  wire _17577_;
  wire _17578_;
  wire _17579_;
  wire _17580_;
  wire _17581_;
  wire _17582_;
  wire _17583_;
  wire _17584_;
  wire _17585_;
  wire _17586_;
  wire _17587_;
  wire _17588_;
  wire _17589_;
  wire _17590_;
  wire _17591_;
  wire _17592_;
  wire _17593_;
  wire _17594_;
  wire _17595_;
  wire _17596_;
  wire _17597_;
  wire _17598_;
  wire _17599_;
  wire _17600_;
  wire _17601_;
  wire _17602_;
  wire _17603_;
  wire _17604_;
  wire _17605_;
  wire _17606_;
  wire _17607_;
  wire _17608_;
  wire _17609_;
  wire _17610_;
  wire _17611_;
  wire _17612_;
  wire _17613_;
  wire _17614_;
  wire _17615_;
  wire _17616_;
  wire _17617_;
  wire _17618_;
  wire _17619_;
  wire _17620_;
  wire _17621_;
  wire _17622_;
  wire _17623_;
  wire _17624_;
  wire _17625_;
  wire _17626_;
  wire _17627_;
  wire _17628_;
  wire _17629_;
  wire _17630_;
  wire _17631_;
  wire _17632_;
  wire _17633_;
  wire _17634_;
  wire _17635_;
  wire _17636_;
  wire _17637_;
  wire _17638_;
  wire _17639_;
  wire _17640_;
  wire _17641_;
  wire _17642_;
  wire _17643_;
  wire _17644_;
  wire _17645_;
  wire _17646_;
  wire _17647_;
  wire _17648_;
  wire _17649_;
  wire _17650_;
  wire _17651_;
  wire _17652_;
  wire _17653_;
  wire _17654_;
  wire _17655_;
  wire _17656_;
  wire _17657_;
  wire _17658_;
  wire _17659_;
  wire _17660_;
  wire _17661_;
  wire _17662_;
  wire _17663_;
  wire _17664_;
  wire _17665_;
  wire _17666_;
  wire _17667_;
  wire _17668_;
  wire _17669_;
  wire _17670_;
  wire _17671_;
  wire _17672_;
  wire _17673_;
  wire _17674_;
  wire _17675_;
  wire _17676_;
  wire _17677_;
  wire _17678_;
  wire _17679_;
  wire _17680_;
  wire _17681_;
  wire _17682_;
  wire _17683_;
  wire _17684_;
  wire _17685_;
  wire _17686_;
  wire _17687_;
  wire _17688_;
  wire _17689_;
  wire _17690_;
  wire _17691_;
  wire _17692_;
  wire _17693_;
  wire _17694_;
  wire _17695_;
  wire _17696_;
  wire _17697_;
  wire _17698_;
  wire _17699_;
  wire _17700_;
  wire _17701_;
  wire _17702_;
  wire _17703_;
  wire _17704_;
  wire _17705_;
  wire _17706_;
  wire _17707_;
  wire _17708_;
  wire _17709_;
  wire _17710_;
  wire _17711_;
  wire _17712_;
  wire _17713_;
  wire _17714_;
  wire _17715_;
  wire _17716_;
  wire _17717_;
  wire _17718_;
  wire _17719_;
  wire _17720_;
  wire _17721_;
  wire _17722_;
  wire _17723_;
  wire _17724_;
  wire _17725_;
  wire _17726_;
  wire _17727_;
  wire _17728_;
  wire _17729_;
  wire _17730_;
  wire _17731_;
  wire _17732_;
  wire _17733_;
  wire _17734_;
  wire _17735_;
  wire _17736_;
  wire _17737_;
  wire _17738_;
  wire _17739_;
  wire _17740_;
  wire _17741_;
  wire _17742_;
  wire _17743_;
  wire _17744_;
  wire _17745_;
  wire _17746_;
  wire _17747_;
  wire _17748_;
  wire _17749_;
  wire _17750_;
  wire _17751_;
  wire _17752_;
  wire _17753_;
  wire _17754_;
  wire _17755_;
  wire _17756_;
  wire _17757_;
  wire _17758_;
  wire _17759_;
  wire _17760_;
  wire _17761_;
  wire _17762_;
  wire _17763_;
  wire _17764_;
  wire _17765_;
  wire _17766_;
  wire _17767_;
  wire _17768_;
  wire _17769_;
  wire _17770_;
  wire _17771_;
  wire _17772_;
  wire _17773_;
  wire _17774_;
  wire _17775_;
  wire _17776_;
  wire _17777_;
  wire _17778_;
  wire _17779_;
  wire _17780_;
  wire _17781_;
  wire _17782_;
  wire _17783_;
  wire _17784_;
  wire _17785_;
  wire _17786_;
  wire _17787_;
  wire _17788_;
  wire _17789_;
  wire _17790_;
  wire _17791_;
  wire _17792_;
  wire _17793_;
  wire _17794_;
  wire _17795_;
  wire _17796_;
  wire _17797_;
  wire _17798_;
  wire _17799_;
  wire _17800_;
  wire _17801_;
  wire _17802_;
  wire _17803_;
  wire _17804_;
  wire _17805_;
  wire _17806_;
  wire _17807_;
  wire _17808_;
  wire _17809_;
  wire _17810_;
  wire _17811_;
  wire _17812_;
  wire _17813_;
  wire _17814_;
  wire _17815_;
  wire _17816_;
  wire _17817_;
  wire _17818_;
  wire _17819_;
  wire _17820_;
  wire _17821_;
  wire _17822_;
  wire _17823_;
  wire _17824_;
  wire _17825_;
  wire _17826_;
  wire _17827_;
  wire _17828_;
  wire _17829_;
  wire _17830_;
  wire _17831_;
  wire _17832_;
  wire _17833_;
  wire _17834_;
  wire _17835_;
  wire _17836_;
  wire _17837_;
  wire _17838_;
  wire _17839_;
  wire _17840_;
  wire _17841_;
  wire _17842_;
  wire _17843_;
  wire _17844_;
  wire _17845_;
  wire _17846_;
  wire _17847_;
  wire _17848_;
  wire _17849_;
  wire _17850_;
  wire _17851_;
  wire _17852_;
  wire _17853_;
  wire _17854_;
  wire _17855_;
  wire _17856_;
  wire _17857_;
  wire _17858_;
  wire _17859_;
  wire _17860_;
  wire _17861_;
  wire _17862_;
  wire _17863_;
  wire _17864_;
  wire _17865_;
  wire _17866_;
  wire _17867_;
  wire _17868_;
  wire _17869_;
  wire _17870_;
  wire _17871_;
  wire _17872_;
  wire _17873_;
  wire _17874_;
  wire _17875_;
  wire _17876_;
  wire _17877_;
  wire _17878_;
  wire _17879_;
  wire _17880_;
  wire _17881_;
  wire _17882_;
  wire _17883_;
  wire _17884_;
  wire _17885_;
  wire _17886_;
  wire _17887_;
  wire _17888_;
  wire _17889_;
  wire _17890_;
  wire _17891_;
  wire _17892_;
  wire _17893_;
  wire _17894_;
  wire _17895_;
  wire _17896_;
  wire _17897_;
  wire _17898_;
  wire _17899_;
  wire _17900_;
  wire _17901_;
  wire _17902_;
  wire _17903_;
  wire _17904_;
  wire _17905_;
  wire _17906_;
  wire _17907_;
  wire _17908_;
  wire _17909_;
  wire _17910_;
  wire _17911_;
  wire _17912_;
  wire _17913_;
  wire _17914_;
  wire _17915_;
  wire _17916_;
  wire _17917_;
  wire _17918_;
  wire _17919_;
  wire _17920_;
  wire _17921_;
  wire _17922_;
  wire _17923_;
  wire _17924_;
  wire _17925_;
  wire _17926_;
  wire _17927_;
  wire _17928_;
  wire _17929_;
  wire _17930_;
  wire _17931_;
  wire _17932_;
  wire _17933_;
  wire _17934_;
  wire _17935_;
  wire _17936_;
  wire _17937_;
  wire _17938_;
  wire _17939_;
  wire _17940_;
  wire _17941_;
  wire _17942_;
  wire _17943_;
  wire _17944_;
  wire _17945_;
  wire _17946_;
  wire _17947_;
  wire _17948_;
  wire _17949_;
  wire _17950_;
  wire _17951_;
  wire _17952_;
  wire _17953_;
  wire _17954_;
  wire _17955_;
  wire _17956_;
  wire _17957_;
  wire _17958_;
  wire _17959_;
  wire _17960_;
  wire _17961_;
  wire _17962_;
  wire _17963_;
  wire _17964_;
  wire _17965_;
  wire _17966_;
  wire _17967_;
  wire _17968_;
  wire _17969_;
  wire _17970_;
  wire _17971_;
  wire _17972_;
  wire _17973_;
  wire _17974_;
  wire _17975_;
  wire _17976_;
  wire _17977_;
  wire _17978_;
  wire _17979_;
  wire _17980_;
  wire _17981_;
  wire _17982_;
  wire _17983_;
  wire _17984_;
  wire _17985_;
  wire _17986_;
  wire _17987_;
  wire _17988_;
  wire _17989_;
  wire _17990_;
  wire _17991_;
  wire _17992_;
  wire _17993_;
  wire _17994_;
  wire _17995_;
  wire _17996_;
  wire _17997_;
  wire _17998_;
  wire _17999_;
  wire _18000_;
  wire _18001_;
  wire _18002_;
  wire _18003_;
  wire _18004_;
  wire _18005_;
  wire _18006_;
  wire _18007_;
  wire _18008_;
  wire _18009_;
  wire _18010_;
  wire _18011_;
  wire _18012_;
  wire _18013_;
  wire _18014_;
  wire _18015_;
  wire _18016_;
  wire _18017_;
  wire _18018_;
  wire _18019_;
  wire _18020_;
  wire _18021_;
  wire _18022_;
  wire _18023_;
  wire _18024_;
  wire _18025_;
  wire _18026_;
  wire _18027_;
  wire _18028_;
  wire _18029_;
  wire _18030_;
  wire _18031_;
  wire _18032_;
  wire _18033_;
  wire _18034_;
  wire _18035_;
  wire _18036_;
  wire _18037_;
  wire _18038_;
  wire _18039_;
  wire _18040_;
  wire _18041_;
  wire _18042_;
  wire _18043_;
  wire _18044_;
  wire _18045_;
  wire _18046_;
  wire _18047_;
  wire _18048_;
  wire _18049_;
  wire _18050_;
  wire _18051_;
  wire _18052_;
  wire _18053_;
  wire _18054_;
  wire _18055_;
  wire _18056_;
  wire _18057_;
  wire _18058_;
  wire _18059_;
  wire _18060_;
  wire _18061_;
  wire _18062_;
  wire _18063_;
  wire _18064_;
  wire _18065_;
  wire _18066_;
  wire _18067_;
  wire _18068_;
  wire _18069_;
  wire _18070_;
  wire _18071_;
  wire _18072_;
  wire _18073_;
  wire _18074_;
  wire _18075_;
  wire _18076_;
  wire _18077_;
  wire _18078_;
  wire _18079_;
  wire _18080_;
  wire _18081_;
  wire _18082_;
  wire _18083_;
  wire _18084_;
  wire _18085_;
  wire _18086_;
  wire _18087_;
  wire _18088_;
  wire _18089_;
  wire _18090_;
  wire _18091_;
  wire _18092_;
  wire _18093_;
  wire _18094_;
  wire _18095_;
  wire _18096_;
  wire _18097_;
  wire _18098_;
  wire _18099_;
  wire _18100_;
  wire _18101_;
  wire _18102_;
  wire _18103_;
  wire _18104_;
  wire _18105_;
  wire _18106_;
  wire _18107_;
  wire _18108_;
  wire _18109_;
  wire _18110_;
  wire _18111_;
  wire _18112_;
  wire _18113_;
  wire _18114_;
  wire _18115_;
  wire _18116_;
  wire _18117_;
  wire _18118_;
  wire _18119_;
  wire _18120_;
  wire _18121_;
  wire _18122_;
  wire _18123_;
  wire _18124_;
  wire _18125_;
  wire _18126_;
  wire _18127_;
  wire _18128_;
  wire _18129_;
  wire _18130_;
  wire _18131_;
  wire _18132_;
  wire _18133_;
  wire _18134_;
  wire _18135_;
  wire _18136_;
  wire _18137_;
  wire _18138_;
  wire _18139_;
  wire _18140_;
  wire _18141_;
  wire _18142_;
  wire _18143_;
  wire _18144_;
  wire _18145_;
  wire _18146_;
  wire _18147_;
  wire _18148_;
  wire _18149_;
  wire _18150_;
  wire _18151_;
  wire _18152_;
  wire _18153_;
  wire _18154_;
  wire _18155_;
  wire _18156_;
  wire _18157_;
  wire _18158_;
  wire _18159_;
  wire _18160_;
  wire _18161_;
  wire _18162_;
  wire _18163_;
  wire _18164_;
  wire _18165_;
  wire _18166_;
  wire _18167_;
  wire _18168_;
  wire _18169_;
  wire _18170_;
  wire _18171_;
  wire _18172_;
  wire _18173_;
  wire _18174_;
  wire _18175_;
  wire _18176_;
  wire _18177_;
  wire _18178_;
  wire _18179_;
  wire _18180_;
  wire _18181_;
  wire _18182_;
  wire _18183_;
  wire _18184_;
  wire _18185_;
  wire _18186_;
  wire _18187_;
  wire _18188_;
  wire _18189_;
  wire _18190_;
  wire _18191_;
  wire _18192_;
  wire _18193_;
  wire _18194_;
  wire _18195_;
  wire _18196_;
  wire _18197_;
  wire _18198_;
  wire _18199_;
  wire _18200_;
  wire _18201_;
  wire _18202_;
  wire _18203_;
  wire _18204_;
  wire _18205_;
  wire _18206_;
  wire _18207_;
  wire _18208_;
  wire _18209_;
  wire _18210_;
  wire _18211_;
  wire _18212_;
  wire _18213_;
  wire _18214_;
  wire _18215_;
  wire _18216_;
  wire _18217_;
  wire _18218_;
  wire _18219_;
  wire _18220_;
  wire _18221_;
  wire _18222_;
  wire _18223_;
  wire _18224_;
  wire _18225_;
  wire _18226_;
  wire _18227_;
  wire _18228_;
  wire _18229_;
  wire _18230_;
  wire _18231_;
  wire _18232_;
  wire _18233_;
  wire _18234_;
  wire _18235_;
  wire _18236_;
  wire _18237_;
  wire _18238_;
  wire _18239_;
  wire _18240_;
  wire _18241_;
  wire _18242_;
  wire _18243_;
  wire _18244_;
  wire _18245_;
  wire _18246_;
  wire _18247_;
  wire _18248_;
  wire _18249_;
  wire _18250_;
  wire _18251_;
  wire _18252_;
  wire _18253_;
  wire _18254_;
  wire _18255_;
  wire _18256_;
  wire _18257_;
  wire _18258_;
  wire _18259_;
  wire _18260_;
  wire _18261_;
  wire _18262_;
  wire _18263_;
  wire _18264_;
  wire _18265_;
  wire _18266_;
  wire _18267_;
  wire _18268_;
  wire _18269_;
  wire _18270_;
  wire _18271_;
  wire _18272_;
  wire _18273_;
  wire _18274_;
  wire _18275_;
  wire _18276_;
  wire _18277_;
  wire _18278_;
  wire _18279_;
  wire _18280_;
  wire _18281_;
  wire _18282_;
  wire _18283_;
  wire _18284_;
  wire _18285_;
  wire _18286_;
  wire _18287_;
  wire _18288_;
  wire _18289_;
  wire _18290_;
  wire _18291_;
  wire _18292_;
  wire _18293_;
  wire _18294_;
  wire _18295_;
  wire _18296_;
  wire _18297_;
  wire _18298_;
  wire _18299_;
  wire _18300_;
  wire _18301_;
  wire _18302_;
  wire _18303_;
  wire _18304_;
  wire _18305_;
  wire _18306_;
  wire _18307_;
  wire _18308_;
  wire _18309_;
  wire _18310_;
  wire _18311_;
  wire _18312_;
  wire _18313_;
  wire _18314_;
  wire _18315_;
  wire _18316_;
  wire _18317_;
  wire _18318_;
  wire _18319_;
  wire _18320_;
  wire _18321_;
  wire _18322_;
  wire _18323_;
  wire _18324_;
  wire _18325_;
  wire _18326_;
  wire _18327_;
  wire _18328_;
  wire _18329_;
  wire _18330_;
  wire _18331_;
  wire _18332_;
  wire _18333_;
  wire _18334_;
  wire _18335_;
  wire _18336_;
  wire _18337_;
  wire _18338_;
  wire _18339_;
  wire _18340_;
  wire _18341_;
  wire _18342_;
  wire _18343_;
  wire _18344_;
  wire _18345_;
  wire _18346_;
  wire _18347_;
  wire _18348_;
  wire _18349_;
  wire _18350_;
  wire _18351_;
  wire _18352_;
  wire _18353_;
  wire _18354_;
  wire _18355_;
  wire _18356_;
  wire _18357_;
  wire _18358_;
  wire _18359_;
  wire _18360_;
  wire _18361_;
  wire _18362_;
  wire _18363_;
  wire _18364_;
  wire _18365_;
  wire _18366_;
  wire _18367_;
  wire _18368_;
  wire _18369_;
  wire _18370_;
  wire _18371_;
  wire _18372_;
  wire _18373_;
  wire _18374_;
  wire _18375_;
  wire _18376_;
  wire _18377_;
  wire _18378_;
  wire _18379_;
  wire _18380_;
  wire _18381_;
  wire _18382_;
  wire _18383_;
  wire _18384_;
  wire _18385_;
  wire _18386_;
  wire _18387_;
  wire _18388_;
  wire _18389_;
  wire _18390_;
  wire _18391_;
  wire _18392_;
  wire _18393_;
  wire _18394_;
  wire _18395_;
  wire _18396_;
  wire _18397_;
  wire _18398_;
  wire _18399_;
  wire _18400_;
  wire _18401_;
  wire _18402_;
  wire _18403_;
  wire _18404_;
  wire _18405_;
  wire _18406_;
  wire _18407_;
  wire _18408_;
  wire _18409_;
  wire _18410_;
  wire _18411_;
  wire _18412_;
  wire _18413_;
  wire _18414_;
  wire _18415_;
  wire _18416_;
  wire _18417_;
  wire _18418_;
  wire _18419_;
  wire _18420_;
  wire _18421_;
  wire _18422_;
  wire _18423_;
  wire _18424_;
  wire _18425_;
  wire _18426_;
  wire _18427_;
  wire _18428_;
  wire _18429_;
  wire _18430_;
  wire _18431_;
  wire _18432_;
  wire _18433_;
  wire _18434_;
  wire _18435_;
  wire _18436_;
  wire _18437_;
  wire _18438_;
  wire _18439_;
  wire _18440_;
  wire _18441_;
  wire _18442_;
  wire _18443_;
  wire _18444_;
  wire _18445_;
  wire _18446_;
  wire _18447_;
  wire _18448_;
  wire _18449_;
  wire _18450_;
  wire _18451_;
  wire _18452_;
  wire _18453_;
  wire _18454_;
  wire _18455_;
  wire _18456_;
  wire _18457_;
  wire _18458_;
  wire _18459_;
  wire _18460_;
  wire _18461_;
  wire _18462_;
  wire _18463_;
  wire _18464_;
  wire _18465_;
  wire _18466_;
  wire _18467_;
  wire _18468_;
  wire _18469_;
  wire _18470_;
  wire _18471_;
  wire _18472_;
  wire _18473_;
  wire _18474_;
  wire _18475_;
  wire _18476_;
  wire _18477_;
  wire _18478_;
  wire _18479_;
  wire _18480_;
  wire _18481_;
  wire _18482_;
  wire _18483_;
  wire _18484_;
  wire _18485_;
  wire _18486_;
  wire _18487_;
  wire _18488_;
  wire _18489_;
  wire _18490_;
  wire _18491_;
  wire _18492_;
  wire _18493_;
  wire _18494_;
  wire _18495_;
  wire _18496_;
  wire _18497_;
  wire _18498_;
  wire _18499_;
  wire _18500_;
  wire _18501_;
  wire _18502_;
  wire _18503_;
  wire _18504_;
  wire _18505_;
  wire _18506_;
  wire _18507_;
  wire _18508_;
  wire _18509_;
  wire _18510_;
  wire _18511_;
  wire _18512_;
  wire _18513_;
  wire _18514_;
  wire _18515_;
  wire _18516_;
  wire _18517_;
  wire _18518_;
  wire _18519_;
  wire _18520_;
  wire _18521_;
  wire _18522_;
  wire _18523_;
  wire _18524_;
  wire _18525_;
  wire _18526_;
  wire _18527_;
  wire _18528_;
  wire _18529_;
  wire _18530_;
  wire _18531_;
  wire _18532_;
  wire _18533_;
  wire _18534_;
  wire _18535_;
  wire _18536_;
  wire _18537_;
  wire _18538_;
  wire _18539_;
  wire _18540_;
  wire _18541_;
  wire _18542_;
  wire _18543_;
  wire _18544_;
  wire _18545_;
  wire _18546_;
  wire _18547_;
  wire _18548_;
  wire _18549_;
  wire _18550_;
  wire _18551_;
  wire _18552_;
  wire _18553_;
  wire _18554_;
  wire _18555_;
  wire _18556_;
  wire _18557_;
  wire _18558_;
  wire _18559_;
  wire _18560_;
  wire _18561_;
  wire _18562_;
  wire _18563_;
  wire _18564_;
  wire _18565_;
  wire _18566_;
  wire _18567_;
  wire _18568_;
  wire _18569_;
  wire _18570_;
  wire _18571_;
  wire _18572_;
  wire _18573_;
  wire _18574_;
  wire _18575_;
  wire _18576_;
  wire _18577_;
  wire _18578_;
  wire _18579_;
  wire _18580_;
  wire _18581_;
  wire _18582_;
  wire _18583_;
  wire _18584_;
  wire _18585_;
  wire _18586_;
  wire _18587_;
  wire _18588_;
  wire _18589_;
  wire _18590_;
  wire _18591_;
  wire _18592_;
  wire _18593_;
  wire _18594_;
  wire _18595_;
  wire _18596_;
  wire _18597_;
  wire _18598_;
  wire _18599_;
  wire _18600_;
  wire _18601_;
  wire _18602_;
  wire _18603_;
  wire _18604_;
  wire _18605_;
  wire _18606_;
  wire _18607_;
  wire _18608_;
  wire _18609_;
  wire _18610_;
  wire _18611_;
  wire _18612_;
  wire _18613_;
  wire _18614_;
  wire _18615_;
  wire _18616_;
  wire _18617_;
  wire _18618_;
  wire _18619_;
  wire _18620_;
  wire _18621_;
  wire _18622_;
  wire _18623_;
  wire _18624_;
  wire _18625_;
  wire _18626_;
  wire _18627_;
  wire _18628_;
  wire _18629_;
  wire _18630_;
  wire _18631_;
  wire _18632_;
  wire _18633_;
  wire _18634_;
  wire _18635_;
  wire _18636_;
  wire _18637_;
  wire _18638_;
  wire _18639_;
  wire _18640_;
  wire _18641_;
  wire _18642_;
  wire _18643_;
  wire _18644_;
  wire _18645_;
  wire _18646_;
  wire _18647_;
  wire _18648_;
  wire _18649_;
  wire _18650_;
  wire _18651_;
  wire _18652_;
  wire _18653_;
  wire _18654_;
  wire _18655_;
  wire _18656_;
  wire _18657_;
  wire _18658_;
  wire _18659_;
  wire _18660_;
  wire _18661_;
  wire _18662_;
  wire _18663_;
  wire _18664_;
  wire _18665_;
  wire _18666_;
  wire _18667_;
  wire _18668_;
  wire _18669_;
  wire _18670_;
  wire _18671_;
  wire _18672_;
  wire _18673_;
  wire _18674_;
  wire _18675_;
  wire _18676_;
  wire _18677_;
  wire _18678_;
  wire _18679_;
  wire _18680_;
  wire _18681_;
  wire _18682_;
  wire _18683_;
  wire _18684_;
  wire _18685_;
  wire _18686_;
  wire _18687_;
  wire _18688_;
  wire _18689_;
  wire _18690_;
  wire _18691_;
  wire _18692_;
  wire _18693_;
  wire _18694_;
  wire _18695_;
  wire _18696_;
  wire _18697_;
  wire _18698_;
  wire _18699_;
  wire _18700_;
  wire _18701_;
  wire _18702_;
  wire _18703_;
  wire _18704_;
  wire _18705_;
  wire _18706_;
  wire _18707_;
  wire _18708_;
  wire _18709_;
  wire _18710_;
  wire _18711_;
  wire _18712_;
  wire _18713_;
  wire _18714_;
  wire _18715_;
  wire _18716_;
  wire _18717_;
  wire _18718_;
  wire _18719_;
  wire _18720_;
  wire _18721_;
  wire _18722_;
  wire _18723_;
  wire _18724_;
  wire _18725_;
  wire _18726_;
  wire _18727_;
  wire _18728_;
  wire _18729_;
  wire _18730_;
  wire _18731_;
  wire _18732_;
  wire _18733_;
  wire _18734_;
  wire _18735_;
  wire _18736_;
  wire _18737_;
  wire _18738_;
  wire _18739_;
  wire _18740_;
  wire _18741_;
  wire _18742_;
  wire _18743_;
  wire _18744_;
  wire _18745_;
  wire _18746_;
  wire _18747_;
  wire _18748_;
  wire _18749_;
  wire _18750_;
  wire _18751_;
  wire _18752_;
  wire _18753_;
  wire _18754_;
  wire _18755_;
  wire _18756_;
  wire _18757_;
  wire _18758_;
  wire _18759_;
  wire _18760_;
  wire _18761_;
  wire _18762_;
  wire _18763_;
  wire _18764_;
  wire _18765_;
  wire _18766_;
  wire _18767_;
  wire _18768_;
  wire _18769_;
  wire _18770_;
  wire _18771_;
  wire _18772_;
  wire _18773_;
  wire _18774_;
  wire _18775_;
  wire _18776_;
  wire _18777_;
  wire _18778_;
  wire _18779_;
  wire _18780_;
  wire _18781_;
  wire _18782_;
  wire _18783_;
  wire _18784_;
  wire _18785_;
  wire _18786_;
  wire _18787_;
  wire _18788_;
  wire _18789_;
  wire _18790_;
  wire _18791_;
  wire _18792_;
  wire _18793_;
  wire _18794_;
  wire _18795_;
  wire _18796_;
  wire _18797_;
  wire _18798_;
  wire _18799_;
  wire _18800_;
  wire _18801_;
  wire _18802_;
  wire _18803_;
  wire _18804_;
  wire _18805_;
  wire _18806_;
  wire _18807_;
  wire _18808_;
  wire _18809_;
  wire _18810_;
  wire _18811_;
  wire _18812_;
  wire _18813_;
  wire _18814_;
  wire _18815_;
  wire _18816_;
  wire _18817_;
  wire _18818_;
  wire _18819_;
  wire _18820_;
  wire _18821_;
  wire _18822_;
  wire _18823_;
  wire _18824_;
  wire _18825_;
  wire _18826_;
  wire _18827_;
  wire _18828_;
  wire _18829_;
  wire _18830_;
  wire _18831_;
  wire _18832_;
  wire _18833_;
  wire _18834_;
  wire _18835_;
  wire _18836_;
  wire _18837_;
  wire _18838_;
  wire _18839_;
  wire _18840_;
  wire _18841_;
  wire _18842_;
  wire _18843_;
  wire _18844_;
  wire _18845_;
  wire _18846_;
  wire _18847_;
  wire _18848_;
  wire _18849_;
  wire _18850_;
  wire _18851_;
  wire _18852_;
  wire _18853_;
  wire _18854_;
  wire _18855_;
  wire _18856_;
  wire _18857_;
  wire _18858_;
  wire _18859_;
  wire _18860_;
  wire _18861_;
  wire _18862_;
  wire _18863_;
  wire _18864_;
  wire _18865_;
  wire _18866_;
  wire _18867_;
  wire _18868_;
  wire _18869_;
  wire _18870_;
  wire _18871_;
  wire _18872_;
  wire _18873_;
  wire _18874_;
  wire _18875_;
  wire _18876_;
  wire _18877_;
  wire _18878_;
  wire _18879_;
  wire _18880_;
  wire _18881_;
  wire _18882_;
  wire _18883_;
  wire _18884_;
  wire _18885_;
  wire _18886_;
  wire _18887_;
  wire _18888_;
  wire _18889_;
  wire _18890_;
  wire _18891_;
  wire _18892_;
  wire _18893_;
  wire _18894_;
  wire _18895_;
  wire _18896_;
  wire _18897_;
  wire _18898_;
  wire _18899_;
  wire _18900_;
  wire _18901_;
  wire _18902_;
  wire _18903_;
  wire _18904_;
  wire _18905_;
  wire _18906_;
  wire _18907_;
  wire _18908_;
  wire _18909_;
  wire _18910_;
  wire _18911_;
  wire _18912_;
  wire _18913_;
  wire _18914_;
  wire _18915_;
  wire _18916_;
  wire _18917_;
  wire _18918_;
  wire _18919_;
  wire _18920_;
  wire _18921_;
  wire _18922_;
  wire _18923_;
  wire _18924_;
  wire _18925_;
  wire _18926_;
  wire _18927_;
  wire _18928_;
  wire _18929_;
  wire _18930_;
  wire _18931_;
  wire _18932_;
  wire _18933_;
  wire _18934_;
  wire _18935_;
  wire _18936_;
  wire _18937_;
  wire _18938_;
  wire _18939_;
  wire _18940_;
  wire _18941_;
  wire _18942_;
  wire _18943_;
  wire _18944_;
  wire _18945_;
  wire _18946_;
  wire _18947_;
  wire _18948_;
  wire _18949_;
  wire _18950_;
  wire _18951_;
  wire _18952_;
  wire _18953_;
  wire _18954_;
  wire _18955_;
  wire _18956_;
  wire _18957_;
  wire _18958_;
  wire _18959_;
  wire _18960_;
  wire _18961_;
  wire _18962_;
  wire _18963_;
  wire _18964_;
  wire _18965_;
  wire _18966_;
  wire _18967_;
  wire _18968_;
  wire _18969_;
  wire _18970_;
  wire _18971_;
  wire _18972_;
  wire _18973_;
  wire _18974_;
  wire _18975_;
  wire _18976_;
  wire _18977_;
  wire _18978_;
  wire _18979_;
  wire _18980_;
  wire _18981_;
  wire _18982_;
  wire _18983_;
  wire _18984_;
  wire _18985_;
  wire _18986_;
  wire _18987_;
  wire _18988_;
  wire _18989_;
  wire _18990_;
  wire _18991_;
  wire _18992_;
  wire _18993_;
  wire _18994_;
  wire _18995_;
  wire _18996_;
  wire _18997_;
  wire _18998_;
  wire _18999_;
  wire _19000_;
  wire _19001_;
  wire _19002_;
  wire _19003_;
  wire _19004_;
  wire _19005_;
  wire _19006_;
  wire _19007_;
  wire _19008_;
  wire _19009_;
  wire _19010_;
  wire _19011_;
  wire _19012_;
  wire _19013_;
  wire _19014_;
  wire _19015_;
  wire _19016_;
  wire _19017_;
  wire _19018_;
  wire _19019_;
  wire _19020_;
  wire _19021_;
  wire _19022_;
  wire _19023_;
  wire _19024_;
  wire _19025_;
  wire _19026_;
  wire _19027_;
  wire _19028_;
  wire _19029_;
  wire _19030_;
  wire _19031_;
  wire _19032_;
  wire _19033_;
  wire _19034_;
  wire _19035_;
  wire _19036_;
  wire _19037_;
  wire _19038_;
  wire _19039_;
  wire _19040_;
  wire _19041_;
  wire _19042_;
  wire _19043_;
  wire _19044_;
  wire _19045_;
  wire _19046_;
  wire _19047_;
  wire _19048_;
  wire _19049_;
  wire _19050_;
  wire _19051_;
  wire _19052_;
  wire _19053_;
  wire _19054_;
  wire _19055_;
  wire _19056_;
  wire _19057_;
  wire _19058_;
  wire _19059_;
  wire _19060_;
  wire _19061_;
  wire _19062_;
  wire _19063_;
  wire _19064_;
  wire _19065_;
  wire _19066_;
  wire _19067_;
  wire _19068_;
  wire _19069_;
  wire _19070_;
  wire _19071_;
  wire _19072_;
  wire _19073_;
  wire _19074_;
  wire _19075_;
  wire _19076_;
  wire _19077_;
  wire _19078_;
  wire _19079_;
  wire _19080_;
  wire _19081_;
  wire _19082_;
  wire _19083_;
  wire _19084_;
  wire _19085_;
  wire _19086_;
  wire _19087_;
  wire _19088_;
  wire _19089_;
  wire _19090_;
  wire _19091_;
  wire _19092_;
  wire _19093_;
  wire _19094_;
  wire _19095_;
  wire _19096_;
  wire _19097_;
  wire _19098_;
  wire _19099_;
  wire _19100_;
  wire _19101_;
  wire _19102_;
  wire _19103_;
  wire _19104_;
  wire _19105_;
  wire _19106_;
  wire _19107_;
  wire _19108_;
  wire _19109_;
  wire _19110_;
  wire _19111_;
  wire _19112_;
  wire _19113_;
  wire _19114_;
  wire _19115_;
  wire _19116_;
  wire _19117_;
  wire _19118_;
  wire _19119_;
  wire _19120_;
  wire _19121_;
  wire _19122_;
  wire _19123_;
  wire _19124_;
  wire _19125_;
  wire _19126_;
  wire _19127_;
  wire _19128_;
  wire _19129_;
  wire _19130_;
  wire _19131_;
  wire _19132_;
  wire _19133_;
  wire _19134_;
  wire _19135_;
  wire _19136_;
  wire _19137_;
  wire _19138_;
  wire _19139_;
  wire _19140_;
  wire _19141_;
  wire _19142_;
  wire _19143_;
  wire _19144_;
  wire _19145_;
  wire _19146_;
  wire _19147_;
  wire _19148_;
  wire _19149_;
  wire _19150_;
  wire _19151_;
  wire _19152_;
  wire _19153_;
  wire _19154_;
  wire _19155_;
  wire _19156_;
  wire _19157_;
  wire _19158_;
  wire _19159_;
  wire _19160_;
  wire _19161_;
  wire _19162_;
  wire _19163_;
  wire _19164_;
  wire _19165_;
  wire _19166_;
  wire _19167_;
  wire _19168_;
  wire _19169_;
  wire _19170_;
  wire _19171_;
  wire _19172_;
  wire _19173_;
  wire _19174_;
  wire _19175_;
  wire _19176_;
  wire _19177_;
  wire _19178_;
  wire _19179_;
  wire _19180_;
  wire _19181_;
  wire _19182_;
  wire _19183_;
  wire _19184_;
  wire _19185_;
  wire _19186_;
  wire _19187_;
  wire _19188_;
  wire _19189_;
  wire _19190_;
  wire _19191_;
  wire _19192_;
  wire _19193_;
  wire _19194_;
  wire _19195_;
  wire _19196_;
  wire _19197_;
  wire _19198_;
  wire _19199_;
  wire _19200_;
  wire _19201_;
  wire _19202_;
  wire _19203_;
  wire _19204_;
  wire _19205_;
  wire _19206_;
  wire _19207_;
  wire _19208_;
  wire _19209_;
  wire _19210_;
  wire _19211_;
  wire _19212_;
  wire _19213_;
  wire _19214_;
  wire _19215_;
  wire _19216_;
  wire _19217_;
  wire _19218_;
  wire _19219_;
  wire _19220_;
  wire _19221_;
  wire _19222_;
  wire _19223_;
  wire _19224_;
  wire _19225_;
  wire _19226_;
  wire _19227_;
  wire _19228_;
  wire _19229_;
  wire _19230_;
  wire _19231_;
  wire _19232_;
  wire _19233_;
  wire _19234_;
  wire _19235_;
  wire _19236_;
  wire _19237_;
  wire _19238_;
  wire _19239_;
  wire _19240_;
  wire _19241_;
  wire _19242_;
  wire _19243_;
  wire _19244_;
  wire _19245_;
  wire _19246_;
  wire _19247_;
  wire _19248_;
  wire _19249_;
  wire _19250_;
  wire _19251_;
  wire _19252_;
  wire _19253_;
  wire _19254_;
  wire _19255_;
  wire _19256_;
  wire _19257_;
  wire _19258_;
  wire _19259_;
  wire _19260_;
  wire _19261_;
  wire _19262_;
  wire _19263_;
  wire _19264_;
  wire _19265_;
  wire _19266_;
  wire _19267_;
  wire _19268_;
  wire _19269_;
  wire _19270_;
  wire _19271_;
  wire _19272_;
  wire _19273_;
  wire _19274_;
  wire _19275_;
  wire _19276_;
  wire _19277_;
  wire _19278_;
  wire _19279_;
  wire _19280_;
  wire _19281_;
  wire _19282_;
  wire _19283_;
  wire _19284_;
  wire _19285_;
  wire _19286_;
  wire _19287_;
  wire _19288_;
  wire _19289_;
  wire _19290_;
  wire _19291_;
  wire _19292_;
  wire _19293_;
  wire _19294_;
  wire _19295_;
  wire _19296_;
  wire _19297_;
  wire _19298_;
  wire _19299_;
  wire _19300_;
  wire _19301_;
  wire _19302_;
  wire _19303_;
  wire _19304_;
  wire _19305_;
  wire _19306_;
  wire _19307_;
  wire _19308_;
  wire _19309_;
  wire _19310_;
  wire _19311_;
  wire _19312_;
  wire _19313_;
  wire _19314_;
  wire _19315_;
  wire _19316_;
  wire _19317_;
  wire _19318_;
  wire _19319_;
  wire _19320_;
  wire _19321_;
  wire _19322_;
  wire _19323_;
  wire _19324_;
  wire _19325_;
  wire _19326_;
  wire _19327_;
  wire _19328_;
  wire _19329_;
  wire _19330_;
  wire _19331_;
  wire _19332_;
  wire _19333_;
  wire _19334_;
  wire _19335_;
  wire _19336_;
  wire _19337_;
  wire _19338_;
  wire _19339_;
  wire _19340_;
  wire _19341_;
  wire _19342_;
  wire _19343_;
  wire _19344_;
  wire _19345_;
  wire _19346_;
  wire _19347_;
  wire _19348_;
  wire _19349_;
  wire _19350_;
  wire _19351_;
  wire _19352_;
  wire _19353_;
  wire _19354_;
  wire _19355_;
  wire _19356_;
  wire _19357_;
  wire _19358_;
  wire _19359_;
  wire _19360_;
  wire _19361_;
  wire _19362_;
  wire _19363_;
  wire _19364_;
  wire _19365_;
  wire _19366_;
  wire _19367_;
  wire _19368_;
  wire _19369_;
  wire _19370_;
  wire _19371_;
  wire _19372_;
  wire _19373_;
  wire _19374_;
  wire _19375_;
  wire _19376_;
  wire _19377_;
  wire _19378_;
  wire _19379_;
  wire _19380_;
  wire _19381_;
  wire _19382_;
  wire _19383_;
  wire _19384_;
  wire _19385_;
  wire _19386_;
  wire _19387_;
  wire _19388_;
  wire _19389_;
  wire _19390_;
  wire _19391_;
  wire _19392_;
  wire _19393_;
  wire _19394_;
  wire _19395_;
  wire _19396_;
  wire _19397_;
  wire _19398_;
  wire _19399_;
  wire _19400_;
  wire _19401_;
  wire _19402_;
  wire _19403_;
  wire _19404_;
  wire _19405_;
  wire _19406_;
  wire _19407_;
  wire _19408_;
  wire _19409_;
  wire _19410_;
  wire _19411_;
  wire _19412_;
  wire _19413_;
  wire _19414_;
  wire _19415_;
  wire _19416_;
  wire _19417_;
  wire _19418_;
  wire _19419_;
  wire _19420_;
  wire _19421_;
  wire _19422_;
  wire _19423_;
  wire _19424_;
  wire _19425_;
  wire _19426_;
  wire _19427_;
  wire _19428_;
  wire _19429_;
  wire _19430_;
  wire _19431_;
  wire _19432_;
  wire _19433_;
  wire _19434_;
  wire _19435_;
  wire _19436_;
  wire _19437_;
  wire _19438_;
  wire _19439_;
  wire _19440_;
  wire _19441_;
  wire _19442_;
  wire _19443_;
  wire _19444_;
  wire _19445_;
  wire _19446_;
  wire _19447_;
  wire _19448_;
  wire _19449_;
  wire _19450_;
  wire _19451_;
  wire _19452_;
  wire _19453_;
  wire _19454_;
  wire _19455_;
  wire _19456_;
  wire _19457_;
  wire _19458_;
  wire _19459_;
  wire _19460_;
  wire _19461_;
  wire _19462_;
  wire _19463_;
  wire _19464_;
  wire _19465_;
  wire _19466_;
  wire _19467_;
  wire _19468_;
  wire _19469_;
  wire _19470_;
  wire _19471_;
  wire _19472_;
  wire _19473_;
  wire _19474_;
  wire _19475_;
  wire _19476_;
  wire _19477_;
  wire _19478_;
  wire _19479_;
  wire _19480_;
  wire _19481_;
  wire _19482_;
  wire _19483_;
  wire _19484_;
  wire _19485_;
  wire _19486_;
  wire _19487_;
  wire _19488_;
  wire _19489_;
  wire _19490_;
  wire _19491_;
  wire _19492_;
  wire _19493_;
  wire _19494_;
  wire _19495_;
  wire _19496_;
  wire _19497_;
  wire _19498_;
  wire _19499_;
  wire _19500_;
  wire _19501_;
  wire _19502_;
  wire _19503_;
  wire _19504_;
  wire _19505_;
  wire _19506_;
  wire _19507_;
  wire _19508_;
  wire _19509_;
  wire _19510_;
  wire _19511_;
  wire _19512_;
  wire _19513_;
  wire _19514_;
  wire _19515_;
  wire _19516_;
  wire _19517_;
  wire _19518_;
  wire _19519_;
  wire _19520_;
  wire _19521_;
  wire _19522_;
  wire _19523_;
  wire _19524_;
  wire _19525_;
  wire _19526_;
  wire _19527_;
  wire _19528_;
  wire _19529_;
  wire _19530_;
  wire _19531_;
  wire _19532_;
  wire _19533_;
  wire _19534_;
  wire _19535_;
  wire _19536_;
  wire _19537_;
  wire _19538_;
  wire _19539_;
  wire _19540_;
  wire _19541_;
  wire _19542_;
  wire _19543_;
  wire _19544_;
  wire _19545_;
  wire _19546_;
  wire _19547_;
  wire _19548_;
  wire _19549_;
  wire _19550_;
  wire _19551_;
  wire _19552_;
  wire _19553_;
  wire _19554_;
  wire _19555_;
  wire _19556_;
  wire _19557_;
  wire _19558_;
  wire _19559_;
  wire _19560_;
  wire _19561_;
  wire _19562_;
  wire _19563_;
  wire _19564_;
  wire _19565_;
  wire _19566_;
  wire _19567_;
  wire _19568_;
  wire _19569_;
  wire _19570_;
  wire _19571_;
  wire _19572_;
  wire _19573_;
  wire _19574_;
  wire _19575_;
  wire _19576_;
  wire _19577_;
  wire _19578_;
  wire _19579_;
  wire _19580_;
  wire _19581_;
  wire _19582_;
  wire _19583_;
  wire _19584_;
  wire _19585_;
  wire _19586_;
  wire _19587_;
  wire _19588_;
  wire _19589_;
  wire _19590_;
  wire _19591_;
  wire _19592_;
  wire _19593_;
  wire _19594_;
  wire _19595_;
  wire _19596_;
  wire _19597_;
  wire _19598_;
  wire _19599_;
  wire _19600_;
  wire _19601_;
  wire _19602_;
  wire _19603_;
  wire _19604_;
  wire _19605_;
  wire _19606_;
  wire _19607_;
  wire _19608_;
  wire _19609_;
  wire _19610_;
  wire _19611_;
  wire _19612_;
  wire _19613_;
  wire _19614_;
  wire _19615_;
  wire _19616_;
  wire _19617_;
  wire _19618_;
  wire _19619_;
  wire _19620_;
  wire _19621_;
  wire _19622_;
  wire _19623_;
  wire _19624_;
  wire _19625_;
  wire _19626_;
  wire _19627_;
  wire _19628_;
  wire _19629_;
  wire _19630_;
  wire _19631_;
  wire _19632_;
  wire _19633_;
  wire _19634_;
  wire _19635_;
  wire _19636_;
  wire _19637_;
  wire _19638_;
  wire _19639_;
  wire _19640_;
  wire _19641_;
  wire _19642_;
  wire _19643_;
  wire _19644_;
  wire _19645_;
  wire _19646_;
  wire _19647_;
  wire _19648_;
  wire _19649_;
  wire _19650_;
  wire _19651_;
  wire _19652_;
  wire _19653_;
  wire _19654_;
  wire _19655_;
  wire _19656_;
  wire _19657_;
  wire _19658_;
  wire _19659_;
  wire _19660_;
  wire _19661_;
  wire _19662_;
  wire _19663_;
  wire _19664_;
  wire _19665_;
  wire _19666_;
  wire _19667_;
  wire _19668_;
  wire _19669_;
  wire _19670_;
  wire _19671_;
  wire _19672_;
  wire _19673_;
  wire _19674_;
  wire _19675_;
  wire _19676_;
  wire _19677_;
  wire _19678_;
  wire _19679_;
  wire _19680_;
  wire _19681_;
  wire _19682_;
  wire _19683_;
  wire _19684_;
  wire _19685_;
  wire _19686_;
  wire _19687_;
  wire _19688_;
  wire _19689_;
  wire _19690_;
  wire _19691_;
  wire _19692_;
  wire _19693_;
  wire _19694_;
  wire _19695_;
  wire _19696_;
  wire _19697_;
  wire _19698_;
  wire _19699_;
  wire _19700_;
  wire _19701_;
  wire _19702_;
  wire _19703_;
  wire _19704_;
  wire _19705_;
  wire _19706_;
  wire _19707_;
  wire _19708_;
  wire _19709_;
  wire _19710_;
  wire _19711_;
  wire _19712_;
  wire _19713_;
  wire _19714_;
  wire _19715_;
  wire _19716_;
  wire _19717_;
  wire _19718_;
  wire _19719_;
  wire _19720_;
  wire _19721_;
  wire _19722_;
  wire _19723_;
  wire _19724_;
  wire _19725_;
  wire _19726_;
  wire _19727_;
  wire _19728_;
  wire _19729_;
  wire _19730_;
  wire _19731_;
  wire _19732_;
  wire _19733_;
  wire _19734_;
  wire _19735_;
  wire _19736_;
  wire _19737_;
  wire _19738_;
  wire _19739_;
  wire _19740_;
  wire _19741_;
  wire _19742_;
  wire _19743_;
  wire _19744_;
  wire _19745_;
  wire _19746_;
  wire _19747_;
  wire _19748_;
  wire _19749_;
  wire _19750_;
  wire _19751_;
  wire _19752_;
  wire _19753_;
  wire _19754_;
  wire _19755_;
  wire _19756_;
  wire _19757_;
  wire _19758_;
  wire _19759_;
  wire _19760_;
  wire _19761_;
  wire _19762_;
  wire _19763_;
  wire _19764_;
  wire _19765_;
  wire _19766_;
  wire _19767_;
  wire _19768_;
  wire _19769_;
  wire _19770_;
  wire _19771_;
  wire _19772_;
  wire _19773_;
  wire _19774_;
  wire _19775_;
  wire _19776_;
  wire _19777_;
  wire _19778_;
  wire _19779_;
  wire _19780_;
  wire _19781_;
  wire _19782_;
  wire _19783_;
  wire _19784_;
  wire _19785_;
  wire _19786_;
  wire _19787_;
  wire _19788_;
  wire _19789_;
  wire _19790_;
  wire _19791_;
  wire _19792_;
  wire _19793_;
  wire _19794_;
  wire _19795_;
  wire _19796_;
  wire _19797_;
  wire _19798_;
  wire _19799_;
  wire _19800_;
  wire _19801_;
  wire _19802_;
  wire _19803_;
  wire _19804_;
  wire _19805_;
  wire _19806_;
  wire _19807_;
  wire _19808_;
  wire _19809_;
  wire _19810_;
  wire _19811_;
  wire _19812_;
  wire _19813_;
  wire _19814_;
  wire _19815_;
  wire _19816_;
  wire _19817_;
  wire _19818_;
  wire _19819_;
  wire _19820_;
  wire _19821_;
  wire _19822_;
  wire _19823_;
  wire _19824_;
  wire _19825_;
  wire _19826_;
  wire _19827_;
  wire _19828_;
  wire _19829_;
  wire _19830_;
  wire _19831_;
  wire _19832_;
  wire _19833_;
  wire _19834_;
  wire _19835_;
  wire _19836_;
  wire _19837_;
  wire _19838_;
  wire _19839_;
  wire _19840_;
  wire _19841_;
  wire _19842_;
  wire _19843_;
  wire _19844_;
  wire _19845_;
  wire _19846_;
  wire _19847_;
  wire _19848_;
  wire _19849_;
  wire _19850_;
  wire _19851_;
  wire _19852_;
  wire _19853_;
  wire _19854_;
  wire _19855_;
  wire _19856_;
  wire _19857_;
  wire _19858_;
  wire _19859_;
  wire _19860_;
  wire _19861_;
  wire _19862_;
  wire _19863_;
  wire _19864_;
  wire _19865_;
  wire _19866_;
  wire _19867_;
  wire _19868_;
  wire _19869_;
  wire _19870_;
  wire _19871_;
  wire _19872_;
  wire _19873_;
  wire _19874_;
  wire _19875_;
  wire _19876_;
  wire _19877_;
  wire _19878_;
  wire _19879_;
  wire _19880_;
  wire _19881_;
  wire _19882_;
  wire _19883_;
  wire _19884_;
  wire _19885_;
  wire _19886_;
  wire _19887_;
  wire _19888_;
  wire _19889_;
  wire _19890_;
  wire _19891_;
  wire _19892_;
  wire _19893_;
  wire _19894_;
  wire _19895_;
  wire _19896_;
  wire _19897_;
  wire _19898_;
  wire _19899_;
  wire _19900_;
  wire _19901_;
  wire _19902_;
  wire _19903_;
  wire _19904_;
  wire _19905_;
  wire _19906_;
  wire _19907_;
  wire _19908_;
  wire _19909_;
  wire _19910_;
  wire _19911_;
  wire _19912_;
  wire _19913_;
  wire _19914_;
  wire _19915_;
  wire _19916_;
  wire _19917_;
  wire _19918_;
  wire _19919_;
  wire _19920_;
  wire _19921_;
  wire _19922_;
  wire _19923_;
  wire _19924_;
  wire _19925_;
  wire _19926_;
  wire _19927_;
  wire _19928_;
  wire _19929_;
  wire _19930_;
  wire _19931_;
  wire _19932_;
  wire _19933_;
  wire _19934_;
  wire _19935_;
  wire _19936_;
  wire _19937_;
  wire _19938_;
  wire _19939_;
  wire _19940_;
  wire _19941_;
  wire _19942_;
  wire _19943_;
  wire _19944_;
  wire _19945_;
  wire _19946_;
  wire _19947_;
  wire _19948_;
  wire _19949_;
  wire _19950_;
  wire _19951_;
  wire _19952_;
  wire _19953_;
  wire _19954_;
  wire _19955_;
  wire _19956_;
  wire _19957_;
  wire _19958_;
  wire _19959_;
  wire _19960_;
  wire _19961_;
  wire _19962_;
  wire _19963_;
  wire _19964_;
  wire _19965_;
  wire _19966_;
  wire _19967_;
  wire _19968_;
  wire _19969_;
  wire _19970_;
  wire _19971_;
  wire _19972_;
  wire _19973_;
  wire _19974_;
  wire _19975_;
  wire _19976_;
  wire _19977_;
  wire _19978_;
  wire _19979_;
  wire _19980_;
  wire _19981_;
  wire _19982_;
  wire _19983_;
  wire _19984_;
  wire _19985_;
  wire _19986_;
  wire _19987_;
  wire _19988_;
  wire _19989_;
  wire _19990_;
  wire _19991_;
  wire _19992_;
  wire _19993_;
  wire _19994_;
  wire _19995_;
  wire _19996_;
  wire _19997_;
  wire _19998_;
  wire _19999_;
  wire _20000_;
  wire _20001_;
  wire _20002_;
  wire _20003_;
  wire _20004_;
  wire _20005_;
  wire _20006_;
  wire _20007_;
  wire _20008_;
  wire _20009_;
  wire _20010_;
  wire _20011_;
  wire _20012_;
  wire _20013_;
  wire _20014_;
  wire _20015_;
  wire _20016_;
  wire _20017_;
  wire _20018_;
  wire _20019_;
  wire _20020_;
  wire _20021_;
  wire _20022_;
  wire _20023_;
  wire _20024_;
  wire _20025_;
  wire _20026_;
  wire _20027_;
  wire _20028_;
  wire _20029_;
  wire _20030_;
  wire _20031_;
  wire _20032_;
  wire _20033_;
  wire _20034_;
  wire _20035_;
  wire _20036_;
  wire _20037_;
  wire _20038_;
  wire _20039_;
  wire _20040_;
  wire _20041_;
  wire _20042_;
  wire _20043_;
  wire _20044_;
  wire _20045_;
  wire _20046_;
  wire _20047_;
  wire _20048_;
  wire _20049_;
  wire _20050_;
  wire _20051_;
  wire _20052_;
  wire _20053_;
  wire _20054_;
  wire _20055_;
  wire _20056_;
  wire _20057_;
  wire _20058_;
  wire _20059_;
  wire _20060_;
  wire _20061_;
  wire _20062_;
  wire _20063_;
  wire _20064_;
  wire _20065_;
  wire _20066_;
  wire _20067_;
  wire _20068_;
  wire _20069_;
  wire _20070_;
  wire _20071_;
  wire _20072_;
  wire _20073_;
  wire _20074_;
  wire _20075_;
  wire _20076_;
  wire _20077_;
  wire _20078_;
  wire _20079_;
  wire _20080_;
  wire _20081_;
  wire _20082_;
  wire _20083_;
  wire _20084_;
  wire _20085_;
  wire _20086_;
  wire _20087_;
  wire _20088_;
  wire _20089_;
  wire _20090_;
  wire _20091_;
  wire _20092_;
  wire _20093_;
  wire _20094_;
  wire _20095_;
  wire _20096_;
  wire _20097_;
  wire _20098_;
  wire _20099_;
  wire _20100_;
  wire _20101_;
  wire _20102_;
  wire _20103_;
  wire _20104_;
  wire _20105_;
  wire _20106_;
  wire _20107_;
  wire _20108_;
  wire _20109_;
  wire _20110_;
  wire _20111_;
  wire _20112_;
  wire _20113_;
  wire _20114_;
  wire _20115_;
  wire _20116_;
  wire _20117_;
  wire _20118_;
  wire _20119_;
  wire _20120_;
  wire _20121_;
  wire _20122_;
  wire _20123_;
  wire _20124_;
  wire _20125_;
  wire _20126_;
  wire _20127_;
  wire _20128_;
  wire _20129_;
  wire _20130_;
  wire _20131_;
  wire _20132_;
  wire _20133_;
  wire _20134_;
  wire _20135_;
  wire _20136_;
  wire _20137_;
  wire _20138_;
  wire _20139_;
  wire _20140_;
  wire _20141_;
  wire _20142_;
  wire _20143_;
  wire _20144_;
  wire _20145_;
  wire _20146_;
  wire _20147_;
  wire _20148_;
  wire _20149_;
  wire _20150_;
  wire _20151_;
  wire _20152_;
  wire _20153_;
  wire _20154_;
  wire _20155_;
  wire _20156_;
  wire _20157_;
  wire _20158_;
  wire _20159_;
  wire _20160_;
  wire _20161_;
  wire _20162_;
  wire _20163_;
  wire _20164_;
  wire _20165_;
  wire _20166_;
  wire _20167_;
  wire _20168_;
  wire _20169_;
  wire _20170_;
  wire _20171_;
  wire _20172_;
  wire _20173_;
  wire _20174_;
  wire _20175_;
  wire _20176_;
  wire _20177_;
  wire _20178_;
  wire _20179_;
  wire _20180_;
  wire _20181_;
  wire _20182_;
  wire _20183_;
  wire _20184_;
  wire _20185_;
  wire _20186_;
  wire _20187_;
  wire _20188_;
  wire _20189_;
  wire _20190_;
  wire _20191_;
  wire _20192_;
  wire _20193_;
  wire _20194_;
  wire _20195_;
  wire _20196_;
  wire _20197_;
  wire _20198_;
  wire _20199_;
  wire _20200_;
  wire _20201_;
  wire _20202_;
  wire _20203_;
  wire _20204_;
  wire _20205_;
  wire _20206_;
  wire _20207_;
  wire _20208_;
  wire _20209_;
  wire _20210_;
  wire _20211_;
  wire _20212_;
  wire _20213_;
  wire _20214_;
  wire _20215_;
  wire _20216_;
  wire _20217_;
  wire _20218_;
  wire _20219_;
  wire _20220_;
  wire _20221_;
  wire _20222_;
  wire _20223_;
  wire _20224_;
  wire _20225_;
  wire _20226_;
  wire _20227_;
  wire _20228_;
  wire _20229_;
  wire _20230_;
  wire _20231_;
  wire _20232_;
  wire _20233_;
  wire _20234_;
  wire _20235_;
  wire _20236_;
  wire _20237_;
  wire _20238_;
  wire _20239_;
  wire _20240_;
  wire _20241_;
  wire _20242_;
  wire _20243_;
  wire _20244_;
  wire _20245_;
  wire _20246_;
  wire _20247_;
  wire _20248_;
  wire _20249_;
  wire _20250_;
  wire _20251_;
  wire _20252_;
  wire _20253_;
  wire _20254_;
  wire _20255_;
  wire _20256_;
  wire _20257_;
  wire _20258_;
  wire _20259_;
  wire _20260_;
  wire _20261_;
  wire _20262_;
  wire _20263_;
  wire _20264_;
  wire _20265_;
  wire _20266_;
  wire _20267_;
  wire _20268_;
  wire _20269_;
  wire _20270_;
  wire _20271_;
  wire _20272_;
  wire _20273_;
  wire _20274_;
  wire _20275_;
  wire _20276_;
  wire _20277_;
  wire _20278_;
  wire _20279_;
  wire _20280_;
  wire _20281_;
  wire _20282_;
  wire _20283_;
  wire _20284_;
  wire _20285_;
  wire _20286_;
  wire _20287_;
  wire _20288_;
  wire _20289_;
  wire _20290_;
  wire _20291_;
  wire _20292_;
  wire _20293_;
  wire _20294_;
  wire _20295_;
  wire _20296_;
  wire _20297_;
  wire _20298_;
  wire _20299_;
  wire _20300_;
  wire _20301_;
  wire _20302_;
  wire _20303_;
  wire _20304_;
  wire _20305_;
  wire _20306_;
  wire _20307_;
  wire _20308_;
  wire _20309_;
  wire _20310_;
  wire _20311_;
  wire _20312_;
  wire _20313_;
  wire _20314_;
  wire _20315_;
  wire _20316_;
  wire _20317_;
  wire _20318_;
  wire _20319_;
  wire _20320_;
  wire _20321_;
  wire _20322_;
  wire _20323_;
  wire _20324_;
  wire _20325_;
  wire _20326_;
  wire _20327_;
  wire _20328_;
  wire _20329_;
  wire _20330_;
  wire _20331_;
  wire _20332_;
  wire _20333_;
  wire _20334_;
  wire _20335_;
  wire _20336_;
  wire _20337_;
  wire _20338_;
  wire _20339_;
  wire _20340_;
  wire _20341_;
  wire _20342_;
  wire _20343_;
  wire _20344_;
  wire _20345_;
  wire _20346_;
  wire _20347_;
  wire _20348_;
  wire _20349_;
  wire _20350_;
  wire _20351_;
  wire _20352_;
  wire _20353_;
  wire _20354_;
  wire _20355_;
  wire _20356_;
  wire _20357_;
  wire _20358_;
  wire _20359_;
  wire _20360_;
  wire _20361_;
  wire _20362_;
  wire _20363_;
  wire _20364_;
  wire _20365_;
  wire _20366_;
  wire _20367_;
  wire _20368_;
  wire _20369_;
  wire _20370_;
  wire _20371_;
  wire _20372_;
  wire _20373_;
  wire _20374_;
  wire _20375_;
  wire _20376_;
  wire _20377_;
  wire _20378_;
  wire _20379_;
  wire _20380_;
  wire _20381_;
  wire _20382_;
  wire _20383_;
  wire _20384_;
  wire _20385_;
  wire _20386_;
  wire _20387_;
  wire _20388_;
  wire _20389_;
  wire _20390_;
  wire _20391_;
  wire _20392_;
  wire _20393_;
  wire _20394_;
  wire _20395_;
  wire _20396_;
  wire _20397_;
  wire _20398_;
  wire _20399_;
  wire _20400_;
  wire _20401_;
  wire _20402_;
  wire _20403_;
  wire _20404_;
  wire _20405_;
  wire _20406_;
  wire _20407_;
  wire _20408_;
  wire _20409_;
  wire _20410_;
  wire _20411_;
  wire _20412_;
  wire _20413_;
  wire _20414_;
  wire _20415_;
  wire _20416_;
  wire _20417_;
  wire _20418_;
  wire _20419_;
  wire _20420_;
  wire _20421_;
  wire _20422_;
  wire _20423_;
  wire _20424_;
  wire _20425_;
  wire _20426_;
  wire _20427_;
  wire _20428_;
  wire _20429_;
  wire _20430_;
  wire _20431_;
  wire _20432_;
  wire _20433_;
  wire _20434_;
  wire _20435_;
  wire _20436_;
  wire _20437_;
  wire _20438_;
  wire _20439_;
  wire _20440_;
  wire _20441_;
  wire _20442_;
  wire _20443_;
  wire _20444_;
  wire _20445_;
  wire _20446_;
  wire _20447_;
  wire _20448_;
  wire _20449_;
  wire _20450_;
  wire _20451_;
  wire _20452_;
  wire _20453_;
  wire _20454_;
  wire _20455_;
  wire _20456_;
  wire _20457_;
  wire _20458_;
  wire _20459_;
  wire _20460_;
  wire _20461_;
  wire _20462_;
  wire _20463_;
  wire _20464_;
  wire _20465_;
  wire _20466_;
  wire _20467_;
  wire _20468_;
  wire _20469_;
  wire _20470_;
  wire _20471_;
  wire _20472_;
  wire _20473_;
  wire _20474_;
  wire _20475_;
  wire _20476_;
  wire _20477_;
  wire _20478_;
  wire _20479_;
  wire _20480_;
  wire _20481_;
  wire _20482_;
  wire _20483_;
  wire _20484_;
  wire _20485_;
  wire _20486_;
  wire _20487_;
  wire _20488_;
  wire _20489_;
  wire _20490_;
  wire _20491_;
  wire _20492_;
  wire _20493_;
  wire _20494_;
  wire _20495_;
  wire _20496_;
  wire _20497_;
  wire _20498_;
  wire _20499_;
  wire _20500_;
  wire _20501_;
  wire _20502_;
  wire _20503_;
  wire _20504_;
  wire _20505_;
  wire _20506_;
  wire _20507_;
  wire _20508_;
  wire _20509_;
  wire _20510_;
  wire _20511_;
  wire _20512_;
  wire _20513_;
  wire _20514_;
  wire _20515_;
  wire _20516_;
  wire _20517_;
  wire _20518_;
  wire _20519_;
  wire _20520_;
  wire _20521_;
  wire _20522_;
  wire _20523_;
  wire _20524_;
  wire _20525_;
  wire _20526_;
  wire _20527_;
  wire _20528_;
  wire _20529_;
  wire _20530_;
  wire _20531_;
  wire _20532_;
  wire _20533_;
  wire _20534_;
  wire _20535_;
  wire _20536_;
  wire _20537_;
  wire _20538_;
  wire _20539_;
  wire _20540_;
  wire _20541_;
  wire _20542_;
  wire _20543_;
  wire _20544_;
  wire _20545_;
  wire _20546_;
  wire _20547_;
  wire _20548_;
  wire _20549_;
  wire _20550_;
  wire _20551_;
  wire _20552_;
  wire _20553_;
  wire _20554_;
  wire _20555_;
  wire _20556_;
  wire _20557_;
  wire _20558_;
  wire _20559_;
  wire _20560_;
  wire _20561_;
  wire _20562_;
  wire _20563_;
  wire _20564_;
  wire _20565_;
  wire _20566_;
  wire _20567_;
  wire _20568_;
  wire _20569_;
  wire _20570_;
  wire _20571_;
  wire _20572_;
  wire _20573_;
  wire _20574_;
  wire _20575_;
  wire _20576_;
  wire _20577_;
  wire _20578_;
  wire _20579_;
  wire _20580_;
  wire _20581_;
  wire _20582_;
  wire _20583_;
  wire _20584_;
  wire _20585_;
  wire _20586_;
  wire _20587_;
  wire _20588_;
  wire _20589_;
  wire _20590_;
  wire _20591_;
  wire _20592_;
  wire _20593_;
  wire _20594_;
  wire _20595_;
  wire _20596_;
  wire _20597_;
  wire _20598_;
  wire _20599_;
  wire _20600_;
  wire _20601_;
  wire _20602_;
  wire _20603_;
  wire _20604_;
  wire _20605_;
  wire _20606_;
  wire _20607_;
  wire _20608_;
  wire _20609_;
  wire _20610_;
  wire _20611_;
  wire _20612_;
  wire _20613_;
  wire _20614_;
  wire _20615_;
  wire _20616_;
  wire _20617_;
  wire _20618_;
  wire _20619_;
  wire _20620_;
  wire _20621_;
  wire _20622_;
  wire _20623_;
  wire _20624_;
  wire _20625_;
  wire _20626_;
  wire _20627_;
  wire _20628_;
  wire _20629_;
  wire _20630_;
  wire _20631_;
  wire _20632_;
  wire _20633_;
  wire _20634_;
  wire _20635_;
  wire _20636_;
  wire _20637_;
  wire _20638_;
  wire _20639_;
  wire _20640_;
  wire _20641_;
  wire _20642_;
  wire _20643_;
  wire _20644_;
  wire _20645_;
  wire _20646_;
  wire _20647_;
  wire _20648_;
  wire _20649_;
  wire _20650_;
  wire _20651_;
  wire _20652_;
  wire _20653_;
  wire _20654_;
  wire _20655_;
  wire _20656_;
  wire _20657_;
  wire _20658_;
  wire _20659_;
  wire _20660_;
  wire _20661_;
  wire _20662_;
  wire _20663_;
  wire _20664_;
  wire _20665_;
  wire _20666_;
  wire _20667_;
  wire _20668_;
  wire _20669_;
  wire _20670_;
  wire _20671_;
  wire _20672_;
  wire _20673_;
  wire _20674_;
  wire _20675_;
  wire _20676_;
  wire _20677_;
  wire _20678_;
  wire _20679_;
  wire _20680_;
  wire _20681_;
  wire _20682_;
  wire _20683_;
  wire _20684_;
  wire _20685_;
  wire _20686_;
  wire _20687_;
  wire _20688_;
  wire _20689_;
  wire _20690_;
  wire _20691_;
  wire _20692_;
  wire _20693_;
  wire _20694_;
  wire _20695_;
  wire _20696_;
  wire _20697_;
  wire _20698_;
  wire _20699_;
  wire _20700_;
  wire _20701_;
  wire _20702_;
  wire _20703_;
  wire _20704_;
  wire _20705_;
  wire _20706_;
  wire _20707_;
  wire _20708_;
  wire _20709_;
  wire _20710_;
  wire _20711_;
  wire _20712_;
  wire _20713_;
  wire _20714_;
  wire _20715_;
  wire _20716_;
  wire _20717_;
  wire _20718_;
  wire _20719_;
  wire _20720_;
  wire _20721_;
  wire _20722_;
  wire _20723_;
  wire _20724_;
  wire _20725_;
  wire _20726_;
  wire _20727_;
  wire _20728_;
  wire _20729_;
  wire _20730_;
  wire _20731_;
  wire _20732_;
  wire _20733_;
  wire _20734_;
  wire _20735_;
  wire _20736_;
  wire _20737_;
  wire _20738_;
  wire _20739_;
  wire _20740_;
  wire _20741_;
  wire _20742_;
  wire _20743_;
  wire _20744_;
  wire _20745_;
  wire _20746_;
  wire _20747_;
  wire _20748_;
  wire _20749_;
  wire _20750_;
  wire _20751_;
  wire _20752_;
  wire _20753_;
  wire _20754_;
  wire _20755_;
  wire _20756_;
  wire _20757_;
  wire _20758_;
  wire _20759_;
  wire _20760_;
  wire _20761_;
  wire _20762_;
  wire _20763_;
  wire _20764_;
  wire _20765_;
  wire _20766_;
  wire _20767_;
  wire _20768_;
  wire _20769_;
  wire _20770_;
  wire _20771_;
  wire _20772_;
  wire _20773_;
  wire _20774_;
  wire _20775_;
  wire _20776_;
  wire _20777_;
  wire _20778_;
  wire _20779_;
  wire _20780_;
  wire _20781_;
  wire _20782_;
  wire _20783_;
  wire _20784_;
  wire _20785_;
  wire _20786_;
  wire _20787_;
  wire _20788_;
  wire _20789_;
  wire _20790_;
  wire _20791_;
  wire _20792_;
  wire _20793_;
  wire _20794_;
  wire _20795_;
  wire _20796_;
  wire _20797_;
  wire _20798_;
  wire _20799_;
  wire _20800_;
  wire _20801_;
  wire _20802_;
  wire _20803_;
  wire _20804_;
  wire _20805_;
  wire _20806_;
  wire _20807_;
  wire _20808_;
  wire _20809_;
  wire _20810_;
  wire _20811_;
  wire _20812_;
  wire _20813_;
  wire _20814_;
  wire _20815_;
  wire _20816_;
  wire _20817_;
  wire _20818_;
  wire _20819_;
  wire _20820_;
  wire _20821_;
  wire _20822_;
  wire _20823_;
  wire _20824_;
  wire _20825_;
  wire _20826_;
  wire _20827_;
  wire _20828_;
  wire _20829_;
  wire _20830_;
  wire _20831_;
  wire _20832_;
  wire _20833_;
  wire _20834_;
  wire _20835_;
  wire _20836_;
  wire _20837_;
  wire _20838_;
  wire _20839_;
  wire _20840_;
  wire _20841_;
  wire _20842_;
  wire _20843_;
  wire _20844_;
  wire _20845_;
  wire _20846_;
  wire _20847_;
  wire _20848_;
  wire _20849_;
  wire _20850_;
  wire _20851_;
  wire _20852_;
  wire _20853_;
  wire _20854_;
  wire _20855_;
  wire _20856_;
  wire _20857_;
  wire _20858_;
  wire _20859_;
  wire _20860_;
  wire _20861_;
  wire _20862_;
  wire _20863_;
  wire _20864_;
  wire _20865_;
  wire _20866_;
  wire _20867_;
  wire _20868_;
  wire _20869_;
  wire _20870_;
  wire _20871_;
  wire _20872_;
  wire _20873_;
  wire _20874_;
  wire _20875_;
  wire _20876_;
  wire _20877_;
  wire _20878_;
  wire _20879_;
  wire _20880_;
  wire _20881_;
  wire _20882_;
  wire _20883_;
  wire _20884_;
  wire _20885_;
  wire _20886_;
  wire _20887_;
  wire _20888_;
  wire _20889_;
  wire _20890_;
  wire _20891_;
  wire _20892_;
  wire _20893_;
  wire _20894_;
  wire _20895_;
  wire _20896_;
  wire _20897_;
  wire _20898_;
  wire _20899_;
  wire _20900_;
  wire _20901_;
  wire _20902_;
  wire _20903_;
  wire _20904_;
  wire _20905_;
  wire _20906_;
  wire _20907_;
  wire _20908_;
  wire _20909_;
  wire _20910_;
  wire _20911_;
  wire _20912_;
  wire _20913_;
  wire _20914_;
  wire _20915_;
  wire _20916_;
  wire _20917_;
  wire _20918_;
  wire _20919_;
  wire _20920_;
  wire _20921_;
  wire _20922_;
  wire _20923_;
  wire _20924_;
  wire _20925_;
  wire _20926_;
  wire _20927_;
  wire _20928_;
  wire _20929_;
  wire _20930_;
  wire _20931_;
  wire _20932_;
  wire _20933_;
  wire _20934_;
  wire _20935_;
  wire _20936_;
  wire _20937_;
  wire _20938_;
  wire _20939_;
  wire _20940_;
  wire _20941_;
  wire _20942_;
  wire _20943_;
  wire _20944_;
  wire _20945_;
  wire _20946_;
  wire _20947_;
  wire _20948_;
  wire _20949_;
  wire _20950_;
  wire _20951_;
  wire _20952_;
  wire _20953_;
  wire _20954_;
  wire _20955_;
  wire _20956_;
  wire _20957_;
  wire _20958_;
  wire _20959_;
  wire _20960_;
  wire _20961_;
  wire _20962_;
  wire _20963_;
  wire _20964_;
  wire _20965_;
  wire _20966_;
  wire _20967_;
  wire _20968_;
  wire _20969_;
  wire _20970_;
  wire _20971_;
  wire _20972_;
  wire _20973_;
  wire _20974_;
  wire _20975_;
  wire _20976_;
  wire _20977_;
  wire _20978_;
  wire _20979_;
  wire _20980_;
  wire _20981_;
  wire _20982_;
  wire _20983_;
  wire _20984_;
  wire _20985_;
  wire _20986_;
  wire _20987_;
  wire _20988_;
  wire _20989_;
  wire _20990_;
  wire _20991_;
  wire _20992_;
  wire _20993_;
  wire _20994_;
  wire _20995_;
  wire _20996_;
  wire _20997_;
  wire _20998_;
  wire _20999_;
  wire _21000_;
  wire _21001_;
  wire _21002_;
  wire _21003_;
  wire _21004_;
  wire _21005_;
  wire _21006_;
  wire _21007_;
  wire _21008_;
  wire _21009_;
  wire _21010_;
  wire _21011_;
  wire _21012_;
  wire _21013_;
  wire _21014_;
  wire _21015_;
  wire _21016_;
  wire _21017_;
  wire _21018_;
  wire _21019_;
  wire _21020_;
  wire _21021_;
  wire _21022_;
  wire _21023_;
  wire _21024_;
  wire _21025_;
  wire _21026_;
  wire _21027_;
  wire _21028_;
  wire _21029_;
  wire _21030_;
  wire _21031_;
  wire _21032_;
  wire _21033_;
  wire _21034_;
  wire _21035_;
  wire _21036_;
  wire _21037_;
  wire _21038_;
  wire _21039_;
  wire _21040_;
  wire _21041_;
  wire _21042_;
  wire _21043_;
  wire _21044_;
  wire _21045_;
  wire _21046_;
  wire _21047_;
  wire _21048_;
  wire _21049_;
  wire _21050_;
  wire _21051_;
  wire _21052_;
  wire _21053_;
  wire _21054_;
  wire _21055_;
  wire _21056_;
  wire _21057_;
  wire _21058_;
  wire _21059_;
  wire _21060_;
  wire _21061_;
  wire _21062_;
  wire _21063_;
  wire _21064_;
  wire _21065_;
  wire _21066_;
  wire _21067_;
  wire _21068_;
  wire _21069_;
  wire _21070_;
  wire _21071_;
  wire _21072_;
  wire _21073_;
  wire _21074_;
  wire _21075_;
  wire _21076_;
  wire _21077_;
  wire _21078_;
  wire _21079_;
  wire _21080_;
  wire _21081_;
  wire _21082_;
  wire _21083_;
  wire _21084_;
  wire _21085_;
  wire _21086_;
  wire _21087_;
  wire _21088_;
  wire _21089_;
  wire _21090_;
  wire _21091_;
  wire _21092_;
  wire _21093_;
  wire _21094_;
  wire _21095_;
  wire _21096_;
  wire _21097_;
  wire _21098_;
  wire _21099_;
  wire _21100_;
  wire _21101_;
  wire _21102_;
  wire _21103_;
  wire _21104_;
  wire _21105_;
  wire _21106_;
  wire _21107_;
  wire _21108_;
  wire _21109_;
  wire _21110_;
  wire _21111_;
  wire _21112_;
  wire _21113_;
  wire _21114_;
  wire _21115_;
  wire _21116_;
  wire _21117_;
  wire _21118_;
  wire _21119_;
  wire _21120_;
  wire _21121_;
  wire _21122_;
  wire _21123_;
  wire _21124_;
  wire _21125_;
  wire _21126_;
  wire _21127_;
  wire _21128_;
  wire _21129_;
  wire _21130_;
  wire _21131_;
  wire _21132_;
  wire _21133_;
  wire _21134_;
  wire _21135_;
  wire _21136_;
  wire _21137_;
  wire _21138_;
  wire _21139_;
  wire _21140_;
  wire _21141_;
  wire _21142_;
  wire _21143_;
  wire _21144_;
  wire _21145_;
  wire _21146_;
  wire _21147_;
  wire _21148_;
  wire _21149_;
  wire _21150_;
  wire _21151_;
  wire _21152_;
  wire _21153_;
  wire _21154_;
  wire _21155_;
  wire _21156_;
  wire _21157_;
  wire _21158_;
  wire _21159_;
  wire _21160_;
  wire _21161_;
  wire _21162_;
  wire _21163_;
  wire _21164_;
  wire _21165_;
  wire _21166_;
  wire _21167_;
  wire _21168_;
  wire _21169_;
  wire _21170_;
  wire _21171_;
  wire _21172_;
  wire _21173_;
  wire _21174_;
  wire _21175_;
  wire _21176_;
  wire _21177_;
  wire _21178_;
  wire _21179_;
  wire _21180_;
  wire _21181_;
  wire _21182_;
  wire _21183_;
  wire _21184_;
  wire _21185_;
  wire _21186_;
  wire _21187_;
  wire _21188_;
  wire _21189_;
  wire _21190_;
  wire _21191_;
  wire _21192_;
  wire _21193_;
  wire _21194_;
  wire _21195_;
  wire _21196_;
  wire _21197_;
  wire _21198_;
  wire _21199_;
  wire _21200_;
  wire _21201_;
  wire _21202_;
  wire _21203_;
  wire _21204_;
  wire _21205_;
  wire _21206_;
  wire _21207_;
  wire _21208_;
  wire _21209_;
  wire _21210_;
  wire _21211_;
  wire _21212_;
  wire _21213_;
  wire _21214_;
  wire _21215_;
  wire _21216_;
  wire _21217_;
  wire _21218_;
  wire _21219_;
  wire _21220_;
  wire _21221_;
  wire _21222_;
  wire _21223_;
  wire _21224_;
  wire _21225_;
  wire _21226_;
  wire _21227_;
  wire _21228_;
  wire _21229_;
  wire _21230_;
  wire _21231_;
  wire _21232_;
  wire _21233_;
  wire _21234_;
  wire _21235_;
  wire _21236_;
  wire _21237_;
  wire _21238_;
  wire _21239_;
  wire _21240_;
  wire _21241_;
  wire _21242_;
  wire _21243_;
  wire _21244_;
  wire _21245_;
  wire _21246_;
  wire _21247_;
  wire _21248_;
  wire _21249_;
  wire _21250_;
  wire _21251_;
  wire _21252_;
  wire _21253_;
  wire _21254_;
  wire _21255_;
  wire _21256_;
  wire _21257_;
  wire _21258_;
  wire _21259_;
  wire _21260_;
  wire _21261_;
  wire _21262_;
  wire _21263_;
  wire _21264_;
  wire _21265_;
  wire _21266_;
  wire _21267_;
  wire _21268_;
  wire _21269_;
  wire _21270_;
  wire _21271_;
  wire _21272_;
  wire _21273_;
  wire _21274_;
  wire _21275_;
  wire _21276_;
  wire _21277_;
  wire _21278_;
  wire _21279_;
  wire _21280_;
  wire _21281_;
  wire _21282_;
  wire _21283_;
  wire _21284_;
  wire _21285_;
  wire _21286_;
  wire _21287_;
  wire _21288_;
  wire _21289_;
  wire _21290_;
  wire _21291_;
  wire _21292_;
  wire _21293_;
  wire _21294_;
  wire _21295_;
  wire _21296_;
  wire _21297_;
  wire _21298_;
  wire _21299_;
  wire _21300_;
  wire _21301_;
  wire _21302_;
  wire _21303_;
  wire _21304_;
  wire _21305_;
  wire _21306_;
  wire _21307_;
  wire _21308_;
  wire _21309_;
  wire _21310_;
  wire _21311_;
  wire _21312_;
  wire _21313_;
  wire _21314_;
  wire _21315_;
  wire _21316_;
  wire _21317_;
  wire _21318_;
  wire _21319_;
  wire _21320_;
  wire _21321_;
  wire _21322_;
  wire _21323_;
  wire _21324_;
  wire _21325_;
  wire _21326_;
  wire _21327_;
  wire _21328_;
  wire _21329_;
  wire _21330_;
  wire _21331_;
  wire _21332_;
  wire _21333_;
  wire _21334_;
  wire _21335_;
  wire _21336_;
  wire _21337_;
  wire _21338_;
  wire _21339_;
  wire _21340_;
  wire _21341_;
  wire _21342_;
  wire _21343_;
  wire _21344_;
  wire _21345_;
  wire _21346_;
  wire _21347_;
  wire _21348_;
  wire _21349_;
  wire _21350_;
  wire _21351_;
  wire _21352_;
  wire _21353_;
  wire _21354_;
  wire _21355_;
  wire _21356_;
  wire _21357_;
  wire _21358_;
  wire _21359_;
  wire _21360_;
  wire _21361_;
  wire _21362_;
  wire _21363_;
  wire _21364_;
  wire _21365_;
  wire _21366_;
  wire _21367_;
  wire _21368_;
  wire _21369_;
  wire _21370_;
  wire _21371_;
  wire _21372_;
  wire _21373_;
  wire _21374_;
  wire _21375_;
  wire _21376_;
  wire _21377_;
  wire _21378_;
  wire _21379_;
  wire _21380_;
  wire _21381_;
  wire _21382_;
  wire _21383_;
  wire _21384_;
  wire _21385_;
  wire _21386_;
  wire _21387_;
  wire _21388_;
  wire _21389_;
  wire _21390_;
  wire _21391_;
  wire _21392_;
  wire _21393_;
  wire _21394_;
  wire _21395_;
  wire _21396_;
  wire _21397_;
  wire _21398_;
  wire _21399_;
  wire _21400_;
  wire _21401_;
  wire _21402_;
  wire _21403_;
  wire _21404_;
  wire _21405_;
  wire _21406_;
  wire _21407_;
  wire _21408_;
  wire _21409_;
  wire _21410_;
  wire _21411_;
  wire _21412_;
  wire _21413_;
  wire _21414_;
  wire _21415_;
  wire _21416_;
  wire _21417_;
  wire _21418_;
  wire _21419_;
  wire _21420_;
  wire _21421_;
  wire _21422_;
  wire _21423_;
  wire _21424_;
  wire _21425_;
  wire _21426_;
  wire _21427_;
  wire _21428_;
  wire _21429_;
  wire _21430_;
  wire _21431_;
  wire _21432_;
  wire _21433_;
  wire _21434_;
  wire _21435_;
  wire _21436_;
  wire _21437_;
  wire _21438_;
  wire _21439_;
  wire _21440_;
  wire _21441_;
  wire _21442_;
  wire _21443_;
  wire _21444_;
  wire _21445_;
  wire _21446_;
  wire _21447_;
  wire _21448_;
  wire _21449_;
  wire _21450_;
  wire _21451_;
  wire _21452_;
  wire _21453_;
  wire _21454_;
  wire _21455_;
  wire _21456_;
  wire _21457_;
  wire _21458_;
  wire _21459_;
  wire _21460_;
  wire _21461_;
  wire _21462_;
  wire _21463_;
  wire _21464_;
  wire _21465_;
  wire _21466_;
  wire _21467_;
  wire _21468_;
  wire _21469_;
  wire _21470_;
  wire _21471_;
  wire _21472_;
  wire _21473_;
  wire _21474_;
  wire _21475_;
  wire _21476_;
  wire _21477_;
  wire _21478_;
  wire _21479_;
  wire _21480_;
  wire _21481_;
  wire _21482_;
  wire _21483_;
  wire _21484_;
  wire _21485_;
  wire _21486_;
  wire _21487_;
  wire _21488_;
  wire _21489_;
  wire _21490_;
  wire _21491_;
  wire _21492_;
  wire _21493_;
  wire _21494_;
  wire _21495_;
  wire _21496_;
  wire _21497_;
  wire _21498_;
  wire _21499_;
  wire _21500_;
  wire _21501_;
  wire _21502_;
  wire _21503_;
  wire _21504_;
  wire _21505_;
  wire _21506_;
  wire _21507_;
  wire _21508_;
  wire _21509_;
  wire _21510_;
  wire _21511_;
  wire _21512_;
  wire _21513_;
  wire _21514_;
  wire _21515_;
  wire _21516_;
  wire _21517_;
  wire _21518_;
  wire _21519_;
  wire _21520_;
  wire _21521_;
  wire _21522_;
  wire _21523_;
  wire _21524_;
  wire _21525_;
  wire _21526_;
  wire _21527_;
  wire _21528_;
  wire _21529_;
  wire _21530_;
  wire _21531_;
  wire _21532_;
  wire _21533_;
  wire _21534_;
  wire _21535_;
  wire _21536_;
  wire _21537_;
  wire _21538_;
  wire _21539_;
  wire _21540_;
  wire _21541_;
  wire _21542_;
  wire _21543_;
  wire _21544_;
  wire _21545_;
  wire _21546_;
  wire _21547_;
  wire _21548_;
  wire _21549_;
  wire _21550_;
  wire _21551_;
  wire _21552_;
  wire _21553_;
  wire _21554_;
  wire _21555_;
  wire _21556_;
  wire _21557_;
  wire _21558_;
  wire _21559_;
  wire _21560_;
  wire _21561_;
  wire _21562_;
  wire _21563_;
  wire _21564_;
  wire _21565_;
  wire _21566_;
  wire _21567_;
  wire _21568_;
  wire _21569_;
  wire _21570_;
  wire _21571_;
  wire _21572_;
  wire _21573_;
  wire _21574_;
  wire _21575_;
  wire _21576_;
  wire _21577_;
  wire _21578_;
  wire _21579_;
  wire _21580_;
  wire _21581_;
  wire _21582_;
  wire _21583_;
  wire _21584_;
  wire _21585_;
  wire _21586_;
  wire _21587_;
  wire _21588_;
  wire _21589_;
  wire _21590_;
  wire _21591_;
  wire _21592_;
  wire _21593_;
  wire _21594_;
  wire _21595_;
  wire _21596_;
  wire _21597_;
  wire _21598_;
  wire _21599_;
  wire _21600_;
  wire _21601_;
  wire _21602_;
  wire _21603_;
  wire _21604_;
  wire _21605_;
  wire _21606_;
  wire _21607_;
  wire _21608_;
  wire _21609_;
  wire _21610_;
  wire _21611_;
  wire _21612_;
  wire _21613_;
  wire _21614_;
  wire _21615_;
  wire _21616_;
  wire _21617_;
  wire _21618_;
  wire _21619_;
  wire _21620_;
  wire _21621_;
  wire _21622_;
  wire _21623_;
  wire _21624_;
  wire _21625_;
  wire _21626_;
  wire _21627_;
  wire _21628_;
  wire _21629_;
  wire _21630_;
  wire _21631_;
  wire _21632_;
  wire _21633_;
  wire _21634_;
  wire _21635_;
  wire _21636_;
  wire _21637_;
  wire _21638_;
  wire _21639_;
  wire _21640_;
  wire _21641_;
  wire _21642_;
  wire _21643_;
  wire _21644_;
  wire _21645_;
  wire _21646_;
  wire _21647_;
  wire _21648_;
  wire _21649_;
  wire _21650_;
  wire _21651_;
  wire _21652_;
  wire _21653_;
  wire _21654_;
  wire _21655_;
  wire _21656_;
  wire _21657_;
  wire _21658_;
  wire _21659_;
  wire _21660_;
  wire _21661_;
  wire _21662_;
  wire _21663_;
  wire _21664_;
  wire _21665_;
  wire _21666_;
  wire _21667_;
  wire _21668_;
  wire _21669_;
  wire _21670_;
  wire _21671_;
  wire _21672_;
  wire _21673_;
  wire _21674_;
  wire _21675_;
  wire _21676_;
  wire _21677_;
  wire _21678_;
  wire _21679_;
  wire _21680_;
  wire _21681_;
  wire _21682_;
  wire _21683_;
  wire _21684_;
  wire _21685_;
  wire _21686_;
  wire _21687_;
  wire _21688_;
  wire _21689_;
  wire _21690_;
  wire _21691_;
  wire _21692_;
  wire _21693_;
  wire _21694_;
  wire _21695_;
  wire _21696_;
  wire _21697_;
  wire _21698_;
  wire _21699_;
  wire _21700_;
  wire _21701_;
  wire _21702_;
  wire _21703_;
  wire _21704_;
  wire _21705_;
  wire _21706_;
  wire _21707_;
  wire _21708_;
  wire _21709_;
  wire _21710_;
  wire _21711_;
  wire _21712_;
  wire _21713_;
  wire _21714_;
  wire _21715_;
  wire _21716_;
  wire _21717_;
  wire _21718_;
  wire _21719_;
  wire _21720_;
  wire _21721_;
  wire _21722_;
  wire _21723_;
  wire _21724_;
  wire _21725_;
  wire _21726_;
  wire _21727_;
  wire _21728_;
  wire _21729_;
  wire _21730_;
  wire _21731_;
  wire _21732_;
  wire _21733_;
  wire _21734_;
  wire _21735_;
  wire _21736_;
  wire _21737_;
  wire _21738_;
  wire _21739_;
  wire _21740_;
  wire _21741_;
  wire _21742_;
  wire _21743_;
  wire _21744_;
  wire _21745_;
  wire _21746_;
  wire _21747_;
  wire _21748_;
  wire _21749_;
  wire _21750_;
  wire _21751_;
  wire _21752_;
  wire _21753_;
  wire _21754_;
  wire _21755_;
  wire _21756_;
  wire _21757_;
  wire _21758_;
  wire _21759_;
  wire _21760_;
  wire _21761_;
  wire _21762_;
  wire _21763_;
  wire _21764_;
  wire _21765_;
  wire _21766_;
  wire _21767_;
  wire _21768_;
  wire _21769_;
  wire _21770_;
  wire _21771_;
  wire _21772_;
  wire _21773_;
  wire _21774_;
  wire _21775_;
  wire _21776_;
  wire _21777_;
  wire _21778_;
  wire _21779_;
  wire _21780_;
  wire _21781_;
  wire _21782_;
  wire _21783_;
  wire _21784_;
  wire _21785_;
  wire _21786_;
  wire _21787_;
  wire _21788_;
  wire _21789_;
  wire _21790_;
  wire _21791_;
  wire _21792_;
  wire _21793_;
  wire _21794_;
  wire _21795_;
  wire _21796_;
  wire _21797_;
  wire _21798_;
  wire _21799_;
  wire _21800_;
  wire _21801_;
  wire _21802_;
  wire _21803_;
  wire _21804_;
  wire _21805_;
  wire _21806_;
  wire _21807_;
  wire _21808_;
  wire _21809_;
  wire _21810_;
  wire _21811_;
  wire _21812_;
  wire _21813_;
  wire _21814_;
  wire _21815_;
  wire _21816_;
  wire _21817_;
  wire _21818_;
  wire _21819_;
  wire _21820_;
  wire _21821_;
  wire _21822_;
  wire _21823_;
  wire _21824_;
  wire _21825_;
  wire _21826_;
  wire _21827_;
  wire _21828_;
  wire _21829_;
  wire _21830_;
  wire _21831_;
  wire _21832_;
  wire _21833_;
  wire _21834_;
  wire _21835_;
  wire _21836_;
  wire _21837_;
  wire _21838_;
  wire _21839_;
  wire _21840_;
  wire _21841_;
  wire _21842_;
  wire _21843_;
  wire _21844_;
  wire _21845_;
  wire _21846_;
  wire _21847_;
  wire _21848_;
  wire _21849_;
  wire _21850_;
  wire _21851_;
  wire _21852_;
  wire _21853_;
  wire _21854_;
  wire _21855_;
  wire _21856_;
  wire _21857_;
  wire _21858_;
  wire _21859_;
  wire _21860_;
  wire _21861_;
  wire _21862_;
  wire _21863_;
  wire _21864_;
  wire _21865_;
  wire _21866_;
  wire _21867_;
  wire _21868_;
  wire _21869_;
  wire _21870_;
  wire _21871_;
  wire _21872_;
  wire _21873_;
  wire _21874_;
  wire _21875_;
  wire _21876_;
  wire _21877_;
  wire _21878_;
  wire _21879_;
  wire _21880_;
  wire _21881_;
  wire _21882_;
  wire _21883_;
  wire _21884_;
  wire _21885_;
  wire _21886_;
  wire _21887_;
  wire _21888_;
  wire _21889_;
  wire _21890_;
  wire _21891_;
  wire _21892_;
  wire _21893_;
  wire _21894_;
  wire _21895_;
  wire _21896_;
  wire _21897_;
  wire _21898_;
  wire _21899_;
  wire _21900_;
  wire _21901_;
  wire _21902_;
  wire _21903_;
  wire _21904_;
  wire _21905_;
  wire _21906_;
  wire _21907_;
  wire _21908_;
  wire _21909_;
  wire _21910_;
  wire _21911_;
  wire _21912_;
  wire _21913_;
  wire _21914_;
  wire _21915_;
  wire _21916_;
  wire _21917_;
  wire _21918_;
  wire _21919_;
  wire _21920_;
  wire _21921_;
  wire _21922_;
  wire _21923_;
  wire _21924_;
  wire _21925_;
  wire _21926_;
  wire _21927_;
  wire _21928_;
  wire _21929_;
  wire _21930_;
  wire _21931_;
  wire _21932_;
  wire _21933_;
  wire _21934_;
  wire _21935_;
  wire _21936_;
  wire _21937_;
  wire _21938_;
  wire _21939_;
  wire _21940_;
  wire _21941_;
  wire _21942_;
  wire _21943_;
  wire _21944_;
  wire _21945_;
  wire _21946_;
  wire _21947_;
  wire _21948_;
  wire _21949_;
  wire _21950_;
  wire _21951_;
  wire _21952_;
  wire _21953_;
  wire _21954_;
  wire _21955_;
  wire _21956_;
  wire _21957_;
  wire _21958_;
  wire _21959_;
  wire _21960_;
  wire _21961_;
  wire _21962_;
  wire _21963_;
  wire _21964_;
  wire _21965_;
  wire _21966_;
  wire _21967_;
  wire _21968_;
  wire _21969_;
  wire _21970_;
  wire _21971_;
  wire _21972_;
  wire _21973_;
  wire _21974_;
  wire _21975_;
  wire _21976_;
  wire _21977_;
  wire _21978_;
  wire _21979_;
  wire _21980_;
  wire _21981_;
  wire _21982_;
  wire _21983_;
  wire _21984_;
  wire _21985_;
  wire _21986_;
  wire _21987_;
  wire _21988_;
  wire _21989_;
  wire _21990_;
  wire _21991_;
  wire _21992_;
  wire _21993_;
  wire _21994_;
  wire _21995_;
  wire _21996_;
  wire _21997_;
  wire _21998_;
  wire _21999_;
  wire _22000_;
  wire _22001_;
  wire _22002_;
  wire _22003_;
  wire _22004_;
  wire _22005_;
  wire _22006_;
  wire _22007_;
  wire _22008_;
  wire _22009_;
  wire _22010_;
  wire _22011_;
  wire _22012_;
  wire _22013_;
  wire _22014_;
  wire _22015_;
  wire _22016_;
  wire _22017_;
  wire _22018_;
  wire _22019_;
  wire _22020_;
  wire _22021_;
  wire _22022_;
  wire _22023_;
  wire _22024_;
  wire _22025_;
  wire _22026_;
  wire _22027_;
  wire _22028_;
  wire _22029_;
  wire _22030_;
  wire _22031_;
  wire _22032_;
  wire _22033_;
  wire _22034_;
  wire _22035_;
  wire _22036_;
  wire _22037_;
  wire _22038_;
  wire _22039_;
  wire _22040_;
  wire _22041_;
  wire _22042_;
  wire _22043_;
  wire _22044_;
  wire _22045_;
  wire _22046_;
  wire _22047_;
  wire _22048_;
  wire _22049_;
  wire _22050_;
  wire _22051_;
  wire _22052_;
  wire _22053_;
  wire _22054_;
  wire _22055_;
  wire _22056_;
  wire _22057_;
  wire _22058_;
  wire _22059_;
  wire _22060_;
  wire _22061_;
  wire _22062_;
  wire _22063_;
  wire _22064_;
  wire _22065_;
  wire _22066_;
  wire _22067_;
  wire _22068_;
  wire _22069_;
  wire _22070_;
  wire _22071_;
  wire _22072_;
  wire _22073_;
  wire _22074_;
  wire _22075_;
  wire _22076_;
  wire _22077_;
  wire _22078_;
  wire _22079_;
  wire _22080_;
  wire _22081_;
  wire _22082_;
  wire _22083_;
  wire _22084_;
  wire _22085_;
  wire _22086_;
  wire _22087_;
  wire _22088_;
  wire _22089_;
  wire _22090_;
  wire _22091_;
  wire _22092_;
  wire _22093_;
  wire _22094_;
  wire _22095_;
  wire _22096_;
  wire _22097_;
  wire _22098_;
  wire _22099_;
  wire _22100_;
  wire _22101_;
  wire _22102_;
  wire _22103_;
  wire _22104_;
  wire _22105_;
  wire _22106_;
  wire _22107_;
  wire _22108_;
  wire _22109_;
  wire _22110_;
  wire _22111_;
  wire _22112_;
  wire _22113_;
  wire _22114_;
  wire _22115_;
  wire _22116_;
  wire _22117_;
  wire _22118_;
  wire _22119_;
  wire _22120_;
  wire _22121_;
  wire _22122_;
  wire _22123_;
  wire _22124_;
  wire _22125_;
  wire _22126_;
  wire _22127_;
  wire _22128_;
  wire _22129_;
  wire _22130_;
  wire _22131_;
  wire _22132_;
  wire _22133_;
  wire _22134_;
  wire _22135_;
  wire _22136_;
  wire _22137_;
  wire _22138_;
  wire _22139_;
  wire _22140_;
  wire _22141_;
  wire _22142_;
  wire _22143_;
  wire _22144_;
  wire _22145_;
  wire _22146_;
  wire _22147_;
  wire _22148_;
  wire _22149_;
  wire _22150_;
  wire _22151_;
  wire _22152_;
  wire _22153_;
  wire _22154_;
  wire _22155_;
  wire _22156_;
  wire _22157_;
  wire _22158_;
  wire _22159_;
  wire _22160_;
  wire _22161_;
  wire _22162_;
  wire _22163_;
  wire _22164_;
  wire _22165_;
  wire _22166_;
  wire _22167_;
  wire _22168_;
  wire _22169_;
  wire _22170_;
  wire _22171_;
  wire _22172_;
  wire _22173_;
  wire _22174_;
  wire _22175_;
  wire _22176_;
  wire _22177_;
  wire _22178_;
  wire _22179_;
  wire _22180_;
  wire _22181_;
  wire _22182_;
  wire _22183_;
  wire _22184_;
  wire _22185_;
  wire _22186_;
  wire _22187_;
  wire _22188_;
  wire _22189_;
  wire _22190_;
  wire _22191_;
  wire _22192_;
  wire _22193_;
  wire _22194_;
  wire _22195_;
  wire _22196_;
  wire _22197_;
  wire _22198_;
  wire _22199_;
  wire _22200_;
  wire _22201_;
  wire _22202_;
  wire _22203_;
  wire _22204_;
  wire _22205_;
  wire _22206_;
  wire _22207_;
  wire _22208_;
  wire _22209_;
  wire _22210_;
  wire _22211_;
  wire _22212_;
  wire _22213_;
  wire _22214_;
  wire _22215_;
  wire _22216_;
  wire _22217_;
  wire _22218_;
  wire _22219_;
  wire _22220_;
  wire _22221_;
  wire _22222_;
  wire _22223_;
  wire _22224_;
  wire _22225_;
  wire _22226_;
  wire _22227_;
  wire _22228_;
  wire _22229_;
  wire _22230_;
  wire _22231_;
  wire _22232_;
  wire _22233_;
  wire _22234_;
  wire _22235_;
  wire _22236_;
  wire _22237_;
  wire _22238_;
  wire _22239_;
  wire _22240_;
  wire _22241_;
  wire _22242_;
  wire _22243_;
  wire _22244_;
  wire _22245_;
  wire _22246_;
  wire _22247_;
  wire _22248_;
  wire _22249_;
  wire _22250_;
  wire _22251_;
  wire _22252_;
  wire _22253_;
  wire _22254_;
  wire _22255_;
  wire _22256_;
  wire _22257_;
  wire _22258_;
  wire _22259_;
  wire _22260_;
  wire _22261_;
  wire _22262_;
  wire _22263_;
  wire _22264_;
  wire _22265_;
  wire _22266_;
  wire _22267_;
  wire _22268_;
  wire _22269_;
  wire _22270_;
  wire _22271_;
  wire _22272_;
  wire _22273_;
  wire _22274_;
  wire _22275_;
  wire _22276_;
  wire _22277_;
  wire _22278_;
  wire _22279_;
  wire _22280_;
  wire _22281_;
  wire _22282_;
  wire _22283_;
  wire _22284_;
  wire _22285_;
  wire _22286_;
  wire _22287_;
  wire _22288_;
  wire _22289_;
  wire _22290_;
  wire _22291_;
  wire _22292_;
  wire _22293_;
  wire _22294_;
  wire _22295_;
  wire _22296_;
  wire _22297_;
  wire _22298_;
  wire _22299_;
  wire _22300_;
  wire _22301_;
  wire _22302_;
  wire _22303_;
  wire _22304_;
  wire _22305_;
  wire _22306_;
  wire _22307_;
  wire _22308_;
  wire _22309_;
  wire _22310_;
  wire _22311_;
  wire _22312_;
  wire _22313_;
  wire _22314_;
  wire _22315_;
  wire _22316_;
  wire _22317_;
  wire _22318_;
  wire _22319_;
  wire _22320_;
  wire _22321_;
  wire _22322_;
  wire _22323_;
  wire _22324_;
  wire _22325_;
  wire _22326_;
  wire _22327_;
  wire _22328_;
  wire _22329_;
  wire _22330_;
  wire _22331_;
  wire _22332_;
  wire _22333_;
  wire _22334_;
  wire _22335_;
  wire _22336_;
  wire _22337_;
  wire _22338_;
  wire _22339_;
  wire _22340_;
  wire _22341_;
  wire _22342_;
  wire _22343_;
  wire _22344_;
  wire _22345_;
  wire _22346_;
  wire _22347_;
  wire _22348_;
  wire _22349_;
  wire _22350_;
  wire _22351_;
  wire _22352_;
  wire _22353_;
  wire _22354_;
  wire _22355_;
  wire _22356_;
  wire _22357_;
  wire _22358_;
  wire _22359_;
  wire _22360_;
  wire _22361_;
  wire _22362_;
  wire _22363_;
  wire _22364_;
  wire _22365_;
  wire _22366_;
  wire _22367_;
  wire _22368_;
  wire _22369_;
  wire _22370_;
  wire _22371_;
  wire _22372_;
  wire _22373_;
  wire _22374_;
  wire _22375_;
  wire _22376_;
  wire _22377_;
  wire _22378_;
  wire _22379_;
  wire _22380_;
  wire _22381_;
  wire _22382_;
  wire _22383_;
  wire _22384_;
  wire _22385_;
  wire _22386_;
  wire _22387_;
  wire _22388_;
  wire _22389_;
  wire _22390_;
  wire _22391_;
  wire _22392_;
  wire _22393_;
  wire _22394_;
  wire _22395_;
  wire _22396_;
  wire _22397_;
  wire _22398_;
  wire _22399_;
  wire _22400_;
  wire _22401_;
  wire _22402_;
  wire _22403_;
  wire _22404_;
  wire _22405_;
  wire _22406_;
  wire _22407_;
  wire _22408_;
  wire _22409_;
  wire _22410_;
  wire _22411_;
  wire _22412_;
  wire _22413_;
  wire _22414_;
  wire _22415_;
  wire _22416_;
  wire _22417_;
  wire _22418_;
  wire _22419_;
  wire _22420_;
  wire _22421_;
  wire _22422_;
  wire _22423_;
  wire _22424_;
  wire _22425_;
  wire _22426_;
  wire _22427_;
  wire _22428_;
  wire _22429_;
  wire _22430_;
  wire _22431_;
  wire _22432_;
  wire _22433_;
  wire _22434_;
  wire _22435_;
  wire _22436_;
  wire _22437_;
  wire _22438_;
  wire _22439_;
  wire _22440_;
  wire _22441_;
  wire _22442_;
  wire _22443_;
  wire _22444_;
  wire _22445_;
  wire _22446_;
  wire _22447_;
  wire _22448_;
  wire _22449_;
  wire _22450_;
  wire _22451_;
  wire _22452_;
  wire _22453_;
  wire _22454_;
  wire _22455_;
  wire _22456_;
  wire _22457_;
  wire _22458_;
  wire _22459_;
  wire _22460_;
  wire _22461_;
  wire _22462_;
  wire _22463_;
  wire _22464_;
  wire _22465_;
  wire _22466_;
  wire _22467_;
  wire _22468_;
  wire _22469_;
  wire _22470_;
  wire _22471_;
  wire _22472_;
  wire _22473_;
  wire _22474_;
  wire _22475_;
  wire _22476_;
  wire _22477_;
  wire _22478_;
  wire _22479_;
  wire _22480_;
  wire _22481_;
  wire _22482_;
  wire _22483_;
  wire _22484_;
  wire _22485_;
  wire _22486_;
  wire _22487_;
  wire _22488_;
  wire _22489_;
  wire _22490_;
  wire _22491_;
  wire _22492_;
  wire _22493_;
  wire _22494_;
  wire _22495_;
  wire _22496_;
  wire _22497_;
  wire _22498_;
  wire _22499_;
  wire _22500_;
  wire _22501_;
  wire _22502_;
  wire _22503_;
  wire _22504_;
  wire _22505_;
  wire _22506_;
  wire _22507_;
  wire _22508_;
  wire _22509_;
  wire _22510_;
  wire _22511_;
  wire _22512_;
  wire _22513_;
  wire _22514_;
  wire _22515_;
  wire _22516_;
  wire _22517_;
  wire _22518_;
  wire _22519_;
  wire _22520_;
  wire _22521_;
  wire _22522_;
  wire _22523_;
  wire _22524_;
  wire _22525_;
  wire _22526_;
  wire _22527_;
  wire _22528_;
  wire _22529_;
  wire _22530_;
  wire _22531_;
  wire _22532_;
  wire _22533_;
  wire _22534_;
  wire _22535_;
  wire _22536_;
  wire _22537_;
  wire _22538_;
  wire _22539_;
  wire _22540_;
  wire _22541_;
  wire _22542_;
  wire _22543_;
  wire _22544_;
  wire _22545_;
  wire _22546_;
  wire _22547_;
  wire _22548_;
  wire _22549_;
  wire _22550_;
  wire _22551_;
  wire _22552_;
  wire _22553_;
  wire _22554_;
  wire _22555_;
  wire _22556_;
  wire _22557_;
  wire _22558_;
  wire _22559_;
  wire _22560_;
  wire _22561_;
  wire _22562_;
  wire _22563_;
  wire _22564_;
  wire _22565_;
  wire _22566_;
  wire _22567_;
  wire _22568_;
  wire _22569_;
  wire _22570_;
  wire _22571_;
  wire _22572_;
  wire _22573_;
  wire _22574_;
  wire _22575_;
  wire _22576_;
  wire _22577_;
  wire _22578_;
  wire _22579_;
  wire _22580_;
  wire _22581_;
  wire _22582_;
  wire _22583_;
  wire _22584_;
  wire _22585_;
  wire _22586_;
  wire _22587_;
  wire _22588_;
  wire _22589_;
  wire _22590_;
  wire _22591_;
  wire _22592_;
  wire _22593_;
  wire _22594_;
  wire _22595_;
  wire _22596_;
  wire _22597_;
  wire _22598_;
  wire _22599_;
  wire _22600_;
  wire _22601_;
  wire _22602_;
  wire _22603_;
  wire _22604_;
  wire _22605_;
  wire _22606_;
  wire _22607_;
  wire _22608_;
  wire _22609_;
  wire _22610_;
  wire _22611_;
  wire _22612_;
  wire _22613_;
  wire _22614_;
  wire _22615_;
  wire _22616_;
  wire _22617_;
  wire _22618_;
  wire _22619_;
  wire _22620_;
  wire _22621_;
  wire _22622_;
  wire _22623_;
  wire _22624_;
  wire _22625_;
  wire _22626_;
  wire _22627_;
  wire _22628_;
  wire _22629_;
  wire _22630_;
  wire _22631_;
  wire _22632_;
  wire _22633_;
  wire _22634_;
  wire _22635_;
  wire _22636_;
  wire _22637_;
  wire _22638_;
  wire _22639_;
  wire _22640_;
  wire _22641_;
  wire _22642_;
  wire _22643_;
  wire _22644_;
  wire _22645_;
  wire _22646_;
  wire _22647_;
  wire _22648_;
  wire _22649_;
  wire _22650_;
  wire _22651_;
  wire _22652_;
  wire _22653_;
  wire _22654_;
  wire _22655_;
  wire _22656_;
  wire _22657_;
  wire _22658_;
  wire _22659_;
  wire _22660_;
  wire _22661_;
  wire _22662_;
  wire _22663_;
  wire _22664_;
  wire _22665_;
  wire _22666_;
  wire _22667_;
  wire _22668_;
  wire _22669_;
  wire _22670_;
  wire _22671_;
  wire _22672_;
  wire _22673_;
  wire _22674_;
  wire _22675_;
  wire _22676_;
  wire _22677_;
  wire _22678_;
  wire _22679_;
  wire _22680_;
  wire _22681_;
  wire _22682_;
  wire _22683_;
  wire _22684_;
  wire _22685_;
  wire _22686_;
  wire _22687_;
  wire _22688_;
  wire _22689_;
  wire _22690_;
  wire _22691_;
  wire _22692_;
  wire _22693_;
  wire _22694_;
  wire _22695_;
  wire _22696_;
  wire _22697_;
  wire _22698_;
  wire _22699_;
  wire _22700_;
  wire _22701_;
  wire _22702_;
  wire _22703_;
  wire _22704_;
  wire _22705_;
  wire _22706_;
  wire _22707_;
  wire _22708_;
  wire _22709_;
  wire _22710_;
  wire _22711_;
  wire _22712_;
  wire _22713_;
  wire _22714_;
  wire _22715_;
  wire _22716_;
  wire _22717_;
  wire _22718_;
  wire _22719_;
  wire _22720_;
  wire _22721_;
  wire _22722_;
  wire _22723_;
  wire _22724_;
  wire _22725_;
  wire _22726_;
  wire _22727_;
  wire _22728_;
  wire _22729_;
  wire _22730_;
  wire _22731_;
  wire _22732_;
  wire _22733_;
  wire _22734_;
  wire _22735_;
  wire _22736_;
  wire _22737_;
  wire _22738_;
  wire _22739_;
  wire _22740_;
  wire _22741_;
  wire _22742_;
  wire _22743_;
  wire _22744_;
  wire _22745_;
  wire _22746_;
  wire _22747_;
  wire _22748_;
  wire _22749_;
  wire _22750_;
  wire _22751_;
  wire _22752_;
  wire _22753_;
  wire _22754_;
  wire _22755_;
  wire _22756_;
  wire _22757_;
  wire _22758_;
  wire _22759_;
  wire _22760_;
  wire _22761_;
  wire _22762_;
  wire _22763_;
  wire _22764_;
  wire _22765_;
  wire _22766_;
  wire _22767_;
  wire _22768_;
  wire _22769_;
  wire _22770_;
  wire _22771_;
  wire _22772_;
  wire _22773_;
  wire _22774_;
  wire _22775_;
  wire _22776_;
  wire _22777_;
  wire _22778_;
  wire _22779_;
  wire _22780_;
  wire _22781_;
  wire _22782_;
  wire _22783_;
  wire _22784_;
  wire _22785_;
  wire _22786_;
  wire _22787_;
  wire _22788_;
  wire _22789_;
  wire _22790_;
  wire _22791_;
  wire _22792_;
  wire _22793_;
  wire _22794_;
  wire _22795_;
  wire _22796_;
  wire _22797_;
  wire _22798_;
  wire _22799_;
  wire _22800_;
  wire _22801_;
  wire _22802_;
  wire _22803_;
  wire _22804_;
  wire _22805_;
  wire _22806_;
  wire _22807_;
  wire _22808_;
  wire _22809_;
  wire _22810_;
  wire _22811_;
  wire _22812_;
  wire _22813_;
  wire _22814_;
  wire _22815_;
  wire _22816_;
  wire _22817_;
  wire _22818_;
  wire _22819_;
  wire _22820_;
  wire _22821_;
  wire _22822_;
  wire _22823_;
  wire _22824_;
  wire _22825_;
  wire _22826_;
  wire _22827_;
  wire _22828_;
  wire _22829_;
  wire _22830_;
  wire _22831_;
  wire _22832_;
  wire _22833_;
  wire _22834_;
  wire _22835_;
  wire _22836_;
  wire _22837_;
  wire _22838_;
  wire _22839_;
  wire _22840_;
  wire _22841_;
  wire _22842_;
  wire _22843_;
  wire _22844_;
  wire _22845_;
  wire _22846_;
  wire _22847_;
  wire _22848_;
  wire _22849_;
  wire _22850_;
  wire _22851_;
  wire _22852_;
  wire _22853_;
  wire _22854_;
  wire _22855_;
  wire _22856_;
  wire _22857_;
  wire _22858_;
  wire _22859_;
  wire _22860_;
  wire _22861_;
  wire _22862_;
  wire _22863_;
  wire _22864_;
  wire _22865_;
  wire _22866_;
  wire _22867_;
  wire _22868_;
  wire _22869_;
  wire _22870_;
  wire _22871_;
  wire _22872_;
  wire _22873_;
  wire _22874_;
  wire _22875_;
  wire _22876_;
  wire _22877_;
  wire _22878_;
  wire _22879_;
  wire _22880_;
  wire _22881_;
  wire _22882_;
  wire _22883_;
  wire _22884_;
  wire _22885_;
  wire _22886_;
  wire _22887_;
  wire _22888_;
  wire _22889_;
  wire _22890_;
  wire _22891_;
  wire _22892_;
  wire _22893_;
  wire _22894_;
  wire _22895_;
  wire _22896_;
  wire _22897_;
  wire _22898_;
  wire _22899_;
  wire _22900_;
  wire _22901_;
  wire _22902_;
  wire _22903_;
  wire _22904_;
  wire _22905_;
  wire _22906_;
  wire _22907_;
  wire _22908_;
  wire _22909_;
  wire _22910_;
  wire _22911_;
  wire _22912_;
  wire _22913_;
  wire _22914_;
  wire _22915_;
  wire _22916_;
  wire _22917_;
  wire _22918_;
  wire _22919_;
  wire _22920_;
  wire _22921_;
  wire _22922_;
  wire _22923_;
  wire _22924_;
  wire _22925_;
  wire _22926_;
  wire _22927_;
  wire _22928_;
  wire _22929_;
  wire _22930_;
  wire _22931_;
  wire _22932_;
  wire _22933_;
  wire _22934_;
  wire _22935_;
  wire _22936_;
  wire _22937_;
  wire _22938_;
  wire _22939_;
  wire _22940_;
  wire _22941_;
  wire _22942_;
  wire _22943_;
  wire _22944_;
  wire _22945_;
  wire _22946_;
  wire _22947_;
  wire _22948_;
  wire _22949_;
  wire _22950_;
  wire _22951_;
  wire _22952_;
  wire _22953_;
  wire _22954_;
  wire _22955_;
  wire _22956_;
  wire _22957_;
  wire _22958_;
  wire _22959_;
  wire _22960_;
  wire _22961_;
  wire _22962_;
  wire _22963_;
  wire _22964_;
  wire _22965_;
  wire _22966_;
  wire _22967_;
  wire _22968_;
  wire _22969_;
  wire _22970_;
  wire _22971_;
  wire _22972_;
  wire _22973_;
  wire _22974_;
  wire _22975_;
  wire _22976_;
  wire _22977_;
  wire _22978_;
  wire _22979_;
  wire _22980_;
  wire _22981_;
  wire _22982_;
  wire _22983_;
  wire _22984_;
  wire _22985_;
  wire _22986_;
  wire _22987_;
  wire _22988_;
  wire _22989_;
  wire _22990_;
  wire _22991_;
  wire _22992_;
  wire _22993_;
  wire _22994_;
  wire _22995_;
  wire _22996_;
  wire _22997_;
  wire _22998_;
  wire _22999_;
  wire _23000_;
  wire _23001_;
  wire _23002_;
  wire _23003_;
  wire _23004_;
  wire _23005_;
  wire _23006_;
  wire _23007_;
  wire _23008_;
  wire _23009_;
  wire _23010_;
  wire _23011_;
  wire _23012_;
  wire _23013_;
  wire _23014_;
  wire _23015_;
  wire _23016_;
  wire _23017_;
  wire _23018_;
  wire _23019_;
  wire _23020_;
  wire _23021_;
  wire _23022_;
  wire _23023_;
  wire _23024_;
  wire _23025_;
  wire _23026_;
  wire _23027_;
  wire _23028_;
  wire _23029_;
  wire _23030_;
  wire _23031_;
  wire _23032_;
  wire _23033_;
  wire _23034_;
  wire _23035_;
  wire _23036_;
  wire _23037_;
  wire _23038_;
  wire _23039_;
  wire _23040_;
  wire _23041_;
  wire _23042_;
  wire _23043_;
  wire _23044_;
  wire _23045_;
  wire _23046_;
  wire _23047_;
  wire _23048_;
  wire _23049_;
  wire _23050_;
  wire _23051_;
  wire _23052_;
  wire _23053_;
  wire _23054_;
  wire _23055_;
  wire _23056_;
  wire _23057_;
  wire _23058_;
  wire _23059_;
  wire _23060_;
  wire _23061_;
  wire _23062_;
  wire _23063_;
  wire _23064_;
  wire _23065_;
  wire _23066_;
  wire _23067_;
  wire _23068_;
  wire _23069_;
  wire _23070_;
  wire _23071_;
  wire _23072_;
  wire _23073_;
  wire _23074_;
  wire _23075_;
  wire _23076_;
  wire _23077_;
  wire _23078_;
  wire _23079_;
  wire _23080_;
  wire _23081_;
  wire _23082_;
  wire _23083_;
  wire _23084_;
  wire _23085_;
  wire _23086_;
  wire _23087_;
  wire _23088_;
  wire _23089_;
  wire _23090_;
  wire _23091_;
  wire _23092_;
  wire _23093_;
  wire _23094_;
  wire _23095_;
  wire _23096_;
  wire _23097_;
  wire _23098_;
  wire _23099_;
  wire _23100_;
  wire _23101_;
  wire _23102_;
  wire _23103_;
  wire _23104_;
  wire _23105_;
  wire _23106_;
  wire _23107_;
  wire _23108_;
  wire _23109_;
  wire _23110_;
  wire _23111_;
  wire _23112_;
  wire _23113_;
  wire _23114_;
  wire _23115_;
  wire _23116_;
  wire _23117_;
  wire _23118_;
  wire _23119_;
  wire _23120_;
  wire _23121_;
  wire _23122_;
  wire _23123_;
  wire _23124_;
  wire _23125_;
  wire _23126_;
  wire _23127_;
  wire _23128_;
  wire _23129_;
  wire _23130_;
  wire _23131_;
  wire _23132_;
  wire _23133_;
  wire _23134_;
  wire _23135_;
  wire _23136_;
  wire _23137_;
  wire _23138_;
  wire _23139_;
  wire _23140_;
  wire _23141_;
  wire _23142_;
  wire _23143_;
  wire _23144_;
  wire _23145_;
  wire _23146_;
  wire _23147_;
  wire _23148_;
  wire _23149_;
  wire _23150_;
  wire _23151_;
  wire _23152_;
  wire _23153_;
  wire _23154_;
  wire _23155_;
  wire _23156_;
  wire _23157_;
  wire _23158_;
  wire _23159_;
  wire _23160_;
  wire _23161_;
  wire _23162_;
  wire _23163_;
  wire _23164_;
  wire _23165_;
  wire _23166_;
  wire _23167_;
  wire _23168_;
  wire _23169_;
  wire _23170_;
  wire _23171_;
  wire _23172_;
  wire _23173_;
  wire _23174_;
  wire _23175_;
  wire _23176_;
  wire _23177_;
  wire _23178_;
  wire _23179_;
  wire _23180_;
  wire _23181_;
  wire _23182_;
  wire _23183_;
  wire _23184_;
  wire _23185_;
  wire _23186_;
  wire _23187_;
  wire _23188_;
  wire _23189_;
  wire _23190_;
  wire _23191_;
  wire _23192_;
  wire _23193_;
  wire _23194_;
  wire _23195_;
  wire _23196_;
  wire _23197_;
  wire _23198_;
  wire _23199_;
  wire _23200_;
  wire _23201_;
  wire _23202_;
  wire _23203_;
  wire _23204_;
  wire _23205_;
  wire _23206_;
  wire _23207_;
  wire _23208_;
  wire _23209_;
  wire _23210_;
  wire _23211_;
  wire _23212_;
  wire _23213_;
  wire _23214_;
  wire _23215_;
  wire _23216_;
  wire _23217_;
  wire _23218_;
  wire _23219_;
  wire _23220_;
  wire _23221_;
  wire _23222_;
  wire _23223_;
  wire _23224_;
  wire _23225_;
  wire _23226_;
  wire _23227_;
  wire _23228_;
  wire _23229_;
  wire _23230_;
  wire _23231_;
  wire _23232_;
  wire _23233_;
  wire _23234_;
  wire _23235_;
  wire _23236_;
  wire _23237_;
  wire _23238_;
  wire _23239_;
  wire _23240_;
  wire _23241_;
  wire _23242_;
  wire _23243_;
  wire _23244_;
  wire _23245_;
  wire _23246_;
  wire _23247_;
  wire _23248_;
  wire _23249_;
  wire _23250_;
  wire _23251_;
  wire _23252_;
  wire _23253_;
  wire _23254_;
  wire _23255_;
  wire _23256_;
  wire _23257_;
  wire _23258_;
  wire _23259_;
  wire _23260_;
  wire _23261_;
  wire _23262_;
  wire _23263_;
  wire _23264_;
  wire _23265_;
  wire _23266_;
  wire _23267_;
  wire _23268_;
  wire _23269_;
  wire _23270_;
  wire _23271_;
  wire _23272_;
  wire _23273_;
  wire _23274_;
  wire _23275_;
  wire _23276_;
  wire _23277_;
  wire _23278_;
  wire _23279_;
  wire _23280_;
  wire _23281_;
  wire _23282_;
  wire _23283_;
  wire _23284_;
  wire _23285_;
  wire _23286_;
  wire _23287_;
  wire _23288_;
  wire _23289_;
  wire _23290_;
  wire _23291_;
  wire _23292_;
  wire _23293_;
  wire _23294_;
  wire _23295_;
  wire _23296_;
  wire _23297_;
  wire _23298_;
  wire _23299_;
  wire _23300_;
  wire _23301_;
  wire _23302_;
  wire _23303_;
  wire _23304_;
  wire _23305_;
  wire _23306_;
  wire _23307_;
  wire _23308_;
  wire _23309_;
  wire _23310_;
  wire _23311_;
  wire _23312_;
  wire _23313_;
  wire _23314_;
  wire _23315_;
  wire _23316_;
  wire _23317_;
  wire _23318_;
  wire _23319_;
  wire _23320_;
  wire _23321_;
  wire _23322_;
  wire _23323_;
  wire _23324_;
  wire _23325_;
  wire _23326_;
  wire _23327_;
  wire _23328_;
  wire _23329_;
  wire _23330_;
  wire _23331_;
  wire _23332_;
  wire _23333_;
  wire _23334_;
  wire _23335_;
  wire _23336_;
  wire _23337_;
  wire _23338_;
  wire _23339_;
  wire _23340_;
  wire _23341_;
  wire _23342_;
  wire _23343_;
  wire _23344_;
  wire _23345_;
  wire _23346_;
  wire _23347_;
  wire _23348_;
  wire _23349_;
  wire _23350_;
  wire _23351_;
  wire _23352_;
  wire _23353_;
  wire _23354_;
  wire _23355_;
  wire _23356_;
  wire _23357_;
  wire _23358_;
  wire _23359_;
  wire _23360_;
  wire _23361_;
  wire _23362_;
  wire _23363_;
  wire _23364_;
  wire _23365_;
  wire _23366_;
  wire _23367_;
  wire _23368_;
  wire _23369_;
  wire _23370_;
  wire _23371_;
  wire _23372_;
  wire _23373_;
  wire _23374_;
  wire _23375_;
  wire _23376_;
  wire _23377_;
  wire _23378_;
  wire _23379_;
  wire _23380_;
  wire _23381_;
  wire _23382_;
  wire _23383_;
  wire _23384_;
  wire _23385_;
  wire _23386_;
  wire _23387_;
  wire _23388_;
  wire _23389_;
  wire _23390_;
  wire _23391_;
  wire _23392_;
  wire _23393_;
  wire _23394_;
  wire _23395_;
  wire _23396_;
  wire _23397_;
  wire _23398_;
  wire _23399_;
  wire _23400_;
  wire _23401_;
  wire _23402_;
  wire _23403_;
  wire _23404_;
  wire _23405_;
  wire _23406_;
  wire _23407_;
  wire _23408_;
  wire _23409_;
  wire _23410_;
  wire _23411_;
  wire _23412_;
  wire _23413_;
  wire _23414_;
  wire _23415_;
  wire _23416_;
  wire _23417_;
  wire _23418_;
  wire _23419_;
  wire _23420_;
  wire _23421_;
  wire _23422_;
  wire _23423_;
  wire _23424_;
  wire _23425_;
  wire _23426_;
  wire _23427_;
  wire _23428_;
  wire _23429_;
  wire _23430_;
  wire _23431_;
  wire _23432_;
  wire _23433_;
  wire _23434_;
  wire _23435_;
  wire _23436_;
  wire _23437_;
  wire _23438_;
  wire _23439_;
  wire _23440_;
  wire _23441_;
  wire _23442_;
  wire _23443_;
  wire _23444_;
  wire _23445_;
  wire _23446_;
  wire _23447_;
  wire _23448_;
  wire _23449_;
  wire _23450_;
  wire _23451_;
  wire _23452_;
  wire _23453_;
  wire _23454_;
  wire _23455_;
  wire _23456_;
  wire _23457_;
  wire _23458_;
  wire _23459_;
  wire _23460_;
  wire _23461_;
  wire _23462_;
  wire _23463_;
  wire _23464_;
  wire _23465_;
  wire _23466_;
  wire _23467_;
  wire _23468_;
  wire _23469_;
  wire _23470_;
  wire _23471_;
  wire _23472_;
  wire _23473_;
  wire _23474_;
  wire _23475_;
  wire _23476_;
  wire _23477_;
  wire _23478_;
  wire _23479_;
  wire _23480_;
  wire _23481_;
  wire _23482_;
  wire _23483_;
  wire _23484_;
  wire _23485_;
  wire _23486_;
  wire _23487_;
  wire _23488_;
  wire _23489_;
  wire _23490_;
  wire _23491_;
  wire _23492_;
  wire _23493_;
  wire _23494_;
  wire _23495_;
  wire _23496_;
  wire _23497_;
  wire _23498_;
  wire _23499_;
  wire _23500_;
  wire _23501_;
  wire _23502_;
  wire _23503_;
  wire _23504_;
  wire _23505_;
  wire _23506_;
  wire _23507_;
  wire _23508_;
  wire _23509_;
  wire _23510_;
  wire _23511_;
  wire _23512_;
  wire _23513_;
  wire _23514_;
  wire _23515_;
  wire _23516_;
  wire _23517_;
  wire _23518_;
  wire _23519_;
  wire _23520_;
  wire _23521_;
  wire _23522_;
  wire _23523_;
  wire _23524_;
  wire _23525_;
  wire _23526_;
  wire _23527_;
  wire _23528_;
  wire _23529_;
  wire _23530_;
  wire _23531_;
  wire _23532_;
  wire _23533_;
  wire _23534_;
  wire _23535_;
  wire _23536_;
  wire _23537_;
  wire _23538_;
  wire _23539_;
  wire _23540_;
  wire _23541_;
  wire _23542_;
  wire _23543_;
  wire _23544_;
  wire _23545_;
  wire _23546_;
  wire _23547_;
  wire _23548_;
  wire _23549_;
  wire _23550_;
  wire _23551_;
  wire _23552_;
  wire _23553_;
  wire _23554_;
  wire _23555_;
  wire _23556_;
  wire _23557_;
  wire _23558_;
  wire _23559_;
  wire _23560_;
  wire _23561_;
  wire _23562_;
  wire _23563_;
  wire _23564_;
  wire _23565_;
  wire _23566_;
  wire _23567_;
  wire _23568_;
  wire _23569_;
  wire _23570_;
  wire _23571_;
  wire _23572_;
  wire _23573_;
  wire _23574_;
  wire _23575_;
  wire _23576_;
  wire _23577_;
  wire _23578_;
  wire _23579_;
  wire _23580_;
  wire _23581_;
  wire _23582_;
  wire _23583_;
  wire _23584_;
  wire _23585_;
  wire _23586_;
  wire _23587_;
  wire _23588_;
  wire _23589_;
  wire _23590_;
  wire _23591_;
  wire _23592_;
  wire _23593_;
  wire _23594_;
  wire _23595_;
  wire _23596_;
  wire _23597_;
  wire _23598_;
  wire _23599_;
  wire _23600_;
  wire _23601_;
  wire _23602_;
  wire _23603_;
  wire _23604_;
  wire _23605_;
  wire _23606_;
  wire _23607_;
  wire _23608_;
  wire _23609_;
  wire _23610_;
  wire _23611_;
  wire _23612_;
  wire _23613_;
  wire _23614_;
  wire _23615_;
  wire _23616_;
  wire _23617_;
  wire _23618_;
  wire _23619_;
  wire _23620_;
  wire _23621_;
  wire _23622_;
  wire _23623_;
  wire _23624_;
  wire _23625_;
  wire _23626_;
  wire _23627_;
  wire _23628_;
  wire _23629_;
  wire _23630_;
  wire _23631_;
  wire _23632_;
  wire _23633_;
  wire _23634_;
  wire _23635_;
  wire _23636_;
  wire _23637_;
  wire _23638_;
  wire _23639_;
  wire _23640_;
  wire _23641_;
  wire _23642_;
  wire _23643_;
  wire _23644_;
  wire _23645_;
  wire _23646_;
  wire _23647_;
  wire _23648_;
  wire _23649_;
  wire _23650_;
  wire _23651_;
  wire _23652_;
  wire _23653_;
  wire _23654_;
  wire _23655_;
  wire _23656_;
  wire _23657_;
  wire _23658_;
  wire _23659_;
  wire _23660_;
  wire _23661_;
  wire _23662_;
  wire _23663_;
  wire _23664_;
  wire _23665_;
  wire _23666_;
  wire _23667_;
  wire _23668_;
  wire _23669_;
  wire _23670_;
  wire _23671_;
  wire _23672_;
  wire _23673_;
  wire _23674_;
  wire _23675_;
  wire _23676_;
  wire _23677_;
  wire _23678_;
  wire _23679_;
  wire _23680_;
  wire _23681_;
  wire _23682_;
  wire _23683_;
  wire _23684_;
  wire _23685_;
  wire _23686_;
  wire _23687_;
  wire _23688_;
  wire _23689_;
  wire _23690_;
  wire _23691_;
  wire _23692_;
  wire _23693_;
  wire _23694_;
  wire _23695_;
  wire _23696_;
  wire _23697_;
  wire _23698_;
  wire _23699_;
  wire _23700_;
  wire _23701_;
  wire _23702_;
  wire _23703_;
  wire _23704_;
  wire _23705_;
  wire _23706_;
  wire _23707_;
  wire _23708_;
  wire _23709_;
  wire _23710_;
  wire _23711_;
  wire _23712_;
  wire _23713_;
  wire _23714_;
  wire _23715_;
  wire _23716_;
  wire _23717_;
  wire _23718_;
  wire _23719_;
  wire _23720_;
  wire _23721_;
  wire _23722_;
  wire _23723_;
  wire _23724_;
  wire _23725_;
  wire _23726_;
  wire _23727_;
  wire _23728_;
  wire _23729_;
  wire _23730_;
  wire _23731_;
  wire _23732_;
  wire _23733_;
  wire _23734_;
  wire _23735_;
  wire _23736_;
  wire _23737_;
  wire _23738_;
  wire _23739_;
  wire _23740_;
  wire _23741_;
  wire _23742_;
  wire _23743_;
  wire _23744_;
  wire _23745_;
  wire _23746_;
  wire _23747_;
  wire _23748_;
  wire _23749_;
  wire _23750_;
  wire _23751_;
  wire _23752_;
  wire _23753_;
  wire _23754_;
  wire _23755_;
  wire _23756_;
  wire _23757_;
  wire _23758_;
  wire _23759_;
  wire _23760_;
  wire _23761_;
  wire _23762_;
  wire _23763_;
  wire _23764_;
  wire _23765_;
  wire _23766_;
  wire _23767_;
  wire _23768_;
  wire _23769_;
  wire _23770_;
  wire _23771_;
  wire _23772_;
  wire _23773_;
  wire _23774_;
  wire _23775_;
  wire _23776_;
  wire _23777_;
  wire _23778_;
  wire _23779_;
  wire _23780_;
  wire _23781_;
  wire _23782_;
  wire _23783_;
  wire _23784_;
  wire _23785_;
  wire _23786_;
  wire _23787_;
  wire _23788_;
  wire _23789_;
  wire _23790_;
  wire _23791_;
  wire _23792_;
  wire _23793_;
  wire _23794_;
  wire _23795_;
  wire _23796_;
  wire _23797_;
  wire _23798_;
  wire _23799_;
  wire _23800_;
  wire _23801_;
  wire _23802_;
  wire _23803_;
  wire _23804_;
  wire _23805_;
  wire _23806_;
  wire _23807_;
  wire _23808_;
  wire _23809_;
  wire _23810_;
  wire _23811_;
  wire _23812_;
  wire _23813_;
  wire _23814_;
  wire _23815_;
  wire _23816_;
  wire _23817_;
  wire _23818_;
  wire _23819_;
  wire _23820_;
  wire _23821_;
  wire _23822_;
  wire _23823_;
  wire _23824_;
  wire _23825_;
  wire _23826_;
  wire _23827_;
  wire _23828_;
  wire _23829_;
  wire _23830_;
  wire _23831_;
  wire _23832_;
  wire _23833_;
  wire _23834_;
  wire _23835_;
  wire _23836_;
  wire _23837_;
  wire _23838_;
  wire _23839_;
  wire _23840_;
  wire _23841_;
  wire _23842_;
  wire _23843_;
  wire _23844_;
  wire _23845_;
  wire _23846_;
  wire _23847_;
  wire _23848_;
  wire _23849_;
  wire _23850_;
  wire _23851_;
  wire _23852_;
  wire _23853_;
  wire _23854_;
  wire _23855_;
  wire _23856_;
  wire _23857_;
  wire _23858_;
  wire _23859_;
  wire _23860_;
  wire _23861_;
  wire _23862_;
  wire _23863_;
  wire _23864_;
  wire _23865_;
  wire _23866_;
  wire _23867_;
  wire _23868_;
  wire _23869_;
  wire _23870_;
  wire _23871_;
  wire _23872_;
  wire _23873_;
  wire _23874_;
  wire _23875_;
  wire _23876_;
  wire _23877_;
  wire _23878_;
  wire _23879_;
  wire _23880_;
  wire _23881_;
  wire _23882_;
  wire _23883_;
  wire _23884_;
  wire _23885_;
  wire _23886_;
  wire _23887_;
  wire _23888_;
  wire _23889_;
  wire _23890_;
  wire _23891_;
  wire _23892_;
  wire _23893_;
  wire _23894_;
  wire _23895_;
  wire _23896_;
  wire _23897_;
  wire _23898_;
  wire _23899_;
  wire _23900_;
  wire _23901_;
  wire _23902_;
  wire _23903_;
  wire _23904_;
  wire _23905_;
  wire _23906_;
  wire _23907_;
  wire _23908_;
  wire _23909_;
  wire _23910_;
  wire _23911_;
  wire _23912_;
  wire _23913_;
  wire _23914_;
  wire _23915_;
  wire _23916_;
  wire _23917_;
  wire _23918_;
  wire _23919_;
  wire _23920_;
  wire _23921_;
  wire _23922_;
  wire _23923_;
  wire _23924_;
  wire _23925_;
  wire _23926_;
  wire _23927_;
  wire _23928_;
  wire _23929_;
  wire _23930_;
  wire _23931_;
  wire _23932_;
  wire _23933_;
  wire _23934_;
  wire _23935_;
  wire _23936_;
  wire _23937_;
  wire _23938_;
  wire _23939_;
  wire _23940_;
  wire _23941_;
  wire _23942_;
  wire _23943_;
  wire _23944_;
  wire _23945_;
  wire _23946_;
  wire _23947_;
  wire _23948_;
  wire _23949_;
  wire _23950_;
  wire _23951_;
  wire _23952_;
  wire _23953_;
  wire _23954_;
  wire _23955_;
  wire _23956_;
  wire _23957_;
  wire _23958_;
  wire _23959_;
  wire _23960_;
  wire _23961_;
  wire _23962_;
  wire _23963_;
  wire _23964_;
  wire _23965_;
  wire _23966_;
  wire _23967_;
  wire _23968_;
  wire _23969_;
  wire _23970_;
  wire _23971_;
  wire _23972_;
  wire _23973_;
  wire _23974_;
  wire _23975_;
  wire _23976_;
  wire _23977_;
  wire _23978_;
  wire _23979_;
  wire _23980_;
  wire _23981_;
  wire _23982_;
  wire _23983_;
  wire _23984_;
  wire _23985_;
  wire _23986_;
  wire _23987_;
  wire _23988_;
  wire _23989_;
  wire _23990_;
  wire _23991_;
  wire _23992_;
  wire _23993_;
  wire _23994_;
  wire _23995_;
  wire _23996_;
  wire _23997_;
  wire _23998_;
  wire _23999_;
  wire _24000_;
  wire _24001_;
  wire _24002_;
  wire _24003_;
  wire _24004_;
  wire _24005_;
  wire _24006_;
  wire _24007_;
  wire _24008_;
  wire _24009_;
  wire _24010_;
  wire _24011_;
  wire _24012_;
  wire _24013_;
  wire _24014_;
  wire _24015_;
  wire _24016_;
  wire _24017_;
  wire _24018_;
  wire _24019_;
  wire _24020_;
  wire _24021_;
  wire _24022_;
  wire _24023_;
  wire _24024_;
  wire _24025_;
  wire _24026_;
  wire _24027_;
  wire _24028_;
  wire _24029_;
  wire _24030_;
  wire _24031_;
  wire _24032_;
  wire _24033_;
  wire _24034_;
  wire _24035_;
  wire _24036_;
  wire _24037_;
  wire _24038_;
  wire _24039_;
  wire _24040_;
  wire _24041_;
  wire _24042_;
  wire _24043_;
  wire _24044_;
  wire _24045_;
  wire _24046_;
  wire _24047_;
  wire _24048_;
  wire _24049_;
  wire _24050_;
  wire _24051_;
  wire _24052_;
  wire _24053_;
  wire _24054_;
  wire _24055_;
  wire _24056_;
  wire _24057_;
  wire _24058_;
  wire _24059_;
  wire _24060_;
  wire _24061_;
  wire _24062_;
  wire _24063_;
  wire _24064_;
  wire _24065_;
  wire _24066_;
  wire _24067_;
  wire _24068_;
  wire _24069_;
  wire _24070_;
  wire _24071_;
  wire _24072_;
  wire _24073_;
  wire _24074_;
  wire _24075_;
  wire _24076_;
  wire _24077_;
  wire _24078_;
  wire _24079_;
  wire _24080_;
  wire _24081_;
  wire _24082_;
  wire _24083_;
  wire _24084_;
  wire _24085_;
  wire _24086_;
  wire _24087_;
  wire _24088_;
  wire _24089_;
  wire _24090_;
  wire _24091_;
  wire _24092_;
  wire _24093_;
  wire _24094_;
  wire _24095_;
  wire _24096_;
  wire _24097_;
  wire _24098_;
  wire _24099_;
  wire _24100_;
  wire _24101_;
  wire _24102_;
  wire _24103_;
  wire _24104_;
  wire _24105_;
  wire _24106_;
  wire _24107_;
  wire _24108_;
  wire _24109_;
  wire _24110_;
  wire _24111_;
  wire _24112_;
  wire _24113_;
  wire _24114_;
  wire _24115_;
  wire _24116_;
  wire _24117_;
  wire _24118_;
  wire _24119_;
  wire _24120_;
  wire _24121_;
  wire _24122_;
  wire _24123_;
  wire _24124_;
  wire _24125_;
  wire _24126_;
  wire _24127_;
  wire _24128_;
  wire _24129_;
  wire _24130_;
  wire _24131_;
  wire _24132_;
  wire _24133_;
  wire _24134_;
  wire _24135_;
  wire _24136_;
  wire _24137_;
  wire _24138_;
  wire _24139_;
  wire _24140_;
  wire _24141_;
  wire _24142_;
  wire _24143_;
  wire _24144_;
  wire _24145_;
  wire _24146_;
  wire _24147_;
  wire _24148_;
  wire _24149_;
  wire _24150_;
  wire _24151_;
  wire _24152_;
  wire _24153_;
  wire _24154_;
  wire _24155_;
  wire _24156_;
  wire _24157_;
  wire _24158_;
  wire _24159_;
  wire _24160_;
  wire _24161_;
  wire _24162_;
  wire _24163_;
  wire _24164_;
  wire _24165_;
  wire _24166_;
  wire _24167_;
  wire _24168_;
  wire _24169_;
  wire _24170_;
  wire _24171_;
  wire _24172_;
  wire _24173_;
  wire _24174_;
  wire _24175_;
  wire _24176_;
  wire _24177_;
  wire _24178_;
  wire _24179_;
  wire _24180_;
  wire _24181_;
  wire _24182_;
  wire _24183_;
  wire _24184_;
  wire _24185_;
  wire _24186_;
  wire _24187_;
  wire _24188_;
  wire _24189_;
  wire _24190_;
  wire _24191_;
  wire _24192_;
  wire _24193_;
  wire _24194_;
  wire _24195_;
  wire _24196_;
  wire _24197_;
  wire _24198_;
  wire _24199_;
  wire _24200_;
  wire _24201_;
  wire _24202_;
  wire _24203_;
  wire _24204_;
  wire _24205_;
  wire _24206_;
  wire _24207_;
  wire _24208_;
  wire _24209_;
  wire _24210_;
  wire _24211_;
  wire _24212_;
  wire _24213_;
  wire _24214_;
  wire _24215_;
  wire _24216_;
  wire _24217_;
  wire _24218_;
  wire _24219_;
  wire _24220_;
  wire _24221_;
  wire _24222_;
  wire _24223_;
  wire _24224_;
  wire _24225_;
  wire _24226_;
  wire _24227_;
  wire _24228_;
  wire _24229_;
  wire _24230_;
  wire _24231_;
  wire _24232_;
  wire _24233_;
  wire _24234_;
  wire _24235_;
  wire _24236_;
  wire _24237_;
  wire _24238_;
  wire _24239_;
  wire _24240_;
  wire _24241_;
  wire _24242_;
  wire _24243_;
  wire _24244_;
  wire _24245_;
  wire _24246_;
  wire _24247_;
  wire _24248_;
  wire _24249_;
  wire _24250_;
  wire _24251_;
  wire _24252_;
  wire _24253_;
  wire _24254_;
  wire _24255_;
  wire _24256_;
  wire _24257_;
  wire _24258_;
  wire _24259_;
  wire _24260_;
  wire _24261_;
  wire _24262_;
  wire _24263_;
  wire _24264_;
  wire _24265_;
  wire _24266_;
  wire _24267_;
  wire _24268_;
  wire _24269_;
  wire _24270_;
  wire _24271_;
  wire _24272_;
  wire _24273_;
  wire _24274_;
  wire _24275_;
  wire _24276_;
  wire _24277_;
  wire _24278_;
  wire _24279_;
  wire _24280_;
  wire _24281_;
  wire _24282_;
  wire _24283_;
  wire _24284_;
  wire _24285_;
  wire _24286_;
  wire _24287_;
  wire _24288_;
  wire _24289_;
  wire _24290_;
  wire _24291_;
  wire _24292_;
  wire _24293_;
  wire _24294_;
  wire _24295_;
  wire _24296_;
  wire _24297_;
  wire _24298_;
  wire _24299_;
  wire _24300_;
  wire _24301_;
  wire _24302_;
  wire _24303_;
  wire _24304_;
  wire _24305_;
  wire _24306_;
  wire _24307_;
  wire _24308_;
  wire _24309_;
  wire _24310_;
  wire _24311_;
  wire _24312_;
  wire _24313_;
  wire _24314_;
  wire _24315_;
  wire _24316_;
  wire _24317_;
  wire _24318_;
  wire _24319_;
  wire _24320_;
  wire _24321_;
  wire _24322_;
  wire _24323_;
  wire _24324_;
  wire _24325_;
  wire _24326_;
  wire _24327_;
  wire _24328_;
  wire _24329_;
  wire _24330_;
  wire _24331_;
  wire _24332_;
  wire _24333_;
  wire _24334_;
  wire _24335_;
  wire _24336_;
  wire _24337_;
  wire _24338_;
  wire _24339_;
  wire _24340_;
  wire _24341_;
  wire _24342_;
  wire _24343_;
  wire _24344_;
  wire _24345_;
  wire _24346_;
  wire _24347_;
  wire _24348_;
  wire _24349_;
  wire _24350_;
  wire _24351_;
  wire _24352_;
  wire _24353_;
  wire _24354_;
  wire _24355_;
  wire _24356_;
  wire _24357_;
  wire _24358_;
  wire _24359_;
  wire _24360_;
  wire _24361_;
  wire _24362_;
  wire _24363_;
  wire _24364_;
  wire _24365_;
  wire _24366_;
  wire _24367_;
  wire _24368_;
  wire _24369_;
  wire _24370_;
  wire _24371_;
  wire _24372_;
  wire _24373_;
  wire _24374_;
  wire _24375_;
  wire _24376_;
  wire _24377_;
  wire _24378_;
  wire _24379_;
  wire _24380_;
  wire _24381_;
  wire _24382_;
  wire _24383_;
  wire _24384_;
  wire _24385_;
  wire _24386_;
  wire _24387_;
  wire _24388_;
  wire _24389_;
  wire _24390_;
  wire _24391_;
  wire _24392_;
  wire _24393_;
  wire _24394_;
  wire _24395_;
  wire _24396_;
  wire _24397_;
  wire _24398_;
  wire _24399_;
  wire _24400_;
  wire _24401_;
  wire _24402_;
  wire _24403_;
  wire _24404_;
  wire _24405_;
  wire _24406_;
  wire _24407_;
  wire _24408_;
  wire _24409_;
  wire _24410_;
  wire _24411_;
  wire _24412_;
  wire _24413_;
  wire _24414_;
  wire _24415_;
  wire _24416_;
  wire _24417_;
  wire _24418_;
  wire _24419_;
  wire _24420_;
  wire _24421_;
  wire _24422_;
  wire _24423_;
  wire _24424_;
  wire _24425_;
  wire _24426_;
  wire _24427_;
  wire _24428_;
  wire _24429_;
  wire _24430_;
  wire _24431_;
  wire _24432_;
  wire _24433_;
  wire _24434_;
  wire _24435_;
  wire _24436_;
  wire _24437_;
  wire _24438_;
  wire _24439_;
  wire _24440_;
  wire _24441_;
  wire _24442_;
  wire _24443_;
  wire _24444_;
  wire _24445_;
  wire _24446_;
  wire _24447_;
  wire _24448_;
  wire _24449_;
  wire _24450_;
  wire _24451_;
  wire _24452_;
  wire _24453_;
  wire _24454_;
  wire _24455_;
  wire _24456_;
  wire _24457_;
  wire _24458_;
  wire _24459_;
  wire _24460_;
  wire _24461_;
  wire _24462_;
  wire _24463_;
  wire _24464_;
  wire _24465_;
  wire _24466_;
  wire _24467_;
  wire _24468_;
  wire _24469_;
  wire _24470_;
  wire _24471_;
  wire _24472_;
  wire _24473_;
  wire _24474_;
  wire _24475_;
  wire _24476_;
  wire _24477_;
  wire _24478_;
  wire _24479_;
  wire _24480_;
  wire _24481_;
  wire _24482_;
  wire _24483_;
  wire _24484_;
  wire _24485_;
  wire _24486_;
  wire _24487_;
  wire _24488_;
  wire _24489_;
  wire _24490_;
  wire _24491_;
  wire _24492_;
  wire _24493_;
  wire _24494_;
  wire _24495_;
  wire _24496_;
  wire _24497_;
  wire _24498_;
  wire _24499_;
  wire _24500_;
  wire _24501_;
  wire _24502_;
  wire _24503_;
  wire _24504_;
  wire _24505_;
  wire _24506_;
  wire _24507_;
  wire _24508_;
  wire _24509_;
  wire _24510_;
  wire _24511_;
  wire _24512_;
  wire _24513_;
  wire _24514_;
  wire _24515_;
  wire _24516_;
  wire _24517_;
  wire _24518_;
  wire _24519_;
  wire _24520_;
  wire _24521_;
  wire _24522_;
  wire _24523_;
  wire _24524_;
  wire _24525_;
  wire _24526_;
  wire _24527_;
  wire _24528_;
  wire _24529_;
  wire _24530_;
  wire _24531_;
  wire _24532_;
  wire _24533_;
  wire _24534_;
  wire _24535_;
  wire _24536_;
  wire _24537_;
  wire _24538_;
  wire _24539_;
  wire _24540_;
  wire _24541_;
  wire _24542_;
  wire _24543_;
  wire _24544_;
  wire _24545_;
  wire _24546_;
  wire _24547_;
  wire _24548_;
  wire _24549_;
  wire _24550_;
  wire _24551_;
  wire _24552_;
  wire _24553_;
  wire _24554_;
  wire _24555_;
  wire _24556_;
  wire _24557_;
  wire _24558_;
  wire _24559_;
  wire _24560_;
  wire _24561_;
  wire _24562_;
  wire _24563_;
  wire _24564_;
  wire _24565_;
  wire _24566_;
  wire _24567_;
  wire _24568_;
  wire _24569_;
  wire _24570_;
  wire _24571_;
  wire _24572_;
  wire _24573_;
  wire _24574_;
  wire _24575_;
  wire _24576_;
  wire _24577_;
  wire _24578_;
  wire _24579_;
  wire _24580_;
  wire _24581_;
  wire _24582_;
  wire _24583_;
  wire _24584_;
  wire _24585_;
  wire _24586_;
  wire _24587_;
  wire _24588_;
  wire _24589_;
  wire _24590_;
  wire _24591_;
  wire _24592_;
  wire _24593_;
  wire _24594_;
  wire _24595_;
  wire _24596_;
  wire _24597_;
  wire _24598_;
  wire _24599_;
  wire _24600_;
  wire _24601_;
  wire _24602_;
  wire _24603_;
  wire _24604_;
  wire _24605_;
  wire _24606_;
  wire _24607_;
  wire _24608_;
  wire _24609_;
  wire _24610_;
  wire _24611_;
  wire _24612_;
  wire _24613_;
  wire _24614_;
  wire _24615_;
  wire _24616_;
  wire _24617_;
  wire _24618_;
  wire _24619_;
  wire _24620_;
  wire _24621_;
  wire _24622_;
  wire _24623_;
  wire _24624_;
  wire _24625_;
  wire _24626_;
  wire _24627_;
  wire _24628_;
  wire _24629_;
  wire _24630_;
  wire _24631_;
  wire _24632_;
  wire _24633_;
  wire _24634_;
  wire _24635_;
  wire _24636_;
  wire _24637_;
  wire _24638_;
  wire _24639_;
  wire _24640_;
  wire _24641_;
  wire _24642_;
  wire _24643_;
  wire _24644_;
  wire _24645_;
  wire _24646_;
  wire _24647_;
  wire _24648_;
  wire _24649_;
  wire _24650_;
  wire _24651_;
  wire _24652_;
  wire _24653_;
  wire _24654_;
  wire _24655_;
  wire _24656_;
  wire _24657_;
  wire _24658_;
  wire _24659_;
  wire _24660_;
  wire _24661_;
  wire _24662_;
  wire _24663_;
  wire _24664_;
  wire _24665_;
  wire _24666_;
  wire _24667_;
  wire _24668_;
  wire _24669_;
  wire _24670_;
  wire _24671_;
  wire _24672_;
  wire _24673_;
  wire _24674_;
  wire _24675_;
  wire _24676_;
  wire _24677_;
  wire _24678_;
  wire _24679_;
  wire _24680_;
  wire _24681_;
  wire _24682_;
  wire _24683_;
  wire _24684_;
  wire _24685_;
  wire _24686_;
  wire _24687_;
  wire _24688_;
  wire _24689_;
  wire _24690_;
  wire _24691_;
  wire _24692_;
  wire _24693_;
  wire _24694_;
  wire _24695_;
  wire _24696_;
  wire _24697_;
  wire _24698_;
  wire _24699_;
  wire _24700_;
  wire _24701_;
  wire _24702_;
  wire _24703_;
  wire _24704_;
  wire _24705_;
  wire _24706_;
  wire _24707_;
  wire _24708_;
  wire _24709_;
  wire _24710_;
  wire _24711_;
  wire _24712_;
  wire _24713_;
  wire _24714_;
  wire _24715_;
  wire _24716_;
  wire _24717_;
  wire _24718_;
  wire _24719_;
  wire _24720_;
  wire _24721_;
  wire _24722_;
  wire _24723_;
  wire _24724_;
  wire _24725_;
  wire _24726_;
  wire _24727_;
  wire _24728_;
  wire _24729_;
  wire _24730_;
  wire _24731_;
  wire _24732_;
  wire _24733_;
  wire _24734_;
  wire _24735_;
  wire _24736_;
  wire _24737_;
  wire _24738_;
  wire _24739_;
  wire _24740_;
  wire _24741_;
  wire _24742_;
  wire _24743_;
  wire _24744_;
  wire _24745_;
  wire _24746_;
  wire _24747_;
  wire _24748_;
  wire _24749_;
  wire _24750_;
  wire _24751_;
  wire _24752_;
  wire _24753_;
  wire _24754_;
  wire _24755_;
  wire _24756_;
  wire _24757_;
  wire _24758_;
  wire _24759_;
  wire _24760_;
  wire _24761_;
  wire _24762_;
  wire _24763_;
  wire _24764_;
  wire _24765_;
  wire _24766_;
  wire _24767_;
  wire _24768_;
  wire _24769_;
  wire _24770_;
  wire _24771_;
  wire _24772_;
  wire _24773_;
  wire _24774_;
  wire _24775_;
  wire _24776_;
  wire _24777_;
  wire _24778_;
  wire _24779_;
  wire _24780_;
  wire _24781_;
  wire _24782_;
  wire _24783_;
  wire _24784_;
  wire _24785_;
  wire _24786_;
  wire _24787_;
  wire _24788_;
  wire _24789_;
  wire _24790_;
  wire _24791_;
  wire _24792_;
  wire _24793_;
  wire _24794_;
  wire _24795_;
  wire _24796_;
  wire _24797_;
  wire _24798_;
  wire _24799_;
  wire _24800_;
  wire _24801_;
  wire _24802_;
  wire _24803_;
  wire _24804_;
  wire _24805_;
  wire _24806_;
  wire _24807_;
  wire _24808_;
  wire _24809_;
  wire _24810_;
  wire _24811_;
  wire _24812_;
  wire _24813_;
  wire _24814_;
  wire _24815_;
  wire _24816_;
  wire _24817_;
  wire _24818_;
  wire _24819_;
  wire _24820_;
  wire _24821_;
  wire _24822_;
  wire _24823_;
  wire _24824_;
  wire _24825_;
  wire _24826_;
  wire _24827_;
  wire _24828_;
  wire _24829_;
  wire _24830_;
  wire _24831_;
  wire _24832_;
  wire _24833_;
  wire _24834_;
  wire _24835_;
  wire _24836_;
  wire _24837_;
  wire _24838_;
  wire _24839_;
  wire _24840_;
  wire _24841_;
  wire _24842_;
  wire _24843_;
  wire _24844_;
  wire _24845_;
  wire _24846_;
  wire _24847_;
  wire _24848_;
  wire _24849_;
  wire _24850_;
  wire _24851_;
  wire _24852_;
  wire _24853_;
  wire _24854_;
  wire _24855_;
  wire _24856_;
  wire _24857_;
  wire _24858_;
  wire _24859_;
  wire _24860_;
  wire _24861_;
  wire _24862_;
  wire _24863_;
  wire _24864_;
  wire _24865_;
  wire _24866_;
  wire _24867_;
  wire _24868_;
  wire _24869_;
  wire _24870_;
  wire _24871_;
  wire _24872_;
  wire _24873_;
  wire _24874_;
  wire _24875_;
  wire _24876_;
  wire _24877_;
  wire _24878_;
  wire _24879_;
  wire _24880_;
  wire _24881_;
  wire _24882_;
  wire _24883_;
  wire _24884_;
  wire _24885_;
  wire _24886_;
  wire _24887_;
  wire _24888_;
  wire _24889_;
  wire _24890_;
  wire _24891_;
  wire _24892_;
  wire _24893_;
  wire _24894_;
  wire _24895_;
  wire _24896_;
  wire _24897_;
  wire _24898_;
  wire _24899_;
  wire _24900_;
  wire _24901_;
  wire _24902_;
  wire _24903_;
  wire _24904_;
  wire _24905_;
  wire _24906_;
  wire _24907_;
  wire _24908_;
  wire _24909_;
  wire _24910_;
  wire _24911_;
  wire _24912_;
  wire _24913_;
  wire _24914_;
  wire _24915_;
  wire _24916_;
  wire _24917_;
  wire _24918_;
  wire _24919_;
  wire _24920_;
  wire _24921_;
  wire _24922_;
  wire _24923_;
  wire _24924_;
  wire _24925_;
  wire _24926_;
  wire _24927_;
  wire _24928_;
  wire _24929_;
  wire _24930_;
  wire _24931_;
  wire _24932_;
  wire _24933_;
  wire _24934_;
  wire _24935_;
  wire _24936_;
  wire _24937_;
  wire _24938_;
  wire _24939_;
  wire _24940_;
  wire _24941_;
  wire _24942_;
  wire _24943_;
  wire _24944_;
  wire _24945_;
  wire _24946_;
  wire _24947_;
  wire _24948_;
  wire _24949_;
  wire _24950_;
  wire _24951_;
  wire _24952_;
  wire _24953_;
  wire _24954_;
  wire _24955_;
  wire _24956_;
  wire _24957_;
  wire _24958_;
  wire _24959_;
  wire _24960_;
  wire _24961_;
  wire _24962_;
  wire _24963_;
  wire _24964_;
  wire _24965_;
  wire _24966_;
  wire _24967_;
  wire _24968_;
  wire _24969_;
  wire _24970_;
  wire _24971_;
  wire _24972_;
  wire _24973_;
  wire _24974_;
  wire _24975_;
  wire _24976_;
  wire _24977_;
  wire _24978_;
  wire _24979_;
  wire _24980_;
  wire _24981_;
  wire _24982_;
  wire _24983_;
  wire _24984_;
  wire _24985_;
  wire _24986_;
  wire _24987_;
  wire _24988_;
  wire _24989_;
  wire _24990_;
  wire _24991_;
  wire _24992_;
  wire _24993_;
  wire _24994_;
  wire _24995_;
  wire _24996_;
  wire _24997_;
  wire _24998_;
  wire _24999_;
  wire _25000_;
  wire _25001_;
  wire _25002_;
  wire _25003_;
  wire _25004_;
  wire _25005_;
  wire _25006_;
  wire _25007_;
  wire _25008_;
  wire _25009_;
  wire _25010_;
  wire _25011_;
  wire _25012_;
  wire _25013_;
  wire _25014_;
  wire _25015_;
  wire _25016_;
  wire _25017_;
  wire _25018_;
  wire _25019_;
  wire _25020_;
  wire _25021_;
  wire _25022_;
  wire _25023_;
  wire _25024_;
  wire _25025_;
  wire _25026_;
  wire _25027_;
  wire _25028_;
  wire _25029_;
  wire _25030_;
  wire _25031_;
  wire _25032_;
  wire _25033_;
  wire _25034_;
  wire _25035_;
  wire _25036_;
  wire _25037_;
  wire _25038_;
  wire _25039_;
  wire _25040_;
  wire _25041_;
  wire _25042_;
  wire _25043_;
  wire _25044_;
  wire _25045_;
  wire _25046_;
  wire _25047_;
  wire _25048_;
  wire _25049_;
  wire _25050_;
  wire _25051_;
  wire _25052_;
  wire _25053_;
  wire _25054_;
  wire _25055_;
  wire _25056_;
  wire _25057_;
  wire _25058_;
  wire _25059_;
  wire _25060_;
  wire _25061_;
  wire _25062_;
  wire _25063_;
  wire _25064_;
  wire _25065_;
  wire _25066_;
  wire _25067_;
  wire _25068_;
  wire _25069_;
  wire _25070_;
  wire _25071_;
  wire _25072_;
  wire _25073_;
  wire _25074_;
  wire _25075_;
  wire _25076_;
  wire _25077_;
  wire _25078_;
  wire _25079_;
  wire _25080_;
  wire _25081_;
  wire _25082_;
  wire _25083_;
  wire _25084_;
  wire _25085_;
  wire _25086_;
  wire _25087_;
  wire _25088_;
  wire _25089_;
  wire _25090_;
  wire _25091_;
  wire _25092_;
  wire _25093_;
  wire _25094_;
  wire _25095_;
  wire _25096_;
  wire _25097_;
  wire _25098_;
  wire _25099_;
  wire _25100_;
  wire _25101_;
  wire _25102_;
  wire _25103_;
  wire _25104_;
  wire _25105_;
  wire _25106_;
  wire _25107_;
  wire _25108_;
  wire _25109_;
  wire _25110_;
  wire _25111_;
  wire _25112_;
  wire _25113_;
  wire _25114_;
  wire _25115_;
  wire _25116_;
  wire _25117_;
  wire _25118_;
  wire _25119_;
  wire _25120_;
  wire _25121_;
  wire _25122_;
  wire _25123_;
  wire _25124_;
  wire _25125_;
  wire _25126_;
  wire _25127_;
  wire _25128_;
  wire _25129_;
  wire _25130_;
  wire _25131_;
  wire _25132_;
  wire _25133_;
  wire _25134_;
  wire _25135_;
  wire _25136_;
  wire _25137_;
  wire _25138_;
  wire _25139_;
  wire _25140_;
  wire _25141_;
  wire _25142_;
  wire _25143_;
  wire _25144_;
  wire _25145_;
  wire _25146_;
  wire _25147_;
  wire _25148_;
  wire _25149_;
  wire _25150_;
  wire _25151_;
  wire _25152_;
  wire _25153_;
  wire _25154_;
  wire _25155_;
  wire _25156_;
  wire _25157_;
  wire _25158_;
  wire _25159_;
  wire _25160_;
  wire _25161_;
  wire _25162_;
  wire _25163_;
  wire _25164_;
  wire _25165_;
  wire _25166_;
  wire _25167_;
  wire _25168_;
  wire _25169_;
  wire _25170_;
  wire _25171_;
  wire _25172_;
  wire _25173_;
  wire _25174_;
  wire _25175_;
  wire _25176_;
  wire _25177_;
  wire _25178_;
  wire _25179_;
  wire _25180_;
  wire _25181_;
  wire _25182_;
  wire _25183_;
  wire _25184_;
  wire _25185_;
  wire _25186_;
  wire _25187_;
  wire _25188_;
  wire _25189_;
  wire _25190_;
  wire _25191_;
  wire _25192_;
  wire _25193_;
  wire _25194_;
  wire _25195_;
  wire _25196_;
  wire _25197_;
  wire _25198_;
  wire _25199_;
  wire _25200_;
  wire _25201_;
  wire _25202_;
  wire _25203_;
  wire _25204_;
  wire _25205_;
  wire _25206_;
  wire _25207_;
  wire _25208_;
  wire _25209_;
  wire _25210_;
  wire _25211_;
  wire _25212_;
  wire _25213_;
  wire _25214_;
  wire _25215_;
  wire _25216_;
  wire _25217_;
  wire _25218_;
  wire _25219_;
  wire _25220_;
  wire _25221_;
  wire _25222_;
  wire _25223_;
  wire _25224_;
  wire _25225_;
  wire _25226_;
  wire _25227_;
  wire _25228_;
  wire _25229_;
  wire _25230_;
  wire _25231_;
  wire _25232_;
  wire _25233_;
  wire _25234_;
  wire _25235_;
  wire _25236_;
  wire _25237_;
  wire _25238_;
  wire _25239_;
  wire _25240_;
  wire _25241_;
  wire _25242_;
  wire _25243_;
  wire _25244_;
  wire _25245_;
  wire _25246_;
  wire _25247_;
  wire _25248_;
  wire _25249_;
  wire _25250_;
  wire _25251_;
  wire _25252_;
  wire _25253_;
  wire _25254_;
  wire _25255_;
  wire _25256_;
  wire _25257_;
  wire _25258_;
  wire _25259_;
  wire _25260_;
  wire _25261_;
  wire _25262_;
  wire _25263_;
  wire _25264_;
  wire _25265_;
  wire _25266_;
  wire _25267_;
  wire _25268_;
  wire _25269_;
  wire _25270_;
  wire _25271_;
  wire _25272_;
  wire _25273_;
  wire _25274_;
  wire _25275_;
  wire _25276_;
  wire _25277_;
  wire _25278_;
  wire _25279_;
  wire _25280_;
  wire _25281_;
  wire _25282_;
  wire _25283_;
  wire _25284_;
  wire _25285_;
  wire _25286_;
  wire _25287_;
  wire _25288_;
  wire _25289_;
  wire _25290_;
  wire _25291_;
  wire _25292_;
  wire _25293_;
  wire _25294_;
  wire _25295_;
  wire _25296_;
  wire _25297_;
  wire _25298_;
  wire _25299_;
  wire _25300_;
  wire _25301_;
  wire _25302_;
  wire _25303_;
  wire _25304_;
  wire _25305_;
  wire _25306_;
  wire _25307_;
  wire _25308_;
  wire _25309_;
  wire _25310_;
  wire _25311_;
  wire _25312_;
  wire _25313_;
  wire _25314_;
  wire _25315_;
  wire _25316_;
  wire _25317_;
  wire _25318_;
  wire _25319_;
  wire _25320_;
  wire _25321_;
  wire _25322_;
  wire _25323_;
  wire _25324_;
  wire _25325_;
  wire _25326_;
  wire _25327_;
  wire _25328_;
  wire _25329_;
  wire _25330_;
  wire _25331_;
  wire _25332_;
  wire _25333_;
  wire _25334_;
  wire _25335_;
  wire _25336_;
  wire _25337_;
  wire _25338_;
  wire _25339_;
  wire _25340_;
  wire _25341_;
  wire _25342_;
  wire _25343_;
  wire _25344_;
  wire _25345_;
  wire _25346_;
  wire _25347_;
  wire _25348_;
  wire _25349_;
  wire _25350_;
  wire _25351_;
  wire _25352_;
  wire _25353_;
  wire _25354_;
  wire _25355_;
  wire _25356_;
  wire _25357_;
  wire _25358_;
  wire _25359_;
  wire _25360_;
  wire _25361_;
  wire _25362_;
  wire _25363_;
  wire _25364_;
  wire _25365_;
  wire _25366_;
  wire _25367_;
  wire _25368_;
  wire _25369_;
  wire _25370_;
  wire _25371_;
  wire _25372_;
  wire _25373_;
  wire _25374_;
  wire _25375_;
  wire _25376_;
  wire _25377_;
  wire _25378_;
  wire _25379_;
  wire _25380_;
  wire _25381_;
  wire _25382_;
  wire _25383_;
  wire _25384_;
  wire _25385_;
  wire _25386_;
  wire _25387_;
  wire _25388_;
  wire _25389_;
  wire _25390_;
  wire _25391_;
  wire _25392_;
  wire _25393_;
  wire _25394_;
  wire _25395_;
  wire _25396_;
  wire _25397_;
  wire _25398_;
  wire _25399_;
  wire _25400_;
  wire _25401_;
  wire _25402_;
  wire _25403_;
  wire _25404_;
  wire _25405_;
  wire _25406_;
  wire _25407_;
  wire _25408_;
  wire _25409_;
  wire _25410_;
  wire _25411_;
  wire _25412_;
  wire _25413_;
  wire _25414_;
  wire _25415_;
  wire _25416_;
  wire _25417_;
  wire _25418_;
  wire _25419_;
  wire _25420_;
  wire _25421_;
  wire _25422_;
  wire _25423_;
  wire _25424_;
  wire _25425_;
  wire _25426_;
  wire _25427_;
  wire _25428_;
  wire _25429_;
  wire _25430_;
  wire _25431_;
  wire _25432_;
  wire _25433_;
  wire _25434_;
  wire _25435_;
  wire _25436_;
  wire _25437_;
  wire _25438_;
  wire _25439_;
  wire _25440_;
  wire _25441_;
  wire _25442_;
  wire _25443_;
  wire _25444_;
  wire _25445_;
  wire _25446_;
  wire _25447_;
  wire _25448_;
  wire _25449_;
  wire _25450_;
  wire _25451_;
  wire _25452_;
  wire _25453_;
  wire _25454_;
  wire _25455_;
  wire _25456_;
  wire _25457_;
  wire _25458_;
  wire _25459_;
  wire _25460_;
  wire _25461_;
  wire _25462_;
  wire _25463_;
  wire _25464_;
  wire _25465_;
  wire _25466_;
  wire _25467_;
  wire _25468_;
  wire _25469_;
  wire _25470_;
  wire _25471_;
  wire _25472_;
  wire _25473_;
  wire _25474_;
  wire _25475_;
  wire _25476_;
  wire _25477_;
  wire _25478_;
  wire _25479_;
  wire _25480_;
  wire _25481_;
  wire _25482_;
  wire _25483_;
  wire _25484_;
  wire _25485_;
  wire _25486_;
  wire _25487_;
  wire _25488_;
  wire _25489_;
  wire _25490_;
  wire _25491_;
  wire _25492_;
  wire _25493_;
  wire _25494_;
  wire _25495_;
  wire _25496_;
  wire _25497_;
  wire _25498_;
  wire _25499_;
  wire _25500_;
  wire _25501_;
  wire _25502_;
  wire _25503_;
  wire _25504_;
  wire _25505_;
  wire _25506_;
  wire _25507_;
  wire _25508_;
  wire _25509_;
  wire _25510_;
  wire _25511_;
  wire _25512_;
  wire _25513_;
  wire _25514_;
  wire _25515_;
  wire _25516_;
  wire _25517_;
  wire _25518_;
  wire _25519_;
  wire _25520_;
  wire _25521_;
  wire _25522_;
  wire _25523_;
  wire _25524_;
  wire _25525_;
  wire _25526_;
  wire _25527_;
  wire _25528_;
  wire _25529_;
  wire _25530_;
  wire _25531_;
  wire _25532_;
  wire _25533_;
  wire _25534_;
  wire _25535_;
  wire _25536_;
  wire _25537_;
  wire _25538_;
  wire _25539_;
  wire _25540_;
  wire _25541_;
  wire _25542_;
  wire _25543_;
  wire _25544_;
  wire _25545_;
  wire _25546_;
  wire _25547_;
  wire _25548_;
  wire _25549_;
  wire _25550_;
  wire _25551_;
  wire _25552_;
  wire _25553_;
  wire _25554_;
  wire _25555_;
  wire _25556_;
  wire _25557_;
  wire _25558_;
  wire _25559_;
  wire _25560_;
  wire _25561_;
  wire _25562_;
  wire _25563_;
  wire _25564_;
  wire _25565_;
  wire _25566_;
  wire _25567_;
  wire _25568_;
  wire _25569_;
  wire _25570_;
  wire _25571_;
  wire _25572_;
  wire _25573_;
  wire _25574_;
  wire _25575_;
  wire _25576_;
  wire _25577_;
  wire _25578_;
  wire _25579_;
  wire _25580_;
  wire _25581_;
  wire _25582_;
  wire _25583_;
  wire _25584_;
  wire _25585_;
  wire _25586_;
  wire _25587_;
  wire _25588_;
  wire _25589_;
  wire _25590_;
  wire _25591_;
  wire _25592_;
  wire _25593_;
  wire _25594_;
  wire _25595_;
  wire _25596_;
  wire _25597_;
  wire _25598_;
  wire _25599_;
  wire _25600_;
  wire _25601_;
  wire _25602_;
  wire _25603_;
  wire _25604_;
  wire _25605_;
  wire _25606_;
  wire _25607_;
  wire _25608_;
  wire _25609_;
  wire _25610_;
  wire _25611_;
  wire _25612_;
  wire _25613_;
  wire _25614_;
  wire _25615_;
  wire _25616_;
  wire _25617_;
  wire _25618_;
  wire _25619_;
  wire _25620_;
  wire _25621_;
  wire _25622_;
  wire _25623_;
  wire _25624_;
  wire _25625_;
  wire _25626_;
  wire _25627_;
  wire _25628_;
  wire _25629_;
  wire _25630_;
  wire _25631_;
  wire _25632_;
  wire _25633_;
  wire _25634_;
  wire _25635_;
  wire _25636_;
  wire _25637_;
  wire _25638_;
  wire _25639_;
  wire _25640_;
  wire _25641_;
  wire _25642_;
  wire _25643_;
  wire _25644_;
  wire _25645_;
  wire _25646_;
  wire _25647_;
  wire _25648_;
  wire _25649_;
  wire _25650_;
  wire _25651_;
  wire _25652_;
  wire _25653_;
  wire _25654_;
  wire _25655_;
  wire _25656_;
  wire _25657_;
  wire _25658_;
  wire _25659_;
  wire _25660_;
  wire _25661_;
  wire _25662_;
  wire _25663_;
  wire _25664_;
  wire _25665_;
  wire _25666_;
  wire _25667_;
  wire _25668_;
  wire _25669_;
  wire _25670_;
  wire _25671_;
  wire _25672_;
  wire _25673_;
  wire _25674_;
  wire _25675_;
  wire _25676_;
  wire _25677_;
  wire _25678_;
  wire _25679_;
  wire _25680_;
  wire _25681_;
  wire _25682_;
  wire _25683_;
  wire _25684_;
  wire _25685_;
  wire _25686_;
  wire _25687_;
  wire _25688_;
  wire _25689_;
  wire _25690_;
  wire _25691_;
  wire _25692_;
  wire _25693_;
  wire _25694_;
  wire _25695_;
  wire _25696_;
  wire _25697_;
  wire _25698_;
  wire _25699_;
  wire _25700_;
  wire _25701_;
  wire _25702_;
  wire _25703_;
  wire _25704_;
  wire _25705_;
  wire _25706_;
  wire _25707_;
  wire _25708_;
  wire _25709_;
  wire _25710_;
  wire _25711_;
  wire _25712_;
  wire _25713_;
  wire _25714_;
  wire _25715_;
  wire _25716_;
  wire _25717_;
  wire _25718_;
  wire _25719_;
  wire _25720_;
  wire _25721_;
  wire _25722_;
  wire _25723_;
  wire _25724_;
  wire _25725_;
  wire _25726_;
  wire _25727_;
  wire _25728_;
  wire _25729_;
  wire _25730_;
  wire _25731_;
  wire _25732_;
  wire _25733_;
  wire _25734_;
  wire _25735_;
  wire _25736_;
  wire _25737_;
  wire _25738_;
  wire _25739_;
  wire _25740_;
  wire _25741_;
  wire _25742_;
  wire _25743_;
  wire _25744_;
  wire _25745_;
  wire _25746_;
  wire _25747_;
  wire _25748_;
  wire _25749_;
  wire _25750_;
  wire _25751_;
  wire _25752_;
  wire _25753_;
  wire _25754_;
  wire _25755_;
  wire _25756_;
  wire _25757_;
  wire _25758_;
  wire _25759_;
  wire _25760_;
  wire _25761_;
  wire _25762_;
  wire _25763_;
  wire _25764_;
  wire _25765_;
  wire _25766_;
  wire _25767_;
  wire _25768_;
  wire _25769_;
  wire _25770_;
  wire _25771_;
  wire _25772_;
  wire _25773_;
  wire _25774_;
  wire _25775_;
  wire _25776_;
  wire _25777_;
  wire _25778_;
  wire _25779_;
  wire _25780_;
  wire _25781_;
  wire _25782_;
  wire _25783_;
  wire _25784_;
  wire _25785_;
  wire _25786_;
  wire _25787_;
  wire _25788_;
  wire _25789_;
  wire _25790_;
  wire _25791_;
  wire _25792_;
  wire _25793_;
  wire _25794_;
  wire _25795_;
  wire _25796_;
  wire _25797_;
  wire _25798_;
  wire _25799_;
  wire _25800_;
  wire _25801_;
  wire _25802_;
  wire _25803_;
  wire _25804_;
  wire _25805_;
  wire _25806_;
  wire _25807_;
  wire _25808_;
  wire _25809_;
  wire _25810_;
  wire _25811_;
  wire _25812_;
  wire _25813_;
  wire _25814_;
  wire _25815_;
  wire _25816_;
  wire _25817_;
  wire _25818_;
  wire _25819_;
  wire _25820_;
  wire _25821_;
  wire _25822_;
  wire _25823_;
  wire _25824_;
  wire _25825_;
  wire _25826_;
  wire _25827_;
  wire _25828_;
  wire _25829_;
  wire _25830_;
  wire _25831_;
  wire _25832_;
  wire _25833_;
  wire _25834_;
  wire _25835_;
  wire _25836_;
  wire _25837_;
  wire _25838_;
  wire _25839_;
  wire _25840_;
  wire _25841_;
  wire _25842_;
  wire _25843_;
  wire _25844_;
  wire _25845_;
  wire _25846_;
  wire _25847_;
  wire _25848_;
  wire _25849_;
  wire _25850_;
  wire _25851_;
  wire _25852_;
  wire _25853_;
  wire _25854_;
  wire _25855_;
  wire _25856_;
  wire _25857_;
  wire _25858_;
  wire _25859_;
  wire _25860_;
  wire _25861_;
  wire _25862_;
  wire _25863_;
  wire _25864_;
  wire _25865_;
  wire _25866_;
  wire _25867_;
  wire _25868_;
  wire _25869_;
  wire _25870_;
  wire _25871_;
  wire _25872_;
  wire _25873_;
  wire _25874_;
  wire _25875_;
  wire _25876_;
  wire _25877_;
  wire _25878_;
  wire _25879_;
  wire _25880_;
  wire _25881_;
  wire _25882_;
  wire _25883_;
  wire _25884_;
  wire _25885_;
  wire _25886_;
  wire _25887_;
  wire _25888_;
  wire _25889_;
  wire _25890_;
  wire _25891_;
  wire _25892_;
  wire _25893_;
  wire _25894_;
  wire _25895_;
  wire _25896_;
  wire _25897_;
  wire _25898_;
  wire _25899_;
  wire _25900_;
  wire _25901_;
  wire _25902_;
  wire _25903_;
  wire _25904_;
  wire _25905_;
  wire _25906_;
  wire _25907_;
  wire _25908_;
  wire _25909_;
  wire _25910_;
  wire _25911_;
  wire _25912_;
  wire _25913_;
  wire _25914_;
  wire _25915_;
  wire _25916_;
  wire _25917_;
  wire _25918_;
  wire _25919_;
  wire _25920_;
  wire _25921_;
  wire _25922_;
  wire _25923_;
  wire _25924_;
  wire _25925_;
  wire _25926_;
  wire _25927_;
  wire _25928_;
  wire _25929_;
  wire _25930_;
  wire _25931_;
  wire _25932_;
  wire _25933_;
  wire _25934_;
  wire _25935_;
  wire _25936_;
  wire _25937_;
  wire _25938_;
  wire _25939_;
  wire _25940_;
  wire _25941_;
  wire _25942_;
  wire _25943_;
  wire _25944_;
  wire _25945_;
  wire _25946_;
  wire _25947_;
  wire _25948_;
  wire _25949_;
  wire _25950_;
  wire _25951_;
  wire _25952_;
  wire _25953_;
  wire _25954_;
  wire _25955_;
  wire _25956_;
  wire _25957_;
  wire _25958_;
  wire _25959_;
  wire _25960_;
  wire _25961_;
  wire _25962_;
  wire _25963_;
  wire _25964_;
  wire _25965_;
  wire _25966_;
  wire _25967_;
  wire _25968_;
  wire _25969_;
  wire _25970_;
  wire _25971_;
  wire _25972_;
  wire _25973_;
  wire _25974_;
  wire _25975_;
  wire _25976_;
  wire _25977_;
  wire _25978_;
  wire _25979_;
  wire _25980_;
  wire _25981_;
  wire _25982_;
  wire _25983_;
  wire _25984_;
  wire _25985_;
  wire _25986_;
  wire _25987_;
  wire _25988_;
  wire _25989_;
  wire _25990_;
  wire _25991_;
  wire _25992_;
  wire _25993_;
  wire _25994_;
  wire _25995_;
  wire _25996_;
  wire _25997_;
  wire _25998_;
  wire _25999_;
  wire _26000_;
  wire _26001_;
  wire _26002_;
  wire _26003_;
  wire _26004_;
  wire _26005_;
  wire _26006_;
  wire _26007_;
  wire _26008_;
  wire _26009_;
  wire _26010_;
  wire _26011_;
  wire _26012_;
  wire _26013_;
  wire _26014_;
  wire _26015_;
  wire _26016_;
  wire _26017_;
  wire _26018_;
  wire _26019_;
  wire _26020_;
  wire _26021_;
  wire _26022_;
  wire _26023_;
  wire _26024_;
  wire _26025_;
  wire _26026_;
  wire _26027_;
  wire _26028_;
  wire _26029_;
  wire _26030_;
  wire _26031_;
  wire _26032_;
  wire _26033_;
  wire _26034_;
  wire _26035_;
  wire _26036_;
  wire _26037_;
  wire _26038_;
  wire _26039_;
  wire _26040_;
  wire _26041_;
  wire _26042_;
  wire _26043_;
  wire _26044_;
  wire _26045_;
  wire _26046_;
  wire _26047_;
  wire _26048_;
  wire _26049_;
  wire _26050_;
  wire _26051_;
  wire _26052_;
  wire _26053_;
  wire _26054_;
  wire _26055_;
  wire _26056_;
  wire _26057_;
  wire _26058_;
  wire _26059_;
  wire _26060_;
  wire _26061_;
  wire _26062_;
  wire _26063_;
  wire _26064_;
  wire _26065_;
  wire _26066_;
  wire _26067_;
  wire _26068_;
  wire _26069_;
  wire _26070_;
  wire _26071_;
  wire _26072_;
  wire _26073_;
  wire _26074_;
  wire _26075_;
  wire _26076_;
  wire _26077_;
  wire _26078_;
  wire _26079_;
  wire _26080_;
  wire _26081_;
  wire _26082_;
  wire _26083_;
  wire _26084_;
  wire _26085_;
  wire _26086_;
  wire _26087_;
  wire _26088_;
  wire _26089_;
  wire _26090_;
  wire _26091_;
  wire _26092_;
  wire _26093_;
  wire _26094_;
  wire _26095_;
  wire _26096_;
  wire _26097_;
  wire _26098_;
  wire _26099_;
  wire _26100_;
  wire _26101_;
  wire _26102_;
  wire _26103_;
  wire _26104_;
  wire _26105_;
  wire _26106_;
  wire _26107_;
  wire _26108_;
  wire _26109_;
  wire _26110_;
  wire _26111_;
  wire _26112_;
  wire _26113_;
  wire _26114_;
  wire _26115_;
  wire _26116_;
  wire _26117_;
  wire _26118_;
  wire _26119_;
  wire _26120_;
  wire _26121_;
  wire _26122_;
  wire _26123_;
  wire _26124_;
  wire _26125_;
  wire _26126_;
  wire _26127_;
  wire _26128_;
  wire _26129_;
  wire _26130_;
  wire _26131_;
  wire _26132_;
  wire _26133_;
  wire _26134_;
  wire _26135_;
  wire _26136_;
  wire _26137_;
  wire _26138_;
  wire _26139_;
  wire _26140_;
  wire _26141_;
  wire _26142_;
  wire _26143_;
  wire _26144_;
  wire _26145_;
  wire _26146_;
  wire _26147_;
  wire _26148_;
  wire _26149_;
  wire _26150_;
  wire _26151_;
  wire _26152_;
  wire _26153_;
  wire _26154_;
  wire _26155_;
  wire _26156_;
  wire _26157_;
  wire _26158_;
  wire _26159_;
  wire _26160_;
  wire _26161_;
  wire _26162_;
  wire _26163_;
  wire _26164_;
  wire _26165_;
  wire _26166_;
  wire _26167_;
  wire _26168_;
  wire _26169_;
  wire _26170_;
  wire _26171_;
  wire _26172_;
  wire _26173_;
  wire _26174_;
  wire _26175_;
  wire _26176_;
  wire _26177_;
  wire _26178_;
  wire _26179_;
  wire _26180_;
  wire _26181_;
  wire _26182_;
  wire _26183_;
  wire _26184_;
  wire _26185_;
  wire _26186_;
  wire _26187_;
  wire _26188_;
  wire _26189_;
  wire _26190_;
  wire _26191_;
  wire _26192_;
  wire _26193_;
  wire _26194_;
  wire _26195_;
  wire _26196_;
  wire _26197_;
  wire _26198_;
  wire _26199_;
  wire _26200_;
  wire _26201_;
  wire _26202_;
  wire _26203_;
  wire _26204_;
  wire _26205_;
  wire _26206_;
  wire _26207_;
  wire _26208_;
  wire _26209_;
  wire _26210_;
  wire _26211_;
  wire _26212_;
  wire _26213_;
  wire _26214_;
  wire _26215_;
  wire _26216_;
  wire _26217_;
  wire _26218_;
  wire _26219_;
  wire _26220_;
  wire _26221_;
  wire _26222_;
  wire _26223_;
  wire _26224_;
  wire _26225_;
  wire _26226_;
  wire _26227_;
  wire _26228_;
  wire _26229_;
  wire _26230_;
  wire _26231_;
  wire _26232_;
  wire _26233_;
  wire _26234_;
  wire _26235_;
  wire _26236_;
  wire _26237_;
  wire _26238_;
  wire _26239_;
  wire _26240_;
  wire _26241_;
  wire _26242_;
  wire _26243_;
  wire _26244_;
  wire _26245_;
  wire _26246_;
  wire _26247_;
  wire _26248_;
  wire _26249_;
  wire _26250_;
  wire _26251_;
  wire _26252_;
  wire _26253_;
  wire _26254_;
  wire _26255_;
  wire _26256_;
  wire _26257_;
  wire _26258_;
  wire _26259_;
  wire _26260_;
  wire _26261_;
  wire _26262_;
  wire _26263_;
  wire _26264_;
  wire _26265_;
  wire _26266_;
  wire _26267_;
  wire _26268_;
  wire _26269_;
  wire _26270_;
  wire _26271_;
  wire _26272_;
  wire _26273_;
  wire _26274_;
  wire _26275_;
  wire _26276_;
  wire _26277_;
  wire _26278_;
  wire _26279_;
  wire _26280_;
  wire _26281_;
  wire _26282_;
  wire _26283_;
  wire _26284_;
  wire _26285_;
  wire _26286_;
  wire _26287_;
  wire _26288_;
  wire _26289_;
  wire _26290_;
  wire _26291_;
  wire _26292_;
  wire _26293_;
  wire _26294_;
  wire _26295_;
  wire _26296_;
  wire _26297_;
  wire _26298_;
  wire _26299_;
  wire _26300_;
  wire _26301_;
  wire _26302_;
  wire _26303_;
  wire _26304_;
  wire _26305_;
  wire _26306_;
  wire _26307_;
  wire _26308_;
  wire _26309_;
  wire _26310_;
  wire _26311_;
  wire _26312_;
  wire _26313_;
  wire _26314_;
  wire _26315_;
  wire _26316_;
  wire _26317_;
  wire _26318_;
  wire _26319_;
  wire _26320_;
  wire _26321_;
  wire _26322_;
  wire _26323_;
  wire _26324_;
  wire _26325_;
  wire _26326_;
  wire _26327_;
  wire _26328_;
  wire _26329_;
  wire _26330_;
  wire _26331_;
  wire _26332_;
  wire _26333_;
  wire _26334_;
  wire _26335_;
  wire _26336_;
  wire _26337_;
  wire _26338_;
  wire _26339_;
  wire _26340_;
  wire _26341_;
  wire _26342_;
  wire _26343_;
  wire _26344_;
  wire _26345_;
  wire _26346_;
  wire _26347_;
  wire _26348_;
  wire _26349_;
  wire _26350_;
  wire _26351_;
  wire _26352_;
  wire _26353_;
  wire _26354_;
  wire _26355_;
  wire _26356_;
  wire _26357_;
  wire _26358_;
  wire _26359_;
  wire _26360_;
  wire _26361_;
  wire _26362_;
  wire _26363_;
  wire _26364_;
  wire _26365_;
  wire _26366_;
  wire _26367_;
  wire _26368_;
  wire _26369_;
  wire _26370_;
  wire _26371_;
  wire _26372_;
  wire _26373_;
  wire _26374_;
  wire _26375_;
  wire _26376_;
  wire _26377_;
  wire _26378_;
  wire _26379_;
  wire _26380_;
  wire _26381_;
  wire _26382_;
  wire _26383_;
  wire _26384_;
  wire _26385_;
  wire _26386_;
  wire _26387_;
  wire _26388_;
  wire _26389_;
  wire _26390_;
  wire _26391_;
  wire _26392_;
  wire _26393_;
  wire _26394_;
  wire _26395_;
  wire _26396_;
  wire _26397_;
  wire _26398_;
  wire _26399_;
  wire _26400_;
  wire _26401_;
  wire _26402_;
  wire _26403_;
  wire _26404_;
  wire _26405_;
  wire _26406_;
  wire _26407_;
  wire _26408_;
  wire _26409_;
  wire _26410_;
  wire _26411_;
  wire _26412_;
  wire _26413_;
  wire _26414_;
  wire _26415_;
  wire _26416_;
  wire _26417_;
  wire _26418_;
  wire _26419_;
  wire _26420_;
  wire _26421_;
  wire _26422_;
  wire _26423_;
  wire _26424_;
  wire _26425_;
  wire _26426_;
  wire _26427_;
  wire _26428_;
  wire _26429_;
  wire _26430_;
  wire _26431_;
  wire _26432_;
  wire _26433_;
  wire _26434_;
  wire _26435_;
  wire _26436_;
  wire _26437_;
  wire _26438_;
  wire _26439_;
  wire _26440_;
  wire _26441_;
  wire _26442_;
  wire _26443_;
  wire _26444_;
  wire _26445_;
  wire _26446_;
  wire _26447_;
  wire _26448_;
  wire _26449_;
  wire _26450_;
  wire _26451_;
  wire _26452_;
  wire _26453_;
  wire _26454_;
  wire _26455_;
  wire _26456_;
  wire _26457_;
  wire _26458_;
  wire _26459_;
  wire _26460_;
  wire _26461_;
  wire _26462_;
  wire _26463_;
  wire _26464_;
  wire _26465_;
  wire _26466_;
  wire _26467_;
  wire _26468_;
  wire _26469_;
  wire _26470_;
  wire _26471_;
  wire _26472_;
  wire _26473_;
  wire _26474_;
  wire _26475_;
  wire _26476_;
  wire _26477_;
  wire _26478_;
  wire _26479_;
  wire _26480_;
  wire _26481_;
  wire _26482_;
  wire _26483_;
  wire _26484_;
  wire _26485_;
  wire _26486_;
  wire _26487_;
  wire _26488_;
  wire _26489_;
  wire _26490_;
  wire _26491_;
  wire _26492_;
  wire _26493_;
  wire _26494_;
  wire _26495_;
  wire _26496_;
  wire _26497_;
  wire _26498_;
  wire _26499_;
  wire _26500_;
  wire _26501_;
  wire _26502_;
  wire _26503_;
  wire _26504_;
  wire _26505_;
  wire _26506_;
  wire _26507_;
  wire _26508_;
  wire _26509_;
  wire _26510_;
  wire _26511_;
  wire _26512_;
  wire _26513_;
  wire _26514_;
  wire _26515_;
  wire _26516_;
  wire _26517_;
  wire _26518_;
  wire _26519_;
  wire _26520_;
  wire _26521_;
  wire _26522_;
  wire _26523_;
  wire _26524_;
  wire _26525_;
  wire _26526_;
  wire _26527_;
  wire _26528_;
  wire _26529_;
  wire _26530_;
  wire _26531_;
  wire _26532_;
  wire _26533_;
  wire _26534_;
  wire _26535_;
  wire _26536_;
  wire _26537_;
  wire _26538_;
  wire _26539_;
  wire _26540_;
  wire _26541_;
  wire _26542_;
  wire _26543_;
  wire _26544_;
  wire _26545_;
  wire _26546_;
  wire _26547_;
  wire _26548_;
  wire _26549_;
  wire _26550_;
  wire _26551_;
  wire _26552_;
  wire _26553_;
  wire _26554_;
  wire _26555_;
  wire _26556_;
  wire _26557_;
  wire _26558_;
  wire _26559_;
  wire _26560_;
  wire _26561_;
  wire _26562_;
  wire _26563_;
  wire _26564_;
  wire _26565_;
  wire _26566_;
  wire _26567_;
  wire _26568_;
  wire _26569_;
  wire _26570_;
  wire _26571_;
  wire _26572_;
  wire _26573_;
  wire _26574_;
  wire _26575_;
  wire _26576_;
  wire _26577_;
  wire _26578_;
  wire _26579_;
  wire _26580_;
  wire _26581_;
  wire _26582_;
  wire _26583_;
  wire _26584_;
  wire _26585_;
  wire _26586_;
  wire _26587_;
  wire _26588_;
  wire _26589_;
  wire _26590_;
  wire _26591_;
  wire _26592_;
  wire _26593_;
  wire _26594_;
  wire _26595_;
  wire _26596_;
  wire _26597_;
  wire _26598_;
  wire _26599_;
  wire _26600_;
  wire _26601_;
  wire _26602_;
  wire _26603_;
  wire _26604_;
  wire _26605_;
  wire _26606_;
  wire _26607_;
  wire _26608_;
  wire _26609_;
  wire _26610_;
  wire _26611_;
  wire _26612_;
  wire _26613_;
  wire _26614_;
  wire _26615_;
  wire _26616_;
  wire _26617_;
  wire _26618_;
  wire _26619_;
  wire _26620_;
  wire _26621_;
  wire _26622_;
  wire _26623_;
  wire _26624_;
  wire _26625_;
  wire _26626_;
  wire _26627_;
  wire _26628_;
  wire _26629_;
  wire _26630_;
  wire _26631_;
  wire _26632_;
  wire _26633_;
  wire _26634_;
  wire _26635_;
  wire _26636_;
  wire _26637_;
  wire _26638_;
  wire _26639_;
  wire _26640_;
  wire _26641_;
  wire _26642_;
  wire _26643_;
  wire _26644_;
  wire _26645_;
  wire _26646_;
  wire _26647_;
  wire _26648_;
  wire _26649_;
  wire _26650_;
  wire _26651_;
  wire _26652_;
  wire _26653_;
  wire _26654_;
  wire _26655_;
  wire _26656_;
  wire _26657_;
  wire _26658_;
  wire _26659_;
  wire _26660_;
  wire _26661_;
  wire _26662_;
  wire _26663_;
  wire _26664_;
  wire _26665_;
  wire _26666_;
  wire _26667_;
  wire _26668_;
  wire _26669_;
  wire _26670_;
  wire _26671_;
  wire _26672_;
  wire _26673_;
  wire _26674_;
  wire _26675_;
  wire _26676_;
  wire _26677_;
  wire _26678_;
  wire _26679_;
  wire _26680_;
  wire _26681_;
  wire _26682_;
  wire _26683_;
  wire _26684_;
  wire _26685_;
  wire _26686_;
  wire _26687_;
  wire _26688_;
  wire _26689_;
  wire _26690_;
  wire _26691_;
  wire _26692_;
  wire _26693_;
  wire _26694_;
  wire _26695_;
  wire _26696_;
  wire _26697_;
  wire _26698_;
  wire _26699_;
  wire _26700_;
  wire _26701_;
  wire _26702_;
  wire _26703_;
  wire _26704_;
  wire _26705_;
  wire _26706_;
  wire _26707_;
  wire _26708_;
  wire _26709_;
  wire _26710_;
  wire _26711_;
  wire _26712_;
  wire _26713_;
  wire _26714_;
  wire _26715_;
  wire _26716_;
  wire _26717_;
  wire _26718_;
  wire _26719_;
  wire _26720_;
  wire _26721_;
  wire _26722_;
  wire _26723_;
  wire _26724_;
  wire _26725_;
  wire _26726_;
  wire _26727_;
  wire _26728_;
  wire _26729_;
  wire _26730_;
  wire _26731_;
  wire _26732_;
  wire _26733_;
  wire _26734_;
  wire _26735_;
  wire _26736_;
  wire _26737_;
  wire _26738_;
  wire _26739_;
  wire _26740_;
  wire _26741_;
  wire _26742_;
  wire _26743_;
  wire _26744_;
  wire _26745_;
  wire _26746_;
  wire _26747_;
  wire _26748_;
  wire _26749_;
  wire _26750_;
  wire _26751_;
  wire _26752_;
  wire _26753_;
  wire _26754_;
  wire _26755_;
  wire _26756_;
  wire _26757_;
  wire _26758_;
  wire _26759_;
  wire _26760_;
  wire _26761_;
  wire _26762_;
  wire _26763_;
  wire _26764_;
  wire _26765_;
  wire _26766_;
  wire _26767_;
  wire _26768_;
  wire _26769_;
  wire _26770_;
  wire _26771_;
  wire _26772_;
  wire _26773_;
  wire _26774_;
  wire _26775_;
  wire _26776_;
  wire _26777_;
  wire _26778_;
  wire _26779_;
  wire _26780_;
  wire _26781_;
  wire _26782_;
  wire _26783_;
  wire _26784_;
  wire _26785_;
  wire _26786_;
  wire _26787_;
  wire _26788_;
  wire _26789_;
  wire _26790_;
  wire _26791_;
  wire _26792_;
  wire _26793_;
  wire _26794_;
  wire _26795_;
  wire _26796_;
  wire _26797_;
  wire _26798_;
  wire _26799_;
  wire _26800_;
  wire _26801_;
  wire _26802_;
  wire _26803_;
  wire _26804_;
  wire _26805_;
  wire _26806_;
  wire _26807_;
  wire _26808_;
  wire _26809_;
  wire _26810_;
  wire _26811_;
  wire _26812_;
  wire _26813_;
  wire _26814_;
  wire _26815_;
  wire _26816_;
  wire _26817_;
  wire _26818_;
  wire _26819_;
  wire _26820_;
  wire _26821_;
  wire _26822_;
  wire _26823_;
  wire _26824_;
  wire _26825_;
  wire _26826_;
  wire _26827_;
  wire _26828_;
  wire _26829_;
  wire _26830_;
  wire _26831_;
  wire _26832_;
  wire _26833_;
  wire _26834_;
  wire _26835_;
  wire _26836_;
  wire _26837_;
  wire _26838_;
  wire _26839_;
  wire _26840_;
  wire _26841_;
  wire _26842_;
  wire _26843_;
  wire _26844_;
  wire _26845_;
  wire _26846_;
  wire _26847_;
  wire _26848_;
  wire _26849_;
  wire _26850_;
  wire _26851_;
  wire _26852_;
  wire _26853_;
  wire _26854_;
  wire _26855_;
  wire _26856_;
  wire _26857_;
  wire _26858_;
  wire _26859_;
  wire _26860_;
  wire _26861_;
  wire _26862_;
  wire _26863_;
  wire _26864_;
  wire _26865_;
  wire _26866_;
  wire _26867_;
  wire _26868_;
  wire _26869_;
  wire _26870_;
  wire _26871_;
  wire _26872_;
  wire _26873_;
  wire _26874_;
  wire _26875_;
  wire _26876_;
  wire _26877_;
  wire _26878_;
  wire _26879_;
  wire _26880_;
  wire _26881_;
  wire _26882_;
  wire _26883_;
  wire _26884_;
  wire _26885_;
  wire _26886_;
  wire _26887_;
  wire _26888_;
  wire _26889_;
  wire _26890_;
  wire _26891_;
  wire _26892_;
  wire _26893_;
  wire _26894_;
  wire _26895_;
  wire _26896_;
  wire _26897_;
  wire _26898_;
  wire _26899_;
  wire _26900_;
  wire _26901_;
  wire _26902_;
  wire _26903_;
  wire _26904_;
  wire _26905_;
  wire _26906_;
  wire _26907_;
  wire _26908_;
  wire _26909_;
  wire _26910_;
  wire _26911_;
  wire _26912_;
  wire _26913_;
  wire _26914_;
  wire _26915_;
  wire _26916_;
  wire _26917_;
  wire _26918_;
  wire _26919_;
  wire _26920_;
  wire _26921_;
  wire _26922_;
  wire _26923_;
  wire _26924_;
  wire _26925_;
  wire _26926_;
  wire _26927_;
  wire _26928_;
  wire _26929_;
  wire _26930_;
  wire _26931_;
  wire _26932_;
  wire _26933_;
  wire _26934_;
  wire _26935_;
  wire _26936_;
  wire _26937_;
  wire _26938_;
  wire _26939_;
  wire _26940_;
  wire _26941_;
  wire _26942_;
  wire _26943_;
  wire _26944_;
  wire _26945_;
  wire _26946_;
  wire _26947_;
  wire _26948_;
  wire _26949_;
  wire _26950_;
  wire _26951_;
  wire _26952_;
  wire _26953_;
  wire _26954_;
  wire _26955_;
  wire _26956_;
  wire _26957_;
  wire _26958_;
  wire _26959_;
  wire _26960_;
  wire _26961_;
  wire _26962_;
  wire _26963_;
  wire _26964_;
  wire _26965_;
  wire _26966_;
  wire _26967_;
  wire _26968_;
  wire _26969_;
  wire _26970_;
  wire _26971_;
  wire _26972_;
  wire _26973_;
  wire _26974_;
  wire _26975_;
  wire _26976_;
  wire _26977_;
  wire _26978_;
  wire _26979_;
  wire _26980_;
  wire _26981_;
  wire _26982_;
  wire _26983_;
  wire _26984_;
  wire _26985_;
  wire _26986_;
  wire _26987_;
  wire _26988_;
  wire _26989_;
  wire _26990_;
  wire _26991_;
  wire _26992_;
  wire _26993_;
  wire _26994_;
  wire _26995_;
  wire _26996_;
  wire _26997_;
  wire _26998_;
  wire _26999_;
  wire _27000_;
  wire _27001_;
  wire _27002_;
  wire _27003_;
  wire _27004_;
  wire _27005_;
  wire _27006_;
  wire _27007_;
  wire _27008_;
  wire _27009_;
  wire _27010_;
  wire _27011_;
  wire _27012_;
  wire _27013_;
  wire _27014_;
  wire _27015_;
  wire _27016_;
  wire _27017_;
  wire _27018_;
  wire _27019_;
  wire _27020_;
  wire _27021_;
  wire _27022_;
  wire _27023_;
  wire _27024_;
  wire _27025_;
  wire _27026_;
  wire _27027_;
  wire _27028_;
  wire _27029_;
  wire _27030_;
  wire _27031_;
  wire _27032_;
  wire _27033_;
  wire _27034_;
  wire _27035_;
  wire _27036_;
  wire _27037_;
  wire _27038_;
  wire _27039_;
  wire _27040_;
  wire _27041_;
  wire _27042_;
  wire _27043_;
  wire _27044_;
  wire _27045_;
  wire _27046_;
  wire _27047_;
  wire _27048_;
  wire _27049_;
  wire _27050_;
  wire _27051_;
  wire _27052_;
  wire _27053_;
  wire _27054_;
  wire _27055_;
  wire _27056_;
  wire _27057_;
  wire _27058_;
  wire _27059_;
  wire _27060_;
  wire _27061_;
  wire _27062_;
  wire _27063_;
  wire _27064_;
  wire _27065_;
  wire _27066_;
  wire _27067_;
  wire _27068_;
  wire _27069_;
  wire _27070_;
  wire _27071_;
  wire _27072_;
  wire _27073_;
  wire _27074_;
  wire _27075_;
  wire _27076_;
  wire _27077_;
  wire _27078_;
  wire _27079_;
  wire _27080_;
  wire _27081_;
  wire _27082_;
  wire _27083_;
  wire _27084_;
  wire _27085_;
  wire _27086_;
  wire _27087_;
  wire _27088_;
  wire _27089_;
  wire _27090_;
  wire _27091_;
  wire _27092_;
  wire _27093_;
  wire _27094_;
  wire _27095_;
  wire _27096_;
  wire _27097_;
  wire _27098_;
  wire _27099_;
  wire _27100_;
  wire _27101_;
  wire _27102_;
  wire _27103_;
  wire _27104_;
  wire _27105_;
  wire _27106_;
  wire _27107_;
  wire _27108_;
  wire _27109_;
  wire _27110_;
  wire _27111_;
  wire _27112_;
  wire _27113_;
  wire _27114_;
  wire _27115_;
  wire _27116_;
  wire _27117_;
  wire _27118_;
  wire _27119_;
  wire _27120_;
  wire _27121_;
  wire _27122_;
  wire _27123_;
  wire _27124_;
  wire _27125_;
  wire _27126_;
  wire _27127_;
  wire _27128_;
  wire _27129_;
  wire _27130_;
  wire _27131_;
  wire _27132_;
  wire _27133_;
  wire _27134_;
  wire _27135_;
  wire _27136_;
  wire _27137_;
  wire _27138_;
  wire _27139_;
  wire _27140_;
  wire _27141_;
  wire _27142_;
  wire _27143_;
  wire _27144_;
  wire _27145_;
  wire _27146_;
  wire _27147_;
  wire _27148_;
  wire _27149_;
  wire _27150_;
  wire _27151_;
  wire _27152_;
  wire _27153_;
  wire _27154_;
  wire _27155_;
  wire _27156_;
  wire _27157_;
  wire _27158_;
  wire _27159_;
  wire _27160_;
  wire _27161_;
  wire _27162_;
  wire _27163_;
  wire _27164_;
  wire _27165_;
  wire _27166_;
  wire _27167_;
  wire _27168_;
  wire _27169_;
  wire _27170_;
  wire _27171_;
  wire _27172_;
  wire _27173_;
  wire _27174_;
  wire _27175_;
  wire _27176_;
  wire _27177_;
  wire _27178_;
  wire _27179_;
  wire _27180_;
  wire _27181_;
  wire _27182_;
  wire _27183_;
  wire _27184_;
  wire _27185_;
  wire _27186_;
  wire _27187_;
  wire _27188_;
  wire _27189_;
  wire _27190_;
  wire _27191_;
  wire _27192_;
  wire _27193_;
  wire _27194_;
  wire _27195_;
  wire _27196_;
  wire _27197_;
  wire _27198_;
  wire _27199_;
  wire _27200_;
  wire _27201_;
  wire _27202_;
  wire _27203_;
  wire _27204_;
  wire _27205_;
  wire _27206_;
  wire _27207_;
  wire _27208_;
  wire _27209_;
  wire _27210_;
  wire _27211_;
  wire _27212_;
  wire _27213_;
  wire _27214_;
  wire _27215_;
  wire _27216_;
  wire _27217_;
  wire _27218_;
  wire _27219_;
  wire _27220_;
  wire _27221_;
  wire _27222_;
  wire _27223_;
  wire _27224_;
  wire _27225_;
  wire _27226_;
  wire _27227_;
  wire _27228_;
  wire _27229_;
  wire _27230_;
  wire _27231_;
  wire _27232_;
  wire _27233_;
  wire _27234_;
  wire _27235_;
  wire _27236_;
  wire _27237_;
  wire _27238_;
  wire _27239_;
  wire _27240_;
  wire _27241_;
  wire _27242_;
  wire _27243_;
  wire _27244_;
  wire _27245_;
  wire _27246_;
  wire _27247_;
  wire _27248_;
  wire _27249_;
  wire _27250_;
  wire _27251_;
  wire _27252_;
  wire _27253_;
  wire _27254_;
  wire _27255_;
  wire _27256_;
  wire _27257_;
  wire _27258_;
  wire _27259_;
  wire _27260_;
  wire _27261_;
  wire _27262_;
  wire _27263_;
  wire _27264_;
  wire _27265_;
  wire _27266_;
  wire _27267_;
  wire _27268_;
  wire _27269_;
  wire _27270_;
  wire _27271_;
  wire _27272_;
  wire _27273_;
  wire _27274_;
  wire _27275_;
  wire _27276_;
  wire _27277_;
  wire _27278_;
  wire _27279_;
  wire _27280_;
  wire _27281_;
  wire _27282_;
  wire _27283_;
  wire _27284_;
  wire _27285_;
  wire _27286_;
  wire _27287_;
  wire _27288_;
  wire _27289_;
  wire _27290_;
  wire _27291_;
  wire _27292_;
  wire _27293_;
  wire _27294_;
  wire _27295_;
  wire _27296_;
  wire _27297_;
  wire _27298_;
  wire _27299_;
  wire _27300_;
  wire _27301_;
  wire _27302_;
  wire _27303_;
  wire _27304_;
  wire _27305_;
  wire _27306_;
  wire _27307_;
  wire _27308_;
  wire _27309_;
  wire _27310_;
  wire _27311_;
  wire _27312_;
  wire _27313_;
  wire _27314_;
  wire _27315_;
  wire _27316_;
  wire _27317_;
  wire _27318_;
  wire _27319_;
  wire _27320_;
  wire _27321_;
  wire _27322_;
  wire _27323_;
  wire _27324_;
  wire _27325_;
  wire _27326_;
  wire _27327_;
  wire _27328_;
  wire _27329_;
  wire _27330_;
  wire _27331_;
  wire _27332_;
  wire _27333_;
  wire _27334_;
  wire _27335_;
  wire _27336_;
  wire _27337_;
  wire _27338_;
  wire _27339_;
  wire _27340_;
  wire _27341_;
  wire _27342_;
  wire _27343_;
  wire _27344_;
  wire _27345_;
  wire _27346_;
  wire _27347_;
  wire _27348_;
  wire _27349_;
  wire _27350_;
  wire _27351_;
  wire _27352_;
  wire _27353_;
  wire _27354_;
  wire _27355_;
  wire _27356_;
  wire _27357_;
  wire _27358_;
  wire _27359_;
  wire _27360_;
  wire _27361_;
  wire _27362_;
  wire _27363_;
  wire _27364_;
  wire _27365_;
  wire _27366_;
  wire _27367_;
  wire _27368_;
  wire _27369_;
  wire _27370_;
  wire _27371_;
  wire _27372_;
  wire _27373_;
  wire _27374_;
  wire _27375_;
  wire _27376_;
  wire _27377_;
  wire _27378_;
  wire _27379_;
  wire _27380_;
  wire _27381_;
  wire _27382_;
  wire _27383_;
  wire _27384_;
  wire _27385_;
  wire _27386_;
  wire _27387_;
  wire _27388_;
  wire _27389_;
  wire _27390_;
  wire _27391_;
  wire _27392_;
  wire _27393_;
  wire _27394_;
  wire _27395_;
  wire _27396_;
  wire _27397_;
  wire _27398_;
  wire _27399_;
  wire _27400_;
  wire _27401_;
  wire _27402_;
  wire _27403_;
  wire _27404_;
  wire _27405_;
  wire _27406_;
  wire _27407_;
  wire _27408_;
  wire _27409_;
  wire _27410_;
  wire _27411_;
  wire _27412_;
  wire _27413_;
  wire _27414_;
  wire _27415_;
  wire _27416_;
  wire _27417_;
  wire _27418_;
  wire _27419_;
  wire _27420_;
  wire _27421_;
  wire _27422_;
  wire _27423_;
  wire _27424_;
  wire _27425_;
  wire _27426_;
  wire _27427_;
  wire _27428_;
  wire _27429_;
  wire _27430_;
  wire _27431_;
  wire _27432_;
  wire _27433_;
  wire _27434_;
  wire _27435_;
  wire _27436_;
  wire _27437_;
  wire _27438_;
  wire _27439_;
  wire _27440_;
  wire _27441_;
  wire _27442_;
  wire _27443_;
  wire _27444_;
  wire _27445_;
  wire _27446_;
  wire _27447_;
  wire _27448_;
  wire _27449_;
  wire _27450_;
  wire _27451_;
  wire _27452_;
  wire _27453_;
  wire _27454_;
  wire _27455_;
  wire _27456_;
  wire _27457_;
  wire _27458_;
  wire _27459_;
  wire _27460_;
  wire _27461_;
  wire _27462_;
  wire _27463_;
  wire _27464_;
  wire _27465_;
  wire _27466_;
  wire _27467_;
  wire _27468_;
  wire _27469_;
  wire _27470_;
  wire _27471_;
  wire _27472_;
  wire _27473_;
  wire _27474_;
  wire _27475_;
  wire _27476_;
  wire _27477_;
  wire _27478_;
  wire _27479_;
  wire _27480_;
  wire _27481_;
  wire _27482_;
  wire _27483_;
  wire _27484_;
  wire _27485_;
  wire _27486_;
  wire _27487_;
  wire _27488_;
  wire _27489_;
  wire _27490_;
  wire _27491_;
  wire _27492_;
  wire _27493_;
  wire _27494_;
  wire _27495_;
  wire _27496_;
  wire _27497_;
  wire _27498_;
  wire _27499_;
  wire _27500_;
  wire _27501_;
  wire _27502_;
  wire _27503_;
  wire _27504_;
  wire _27505_;
  wire _27506_;
  wire _27507_;
  wire _27508_;
  wire _27509_;
  wire _27510_;
  wire _27511_;
  wire _27512_;
  wire _27513_;
  wire _27514_;
  wire _27515_;
  wire _27516_;
  wire _27517_;
  wire _27518_;
  wire _27519_;
  wire _27520_;
  wire _27521_;
  wire _27522_;
  wire _27523_;
  wire _27524_;
  wire _27525_;
  wire _27526_;
  wire _27527_;
  wire _27528_;
  wire _27529_;
  wire _27530_;
  wire _27531_;
  wire _27532_;
  wire _27533_;
  wire _27534_;
  wire _27535_;
  wire _27536_;
  wire _27537_;
  wire _27538_;
  wire _27539_;
  wire _27540_;
  wire _27541_;
  wire _27542_;
  wire _27543_;
  wire _27544_;
  wire _27545_;
  wire _27546_;
  wire _27547_;
  wire _27548_;
  wire _27549_;
  wire _27550_;
  wire _27551_;
  wire _27552_;
  wire _27553_;
  wire _27554_;
  wire _27555_;
  wire _27556_;
  wire _27557_;
  wire _27558_;
  wire _27559_;
  wire _27560_;
  wire _27561_;
  wire _27562_;
  wire _27563_;
  wire _27564_;
  wire _27565_;
  wire _27566_;
  wire _27567_;
  wire _27568_;
  wire _27569_;
  wire _27570_;
  wire _27571_;
  wire _27572_;
  wire _27573_;
  wire _27574_;
  wire _27575_;
  wire _27576_;
  wire _27577_;
  wire _27578_;
  wire _27579_;
  wire _27580_;
  wire _27581_;
  wire _27582_;
  wire _27583_;
  wire _27584_;
  wire _27585_;
  wire _27586_;
  wire _27587_;
  wire _27588_;
  wire _27589_;
  wire _27590_;
  wire _27591_;
  wire _27592_;
  wire _27593_;
  wire _27594_;
  wire _27595_;
  wire _27596_;
  wire _27597_;
  wire _27598_;
  wire _27599_;
  wire _27600_;
  wire _27601_;
  wire _27602_;
  wire _27603_;
  wire _27604_;
  wire _27605_;
  wire _27606_;
  wire _27607_;
  wire _27608_;
  wire _27609_;
  wire _27610_;
  wire _27611_;
  wire _27612_;
  wire _27613_;
  wire _27614_;
  wire _27615_;
  wire _27616_;
  wire _27617_;
  wire _27618_;
  wire _27619_;
  wire _27620_;
  wire _27621_;
  wire _27622_;
  wire _27623_;
  wire _27624_;
  wire _27625_;
  wire _27626_;
  wire _27627_;
  wire _27628_;
  wire _27629_;
  wire _27630_;
  wire _27631_;
  wire _27632_;
  wire _27633_;
  wire _27634_;
  wire _27635_;
  wire _27636_;
  wire _27637_;
  wire _27638_;
  wire _27639_;
  wire _27640_;
  wire _27641_;
  wire _27642_;
  wire _27643_;
  wire _27644_;
  wire _27645_;
  wire _27646_;
  wire _27647_;
  wire _27648_;
  wire _27649_;
  wire _27650_;
  wire _27651_;
  wire _27652_;
  wire _27653_;
  wire _27654_;
  wire _27655_;
  wire _27656_;
  wire _27657_;
  wire _27658_;
  wire _27659_;
  wire _27660_;
  wire _27661_;
  wire _27662_;
  wire _27663_;
  wire _27664_;
  wire _27665_;
  wire _27666_;
  wire _27667_;
  wire _27668_;
  wire _27669_;
  wire _27670_;
  wire _27671_;
  wire _27672_;
  wire _27673_;
  wire _27674_;
  wire _27675_;
  wire _27676_;
  wire _27677_;
  wire _27678_;
  wire _27679_;
  wire _27680_;
  wire _27681_;
  wire _27682_;
  wire _27683_;
  wire _27684_;
  wire _27685_;
  wire _27686_;
  wire _27687_;
  wire _27688_;
  wire _27689_;
  wire _27690_;
  wire _27691_;
  wire _27692_;
  wire _27693_;
  wire _27694_;
  wire _27695_;
  wire _27696_;
  wire _27697_;
  wire _27698_;
  wire _27699_;
  wire _27700_;
  wire _27701_;
  wire _27702_;
  wire _27703_;
  wire _27704_;
  wire _27705_;
  wire _27706_;
  wire _27707_;
  wire _27708_;
  wire _27709_;
  wire _27710_;
  wire _27711_;
  wire _27712_;
  wire _27713_;
  wire _27714_;
  wire _27715_;
  wire _27716_;
  wire _27717_;
  wire _27718_;
  wire _27719_;
  wire _27720_;
  wire _27721_;
  wire _27722_;
  wire _27723_;
  wire _27724_;
  wire _27725_;
  wire _27726_;
  wire _27727_;
  wire _27728_;
  wire _27729_;
  wire _27730_;
  wire _27731_;
  wire _27732_;
  wire _27733_;
  wire _27734_;
  wire _27735_;
  wire _27736_;
  wire _27737_;
  wire _27738_;
  wire _27739_;
  wire _27740_;
  wire _27741_;
  wire _27742_;
  wire _27743_;
  wire _27744_;
  wire _27745_;
  wire _27746_;
  wire _27747_;
  wire _27748_;
  wire _27749_;
  wire _27750_;
  wire _27751_;
  wire _27752_;
  wire _27753_;
  wire _27754_;
  wire _27755_;
  wire _27756_;
  wire _27757_;
  wire _27758_;
  wire _27759_;
  wire _27760_;
  wire _27761_;
  wire _27762_;
  wire _27763_;
  wire _27764_;
  wire _27765_;
  wire _27766_;
  wire _27767_;
  wire _27768_;
  wire _27769_;
  wire _27770_;
  wire _27771_;
  wire _27772_;
  wire _27773_;
  wire _27774_;
  wire _27775_;
  wire _27776_;
  wire _27777_;
  wire _27778_;
  wire _27779_;
  wire _27780_;
  wire _27781_;
  wire _27782_;
  wire _27783_;
  wire _27784_;
  wire _27785_;
  wire _27786_;
  wire _27787_;
  wire _27788_;
  wire _27789_;
  wire _27790_;
  wire _27791_;
  wire _27792_;
  wire _27793_;
  wire _27794_;
  wire _27795_;
  wire _27796_;
  wire _27797_;
  wire _27798_;
  wire _27799_;
  wire _27800_;
  wire _27801_;
  wire _27802_;
  wire _27803_;
  wire _27804_;
  wire _27805_;
  wire _27806_;
  wire _27807_;
  wire _27808_;
  wire _27809_;
  wire _27810_;
  wire _27811_;
  wire _27812_;
  wire _27813_;
  wire _27814_;
  wire _27815_;
  wire _27816_;
  wire _27817_;
  wire _27818_;
  wire _27819_;
  wire _27820_;
  wire _27821_;
  wire _27822_;
  wire _27823_;
  wire _27824_;
  wire _27825_;
  wire _27826_;
  wire _27827_;
  wire _27828_;
  wire _27829_;
  wire _27830_;
  wire _27831_;
  wire _27832_;
  wire _27833_;
  wire _27834_;
  wire _27835_;
  wire _27836_;
  wire _27837_;
  wire _27838_;
  wire _27839_;
  wire _27840_;
  wire _27841_;
  wire _27842_;
  wire _27843_;
  wire _27844_;
  wire _27845_;
  wire _27846_;
  wire _27847_;
  wire _27848_;
  wire _27849_;
  wire _27850_;
  wire _27851_;
  wire _27852_;
  wire _27853_;
  wire _27854_;
  wire _27855_;
  wire _27856_;
  wire _27857_;
  wire _27858_;
  wire _27859_;
  wire _27860_;
  wire _27861_;
  wire _27862_;
  wire _27863_;
  wire _27864_;
  wire _27865_;
  wire _27866_;
  wire _27867_;
  wire _27868_;
  wire _27869_;
  wire _27870_;
  wire _27871_;
  wire _27872_;
  wire _27873_;
  wire _27874_;
  wire _27875_;
  wire _27876_;
  wire _27877_;
  wire _27878_;
  wire _27879_;
  wire _27880_;
  wire _27881_;
  wire _27882_;
  wire _27883_;
  wire _27884_;
  wire _27885_;
  wire _27886_;
  wire _27887_;
  wire _27888_;
  wire _27889_;
  wire _27890_;
  wire _27891_;
  wire _27892_;
  wire _27893_;
  wire _27894_;
  wire _27895_;
  wire _27896_;
  wire _27897_;
  wire _27898_;
  wire _27899_;
  wire _27900_;
  wire _27901_;
  wire _27902_;
  wire _27903_;
  wire _27904_;
  wire _27905_;
  wire _27906_;
  wire _27907_;
  wire _27908_;
  wire _27909_;
  wire _27910_;
  wire _27911_;
  wire _27912_;
  wire _27913_;
  wire _27914_;
  wire _27915_;
  wire _27916_;
  wire _27917_;
  wire _27918_;
  wire _27919_;
  wire _27920_;
  wire _27921_;
  wire _27922_;
  wire _27923_;
  wire _27924_;
  wire _27925_;
  wire _27926_;
  wire _27927_;
  wire _27928_;
  wire _27929_;
  wire _27930_;
  wire _27931_;
  wire _27932_;
  wire _27933_;
  wire _27934_;
  wire _27935_;
  wire _27936_;
  wire _27937_;
  wire _27938_;
  wire _27939_;
  wire _27940_;
  wire _27941_;
  wire _27942_;
  wire _27943_;
  wire _27944_;
  wire _27945_;
  wire _27946_;
  wire _27947_;
  wire _27948_;
  wire _27949_;
  wire _27950_;
  wire _27951_;
  wire _27952_;
  wire _27953_;
  wire _27954_;
  wire _27955_;
  wire _27956_;
  wire _27957_;
  wire _27958_;
  wire _27959_;
  wire _27960_;
  wire _27961_;
  wire _27962_;
  wire _27963_;
  wire _27964_;
  wire _27965_;
  wire _27966_;
  wire _27967_;
  wire _27968_;
  wire _27969_;
  wire _27970_;
  wire _27971_;
  wire _27972_;
  wire _27973_;
  wire _27974_;
  wire _27975_;
  wire _27976_;
  wire _27977_;
  wire _27978_;
  wire _27979_;
  wire _27980_;
  wire _27981_;
  wire _27982_;
  wire _27983_;
  wire _27984_;
  wire _27985_;
  wire _27986_;
  wire _27987_;
  wire _27988_;
  wire _27989_;
  wire _27990_;
  wire _27991_;
  wire _27992_;
  wire _27993_;
  wire _27994_;
  wire _27995_;
  wire _27996_;
  wire _27997_;
  wire _27998_;
  wire _27999_;
  wire _28000_;
  wire _28001_;
  wire _28002_;
  wire _28003_;
  wire _28004_;
  wire _28005_;
  wire _28006_;
  wire _28007_;
  wire _28008_;
  wire _28009_;
  wire _28010_;
  wire _28011_;
  wire _28012_;
  wire _28013_;
  wire _28014_;
  wire _28015_;
  wire _28016_;
  wire _28017_;
  wire _28018_;
  wire _28019_;
  wire _28020_;
  wire _28021_;
  wire _28022_;
  wire _28023_;
  wire _28024_;
  wire _28025_;
  wire _28026_;
  wire _28027_;
  wire _28028_;
  wire _28029_;
  wire _28030_;
  wire _28031_;
  wire _28032_;
  wire _28033_;
  wire _28034_;
  wire _28035_;
  wire _28036_;
  wire _28037_;
  wire _28038_;
  wire _28039_;
  wire _28040_;
  wire _28041_;
  wire _28042_;
  wire _28043_;
  wire _28044_;
  wire _28045_;
  wire _28046_;
  wire _28047_;
  wire _28048_;
  wire _28049_;
  wire _28050_;
  wire _28051_;
  wire _28052_;
  wire _28053_;
  wire _28054_;
  wire _28055_;
  wire _28056_;
  wire _28057_;
  wire _28058_;
  wire _28059_;
  wire _28060_;
  wire _28061_;
  wire _28062_;
  wire _28063_;
  wire _28064_;
  wire _28065_;
  wire _28066_;
  wire _28067_;
  wire _28068_;
  wire _28069_;
  wire _28070_;
  wire _28071_;
  wire _28072_;
  wire _28073_;
  wire _28074_;
  wire _28075_;
  wire _28076_;
  wire _28077_;
  wire _28078_;
  wire _28079_;
  wire _28080_;
  wire _28081_;
  wire _28082_;
  wire _28083_;
  wire _28084_;
  wire _28085_;
  wire _28086_;
  wire _28087_;
  wire _28088_;
  wire _28089_;
  wire _28090_;
  wire _28091_;
  wire _28092_;
  wire _28093_;
  wire _28094_;
  wire _28095_;
  wire _28096_;
  wire _28097_;
  wire _28098_;
  wire _28099_;
  wire _28100_;
  wire _28101_;
  wire _28102_;
  wire _28103_;
  wire _28104_;
  wire _28105_;
  wire _28106_;
  wire _28107_;
  wire _28108_;
  wire _28109_;
  wire _28110_;
  wire _28111_;
  wire _28112_;
  wire _28113_;
  wire _28114_;
  wire _28115_;
  wire _28116_;
  wire _28117_;
  wire _28118_;
  wire _28119_;
  wire _28120_;
  wire _28121_;
  wire _28122_;
  wire _28123_;
  wire _28124_;
  wire _28125_;
  wire _28126_;
  wire _28127_;
  wire _28128_;
  wire _28129_;
  wire _28130_;
  wire _28131_;
  wire _28132_;
  wire _28133_;
  wire _28134_;
  wire _28135_;
  wire _28136_;
  wire _28137_;
  wire _28138_;
  wire _28139_;
  wire _28140_;
  wire _28141_;
  wire _28142_;
  wire _28143_;
  wire _28144_;
  wire _28145_;
  wire _28146_;
  wire _28147_;
  wire _28148_;
  wire _28149_;
  wire _28150_;
  wire _28151_;
  wire _28152_;
  wire _28153_;
  wire _28154_;
  wire _28155_;
  wire _28156_;
  wire _28157_;
  wire _28158_;
  wire _28159_;
  wire _28160_;
  wire _28161_;
  wire _28162_;
  wire _28163_;
  wire _28164_;
  wire _28165_;
  wire _28166_;
  wire _28167_;
  wire _28168_;
  wire _28169_;
  wire _28170_;
  wire _28171_;
  wire _28172_;
  wire _28173_;
  wire _28174_;
  wire _28175_;
  wire _28176_;
  wire _28177_;
  wire _28178_;
  wire _28179_;
  wire _28180_;
  wire _28181_;
  wire _28182_;
  wire _28183_;
  wire _28184_;
  wire _28185_;
  wire _28186_;
  wire _28187_;
  wire _28188_;
  wire _28189_;
  wire _28190_;
  wire _28191_;
  wire _28192_;
  wire _28193_;
  wire _28194_;
  wire _28195_;
  wire _28196_;
  wire _28197_;
  wire _28198_;
  wire _28199_;
  wire _28200_;
  wire _28201_;
  wire _28202_;
  wire _28203_;
  wire _28204_;
  wire _28205_;
  wire _28206_;
  wire _28207_;
  wire _28208_;
  wire _28209_;
  wire _28210_;
  wire _28211_;
  wire _28212_;
  wire _28213_;
  wire _28214_;
  wire _28215_;
  wire _28216_;
  wire _28217_;
  wire _28218_;
  wire _28219_;
  wire _28220_;
  wire _28221_;
  wire _28222_;
  wire _28223_;
  wire _28224_;
  wire _28225_;
  wire _28226_;
  wire _28227_;
  wire _28228_;
  wire _28229_;
  wire _28230_;
  wire _28231_;
  wire _28232_;
  wire _28233_;
  wire _28234_;
  wire _28235_;
  wire _28236_;
  wire _28237_;
  wire _28238_;
  wire _28239_;
  wire _28240_;
  wire _28241_;
  wire _28242_;
  wire _28243_;
  wire _28244_;
  wire _28245_;
  wire _28246_;
  wire _28247_;
  wire _28248_;
  wire _28249_;
  wire _28250_;
  wire _28251_;
  wire _28252_;
  wire _28253_;
  wire _28254_;
  wire _28255_;
  wire _28256_;
  wire _28257_;
  wire _28258_;
  wire _28259_;
  wire _28260_;
  wire _28261_;
  wire _28262_;
  wire _28263_;
  wire _28264_;
  wire _28265_;
  wire _28266_;
  wire _28267_;
  wire _28268_;
  wire _28269_;
  wire _28270_;
  wire _28271_;
  wire _28272_;
  wire _28273_;
  wire _28274_;
  wire _28275_;
  wire _28276_;
  wire _28277_;
  wire _28278_;
  wire _28279_;
  wire _28280_;
  wire _28281_;
  wire _28282_;
  wire _28283_;
  wire _28284_;
  wire _28285_;
  wire _28286_;
  wire _28287_;
  wire _28288_;
  wire _28289_;
  wire _28290_;
  wire _28291_;
  wire _28292_;
  wire _28293_;
  wire _28294_;
  wire _28295_;
  wire _28296_;
  wire _28297_;
  wire _28298_;
  wire _28299_;
  wire _28300_;
  wire _28301_;
  wire _28302_;
  wire _28303_;
  wire _28304_;
  wire _28305_;
  wire _28306_;
  wire _28307_;
  wire _28308_;
  wire _28309_;
  wire _28310_;
  wire _28311_;
  wire _28312_;
  wire _28313_;
  wire _28314_;
  wire _28315_;
  wire _28316_;
  wire _28317_;
  wire _28318_;
  wire _28319_;
  wire _28320_;
  wire _28321_;
  wire _28322_;
  wire _28323_;
  wire _28324_;
  wire _28325_;
  wire _28326_;
  wire _28327_;
  wire _28328_;
  wire _28329_;
  wire _28330_;
  wire _28331_;
  wire _28332_;
  wire _28333_;
  wire _28334_;
  wire _28335_;
  wire _28336_;
  wire _28337_;
  wire _28338_;
  wire _28339_;
  wire _28340_;
  wire _28341_;
  wire _28342_;
  wire _28343_;
  wire _28344_;
  wire _28345_;
  wire _28346_;
  wire _28347_;
  wire _28348_;
  wire _28349_;
  wire _28350_;
  wire _28351_;
  wire _28352_;
  wire _28353_;
  wire _28354_;
  wire _28355_;
  wire _28356_;
  wire _28357_;
  wire _28358_;
  wire _28359_;
  wire _28360_;
  wire _28361_;
  wire _28362_;
  wire _28363_;
  wire _28364_;
  wire _28365_;
  wire _28366_;
  wire _28367_;
  wire _28368_;
  wire _28369_;
  wire _28370_;
  wire _28371_;
  wire _28372_;
  wire _28373_;
  wire _28374_;
  wire _28375_;
  wire _28376_;
  wire _28377_;
  wire _28378_;
  wire _28379_;
  wire _28380_;
  wire _28381_;
  wire _28382_;
  wire _28383_;
  wire _28384_;
  wire _28385_;
  wire _28386_;
  wire _28387_;
  wire _28388_;
  wire _28389_;
  wire _28390_;
  wire _28391_;
  wire _28392_;
  wire _28393_;
  wire _28394_;
  wire _28395_;
  wire _28396_;
  wire _28397_;
  wire _28398_;
  wire _28399_;
  wire _28400_;
  wire _28401_;
  wire _28402_;
  wire _28403_;
  wire _28404_;
  wire _28405_;
  wire _28406_;
  wire _28407_;
  wire _28408_;
  wire _28409_;
  wire _28410_;
  wire _28411_;
  wire _28412_;
  wire _28413_;
  wire _28414_;
  wire _28415_;
  wire _28416_;
  wire _28417_;
  wire _28418_;
  wire _28419_;
  wire _28420_;
  wire _28421_;
  wire _28422_;
  wire _28423_;
  wire _28424_;
  wire _28425_;
  wire _28426_;
  wire _28427_;
  wire _28428_;
  wire _28429_;
  wire _28430_;
  wire _28431_;
  wire _28432_;
  wire _28433_;
  wire _28434_;
  wire _28435_;
  wire _28436_;
  wire _28437_;
  wire _28438_;
  wire _28439_;
  wire _28440_;
  wire _28441_;
  wire _28442_;
  wire _28443_;
  wire _28444_;
  wire _28445_;
  wire _28446_;
  wire _28447_;
  wire _28448_;
  wire _28449_;
  wire _28450_;
  wire _28451_;
  wire _28452_;
  wire _28453_;
  wire _28454_;
  wire _28455_;
  wire _28456_;
  wire _28457_;
  wire _28458_;
  wire _28459_;
  wire _28460_;
  wire _28461_;
  wire _28462_;
  wire _28463_;
  wire _28464_;
  wire _28465_;
  wire _28466_;
  wire _28467_;
  wire _28468_;
  wire _28469_;
  wire _28470_;
  wire _28471_;
  wire _28472_;
  wire _28473_;
  wire _28474_;
  wire _28475_;
  wire _28476_;
  wire _28477_;
  wire _28478_;
  wire _28479_;
  wire _28480_;
  wire _28481_;
  wire _28482_;
  wire _28483_;
  wire _28484_;
  wire _28485_;
  wire _28486_;
  wire _28487_;
  wire _28488_;
  wire _28489_;
  wire _28490_;
  wire _28491_;
  wire _28492_;
  wire _28493_;
  wire _28494_;
  wire _28495_;
  wire _28496_;
  wire _28497_;
  wire _28498_;
  wire _28499_;
  wire _28500_;
  wire _28501_;
  wire _28502_;
  wire _28503_;
  wire _28504_;
  wire _28505_;
  wire _28506_;
  wire _28507_;
  wire _28508_;
  wire _28509_;
  wire _28510_;
  wire _28511_;
  wire _28512_;
  wire _28513_;
  wire _28514_;
  wire _28515_;
  wire _28516_;
  wire _28517_;
  wire _28518_;
  wire _28519_;
  wire _28520_;
  wire _28521_;
  wire _28522_;
  wire _28523_;
  wire _28524_;
  wire _28525_;
  wire _28526_;
  wire _28527_;
  wire _28528_;
  wire _28529_;
  wire _28530_;
  wire _28531_;
  wire _28532_;
  wire _28533_;
  wire _28534_;
  wire _28535_;
  wire _28536_;
  wire _28537_;
  wire _28538_;
  wire _28539_;
  wire _28540_;
  wire _28541_;
  wire _28542_;
  wire _28543_;
  wire _28544_;
  wire _28545_;
  wire _28546_;
  wire _28547_;
  wire _28548_;
  wire _28549_;
  wire _28550_;
  wire _28551_;
  wire _28552_;
  wire _28553_;
  wire _28554_;
  wire _28555_;
  wire _28556_;
  wire _28557_;
  wire _28558_;
  wire _28559_;
  wire _28560_;
  wire _28561_;
  wire _28562_;
  wire _28563_;
  wire _28564_;
  wire _28565_;
  wire _28566_;
  wire _28567_;
  wire _28568_;
  wire _28569_;
  wire _28570_;
  wire _28571_;
  wire _28572_;
  wire _28573_;
  wire _28574_;
  wire _28575_;
  wire _28576_;
  wire _28577_;
  wire _28578_;
  wire _28579_;
  wire _28580_;
  wire _28581_;
  wire _28582_;
  wire _28583_;
  wire _28584_;
  wire _28585_;
  wire _28586_;
  wire _28587_;
  wire _28588_;
  wire _28589_;
  wire _28590_;
  wire _28591_;
  wire _28592_;
  wire _28593_;
  wire _28594_;
  wire _28595_;
  wire _28596_;
  wire _28597_;
  wire _28598_;
  wire _28599_;
  wire _28600_;
  wire _28601_;
  wire _28602_;
  wire _28603_;
  wire _28604_;
  wire _28605_;
  wire _28606_;
  wire _28607_;
  wire _28608_;
  wire _28609_;
  wire _28610_;
  wire _28611_;
  wire _28612_;
  wire _28613_;
  wire _28614_;
  wire _28615_;
  wire _28616_;
  wire _28617_;
  wire _28618_;
  wire _28619_;
  wire _28620_;
  wire _28621_;
  wire _28622_;
  wire _28623_;
  wire _28624_;
  wire _28625_;
  wire _28626_;
  wire _28627_;
  wire _28628_;
  wire _28629_;
  wire _28630_;
  wire _28631_;
  wire _28632_;
  wire _28633_;
  wire _28634_;
  wire _28635_;
  wire _28636_;
  wire _28637_;
  wire _28638_;
  wire _28639_;
  wire _28640_;
  wire _28641_;
  wire _28642_;
  wire _28643_;
  wire _28644_;
  wire _28645_;
  wire _28646_;
  wire _28647_;
  wire _28648_;
  wire _28649_;
  wire _28650_;
  wire _28651_;
  wire _28652_;
  wire _28653_;
  wire _28654_;
  wire _28655_;
  wire _28656_;
  wire _28657_;
  wire _28658_;
  wire _28659_;
  wire _28660_;
  wire _28661_;
  wire _28662_;
  wire _28663_;
  wire _28664_;
  wire _28665_;
  wire _28666_;
  wire _28667_;
  wire _28668_;
  wire _28669_;
  wire _28670_;
  wire _28671_;
  wire _28672_;
  wire _28673_;
  wire _28674_;
  wire _28675_;
  wire _28676_;
  wire _28677_;
  wire _28678_;
  wire _28679_;
  wire _28680_;
  wire _28681_;
  wire _28682_;
  wire _28683_;
  wire _28684_;
  wire _28685_;
  wire _28686_;
  wire _28687_;
  wire _28688_;
  wire _28689_;
  wire _28690_;
  wire _28691_;
  wire _28692_;
  wire _28693_;
  wire _28694_;
  wire _28695_;
  wire _28696_;
  wire _28697_;
  wire _28698_;
  wire _28699_;
  wire _28700_;
  wire _28701_;
  wire _28702_;
  wire _28703_;
  wire _28704_;
  wire _28705_;
  wire _28706_;
  wire _28707_;
  wire _28708_;
  wire _28709_;
  wire _28710_;
  wire _28711_;
  wire _28712_;
  wire _28713_;
  wire _28714_;
  wire _28715_;
  wire _28716_;
  wire _28717_;
  wire _28718_;
  wire _28719_;
  wire _28720_;
  wire _28721_;
  wire _28722_;
  wire _28723_;
  wire _28724_;
  wire _28725_;
  wire _28726_;
  wire _28727_;
  wire _28728_;
  wire _28729_;
  wire _28730_;
  wire _28731_;
  wire _28732_;
  wire _28733_;
  wire _28734_;
  wire _28735_;
  wire _28736_;
  wire _28737_;
  wire _28738_;
  wire _28739_;
  wire _28740_;
  wire _28741_;
  wire _28742_;
  wire _28743_;
  wire _28744_;
  wire _28745_;
  wire _28746_;
  wire _28747_;
  wire _28748_;
  wire _28749_;
  wire _28750_;
  wire _28751_;
  wire _28752_;
  wire _28753_;
  wire _28754_;
  wire _28755_;
  wire _28756_;
  wire _28757_;
  wire _28758_;
  wire _28759_;
  wire _28760_;
  wire _28761_;
  wire _28762_;
  wire _28763_;
  wire _28764_;
  wire _28765_;
  wire _28766_;
  wire _28767_;
  wire _28768_;
  wire _28769_;
  wire _28770_;
  wire _28771_;
  wire _28772_;
  wire _28773_;
  wire _28774_;
  wire _28775_;
  wire _28776_;
  wire _28777_;
  wire _28778_;
  wire _28779_;
  wire _28780_;
  wire _28781_;
  wire _28782_;
  wire _28783_;
  wire _28784_;
  wire _28785_;
  wire _28786_;
  wire _28787_;
  wire _28788_;
  wire _28789_;
  wire _28790_;
  wire _28791_;
  wire _28792_;
  wire _28793_;
  wire _28794_;
  wire _28795_;
  wire _28796_;
  wire _28797_;
  wire _28798_;
  wire _28799_;
  wire _28800_;
  wire _28801_;
  wire _28802_;
  wire _28803_;
  wire _28804_;
  wire _28805_;
  wire _28806_;
  wire _28807_;
  wire _28808_;
  wire _28809_;
  wire _28810_;
  wire _28811_;
  wire _28812_;
  wire _28813_;
  wire _28814_;
  wire _28815_;
  wire _28816_;
  wire _28817_;
  wire _28818_;
  wire _28819_;
  wire _28820_;
  wire _28821_;
  wire _28822_;
  wire _28823_;
  wire _28824_;
  wire _28825_;
  wire _28826_;
  wire _28827_;
  wire _28828_;
  wire _28829_;
  wire _28830_;
  wire _28831_;
  wire _28832_;
  wire _28833_;
  wire _28834_;
  wire _28835_;
  wire _28836_;
  wire _28837_;
  wire _28838_;
  wire _28839_;
  wire _28840_;
  wire _28841_;
  wire _28842_;
  wire _28843_;
  wire _28844_;
  wire _28845_;
  wire _28846_;
  wire _28847_;
  wire _28848_;
  wire _28849_;
  wire _28850_;
  wire _28851_;
  wire _28852_;
  wire _28853_;
  wire _28854_;
  wire _28855_;
  wire _28856_;
  wire _28857_;
  wire _28858_;
  wire _28859_;
  wire _28860_;
  wire _28861_;
  wire _28862_;
  wire _28863_;
  wire _28864_;
  wire _28865_;
  wire _28866_;
  wire _28867_;
  wire _28868_;
  wire _28869_;
  wire _28870_;
  wire _28871_;
  wire _28872_;
  wire _28873_;
  wire _28874_;
  wire _28875_;
  wire _28876_;
  wire _28877_;
  wire _28878_;
  wire _28879_;
  wire _28880_;
  wire _28881_;
  wire _28882_;
  wire _28883_;
  wire _28884_;
  wire _28885_;
  wire _28886_;
  wire _28887_;
  wire _28888_;
  wire _28889_;
  wire _28890_;
  wire _28891_;
  wire _28892_;
  wire _28893_;
  wire _28894_;
  wire _28895_;
  wire _28896_;
  wire _28897_;
  wire _28898_;
  wire _28899_;
  wire _28900_;
  wire _28901_;
  wire _28902_;
  wire _28903_;
  wire _28904_;
  wire _28905_;
  wire _28906_;
  wire _28907_;
  wire _28908_;
  wire _28909_;
  wire _28910_;
  wire _28911_;
  wire _28912_;
  wire _28913_;
  wire _28914_;
  wire _28915_;
  wire _28916_;
  wire _28917_;
  wire _28918_;
  wire _28919_;
  wire _28920_;
  wire _28921_;
  wire _28922_;
  wire _28923_;
  wire _28924_;
  wire _28925_;
  wire _28926_;
  wire _28927_;
  wire _28928_;
  wire _28929_;
  wire _28930_;
  wire _28931_;
  wire _28932_;
  wire _28933_;
  wire _28934_;
  wire _28935_;
  wire _28936_;
  wire _28937_;
  wire _28938_;
  wire _28939_;
  wire _28940_;
  wire _28941_;
  wire _28942_;
  wire _28943_;
  wire _28944_;
  wire _28945_;
  wire _28946_;
  wire _28947_;
  wire _28948_;
  wire _28949_;
  wire _28950_;
  wire _28951_;
  wire _28952_;
  wire _28953_;
  wire _28954_;
  wire _28955_;
  wire _28956_;
  wire _28957_;
  wire _28958_;
  wire _28959_;
  wire _28960_;
  wire _28961_;
  wire _28962_;
  wire _28963_;
  wire _28964_;
  wire _28965_;
  wire _28966_;
  wire _28967_;
  wire _28968_;
  wire _28969_;
  wire _28970_;
  wire _28971_;
  wire _28972_;
  wire _28973_;
  wire _28974_;
  wire _28975_;
  wire _28976_;
  wire _28977_;
  wire _28978_;
  wire _28979_;
  wire _28980_;
  wire _28981_;
  wire _28982_;
  wire _28983_;
  wire _28984_;
  wire _28985_;
  wire _28986_;
  wire _28987_;
  wire _28988_;
  wire _28989_;
  wire _28990_;
  wire _28991_;
  wire _28992_;
  wire _28993_;
  wire _28994_;
  wire _28995_;
  wire _28996_;
  wire _28997_;
  wire _28998_;
  wire _28999_;
  wire _29000_;
  wire _29001_;
  wire _29002_;
  wire _29003_;
  wire _29004_;
  wire _29005_;
  wire _29006_;
  wire _29007_;
  wire _29008_;
  wire _29009_;
  wire _29010_;
  wire _29011_;
  wire _29012_;
  wire _29013_;
  wire _29014_;
  wire _29015_;
  wire _29016_;
  wire _29017_;
  wire _29018_;
  wire _29019_;
  wire _29020_;
  wire _29021_;
  wire _29022_;
  wire _29023_;
  wire _29024_;
  wire _29025_;
  wire _29026_;
  wire _29027_;
  wire _29028_;
  wire _29029_;
  wire _29030_;
  wire _29031_;
  wire _29032_;
  wire _29033_;
  wire _29034_;
  wire _29035_;
  wire _29036_;
  wire _29037_;
  wire _29038_;
  wire _29039_;
  wire _29040_;
  wire _29041_;
  wire _29042_;
  wire _29043_;
  wire _29044_;
  wire _29045_;
  wire _29046_;
  wire _29047_;
  wire _29048_;
  wire _29049_;
  wire _29050_;
  wire _29051_;
  wire _29052_;
  wire _29053_;
  wire _29054_;
  wire _29055_;
  wire _29056_;
  wire _29057_;
  wire _29058_;
  wire _29059_;
  wire _29060_;
  wire _29061_;
  wire _29062_;
  wire _29063_;
  wire _29064_;
  wire _29065_;
  wire _29066_;
  wire _29067_;
  wire _29068_;
  wire _29069_;
  wire _29070_;
  wire _29071_;
  wire _29072_;
  wire _29073_;
  wire _29074_;
  wire _29075_;
  wire _29076_;
  wire _29077_;
  wire _29078_;
  wire _29079_;
  wire _29080_;
  wire _29081_;
  wire _29082_;
  wire _29083_;
  wire _29084_;
  wire _29085_;
  wire _29086_;
  wire _29087_;
  wire _29088_;
  wire _29089_;
  wire _29090_;
  wire _29091_;
  wire _29092_;
  wire _29093_;
  wire _29094_;
  wire _29095_;
  wire _29096_;
  wire _29097_;
  wire _29098_;
  wire _29099_;
  wire _29100_;
  wire _29101_;
  wire _29102_;
  wire _29103_;
  wire _29104_;
  wire _29105_;
  wire _29106_;
  wire _29107_;
  wire _29108_;
  wire _29109_;
  wire _29110_;
  wire _29111_;
  wire _29112_;
  wire _29113_;
  wire _29114_;
  wire _29115_;
  wire _29116_;
  wire _29117_;
  wire _29118_;
  wire _29119_;
  wire _29120_;
  wire _29121_;
  wire _29122_;
  wire _29123_;
  wire _29124_;
  wire _29125_;
  wire _29126_;
  wire _29127_;
  wire _29128_;
  wire _29129_;
  wire _29130_;
  wire _29131_;
  wire _29132_;
  wire _29133_;
  wire _29134_;
  wire _29135_;
  wire _29136_;
  wire _29137_;
  wire _29138_;
  wire _29139_;
  wire _29140_;
  wire _29141_;
  wire _29142_;
  wire _29143_;
  wire _29144_;
  wire _29145_;
  wire _29146_;
  wire _29147_;
  wire _29148_;
  wire _29149_;
  wire _29150_;
  wire _29151_;
  wire _29152_;
  wire _29153_;
  wire _29154_;
  wire _29155_;
  wire _29156_;
  wire _29157_;
  wire _29158_;
  wire _29159_;
  wire _29160_;
  wire _29161_;
  wire _29162_;
  wire _29163_;
  wire _29164_;
  wire _29165_;
  wire _29166_;
  wire _29167_;
  wire _29168_;
  wire _29169_;
  wire _29170_;
  wire _29171_;
  wire _29172_;
  wire _29173_;
  wire _29174_;
  wire _29175_;
  wire _29176_;
  wire _29177_;
  wire _29178_;
  wire _29179_;
  wire _29180_;
  wire _29181_;
  wire _29182_;
  wire _29183_;
  wire _29184_;
  wire _29185_;
  wire _29186_;
  wire _29187_;
  wire _29188_;
  wire _29189_;
  wire _29190_;
  wire _29191_;
  wire _29192_;
  wire _29193_;
  wire _29194_;
  wire _29195_;
  wire _29196_;
  wire _29197_;
  wire _29198_;
  wire _29199_;
  wire _29200_;
  wire _29201_;
  wire _29202_;
  wire _29203_;
  wire _29204_;
  wire _29205_;
  wire _29206_;
  wire _29207_;
  wire _29208_;
  wire _29209_;
  wire _29210_;
  wire _29211_;
  wire _29212_;
  wire _29213_;
  wire _29214_;
  wire _29215_;
  wire _29216_;
  wire _29217_;
  wire _29218_;
  wire _29219_;
  wire _29220_;
  wire _29221_;
  wire _29222_;
  wire _29223_;
  wire _29224_;
  wire _29225_;
  wire _29226_;
  wire _29227_;
  wire _29228_;
  wire _29229_;
  wire _29230_;
  wire _29231_;
  wire _29232_;
  wire _29233_;
  wire _29234_;
  wire _29235_;
  wire _29236_;
  wire _29237_;
  wire _29238_;
  wire _29239_;
  wire _29240_;
  wire _29241_;
  wire _29242_;
  wire _29243_;
  wire _29244_;
  wire _29245_;
  wire _29246_;
  wire _29247_;
  wire _29248_;
  wire _29249_;
  wire _29250_;
  wire _29251_;
  wire _29252_;
  wire _29253_;
  wire _29254_;
  wire _29255_;
  wire _29256_;
  wire _29257_;
  wire _29258_;
  wire _29259_;
  wire _29260_;
  wire _29261_;
  wire _29262_;
  wire _29263_;
  wire _29264_;
  wire _29265_;
  wire _29266_;
  wire _29267_;
  wire _29268_;
  wire _29269_;
  wire _29270_;
  wire _29271_;
  wire _29272_;
  wire _29273_;
  wire _29274_;
  wire _29275_;
  wire _29276_;
  wire _29277_;
  wire _29278_;
  wire _29279_;
  wire _29280_;
  wire _29281_;
  wire _29282_;
  wire _29283_;
  wire _29284_;
  wire _29285_;
  wire _29286_;
  wire _29287_;
  wire _29288_;
  wire _29289_;
  wire _29290_;
  wire _29291_;
  wire _29292_;
  wire _29293_;
  wire _29294_;
  wire _29295_;
  wire _29296_;
  wire _29297_;
  wire _29298_;
  wire _29299_;
  wire _29300_;
  wire _29301_;
  wire _29302_;
  wire _29303_;
  wire _29304_;
  wire _29305_;
  wire _29306_;
  wire _29307_;
  wire _29308_;
  wire _29309_;
  wire _29310_;
  wire _29311_;
  wire _29312_;
  wire _29313_;
  wire _29314_;
  wire _29315_;
  wire _29316_;
  wire _29317_;
  wire _29318_;
  wire _29319_;
  wire _29320_;
  wire _29321_;
  wire _29322_;
  wire _29323_;
  wire _29324_;
  wire _29325_;
  wire _29326_;
  wire _29327_;
  wire _29328_;
  wire _29329_;
  wire _29330_;
  wire _29331_;
  wire _29332_;
  wire _29333_;
  wire _29334_;
  wire _29335_;
  wire _29336_;
  wire _29337_;
  wire _29338_;
  wire _29339_;
  wire _29340_;
  wire _29341_;
  wire _29342_;
  wire _29343_;
  wire _29344_;
  wire _29345_;
  wire _29346_;
  wire _29347_;
  wire _29348_;
  wire _29349_;
  wire _29350_;
  wire _29351_;
  wire _29352_;
  wire _29353_;
  wire _29354_;
  wire _29355_;
  wire _29356_;
  wire _29357_;
  wire _29358_;
  wire _29359_;
  wire _29360_;
  wire _29361_;
  wire _29362_;
  wire _29363_;
  wire _29364_;
  wire _29365_;
  wire _29366_;
  wire _29367_;
  wire _29368_;
  wire _29369_;
  wire _29370_;
  wire _29371_;
  wire _29372_;
  wire _29373_;
  wire _29374_;
  wire _29375_;
  wire _29376_;
  wire _29377_;
  wire _29378_;
  wire _29379_;
  wire _29380_;
  wire _29381_;
  wire _29382_;
  wire _29383_;
  wire _29384_;
  wire _29385_;
  wire _29386_;
  wire _29387_;
  wire _29388_;
  wire _29389_;
  wire _29390_;
  wire _29391_;
  wire _29392_;
  wire _29393_;
  wire _29394_;
  wire _29395_;
  wire _29396_;
  wire _29397_;
  wire _29398_;
  wire _29399_;
  wire _29400_;
  wire _29401_;
  wire _29402_;
  wire _29403_;
  wire _29404_;
  wire _29405_;
  wire _29406_;
  wire _29407_;
  wire _29408_;
  wire _29409_;
  wire _29410_;
  wire _29411_;
  wire _29412_;
  wire _29413_;
  wire _29414_;
  wire _29415_;
  wire _29416_;
  wire _29417_;
  wire _29418_;
  wire _29419_;
  wire _29420_;
  wire _29421_;
  wire _29422_;
  wire _29423_;
  wire _29424_;
  wire _29425_;
  wire _29426_;
  wire _29427_;
  wire _29428_;
  wire _29429_;
  wire _29430_;
  wire _29431_;
  wire _29432_;
  wire _29433_;
  wire _29434_;
  wire _29435_;
  wire _29436_;
  wire _29437_;
  wire _29438_;
  wire _29439_;
  wire _29440_;
  wire _29441_;
  wire _29442_;
  wire _29443_;
  wire _29444_;
  wire _29445_;
  wire _29446_;
  wire _29447_;
  wire _29448_;
  wire _29449_;
  wire _29450_;
  wire _29451_;
  wire _29452_;
  wire _29453_;
  wire _29454_;
  wire _29455_;
  wire _29456_;
  wire _29457_;
  wire _29458_;
  wire _29459_;
  wire _29460_;
  wire _29461_;
  wire _29462_;
  wire _29463_;
  wire _29464_;
  wire _29465_;
  wire _29466_;
  wire _29467_;
  wire _29468_;
  wire _29469_;
  wire _29470_;
  wire _29471_;
  wire _29472_;
  wire _29473_;
  wire _29474_;
  wire _29475_;
  wire _29476_;
  wire _29477_;
  wire _29478_;
  wire _29479_;
  wire _29480_;
  wire _29481_;
  wire _29482_;
  wire _29483_;
  wire _29484_;
  wire _29485_;
  wire _29486_;
  wire _29487_;
  wire _29488_;
  wire _29489_;
  wire _29490_;
  wire _29491_;
  wire _29492_;
  wire _29493_;
  wire _29494_;
  wire _29495_;
  wire _29496_;
  wire _29497_;
  wire _29498_;
  wire _29499_;
  wire _29500_;
  wire _29501_;
  wire _29502_;
  wire _29503_;
  wire _29504_;
  wire _29505_;
  wire _29506_;
  wire _29507_;
  wire _29508_;
  wire _29509_;
  wire _29510_;
  wire _29511_;
  wire _29512_;
  wire _29513_;
  wire _29514_;
  wire _29515_;
  wire _29516_;
  wire _29517_;
  wire _29518_;
  wire _29519_;
  wire _29520_;
  wire _29521_;
  wire _29522_;
  wire _29523_;
  wire _29524_;
  wire _29525_;
  wire _29526_;
  wire _29527_;
  wire _29528_;
  wire _29529_;
  wire _29530_;
  wire _29531_;
  wire _29532_;
  wire _29533_;
  wire _29534_;
  wire _29535_;
  wire _29536_;
  wire _29537_;
  wire _29538_;
  wire _29539_;
  wire _29540_;
  wire _29541_;
  wire _29542_;
  wire _29543_;
  wire _29544_;
  wire _29545_;
  wire _29546_;
  wire _29547_;
  wire _29548_;
  wire _29549_;
  wire _29550_;
  wire _29551_;
  wire _29552_;
  wire _29553_;
  wire _29554_;
  wire _29555_;
  wire _29556_;
  wire _29557_;
  wire _29558_;
  wire _29559_;
  wire _29560_;
  wire _29561_;
  wire _29562_;
  wire _29563_;
  wire _29564_;
  wire _29565_;
  wire _29566_;
  wire _29567_;
  wire _29568_;
  wire _29569_;
  wire _29570_;
  wire _29571_;
  wire _29572_;
  wire _29573_;
  wire _29574_;
  wire _29575_;
  wire _29576_;
  wire _29577_;
  wire _29578_;
  wire _29579_;
  wire _29580_;
  wire _29581_;
  wire _29582_;
  wire _29583_;
  wire _29584_;
  wire _29585_;
  wire _29586_;
  wire _29587_;
  wire _29588_;
  wire _29589_;
  wire _29590_;
  wire _29591_;
  wire _29592_;
  wire _29593_;
  wire _29594_;
  wire _29595_;
  wire _29596_;
  wire _29597_;
  wire _29598_;
  wire _29599_;
  wire _29600_;
  wire _29601_;
  wire _29602_;
  wire _29603_;
  wire _29604_;
  wire _29605_;
  wire _29606_;
  wire _29607_;
  wire _29608_;
  wire _29609_;
  wire _29610_;
  wire _29611_;
  wire _29612_;
  wire _29613_;
  wire _29614_;
  wire _29615_;
  wire _29616_;
  wire _29617_;
  wire _29618_;
  wire _29619_;
  wire _29620_;
  wire _29621_;
  wire _29622_;
  wire _29623_;
  wire _29624_;
  wire _29625_;
  wire _29626_;
  wire _29627_;
  wire _29628_;
  wire _29629_;
  wire _29630_;
  wire _29631_;
  wire _29632_;
  wire _29633_;
  wire _29634_;
  wire _29635_;
  wire _29636_;
  wire _29637_;
  wire _29638_;
  wire _29639_;
  wire _29640_;
  wire _29641_;
  wire _29642_;
  wire _29643_;
  wire _29644_;
  wire _29645_;
  wire _29646_;
  wire _29647_;
  wire _29648_;
  wire _29649_;
  wire _29650_;
  wire _29651_;
  wire _29652_;
  wire _29653_;
  wire _29654_;
  wire _29655_;
  wire _29656_;
  wire _29657_;
  wire _29658_;
  wire _29659_;
  wire _29660_;
  wire _29661_;
  wire _29662_;
  wire _29663_;
  wire _29664_;
  wire _29665_;
  wire _29666_;
  wire _29667_;
  wire _29668_;
  wire _29669_;
  wire _29670_;
  wire _29671_;
  wire _29672_;
  wire _29673_;
  wire _29674_;
  wire _29675_;
  wire _29676_;
  wire _29677_;
  wire _29678_;
  wire _29679_;
  wire _29680_;
  wire _29681_;
  wire _29682_;
  wire _29683_;
  wire _29684_;
  wire _29685_;
  wire _29686_;
  wire _29687_;
  wire _29688_;
  wire _29689_;
  wire _29690_;
  wire _29691_;
  wire _29692_;
  wire _29693_;
  wire _29694_;
  wire _29695_;
  wire _29696_;
  wire _29697_;
  wire _29698_;
  wire _29699_;
  wire _29700_;
  wire _29701_;
  wire _29702_;
  wire _29703_;
  wire _29704_;
  wire _29705_;
  wire _29706_;
  wire _29707_;
  wire _29708_;
  wire _29709_;
  wire _29710_;
  wire _29711_;
  wire _29712_;
  wire _29713_;
  wire _29714_;
  wire _29715_;
  wire _29716_;
  wire _29717_;
  wire _29718_;
  wire _29719_;
  wire _29720_;
  wire _29721_;
  wire _29722_;
  wire _29723_;
  wire _29724_;
  wire _29725_;
  wire _29726_;
  wire _29727_;
  wire _29728_;
  wire _29729_;
  wire _29730_;
  wire _29731_;
  wire _29732_;
  wire _29733_;
  wire _29734_;
  wire _29735_;
  wire _29736_;
  wire _29737_;
  wire _29738_;
  wire _29739_;
  wire _29740_;
  wire _29741_;
  wire _29742_;
  wire _29743_;
  wire _29744_;
  wire _29745_;
  wire _29746_;
  wire _29747_;
  wire _29748_;
  wire _29749_;
  wire _29750_;
  wire _29751_;
  wire _29752_;
  wire _29753_;
  wire _29754_;
  wire _29755_;
  wire _29756_;
  wire _29757_;
  wire _29758_;
  wire _29759_;
  wire _29760_;
  wire _29761_;
  wire _29762_;
  wire _29763_;
  wire _29764_;
  wire _29765_;
  wire _29766_;
  wire _29767_;
  wire _29768_;
  wire _29769_;
  wire _29770_;
  wire _29771_;
  wire _29772_;
  wire _29773_;
  wire _29774_;
  wire _29775_;
  wire _29776_;
  wire _29777_;
  wire _29778_;
  wire _29779_;
  wire _29780_;
  wire _29781_;
  wire _29782_;
  wire _29783_;
  wire _29784_;
  wire _29785_;
  wire _29786_;
  wire _29787_;
  wire _29788_;
  wire _29789_;
  wire _29790_;
  wire _29791_;
  wire _29792_;
  wire _29793_;
  wire _29794_;
  wire _29795_;
  wire _29796_;
  wire _29797_;
  wire _29798_;
  wire _29799_;
  wire _29800_;
  wire _29801_;
  wire _29802_;
  wire _29803_;
  wire _29804_;
  wire _29805_;
  wire _29806_;
  wire _29807_;
  wire _29808_;
  wire _29809_;
  wire _29810_;
  wire _29811_;
  wire _29812_;
  wire _29813_;
  wire _29814_;
  wire _29815_;
  wire _29816_;
  wire _29817_;
  wire _29818_;
  wire _29819_;
  wire _29820_;
  wire _29821_;
  wire _29822_;
  wire _29823_;
  wire _29824_;
  wire _29825_;
  wire _29826_;
  wire _29827_;
  wire _29828_;
  wire _29829_;
  wire _29830_;
  wire _29831_;
  wire _29832_;
  wire _29833_;
  wire _29834_;
  wire _29835_;
  wire _29836_;
  wire _29837_;
  wire _29838_;
  wire _29839_;
  wire _29840_;
  wire _29841_;
  wire _29842_;
  wire _29843_;
  wire _29844_;
  wire _29845_;
  wire _29846_;
  wire _29847_;
  wire _29848_;
  wire _29849_;
  wire _29850_;
  wire _29851_;
  wire _29852_;
  wire _29853_;
  wire _29854_;
  wire _29855_;
  wire _29856_;
  wire _29857_;
  wire _29858_;
  wire _29859_;
  wire _29860_;
  wire _29861_;
  wire _29862_;
  wire _29863_;
  wire _29864_;
  wire _29865_;
  wire _29866_;
  wire _29867_;
  wire _29868_;
  wire _29869_;
  wire _29870_;
  wire _29871_;
  wire _29872_;
  wire _29873_;
  wire _29874_;
  wire _29875_;
  wire _29876_;
  wire _29877_;
  wire _29878_;
  wire _29879_;
  wire _29880_;
  wire _29881_;
  wire _29882_;
  wire _29883_;
  wire _29884_;
  wire _29885_;
  wire _29886_;
  wire _29887_;
  wire _29888_;
  wire _29889_;
  wire _29890_;
  wire _29891_;
  wire _29892_;
  wire _29893_;
  wire _29894_;
  wire _29895_;
  wire _29896_;
  wire _29897_;
  wire _29898_;
  wire _29899_;
  wire _29900_;
  wire _29901_;
  wire _29902_;
  wire _29903_;
  wire _29904_;
  wire _29905_;
  wire _29906_;
  wire _29907_;
  wire _29908_;
  wire _29909_;
  wire _29910_;
  wire _29911_;
  wire _29912_;
  wire _29913_;
  wire _29914_;
  wire _29915_;
  wire _29916_;
  wire _29917_;
  wire _29918_;
  wire _29919_;
  wire _29920_;
  wire _29921_;
  wire _29922_;
  wire _29923_;
  wire _29924_;
  wire _29925_;
  wire _29926_;
  wire _29927_;
  wire _29928_;
  wire _29929_;
  wire _29930_;
  wire _29931_;
  wire _29932_;
  wire _29933_;
  wire _29934_;
  wire _29935_;
  wire _29936_;
  wire _29937_;
  wire _29938_;
  wire _29939_;
  wire _29940_;
  wire _29941_;
  wire _29942_;
  wire _29943_;
  wire _29944_;
  wire _29945_;
  wire _29946_;
  wire _29947_;
  wire _29948_;
  wire _29949_;
  wire _29950_;
  wire _29951_;
  wire _29952_;
  wire _29953_;
  wire _29954_;
  wire _29955_;
  wire _29956_;
  wire _29957_;
  wire _29958_;
  wire _29959_;
  wire _29960_;
  wire _29961_;
  wire _29962_;
  wire _29963_;
  wire _29964_;
  wire _29965_;
  wire _29966_;
  wire _29967_;
  wire _29968_;
  wire _29969_;
  wire _29970_;
  wire _29971_;
  wire _29972_;
  wire _29973_;
  wire _29974_;
  wire _29975_;
  wire _29976_;
  wire _29977_;
  wire _29978_;
  wire _29979_;
  wire _29980_;
  wire _29981_;
  wire _29982_;
  wire _29983_;
  wire _29984_;
  wire _29985_;
  wire _29986_;
  wire _29987_;
  wire _29988_;
  wire _29989_;
  wire _29990_;
  wire _29991_;
  wire _29992_;
  wire _29993_;
  wire _29994_;
  wire _29995_;
  wire _29996_;
  wire _29997_;
  wire _29998_;
  wire _29999_;
  wire _30000_;
  wire _30001_;
  wire _30002_;
  wire _30003_;
  wire _30004_;
  wire _30005_;
  wire _30006_;
  wire _30007_;
  wire _30008_;
  wire _30009_;
  wire _30010_;
  wire _30011_;
  wire _30012_;
  wire _30013_;
  wire _30014_;
  wire _30015_;
  wire _30016_;
  wire _30017_;
  wire _30018_;
  wire _30019_;
  wire _30020_;
  wire _30021_;
  wire _30022_;
  wire _30023_;
  wire _30024_;
  wire _30025_;
  wire _30026_;
  wire _30027_;
  wire _30028_;
  wire _30029_;
  wire _30030_;
  wire _30031_;
  wire _30032_;
  wire _30033_;
  wire _30034_;
  wire _30035_;
  wire _30036_;
  wire _30037_;
  wire _30038_;
  wire _30039_;
  wire _30040_;
  wire _30041_;
  wire _30042_;
  wire _30043_;
  wire _30044_;
  wire _30045_;
  wire _30046_;
  wire _30047_;
  wire _30048_;
  wire _30049_;
  wire _30050_;
  wire _30051_;
  wire _30052_;
  wire _30053_;
  wire _30054_;
  wire _30055_;
  wire _30056_;
  wire _30057_;
  wire _30058_;
  wire _30059_;
  wire _30060_;
  wire _30061_;
  wire _30062_;
  wire _30063_;
  wire _30064_;
  wire _30065_;
  wire _30066_;
  wire _30067_;
  wire _30068_;
  wire _30069_;
  wire _30070_;
  wire _30071_;
  wire _30072_;
  wire _30073_;
  wire _30074_;
  wire _30075_;
  wire _30076_;
  wire _30077_;
  wire _30078_;
  wire _30079_;
  wire _30080_;
  wire _30081_;
  wire _30082_;
  wire _30083_;
  wire _30084_;
  wire _30085_;
  wire _30086_;
  wire _30087_;
  wire _30088_;
  wire _30089_;
  wire _30090_;
  wire _30091_;
  wire _30092_;
  wire _30093_;
  wire _30094_;
  wire _30095_;
  wire _30096_;
  wire _30097_;
  wire _30098_;
  wire _30099_;
  wire _30100_;
  wire _30101_;
  wire _30102_;
  wire _30103_;
  wire _30104_;
  wire _30105_;
  wire _30106_;
  wire _30107_;
  wire _30108_;
  wire _30109_;
  wire _30110_;
  wire _30111_;
  wire _30112_;
  wire _30113_;
  wire _30114_;
  wire _30115_;
  wire _30116_;
  wire _30117_;
  wire _30118_;
  wire _30119_;
  wire _30120_;
  wire _30121_;
  wire _30122_;
  wire _30123_;
  wire _30124_;
  wire _30125_;
  wire _30126_;
  wire _30127_;
  wire _30128_;
  wire _30129_;
  wire _30130_;
  wire _30131_;
  wire _30132_;
  wire _30133_;
  wire _30134_;
  wire _30135_;
  wire _30136_;
  wire _30137_;
  wire _30138_;
  wire _30139_;
  wire _30140_;
  wire _30141_;
  wire _30142_;
  wire _30143_;
  wire _30144_;
  wire _30145_;
  wire _30146_;
  wire _30147_;
  wire _30148_;
  wire _30149_;
  wire _30150_;
  wire _30151_;
  wire _30152_;
  wire _30153_;
  wire _30154_;
  wire _30155_;
  wire _30156_;
  wire _30157_;
  wire _30158_;
  wire _30159_;
  wire _30160_;
  wire _30161_;
  wire _30162_;
  wire _30163_;
  wire _30164_;
  wire _30165_;
  wire _30166_;
  wire _30167_;
  wire _30168_;
  wire _30169_;
  wire _30170_;
  wire _30171_;
  wire _30172_;
  wire _30173_;
  wire _30174_;
  wire _30175_;
  wire _30176_;
  wire _30177_;
  wire _30178_;
  wire _30179_;
  wire _30180_;
  wire _30181_;
  wire _30182_;
  wire _30183_;
  wire _30184_;
  wire _30185_;
  wire _30186_;
  wire _30187_;
  wire _30188_;
  wire _30189_;
  wire _30190_;
  wire _30191_;
  wire _30192_;
  wire _30193_;
  wire _30194_;
  wire _30195_;
  wire _30196_;
  wire _30197_;
  wire _30198_;
  wire _30199_;
  wire _30200_;
  wire _30201_;
  wire _30202_;
  wire _30203_;
  wire _30204_;
  wire _30205_;
  wire _30206_;
  wire _30207_;
  wire _30208_;
  wire _30209_;
  wire _30210_;
  wire _30211_;
  wire _30212_;
  wire _30213_;
  wire _30214_;
  wire _30215_;
  wire _30216_;
  wire _30217_;
  wire _30218_;
  wire _30219_;
  wire _30220_;
  wire _30221_;
  wire _30222_;
  wire _30223_;
  wire _30224_;
  wire _30225_;
  wire _30226_;
  wire _30227_;
  wire _30228_;
  wire _30229_;
  wire _30230_;
  wire _30231_;
  wire _30232_;
  wire _30233_;
  wire _30234_;
  wire _30235_;
  wire _30236_;
  wire _30237_;
  wire _30238_;
  wire _30239_;
  wire _30240_;
  wire _30241_;
  wire _30242_;
  wire _30243_;
  wire _30244_;
  wire _30245_;
  wire _30246_;
  wire _30247_;
  wire _30248_;
  wire _30249_;
  wire _30250_;
  wire _30251_;
  wire _30252_;
  wire _30253_;
  wire _30254_;
  wire _30255_;
  wire _30256_;
  wire _30257_;
  wire _30258_;
  wire _30259_;
  wire _30260_;
  wire _30261_;
  wire _30262_;
  wire _30263_;
  wire _30264_;
  wire _30265_;
  wire _30266_;
  wire _30267_;
  wire _30268_;
  wire _30269_;
  wire _30270_;
  wire _30271_;
  wire _30272_;
  wire _30273_;
  wire _30274_;
  wire _30275_;
  wire _30276_;
  wire _30277_;
  wire _30278_;
  wire _30279_;
  wire _30280_;
  wire _30281_;
  wire _30282_;
  wire _30283_;
  wire _30284_;
  wire _30285_;
  wire _30286_;
  wire _30287_;
  wire _30288_;
  wire _30289_;
  wire _30290_;
  wire _30291_;
  wire _30292_;
  wire _30293_;
  wire _30294_;
  wire _30295_;
  wire _30296_;
  wire _30297_;
  wire _30298_;
  wire _30299_;
  wire _30300_;
  wire _30301_;
  wire _30302_;
  wire _30303_;
  wire _30304_;
  wire _30305_;
  wire _30306_;
  wire _30307_;
  wire _30308_;
  wire _30309_;
  wire _30310_;
  wire _30311_;
  wire _30312_;
  wire _30313_;
  wire _30314_;
  wire _30315_;
  wire _30316_;
  wire _30317_;
  wire _30318_;
  wire _30319_;
  wire _30320_;
  wire _30321_;
  wire _30322_;
  wire _30323_;
  wire _30324_;
  wire _30325_;
  wire _30326_;
  wire _30327_;
  wire _30328_;
  wire _30329_;
  wire _30330_;
  wire _30331_;
  wire _30332_;
  wire _30333_;
  wire _30334_;
  wire _30335_;
  wire _30336_;
  wire _30337_;
  wire _30338_;
  wire _30339_;
  wire _30340_;
  wire _30341_;
  wire _30342_;
  wire _30343_;
  wire _30344_;
  wire _30345_;
  wire _30346_;
  wire _30347_;
  wire _30348_;
  wire _30349_;
  wire _30350_;
  wire _30351_;
  wire _30352_;
  wire _30353_;
  wire _30354_;
  wire _30355_;
  wire _30356_;
  wire _30357_;
  wire _30358_;
  wire _30359_;
  wire _30360_;
  wire _30361_;
  wire _30362_;
  wire _30363_;
  wire _30364_;
  wire _30365_;
  wire _30366_;
  wire _30367_;
  wire _30368_;
  wire _30369_;
  wire _30370_;
  wire _30371_;
  wire _30372_;
  wire _30373_;
  wire _30374_;
  wire _30375_;
  wire _30376_;
  wire _30377_;
  wire _30378_;
  wire _30379_;
  wire _30380_;
  wire _30381_;
  wire _30382_;
  wire _30383_;
  wire _30384_;
  wire _30385_;
  wire _30386_;
  wire _30387_;
  wire _30388_;
  wire _30389_;
  wire _30390_;
  wire _30391_;
  wire _30392_;
  wire _30393_;
  wire _30394_;
  wire _30395_;
  wire _30396_;
  wire _30397_;
  wire _30398_;
  wire _30399_;
  wire _30400_;
  wire _30401_;
  wire _30402_;
  wire _30403_;
  wire _30404_;
  wire _30405_;
  wire _30406_;
  wire _30407_;
  wire _30408_;
  wire _30409_;
  wire _30410_;
  wire _30411_;
  wire _30412_;
  wire _30413_;
  wire _30414_;
  wire _30415_;
  wire _30416_;
  wire _30417_;
  wire _30418_;
  wire _30419_;
  wire _30420_;
  wire _30421_;
  wire _30422_;
  wire _30423_;
  wire _30424_;
  wire _30425_;
  wire _30426_;
  wire _30427_;
  wire _30428_;
  wire _30429_;
  wire _30430_;
  wire _30431_;
  wire _30432_;
  wire _30433_;
  wire _30434_;
  wire _30435_;
  wire _30436_;
  wire _30437_;
  wire _30438_;
  wire _30439_;
  wire _30440_;
  wire _30441_;
  wire _30442_;
  wire _30443_;
  wire _30444_;
  wire _30445_;
  wire _30446_;
  wire _30447_;
  wire _30448_;
  wire _30449_;
  wire _30450_;
  wire _30451_;
  wire _30452_;
  wire _30453_;
  wire _30454_;
  wire _30455_;
  wire _30456_;
  wire _30457_;
  wire _30458_;
  wire _30459_;
  wire _30460_;
  wire _30461_;
  wire _30462_;
  wire _30463_;
  wire _30464_;
  wire _30465_;
  wire _30466_;
  wire _30467_;
  wire _30468_;
  wire _30469_;
  wire _30470_;
  wire _30471_;
  wire _30472_;
  wire _30473_;
  wire _30474_;
  wire _30475_;
  wire _30476_;
  wire _30477_;
  wire _30478_;
  wire _30479_;
  wire _30480_;
  wire _30481_;
  wire _30482_;
  wire _30483_;
  wire _30484_;
  wire _30485_;
  wire _30486_;
  wire _30487_;
  wire _30488_;
  wire _30489_;
  wire _30490_;
  wire _30491_;
  wire _30492_;
  wire _30493_;
  wire _30494_;
  wire _30495_;
  wire _30496_;
  wire _30497_;
  wire _30498_;
  wire _30499_;
  wire _30500_;
  wire _30501_;
  wire _30502_;
  wire _30503_;
  wire _30504_;
  wire _30505_;
  wire _30506_;
  wire _30507_;
  wire _30508_;
  wire _30509_;
  wire _30510_;
  wire _30511_;
  wire _30512_;
  wire _30513_;
  wire _30514_;
  wire _30515_;
  wire _30516_;
  wire _30517_;
  wire _30518_;
  wire _30519_;
  wire _30520_;
  wire _30521_;
  wire _30522_;
  wire _30523_;
  wire _30524_;
  wire _30525_;
  wire _30526_;
  wire _30527_;
  wire _30528_;
  wire _30529_;
  wire _30530_;
  wire _30531_;
  wire _30532_;
  wire _30533_;
  wire _30534_;
  wire _30535_;
  wire _30536_;
  wire _30537_;
  wire _30538_;
  wire _30539_;
  wire _30540_;
  wire _30541_;
  wire _30542_;
  wire _30543_;
  wire _30544_;
  wire _30545_;
  wire _30546_;
  wire _30547_;
  wire _30548_;
  wire _30549_;
  wire _30550_;
  wire _30551_;
  wire _30552_;
  wire _30553_;
  wire _30554_;
  wire _30555_;
  wire _30556_;
  wire _30557_;
  wire _30558_;
  wire _30559_;
  wire _30560_;
  wire _30561_;
  wire _30562_;
  wire _30563_;
  wire _30564_;
  wire _30565_;
  wire _30566_;
  wire _30567_;
  wire _30568_;
  wire _30569_;
  wire _30570_;
  wire _30571_;
  wire _30572_;
  wire _30573_;
  wire _30574_;
  wire _30575_;
  wire _30576_;
  wire _30577_;
  wire _30578_;
  wire _30579_;
  wire _30580_;
  wire _30581_;
  wire _30582_;
  wire _30583_;
  wire _30584_;
  wire _30585_;
  wire _30586_;
  wire _30587_;
  wire _30588_;
  wire _30589_;
  wire _30590_;
  wire _30591_;
  wire _30592_;
  wire _30593_;
  wire _30594_;
  wire _30595_;
  wire _30596_;
  wire _30597_;
  wire _30598_;
  wire _30599_;
  wire _30600_;
  wire _30601_;
  wire _30602_;
  wire _30603_;
  wire _30604_;
  wire _30605_;
  wire _30606_;
  wire _30607_;
  wire _30608_;
  wire _30609_;
  wire _30610_;
  wire _30611_;
  wire _30612_;
  wire _30613_;
  wire _30614_;
  wire _30615_;
  wire _30616_;
  wire _30617_;
  wire _30618_;
  wire _30619_;
  wire _30620_;
  wire _30621_;
  wire _30622_;
  wire _30623_;
  wire _30624_;
  wire _30625_;
  wire _30626_;
  wire _30627_;
  wire _30628_;
  wire _30629_;
  wire _30630_;
  wire _30631_;
  wire _30632_;
  wire _30633_;
  wire _30634_;
  wire _30635_;
  wire _30636_;
  wire _30637_;
  wire _30638_;
  wire _30639_;
  wire _30640_;
  wire _30641_;
  wire _30642_;
  wire _30643_;
  wire _30644_;
  wire _30645_;
  wire _30646_;
  wire _30647_;
  wire _30648_;
  wire _30649_;
  wire _30650_;
  wire _30651_;
  wire _30652_;
  wire _30653_;
  wire _30654_;
  wire _30655_;
  wire _30656_;
  wire _30657_;
  wire _30658_;
  wire _30659_;
  wire _30660_;
  wire _30661_;
  wire _30662_;
  wire _30663_;
  wire _30664_;
  wire _30665_;
  wire _30666_;
  wire _30667_;
  wire _30668_;
  wire _30669_;
  wire _30670_;
  wire _30671_;
  wire _30672_;
  wire _30673_;
  wire _30674_;
  wire _30675_;
  wire _30676_;
  wire _30677_;
  wire _30678_;
  wire _30679_;
  wire _30680_;
  wire _30681_;
  wire _30682_;
  wire _30683_;
  wire _30684_;
  wire _30685_;
  wire _30686_;
  wire _30687_;
  wire _30688_;
  wire _30689_;
  wire _30690_;
  wire _30691_;
  wire _30692_;
  wire _30693_;
  wire _30694_;
  wire _30695_;
  wire _30696_;
  wire _30697_;
  wire _30698_;
  wire _30699_;
  wire _30700_;
  wire _30701_;
  wire _30702_;
  wire _30703_;
  wire _30704_;
  wire _30705_;
  wire _30706_;
  wire _30707_;
  wire _30708_;
  wire _30709_;
  wire _30710_;
  wire _30711_;
  wire _30712_;
  wire _30713_;
  wire _30714_;
  wire _30715_;
  wire _30716_;
  wire _30717_;
  wire _30718_;
  wire _30719_;
  wire _30720_;
  wire _30721_;
  wire _30722_;
  wire _30723_;
  wire _30724_;
  wire _30725_;
  wire _30726_;
  wire _30727_;
  wire _30728_;
  wire _30729_;
  wire _30730_;
  wire _30731_;
  wire _30732_;
  wire _30733_;
  wire _30734_;
  wire _30735_;
  wire _30736_;
  wire _30737_;
  wire _30738_;
  wire _30739_;
  wire _30740_;
  wire _30741_;
  wire _30742_;
  wire _30743_;
  wire _30744_;
  wire _30745_;
  wire _30746_;
  wire _30747_;
  wire _30748_;
  wire _30749_;
  wire _30750_;
  wire _30751_;
  wire _30752_;
  wire _30753_;
  wire _30754_;
  wire _30755_;
  wire _30756_;
  wire _30757_;
  wire _30758_;
  wire _30759_;
  wire _30760_;
  wire _30761_;
  wire _30762_;
  wire _30763_;
  wire _30764_;
  wire _30765_;
  wire _30766_;
  wire _30767_;
  wire _30768_;
  wire _30769_;
  wire _30770_;
  wire _30771_;
  wire _30772_;
  wire _30773_;
  wire _30774_;
  wire _30775_;
  wire _30776_;
  wire _30777_;
  wire _30778_;
  wire _30779_;
  wire _30780_;
  wire _30781_;
  wire _30782_;
  wire _30783_;
  wire _30784_;
  wire _30785_;
  wire _30786_;
  wire _30787_;
  wire _30788_;
  wire _30789_;
  wire _30790_;
  wire _30791_;
  wire _30792_;
  wire _30793_;
  wire _30794_;
  wire _30795_;
  wire _30796_;
  wire _30797_;
  wire _30798_;
  wire _30799_;
  wire _30800_;
  wire _30801_;
  wire _30802_;
  wire _30803_;
  wire _30804_;
  wire _30805_;
  wire _30806_;
  wire _30807_;
  wire _30808_;
  wire _30809_;
  wire _30810_;
  wire _30811_;
  wire _30812_;
  wire _30813_;
  wire _30814_;
  wire _30815_;
  wire _30816_;
  wire _30817_;
  wire _30818_;
  wire _30819_;
  wire _30820_;
  wire _30821_;
  wire _30822_;
  wire _30823_;
  wire _30824_;
  wire _30825_;
  wire _30826_;
  wire _30827_;
  wire _30828_;
  wire _30829_;
  wire _30830_;
  wire _30831_;
  wire _30832_;
  wire _30833_;
  wire _30834_;
  wire _30835_;
  wire _30836_;
  wire _30837_;
  wire _30838_;
  wire _30839_;
  wire _30840_;
  wire _30841_;
  wire _30842_;
  wire _30843_;
  wire _30844_;
  wire _30845_;
  wire _30846_;
  wire _30847_;
  wire _30848_;
  wire _30849_;
  wire _30850_;
  wire _30851_;
  wire _30852_;
  wire _30853_;
  wire _30854_;
  wire _30855_;
  wire _30856_;
  wire _30857_;
  wire _30858_;
  wire _30859_;
  wire _30860_;
  wire _30861_;
  wire _30862_;
  wire _30863_;
  wire _30864_;
  wire _30865_;
  wire _30866_;
  wire _30867_;
  wire _30868_;
  wire _30869_;
  wire _30870_;
  wire _30871_;
  wire _30872_;
  wire _30873_;
  wire _30874_;
  wire _30875_;
  wire _30876_;
  wire _30877_;
  wire _30878_;
  wire _30879_;
  wire _30880_;
  wire _30881_;
  wire _30882_;
  wire _30883_;
  wire _30884_;
  wire _30885_;
  wire _30886_;
  wire _30887_;
  wire _30888_;
  wire _30889_;
  wire _30890_;
  wire _30891_;
  wire _30892_;
  wire _30893_;
  wire _30894_;
  wire _30895_;
  wire _30896_;
  wire _30897_;
  wire _30898_;
  wire _30899_;
  wire _30900_;
  wire _30901_;
  wire _30902_;
  wire _30903_;
  wire _30904_;
  wire _30905_;
  wire _30906_;
  wire _30907_;
  wire _30908_;
  wire _30909_;
  wire _30910_;
  wire _30911_;
  wire _30912_;
  wire _30913_;
  wire _30914_;
  wire _30915_;
  wire _30916_;
  wire _30917_;
  wire _30918_;
  wire _30919_;
  wire _30920_;
  wire _30921_;
  wire _30922_;
  wire _30923_;
  wire _30924_;
  wire _30925_;
  wire _30926_;
  wire _30927_;
  wire _30928_;
  wire _30929_;
  wire _30930_;
  wire _30931_;
  wire _30932_;
  wire _30933_;
  wire _30934_;
  wire _30935_;
  wire _30936_;
  wire _30937_;
  wire _30938_;
  wire _30939_;
  wire _30940_;
  wire _30941_;
  wire _30942_;
  wire _30943_;
  wire _30944_;
  wire _30945_;
  wire _30946_;
  wire _30947_;
  wire _30948_;
  wire _30949_;
  wire _30950_;
  wire _30951_;
  wire _30952_;
  wire _30953_;
  wire _30954_;
  wire _30955_;
  wire _30956_;
  wire _30957_;
  wire _30958_;
  wire _30959_;
  wire _30960_;
  wire _30961_;
  wire _30962_;
  wire _30963_;
  wire _30964_;
  wire _30965_;
  wire _30966_;
  wire _30967_;
  wire _30968_;
  wire _30969_;
  wire _30970_;
  wire _30971_;
  wire _30972_;
  wire _30973_;
  wire _30974_;
  wire _30975_;
  wire _30976_;
  wire _30977_;
  wire _30978_;
  wire _30979_;
  wire _30980_;
  wire _30981_;
  wire _30982_;
  wire _30983_;
  wire _30984_;
  wire _30985_;
  wire _30986_;
  wire _30987_;
  wire _30988_;
  wire _30989_;
  wire _30990_;
  wire _30991_;
  wire _30992_;
  wire _30993_;
  wire _30994_;
  wire _30995_;
  wire _30996_;
  wire _30997_;
  wire _30998_;
  wire _30999_;
  wire _31000_;
  wire _31001_;
  wire _31002_;
  wire _31003_;
  wire _31004_;
  wire _31005_;
  wire _31006_;
  wire _31007_;
  wire _31008_;
  wire _31009_;
  wire _31010_;
  wire _31011_;
  wire _31012_;
  wire _31013_;
  wire _31014_;
  wire _31015_;
  wire _31016_;
  wire _31017_;
  wire _31018_;
  wire _31019_;
  wire _31020_;
  wire _31021_;
  wire _31022_;
  wire _31023_;
  wire _31024_;
  wire _31025_;
  wire _31026_;
  wire _31027_;
  wire _31028_;
  wire _31029_;
  wire _31030_;
  wire _31031_;
  wire _31032_;
  wire _31033_;
  wire _31034_;
  wire _31035_;
  wire _31036_;
  wire _31037_;
  wire _31038_;
  wire _31039_;
  wire _31040_;
  wire _31041_;
  wire _31042_;
  wire _31043_;
  wire _31044_;
  wire _31045_;
  wire _31046_;
  wire _31047_;
  wire _31048_;
  wire _31049_;
  wire _31050_;
  wire _31051_;
  wire _31052_;
  wire _31053_;
  wire _31054_;
  wire _31055_;
  wire _31056_;
  wire _31057_;
  wire _31058_;
  wire _31059_;
  wire _31060_;
  wire _31061_;
  wire _31062_;
  wire _31063_;
  wire _31064_;
  wire _31065_;
  wire _31066_;
  wire _31067_;
  wire _31068_;
  wire _31069_;
  wire _31070_;
  wire _31071_;
  wire _31072_;
  wire _31073_;
  wire _31074_;
  wire _31075_;
  wire _31076_;
  wire _31077_;
  wire _31078_;
  wire _31079_;
  wire _31080_;
  wire _31081_;
  wire _31082_;
  wire _31083_;
  wire _31084_;
  wire _31085_;
  wire _31086_;
  wire _31087_;
  wire _31088_;
  wire _31089_;
  wire _31090_;
  wire _31091_;
  wire _31092_;
  wire _31093_;
  wire _31094_;
  wire _31095_;
  wire _31096_;
  wire _31097_;
  wire _31098_;
  wire _31099_;
  wire _31100_;
  wire _31101_;
  wire _31102_;
  wire _31103_;
  wire _31104_;
  wire _31105_;
  wire _31106_;
  wire _31107_;
  wire _31108_;
  wire _31109_;
  wire _31110_;
  wire _31111_;
  wire _31112_;
  wire _31113_;
  wire _31114_;
  wire _31115_;
  wire _31116_;
  wire _31117_;
  wire _31118_;
  wire _31119_;
  wire _31120_;
  wire _31121_;
  wire _31122_;
  wire _31123_;
  wire _31124_;
  wire _31125_;
  wire _31126_;
  wire _31127_;
  wire _31128_;
  wire _31129_;
  wire _31130_;
  wire _31131_;
  wire _31132_;
  wire _31133_;
  wire _31134_;
  wire _31135_;
  wire _31136_;
  wire _31137_;
  wire _31138_;
  wire _31139_;
  wire _31140_;
  wire _31141_;
  wire _31142_;
  wire _31143_;
  wire _31144_;
  wire _31145_;
  wire _31146_;
  wire _31147_;
  wire _31148_;
  wire _31149_;
  wire _31150_;
  wire _31151_;
  wire _31152_;
  wire _31153_;
  wire _31154_;
  wire _31155_;
  wire _31156_;
  wire _31157_;
  wire _31158_;
  wire _31159_;
  wire _31160_;
  wire _31161_;
  wire _31162_;
  wire _31163_;
  wire _31164_;
  wire _31165_;
  wire _31166_;
  wire _31167_;
  wire _31168_;
  wire _31169_;
  wire _31170_;
  wire _31171_;
  wire _31172_;
  wire _31173_;
  wire _31174_;
  wire _31175_;
  wire _31176_;
  wire _31177_;
  wire _31178_;
  wire _31179_;
  wire _31180_;
  wire _31181_;
  wire _31182_;
  wire _31183_;
  wire _31184_;
  wire _31185_;
  wire _31186_;
  wire _31187_;
  wire _31188_;
  wire _31189_;
  wire _31190_;
  wire _31191_;
  wire _31192_;
  wire _31193_;
  wire _31194_;
  wire _31195_;
  wire _31196_;
  wire _31197_;
  wire _31198_;
  wire _31199_;
  wire _31200_;
  wire _31201_;
  wire _31202_;
  wire _31203_;
  wire _31204_;
  wire _31205_;
  wire _31206_;
  wire _31207_;
  wire _31208_;
  wire _31209_;
  wire _31210_;
  wire _31211_;
  wire _31212_;
  wire _31213_;
  wire _31214_;
  wire _31215_;
  wire _31216_;
  wire _31217_;
  wire _31218_;
  wire _31219_;
  wire _31220_;
  wire _31221_;
  wire _31222_;
  wire _31223_;
  wire _31224_;
  wire _31225_;
  wire _31226_;
  wire _31227_;
  wire _31228_;
  wire _31229_;
  wire _31230_;
  wire _31231_;
  wire _31232_;
  wire _31233_;
  wire _31234_;
  wire _31235_;
  wire _31236_;
  wire _31237_;
  wire _31238_;
  wire _31239_;
  wire _31240_;
  wire _31241_;
  wire _31242_;
  wire _31243_;
  wire _31244_;
  wire _31245_;
  wire _31246_;
  wire _31247_;
  wire _31248_;
  wire _31249_;
  wire _31250_;
  wire _31251_;
  wire _31252_;
  wire _31253_;
  wire _31254_;
  wire _31255_;
  wire _31256_;
  wire _31257_;
  wire _31258_;
  wire _31259_;
  wire _31260_;
  wire _31261_;
  wire _31262_;
  wire _31263_;
  wire _31264_;
  wire _31265_;
  wire _31266_;
  wire _31267_;
  wire _31268_;
  wire _31269_;
  wire _31270_;
  wire _31271_;
  wire _31272_;
  wire _31273_;
  wire _31274_;
  wire _31275_;
  wire _31276_;
  wire _31277_;
  wire _31278_;
  wire _31279_;
  wire _31280_;
  wire _31281_;
  wire _31282_;
  wire _31283_;
  wire _31284_;
  wire _31285_;
  wire _31286_;
  wire _31287_;
  wire _31288_;
  wire _31289_;
  wire _31290_;
  wire _31291_;
  wire _31292_;
  wire _31293_;
  wire _31294_;
  wire _31295_;
  wire _31296_;
  wire _31297_;
  wire _31298_;
  wire _31299_;
  wire _31300_;
  wire _31301_;
  wire _31302_;
  wire _31303_;
  wire _31304_;
  wire _31305_;
  wire _31306_;
  wire _31307_;
  wire _31308_;
  wire _31309_;
  wire _31310_;
  wire _31311_;
  wire _31312_;
  wire _31313_;
  wire _31314_;
  wire _31315_;
  wire _31316_;
  wire _31317_;
  wire _31318_;
  wire _31319_;
  wire _31320_;
  wire _31321_;
  wire _31322_;
  wire _31323_;
  wire _31324_;
  wire _31325_;
  wire _31326_;
  wire _31327_;
  wire _31328_;
  wire _31329_;
  wire _31330_;
  wire _31331_;
  wire _31332_;
  wire _31333_;
  wire _31334_;
  wire _31335_;
  wire _31336_;
  wire _31337_;
  wire _31338_;
  wire _31339_;
  wire _31340_;
  wire _31341_;
  wire _31342_;
  wire _31343_;
  wire _31344_;
  wire _31345_;
  wire _31346_;
  wire _31347_;
  wire _31348_;
  wire _31349_;
  wire _31350_;
  wire _31351_;
  wire _31352_;
  wire _31353_;
  wire _31354_;
  wire _31355_;
  wire _31356_;
  wire _31357_;
  wire _31358_;
  wire _31359_;
  wire _31360_;
  wire _31361_;
  wire _31362_;
  wire _31363_;
  wire _31364_;
  wire _31365_;
  wire _31366_;
  wire _31367_;
  wire _31368_;
  wire _31369_;
  wire _31370_;
  wire _31371_;
  wire _31372_;
  wire _31373_;
  wire _31374_;
  wire _31375_;
  wire _31376_;
  wire _31377_;
  wire _31378_;
  wire _31379_;
  wire _31380_;
  wire _31381_;
  wire _31382_;
  wire _31383_;
  wire _31384_;
  wire _31385_;
  wire _31386_;
  wire _31387_;
  wire _31388_;
  wire _31389_;
  wire _31390_;
  wire _31391_;
  wire _31392_;
  wire _31393_;
  wire _31394_;
  wire _31395_;
  wire _31396_;
  wire _31397_;
  wire _31398_;
  wire _31399_;
  wire _31400_;
  wire _31401_;
  wire _31402_;
  wire _31403_;
  wire _31404_;
  wire _31405_;
  wire _31406_;
  wire _31407_;
  wire _31408_;
  wire _31409_;
  wire _31410_;
  wire _31411_;
  wire _31412_;
  wire _31413_;
  wire _31414_;
  wire _31415_;
  wire _31416_;
  wire _31417_;
  wire _31418_;
  wire _31419_;
  wire _31420_;
  wire _31421_;
  wire _31422_;
  wire _31423_;
  wire _31424_;
  wire _31425_;
  wire _31426_;
  wire _31427_;
  wire _31428_;
  wire _31429_;
  wire _31430_;
  wire _31431_;
  wire _31432_;
  wire _31433_;
  wire _31434_;
  wire _31435_;
  wire _31436_;
  wire _31437_;
  wire _31438_;
  wire _31439_;
  wire _31440_;
  wire _31441_;
  wire _31442_;
  wire _31443_;
  wire _31444_;
  wire _31445_;
  wire _31446_;
  wire _31447_;
  wire _31448_;
  wire _31449_;
  wire _31450_;
  wire _31451_;
  wire _31452_;
  wire _31453_;
  wire _31454_;
  wire _31455_;
  wire _31456_;
  wire _31457_;
  wire _31458_;
  wire _31459_;
  wire _31460_;
  wire _31461_;
  wire _31462_;
  wire _31463_;
  wire _31464_;
  wire _31465_;
  wire _31466_;
  wire _31467_;
  wire _31468_;
  wire _31469_;
  wire _31470_;
  wire _31471_;
  wire _31472_;
  wire _31473_;
  wire _31474_;
  wire _31475_;
  wire _31476_;
  wire _31477_;
  wire _31478_;
  wire _31479_;
  wire _31480_;
  wire _31481_;
  wire _31482_;
  wire _31483_;
  wire _31484_;
  wire _31485_;
  wire _31486_;
  wire _31487_;
  wire _31488_;
  wire _31489_;
  wire _31490_;
  wire _31491_;
  wire _31492_;
  wire _31493_;
  wire _31494_;
  wire _31495_;
  wire _31496_;
  wire _31497_;
  wire _31498_;
  wire _31499_;
  wire _31500_;
  wire _31501_;
  wire _31502_;
  wire _31503_;
  wire _31504_;
  wire _31505_;
  wire _31506_;
  wire _31507_;
  wire _31508_;
  wire _31509_;
  wire _31510_;
  wire _31511_;
  wire _31512_;
  wire _31513_;
  wire _31514_;
  wire _31515_;
  wire _31516_;
  wire _31517_;
  wire _31518_;
  wire _31519_;
  wire _31520_;
  wire _31521_;
  wire _31522_;
  wire _31523_;
  wire _31524_;
  wire _31525_;
  wire _31526_;
  wire _31527_;
  wire _31528_;
  wire _31529_;
  wire _31530_;
  wire _31531_;
  wire _31532_;
  wire _31533_;
  wire _31534_;
  wire _31535_;
  wire _31536_;
  wire _31537_;
  wire _31538_;
  wire _31539_;
  wire _31540_;
  wire _31541_;
  wire _31542_;
  wire _31543_;
  wire _31544_;
  wire _31545_;
  wire _31546_;
  wire _31547_;
  wire _31548_;
  wire _31549_;
  wire _31550_;
  wire _31551_;
  wire _31552_;
  wire _31553_;
  wire _31554_;
  wire _31555_;
  wire _31556_;
  wire _31557_;
  wire _31558_;
  wire _31559_;
  wire _31560_;
  wire _31561_;
  wire _31562_;
  wire _31563_;
  wire _31564_;
  wire _31565_;
  wire _31566_;
  wire _31567_;
  wire _31568_;
  wire _31569_;
  wire _31570_;
  wire _31571_;
  wire _31572_;
  wire _31573_;
  wire _31574_;
  wire _31575_;
  wire _31576_;
  wire _31577_;
  wire _31578_;
  wire _31579_;
  wire _31580_;
  wire _31581_;
  wire _31582_;
  wire _31583_;
  wire _31584_;
  wire _31585_;
  wire _31586_;
  wire _31587_;
  wire _31588_;
  wire _31589_;
  wire _31590_;
  wire _31591_;
  wire _31592_;
  wire _31593_;
  wire _31594_;
  wire _31595_;
  wire _31596_;
  wire _31597_;
  wire _31598_;
  wire _31599_;
  wire _31600_;
  wire _31601_;
  wire _31602_;
  wire _31603_;
  wire _31604_;
  wire _31605_;
  wire _31606_;
  wire _31607_;
  wire _31608_;
  wire _31609_;
  wire _31610_;
  wire _31611_;
  wire _31612_;
  wire _31613_;
  wire _31614_;
  wire _31615_;
  wire _31616_;
  wire _31617_;
  wire _31618_;
  wire _31619_;
  wire _31620_;
  wire _31621_;
  wire _31622_;
  wire _31623_;
  wire _31624_;
  wire _31625_;
  wire _31626_;
  wire _31627_;
  wire _31628_;
  wire _31629_;
  wire _31630_;
  wire _31631_;
  wire _31632_;
  wire _31633_;
  wire _31634_;
  wire _31635_;
  wire _31636_;
  wire _31637_;
  wire _31638_;
  wire _31639_;
  wire _31640_;
  wire _31641_;
  wire _31642_;
  wire _31643_;
  wire _31644_;
  wire _31645_;
  wire _31646_;
  wire _31647_;
  wire _31648_;
  wire _31649_;
  wire _31650_;
  wire _31651_;
  wire _31652_;
  wire _31653_;
  wire _31654_;
  wire _31655_;
  wire _31656_;
  wire _31657_;
  wire _31658_;
  wire _31659_;
  wire _31660_;
  wire _31661_;
  wire _31662_;
  wire _31663_;
  wire _31664_;
  wire _31665_;
  wire _31666_;
  wire _31667_;
  wire _31668_;
  wire _31669_;
  wire _31670_;
  wire _31671_;
  wire _31672_;
  wire _31673_;
  wire _31674_;
  wire _31675_;
  wire _31676_;
  wire _31677_;
  wire _31678_;
  wire _31679_;
  wire _31680_;
  wire _31681_;
  wire _31682_;
  wire _31683_;
  wire _31684_;
  wire _31685_;
  wire _31686_;
  wire _31687_;
  wire _31688_;
  wire _31689_;
  wire _31690_;
  wire _31691_;
  wire _31692_;
  wire _31693_;
  wire _31694_;
  wire _31695_;
  wire _31696_;
  wire _31697_;
  wire _31698_;
  wire _31699_;
  wire _31700_;
  wire _31701_;
  wire _31702_;
  wire _31703_;
  wire _31704_;
  wire _31705_;
  wire _31706_;
  wire _31707_;
  wire _31708_;
  wire _31709_;
  wire _31710_;
  wire _31711_;
  wire _31712_;
  wire _31713_;
  wire _31714_;
  wire _31715_;
  wire _31716_;
  wire _31717_;
  wire _31718_;
  wire _31719_;
  wire _31720_;
  wire _31721_;
  wire _31722_;
  wire _31723_;
  wire _31724_;
  wire _31725_;
  wire _31726_;
  wire _31727_;
  wire _31728_;
  wire _31729_;
  wire _31730_;
  wire _31731_;
  wire _31732_;
  wire _31733_;
  wire _31734_;
  wire _31735_;
  wire _31736_;
  wire _31737_;
  wire _31738_;
  wire _31739_;
  wire _31740_;
  wire _31741_;
  wire _31742_;
  wire _31743_;
  wire _31744_;
  wire _31745_;
  wire _31746_;
  wire _31747_;
  wire _31748_;
  wire _31749_;
  wire _31750_;
  wire _31751_;
  wire _31752_;
  wire _31753_;
  wire _31754_;
  wire _31755_;
  wire _31756_;
  wire _31757_;
  wire _31758_;
  wire _31759_;
  wire _31760_;
  wire _31761_;
  wire _31762_;
  wire _31763_;
  wire _31764_;
  wire _31765_;
  wire _31766_;
  wire _31767_;
  wire _31768_;
  wire _31769_;
  wire _31770_;
  wire _31771_;
  wire _31772_;
  wire _31773_;
  wire _31774_;
  wire _31775_;
  wire _31776_;
  wire _31777_;
  wire _31778_;
  wire _31779_;
  wire _31780_;
  wire _31781_;
  wire _31782_;
  wire _31783_;
  wire _31784_;
  wire _31785_;
  wire _31786_;
  wire _31787_;
  wire _31788_;
  wire _31789_;
  wire _31790_;
  wire _31791_;
  wire _31792_;
  wire _31793_;
  wire _31794_;
  wire _31795_;
  wire _31796_;
  wire _31797_;
  wire _31798_;
  wire _31799_;
  wire _31800_;
  wire _31801_;
  wire _31802_;
  wire _31803_;
  wire _31804_;
  wire _31805_;
  wire _31806_;
  wire _31807_;
  wire _31808_;
  wire _31809_;
  wire _31810_;
  wire _31811_;
  wire _31812_;
  wire _31813_;
  wire _31814_;
  wire _31815_;
  wire _31816_;
  wire _31817_;
  wire _31818_;
  wire _31819_;
  wire _31820_;
  wire _31821_;
  wire _31822_;
  wire _31823_;
  wire _31824_;
  wire _31825_;
  wire _31826_;
  wire _31827_;
  wire _31828_;
  wire _31829_;
  wire _31830_;
  wire _31831_;
  wire _31832_;
  wire _31833_;
  wire _31834_;
  wire _31835_;
  wire _31836_;
  wire _31837_;
  wire _31838_;
  wire _31839_;
  wire _31840_;
  wire _31841_;
  wire _31842_;
  wire _31843_;
  wire _31844_;
  wire _31845_;
  wire _31846_;
  wire _31847_;
  wire _31848_;
  wire _31849_;
  wire _31850_;
  wire _31851_;
  wire _31852_;
  wire _31853_;
  wire _31854_;
  wire _31855_;
  wire _31856_;
  wire _31857_;
  wire _31858_;
  wire _31859_;
  wire _31860_;
  wire _31861_;
  wire _31862_;
  wire _31863_;
  wire _31864_;
  wire _31865_;
  wire _31866_;
  wire _31867_;
  wire _31868_;
  wire _31869_;
  wire _31870_;
  wire _31871_;
  wire _31872_;
  wire _31873_;
  wire _31874_;
  wire _31875_;
  wire _31876_;
  wire _31877_;
  wire _31878_;
  wire _31879_;
  wire _31880_;
  wire _31881_;
  wire _31882_;
  wire _31883_;
  wire _31884_;
  wire _31885_;
  wire _31886_;
  wire _31887_;
  wire _31888_;
  wire _31889_;
  wire _31890_;
  wire _31891_;
  wire _31892_;
  wire _31893_;
  wire _31894_;
  wire _31895_;
  wire _31896_;
  wire _31897_;
  wire _31898_;
  wire _31899_;
  wire _31900_;
  wire _31901_;
  wire _31902_;
  wire _31903_;
  wire _31904_;
  wire _31905_;
  wire _31906_;
  wire _31907_;
  wire _31908_;
  wire _31909_;
  wire _31910_;
  wire _31911_;
  wire _31912_;
  wire _31913_;
  wire _31914_;
  wire _31915_;
  wire _31916_;
  wire _31917_;
  wire _31918_;
  wire _31919_;
  wire _31920_;
  wire _31921_;
  wire _31922_;
  wire _31923_;
  wire _31924_;
  wire _31925_;
  wire _31926_;
  wire _31927_;
  wire _31928_;
  wire _31929_;
  wire _31930_;
  wire _31931_;
  wire _31932_;
  wire _31933_;
  wire _31934_;
  wire _31935_;
  wire _31936_;
  wire _31937_;
  wire _31938_;
  wire _31939_;
  wire _31940_;
  wire _31941_;
  wire _31942_;
  wire _31943_;
  wire _31944_;
  wire _31945_;
  wire _31946_;
  wire _31947_;
  wire _31948_;
  wire _31949_;
  wire _31950_;
  wire _31951_;
  wire _31952_;
  wire _31953_;
  wire _31954_;
  wire _31955_;
  wire _31956_;
  wire _31957_;
  wire _31958_;
  wire _31959_;
  wire _31960_;
  wire _31961_;
  wire _31962_;
  wire _31963_;
  wire _31964_;
  wire _31965_;
  wire _31966_;
  wire _31967_;
  wire _31968_;
  wire _31969_;
  wire _31970_;
  wire _31971_;
  wire _31972_;
  wire _31973_;
  wire _31974_;
  wire _31975_;
  wire _31976_;
  wire _31977_;
  wire _31978_;
  wire _31979_;
  wire _31980_;
  wire _31981_;
  wire _31982_;
  wire _31983_;
  wire _31984_;
  wire _31985_;
  wire _31986_;
  wire _31987_;
  wire _31988_;
  wire _31989_;
  wire _31990_;
  wire _31991_;
  wire _31992_;
  wire _31993_;
  wire _31994_;
  wire _31995_;
  wire _31996_;
  wire _31997_;
  wire _31998_;
  wire _31999_;
  wire _32000_;
  wire _32001_;
  wire _32002_;
  wire _32003_;
  wire _32004_;
  wire _32005_;
  wire _32006_;
  wire _32007_;
  wire _32008_;
  wire _32009_;
  wire _32010_;
  wire _32011_;
  wire _32012_;
  wire _32013_;
  wire _32014_;
  wire _32015_;
  wire _32016_;
  wire _32017_;
  wire _32018_;
  wire _32019_;
  wire _32020_;
  wire _32021_;
  wire _32022_;
  wire _32023_;
  wire _32024_;
  wire _32025_;
  wire _32026_;
  wire _32027_;
  wire _32028_;
  wire _32029_;
  wire _32030_;
  wire _32031_;
  wire _32032_;
  wire _32033_;
  wire _32034_;
  wire _32035_;
  wire _32036_;
  wire _32037_;
  wire _32038_;
  wire _32039_;
  wire _32040_;
  wire _32041_;
  wire _32042_;
  wire _32043_;
  wire _32044_;
  wire _32045_;
  wire _32046_;
  wire _32047_;
  wire _32048_;
  wire _32049_;
  wire _32050_;
  wire _32051_;
  wire _32052_;
  wire _32053_;
  wire _32054_;
  wire _32055_;
  wire _32056_;
  wire _32057_;
  wire _32058_;
  wire _32059_;
  wire _32060_;
  wire _32061_;
  wire _32062_;
  wire _32063_;
  wire _32064_;
  wire _32065_;
  wire _32066_;
  wire _32067_;
  wire _32068_;
  wire _32069_;
  wire _32070_;
  wire _32071_;
  wire _32072_;
  wire _32073_;
  wire _32074_;
  wire _32075_;
  wire _32076_;
  wire _32077_;
  wire _32078_;
  wire _32079_;
  wire _32080_;
  wire _32081_;
  wire _32082_;
  wire _32083_;
  wire _32084_;
  wire _32085_;
  wire _32086_;
  wire _32087_;
  wire _32088_;
  wire _32089_;
  wire _32090_;
  wire _32091_;
  wire _32092_;
  wire _32093_;
  wire _32094_;
  wire _32095_;
  wire _32096_;
  wire _32097_;
  wire _32098_;
  wire _32099_;
  wire _32100_;
  wire _32101_;
  wire _32102_;
  wire _32103_;
  wire _32104_;
  wire _32105_;
  wire _32106_;
  wire _32107_;
  wire _32108_;
  wire _32109_;
  wire _32110_;
  wire _32111_;
  wire _32112_;
  wire _32113_;
  wire _32114_;
  wire _32115_;
  wire _32116_;
  wire _32117_;
  wire _32118_;
  wire _32119_;
  wire _32120_;
  wire _32121_;
  wire _32122_;
  wire _32123_;
  wire _32124_;
  wire _32125_;
  wire _32126_;
  wire _32127_;
  wire _32128_;
  wire _32129_;
  wire _32130_;
  wire _32131_;
  wire _32132_;
  wire _32133_;
  wire _32134_;
  wire _32135_;
  wire _32136_;
  wire _32137_;
  wire _32138_;
  wire _32139_;
  wire _32140_;
  wire _32141_;
  wire _32142_;
  wire _32143_;
  wire _32144_;
  wire _32145_;
  wire _32146_;
  wire _32147_;
  wire _32148_;
  wire _32149_;
  wire _32150_;
  wire _32151_;
  wire _32152_;
  wire _32153_;
  wire _32154_;
  wire _32155_;
  wire _32156_;
  wire _32157_;
  wire _32158_;
  wire _32159_;
  wire _32160_;
  wire _32161_;
  wire _32162_;
  wire _32163_;
  wire _32164_;
  wire _32165_;
  wire _32166_;
  wire _32167_;
  wire _32168_;
  wire _32169_;
  wire _32170_;
  wire _32171_;
  wire _32172_;
  wire _32173_;
  wire _32174_;
  wire _32175_;
  wire _32176_;
  wire _32177_;
  wire _32178_;
  wire _32179_;
  wire _32180_;
  wire _32181_;
  wire _32182_;
  wire _32183_;
  wire _32184_;
  wire _32185_;
  wire _32186_;
  wire _32187_;
  wire _32188_;
  wire _32189_;
  wire _32190_;
  wire _32191_;
  wire _32192_;
  wire _32193_;
  wire _32194_;
  wire _32195_;
  wire _32196_;
  wire _32197_;
  wire _32198_;
  wire _32199_;
  wire _32200_;
  wire _32201_;
  wire _32202_;
  wire _32203_;
  wire _32204_;
  wire _32205_;
  wire _32206_;
  wire _32207_;
  wire _32208_;
  wire _32209_;
  wire _32210_;
  wire _32211_;
  wire _32212_;
  wire _32213_;
  wire _32214_;
  wire _32215_;
  wire _32216_;
  wire _32217_;
  wire _32218_;
  wire _32219_;
  wire _32220_;
  wire _32221_;
  wire _32222_;
  wire _32223_;
  wire _32224_;
  wire _32225_;
  wire _32226_;
  wire _32227_;
  wire _32228_;
  wire _32229_;
  wire _32230_;
  wire _32231_;
  wire _32232_;
  wire _32233_;
  wire _32234_;
  wire _32235_;
  wire _32236_;
  wire _32237_;
  wire _32238_;
  wire _32239_;
  wire _32240_;
  wire _32241_;
  wire _32242_;
  wire _32243_;
  wire _32244_;
  wire _32245_;
  wire _32246_;
  wire _32247_;
  wire _32248_;
  wire _32249_;
  wire _32250_;
  wire _32251_;
  wire _32252_;
  wire _32253_;
  wire _32254_;
  wire _32255_;
  wire _32256_;
  wire _32257_;
  wire _32258_;
  wire _32259_;
  wire _32260_;
  wire _32261_;
  wire _32262_;
  wire _32263_;
  wire _32264_;
  wire _32265_;
  wire _32266_;
  wire _32267_;
  wire _32268_;
  wire _32269_;
  wire _32270_;
  wire _32271_;
  wire _32272_;
  wire _32273_;
  wire _32274_;
  wire _32275_;
  wire _32276_;
  wire _32277_;
  wire _32278_;
  wire _32279_;
  wire _32280_;
  wire _32281_;
  wire _32282_;
  wire _32283_;
  wire _32284_;
  wire _32285_;
  wire _32286_;
  wire _32287_;
  wire _32288_;
  wire _32289_;
  wire _32290_;
  wire _32291_;
  wire _32292_;
  wire _32293_;
  wire _32294_;
  wire _32295_;
  wire _32296_;
  wire _32297_;
  wire _32298_;
  wire _32299_;
  wire _32300_;
  wire _32301_;
  wire _32302_;
  wire _32303_;
  wire _32304_;
  wire _32305_;
  wire _32306_;
  wire _32307_;
  wire _32308_;
  wire _32309_;
  wire _32310_;
  wire _32311_;
  wire _32312_;
  wire _32313_;
  wire _32314_;
  wire _32315_;
  wire _32316_;
  wire _32317_;
  wire _32318_;
  wire _32319_;
  wire _32320_;
  wire _32321_;
  wire _32322_;
  wire _32323_;
  wire _32324_;
  wire _32325_;
  wire _32326_;
  wire _32327_;
  wire _32328_;
  wire _32329_;
  wire _32330_;
  wire _32331_;
  wire _32332_;
  wire _32333_;
  wire _32334_;
  wire _32335_;
  wire _32336_;
  wire _32337_;
  wire _32338_;
  wire _32339_;
  wire _32340_;
  wire _32341_;
  wire _32342_;
  wire _32343_;
  wire _32344_;
  wire _32345_;
  wire _32346_;
  wire _32347_;
  wire _32348_;
  wire _32349_;
  wire _32350_;
  wire _32351_;
  wire _32352_;
  wire _32353_;
  wire _32354_;
  wire _32355_;
  wire _32356_;
  wire _32357_;
  wire _32358_;
  wire _32359_;
  wire _32360_;
  wire _32361_;
  wire _32362_;
  wire _32363_;
  wire _32364_;
  wire _32365_;
  wire _32366_;
  wire _32367_;
  wire _32368_;
  wire _32369_;
  wire _32370_;
  wire _32371_;
  wire _32372_;
  wire _32373_;
  wire _32374_;
  wire _32375_;
  wire _32376_;
  wire _32377_;
  wire _32378_;
  wire _32379_;
  wire _32380_;
  wire _32381_;
  wire _32382_;
  wire _32383_;
  wire _32384_;
  wire _32385_;
  wire _32386_;
  wire _32387_;
  wire _32388_;
  wire _32389_;
  wire _32390_;
  wire _32391_;
  wire _32392_;
  wire _32393_;
  wire _32394_;
  wire _32395_;
  wire _32396_;
  wire _32397_;
  wire _32398_;
  wire _32399_;
  wire _32400_;
  wire _32401_;
  wire _32402_;
  wire _32403_;
  wire _32404_;
  wire _32405_;
  wire _32406_;
  wire _32407_;
  wire _32408_;
  wire _32409_;
  wire _32410_;
  wire _32411_;
  wire _32412_;
  wire _32413_;
  wire _32414_;
  wire _32415_;
  wire _32416_;
  wire _32417_;
  wire _32418_;
  wire _32419_;
  wire _32420_;
  wire _32421_;
  wire _32422_;
  wire _32423_;
  wire _32424_;
  wire _32425_;
  wire _32426_;
  wire _32427_;
  wire _32428_;
  wire _32429_;
  wire _32430_;
  wire _32431_;
  wire _32432_;
  wire _32433_;
  wire _32434_;
  wire _32435_;
  wire _32436_;
  wire _32437_;
  wire _32438_;
  wire _32439_;
  wire _32440_;
  wire _32441_;
  wire _32442_;
  wire _32443_;
  wire _32444_;
  wire _32445_;
  wire _32446_;
  wire _32447_;
  wire _32448_;
  wire _32449_;
  wire _32450_;
  wire _32451_;
  wire _32452_;
  wire _32453_;
  wire _32454_;
  wire _32455_;
  wire _32456_;
  wire _32457_;
  wire _32458_;
  wire _32459_;
  wire _32460_;
  wire _32461_;
  wire _32462_;
  wire _32463_;
  wire _32464_;
  wire _32465_;
  wire _32466_;
  wire _32467_;
  wire _32468_;
  wire _32469_;
  wire _32470_;
  wire _32471_;
  wire _32472_;
  wire _32473_;
  wire _32474_;
  wire _32475_;
  wire _32476_;
  wire _32477_;
  wire _32478_;
  wire _32479_;
  wire _32480_;
  wire _32481_;
  wire _32482_;
  wire _32483_;
  wire _32484_;
  wire _32485_;
  wire _32486_;
  wire _32487_;
  wire _32488_;
  wire _32489_;
  wire _32490_;
  wire _32491_;
  wire _32492_;
  wire _32493_;
  wire _32494_;
  wire _32495_;
  wire _32496_;
  wire _32497_;
  wire _32498_;
  wire _32499_;
  wire _32500_;
  wire _32501_;
  wire _32502_;
  wire _32503_;
  wire _32504_;
  wire _32505_;
  wire _32506_;
  wire _32507_;
  wire _32508_;
  wire _32509_;
  wire _32510_;
  wire _32511_;
  wire _32512_;
  wire _32513_;
  wire _32514_;
  wire _32515_;
  wire _32516_;
  wire _32517_;
  wire _32518_;
  wire _32519_;
  wire _32520_;
  wire _32521_;
  wire _32522_;
  wire _32523_;
  wire _32524_;
  wire _32525_;
  wire _32526_;
  wire _32527_;
  wire _32528_;
  wire _32529_;
  wire _32530_;
  wire _32531_;
  wire _32532_;
  wire _32533_;
  wire _32534_;
  wire _32535_;
  wire _32536_;
  wire _32537_;
  wire _32538_;
  wire _32539_;
  wire _32540_;
  wire _32541_;
  wire _32542_;
  wire _32543_;
  wire _32544_;
  wire _32545_;
  wire _32546_;
  wire _32547_;
  wire _32548_;
  wire _32549_;
  wire _32550_;
  wire _32551_;
  wire _32552_;
  wire _32553_;
  wire _32554_;
  wire _32555_;
  wire _32556_;
  wire _32557_;
  wire _32558_;
  wire _32559_;
  wire _32560_;
  wire _32561_;
  wire _32562_;
  wire _32563_;
  wire _32564_;
  wire _32565_;
  wire _32566_;
  wire _32567_;
  wire _32568_;
  wire _32569_;
  wire _32570_;
  wire _32571_;
  wire _32572_;
  wire _32573_;
  wire _32574_;
  wire _32575_;
  wire _32576_;
  wire _32577_;
  wire _32578_;
  wire _32579_;
  wire _32580_;
  wire _32581_;
  wire _32582_;
  wire _32583_;
  wire _32584_;
  wire _32585_;
  wire _32586_;
  wire _32587_;
  wire _32588_;
  wire _32589_;
  wire _32590_;
  wire _32591_;
  wire _32592_;
  wire _32593_;
  wire _32594_;
  wire _32595_;
  wire _32596_;
  wire _32597_;
  wire _32598_;
  wire _32599_;
  wire _32600_;
  wire _32601_;
  wire _32602_;
  wire _32603_;
  wire _32604_;
  wire _32605_;
  wire _32606_;
  wire _32607_;
  wire _32608_;
  wire _32609_;
  wire _32610_;
  wire _32611_;
  wire _32612_;
  wire _32613_;
  wire _32614_;
  wire _32615_;
  wire _32616_;
  wire _32617_;
  wire _32618_;
  wire _32619_;
  wire _32620_;
  wire _32621_;
  wire _32622_;
  wire _32623_;
  wire _32624_;
  wire _32625_;
  wire _32626_;
  wire _32627_;
  wire _32628_;
  wire _32629_;
  wire _32630_;
  wire _32631_;
  wire _32632_;
  wire _32633_;
  wire _32634_;
  wire _32635_;
  wire _32636_;
  wire _32637_;
  wire _32638_;
  wire _32639_;
  wire _32640_;
  wire _32641_;
  wire _32642_;
  wire _32643_;
  wire _32644_;
  wire _32645_;
  wire _32646_;
  wire _32647_;
  wire _32648_;
  wire _32649_;
  wire _32650_;
  wire _32651_;
  wire _32652_;
  wire _32653_;
  wire _32654_;
  wire _32655_;
  wire _32656_;
  wire _32657_;
  wire _32658_;
  wire _32659_;
  wire _32660_;
  wire _32661_;
  wire _32662_;
  wire _32663_;
  wire _32664_;
  wire _32665_;
  wire _32666_;
  wire _32667_;
  wire _32668_;
  wire _32669_;
  wire _32670_;
  wire _32671_;
  wire _32672_;
  wire _32673_;
  wire _32674_;
  wire _32675_;
  wire _32676_;
  wire _32677_;
  wire _32678_;
  wire _32679_;
  wire _32680_;
  wire _32681_;
  wire _32682_;
  wire _32683_;
  wire _32684_;
  wire _32685_;
  wire _32686_;
  wire _32687_;
  wire _32688_;
  wire _32689_;
  wire _32690_;
  wire _32691_;
  wire _32692_;
  wire _32693_;
  wire _32694_;
  wire _32695_;
  wire _32696_;
  wire _32697_;
  wire _32698_;
  wire _32699_;
  wire _32700_;
  wire _32701_;
  wire _32702_;
  wire _32703_;
  wire _32704_;
  wire _32705_;
  wire _32706_;
  wire _32707_;
  wire _32708_;
  wire _32709_;
  wire _32710_;
  wire _32711_;
  wire _32712_;
  wire _32713_;
  wire _32714_;
  wire _32715_;
  wire _32716_;
  wire _32717_;
  wire _32718_;
  wire _32719_;
  wire _32720_;
  wire _32721_;
  wire _32722_;
  wire _32723_;
  wire _32724_;
  wire _32725_;
  wire _32726_;
  wire _32727_;
  wire _32728_;
  wire _32729_;
  wire _32730_;
  wire _32731_;
  wire _32732_;
  wire _32733_;
  wire _32734_;
  wire _32735_;
  wire _32736_;
  wire _32737_;
  wire _32738_;
  wire _32739_;
  wire _32740_;
  wire _32741_;
  wire _32742_;
  wire _32743_;
  wire _32744_;
  wire _32745_;
  wire _32746_;
  wire _32747_;
  wire _32748_;
  wire _32749_;
  wire _32750_;
  wire _32751_;
  wire _32752_;
  wire _32753_;
  wire _32754_;
  wire _32755_;
  wire _32756_;
  wire _32757_;
  wire _32758_;
  wire _32759_;
  wire _32760_;
  wire _32761_;
  wire _32762_;
  wire _32763_;
  wire _32764_;
  wire _32765_;
  wire _32766_;
  wire _32767_;
  wire _32768_;
  wire _32769_;
  wire _32770_;
  wire _32771_;
  wire _32772_;
  wire _32773_;
  wire _32774_;
  wire _32775_;
  wire _32776_;
  wire _32777_;
  wire _32778_;
  wire _32779_;
  wire _32780_;
  wire _32781_;
  wire _32782_;
  wire _32783_;
  wire _32784_;
  wire _32785_;
  wire _32786_;
  wire _32787_;
  wire _32788_;
  wire _32789_;
  wire _32790_;
  wire _32791_;
  wire _32792_;
  wire _32793_;
  wire _32794_;
  wire _32795_;
  wire _32796_;
  wire _32797_;
  wire _32798_;
  wire _32799_;
  wire _32800_;
  wire _32801_;
  wire _32802_;
  wire _32803_;
  wire _32804_;
  wire _32805_;
  wire _32806_;
  wire _32807_;
  wire _32808_;
  wire _32809_;
  wire _32810_;
  wire _32811_;
  wire _32812_;
  wire _32813_;
  wire _32814_;
  wire _32815_;
  wire _32816_;
  wire _32817_;
  wire _32818_;
  wire _32819_;
  wire _32820_;
  wire _32821_;
  wire _32822_;
  wire _32823_;
  wire _32824_;
  wire _32825_;
  wire _32826_;
  wire _32827_;
  wire _32828_;
  wire _32829_;
  wire _32830_;
  wire _32831_;
  wire _32832_;
  wire _32833_;
  wire _32834_;
  wire _32835_;
  wire _32836_;
  wire _32837_;
  wire _32838_;
  wire _32839_;
  wire _32840_;
  wire _32841_;
  wire _32842_;
  wire _32843_;
  wire _32844_;
  wire _32845_;
  wire _32846_;
  wire _32847_;
  wire _32848_;
  wire _32849_;
  wire _32850_;
  wire _32851_;
  wire _32852_;
  wire _32853_;
  wire _32854_;
  wire _32855_;
  wire _32856_;
  wire _32857_;
  wire _32858_;
  wire _32859_;
  wire _32860_;
  wire _32861_;
  wire _32862_;
  wire _32863_;
  wire _32864_;
  wire _32865_;
  wire _32866_;
  wire _32867_;
  wire _32868_;
  wire _32869_;
  wire _32870_;
  wire _32871_;
  wire _32872_;
  wire _32873_;
  wire _32874_;
  wire _32875_;
  wire _32876_;
  wire _32877_;
  wire _32878_;
  wire _32879_;
  wire _32880_;
  wire _32881_;
  wire _32882_;
  wire _32883_;
  wire _32884_;
  wire _32885_;
  wire _32886_;
  wire _32887_;
  wire _32888_;
  wire _32889_;
  wire _32890_;
  wire _32891_;
  wire _32892_;
  wire _32893_;
  wire _32894_;
  wire _32895_;
  wire _32896_;
  wire _32897_;
  wire _32898_;
  wire _32899_;
  wire _32900_;
  wire _32901_;
  wire _32902_;
  wire _32903_;
  wire _32904_;
  wire _32905_;
  wire _32906_;
  wire _32907_;
  wire _32908_;
  wire _32909_;
  wire _32910_;
  wire _32911_;
  wire _32912_;
  wire _32913_;
  wire _32914_;
  wire _32915_;
  wire _32916_;
  wire _32917_;
  wire _32918_;
  wire _32919_;
  wire _32920_;
  wire _32921_;
  wire _32922_;
  wire _32923_;
  wire _32924_;
  wire _32925_;
  wire _32926_;
  wire _32927_;
  wire _32928_;
  wire _32929_;
  wire _32930_;
  wire _32931_;
  wire _32932_;
  wire _32933_;
  wire _32934_;
  wire _32935_;
  wire _32936_;
  wire _32937_;
  wire _32938_;
  wire _32939_;
  wire _32940_;
  wire _32941_;
  wire _32942_;
  wire _32943_;
  wire _32944_;
  wire _32945_;
  wire _32946_;
  wire _32947_;
  wire _32948_;
  wire _32949_;
  wire _32950_;
  wire _32951_;
  wire _32952_;
  wire _32953_;
  wire _32954_;
  wire _32955_;
  wire _32956_;
  wire _32957_;
  wire _32958_;
  wire _32959_;
  wire _32960_;
  wire _32961_;
  wire _32962_;
  wire _32963_;
  wire _32964_;
  wire _32965_;
  wire _32966_;
  wire _32967_;
  wire _32968_;
  wire _32969_;
  wire _32970_;
  wire _32971_;
  wire _32972_;
  wire _32973_;
  wire _32974_;
  wire _32975_;
  wire _32976_;
  wire _32977_;
  wire _32978_;
  wire _32979_;
  wire _32980_;
  wire _32981_;
  wire _32982_;
  wire _32983_;
  wire _32984_;
  wire _32985_;
  wire _32986_;
  wire _32987_;
  wire _32988_;
  wire _32989_;
  wire _32990_;
  wire _32991_;
  wire _32992_;
  wire _32993_;
  wire _32994_;
  wire _32995_;
  wire _32996_;
  wire _32997_;
  wire _32998_;
  wire _32999_;
  wire _33000_;
  wire _33001_;
  wire _33002_;
  wire _33003_;
  wire _33004_;
  wire _33005_;
  wire _33006_;
  wire _33007_;
  wire _33008_;
  wire _33009_;
  wire _33010_;
  wire _33011_;
  wire _33012_;
  wire _33013_;
  wire _33014_;
  wire _33015_;
  wire _33016_;
  wire _33017_;
  wire _33018_;
  wire _33019_;
  wire _33020_;
  wire _33021_;
  wire _33022_;
  wire _33023_;
  wire _33024_;
  wire _33025_;
  wire _33026_;
  wire _33027_;
  wire _33028_;
  wire _33029_;
  wire _33030_;
  wire _33031_;
  wire _33032_;
  wire _33033_;
  wire _33034_;
  wire _33035_;
  wire _33036_;
  wire _33037_;
  wire _33038_;
  wire _33039_;
  wire _33040_;
  wire _33041_;
  wire _33042_;
  wire _33043_;
  wire _33044_;
  wire _33045_;
  wire _33046_;
  wire _33047_;
  wire _33048_;
  wire _33049_;
  wire _33050_;
  wire _33051_;
  wire _33052_;
  wire _33053_;
  wire _33054_;
  wire _33055_;
  wire _33056_;
  wire _33057_;
  wire _33058_;
  wire _33059_;
  wire _33060_;
  wire _33061_;
  wire _33062_;
  wire _33063_;
  wire _33064_;
  wire _33065_;
  wire _33066_;
  wire _33067_;
  wire _33068_;
  wire _33069_;
  wire _33070_;
  wire _33071_;
  wire _33072_;
  wire _33073_;
  wire _33074_;
  wire _33075_;
  wire _33076_;
  wire _33077_;
  wire _33078_;
  wire _33079_;
  wire _33080_;
  wire _33081_;
  wire _33082_;
  wire _33083_;
  wire _33084_;
  wire _33085_;
  wire _33086_;
  wire _33087_;
  wire _33088_;
  wire _33089_;
  wire _33090_;
  wire _33091_;
  wire _33092_;
  wire _33093_;
  wire _33094_;
  wire _33095_;
  wire _33096_;
  wire _33097_;
  wire _33098_;
  wire _33099_;
  wire _33100_;
  wire _33101_;
  wire _33102_;
  wire _33103_;
  wire _33104_;
  wire _33105_;
  wire _33106_;
  wire _33107_;
  wire _33108_;
  wire _33109_;
  wire _33110_;
  wire _33111_;
  wire _33112_;
  wire _33113_;
  wire _33114_;
  wire _33115_;
  wire _33116_;
  wire _33117_;
  wire _33118_;
  wire _33119_;
  wire _33120_;
  wire _33121_;
  wire _33122_;
  wire _33123_;
  wire _33124_;
  wire _33125_;
  wire _33126_;
  wire _33127_;
  wire _33128_;
  wire _33129_;
  wire _33130_;
  wire _33131_;
  wire _33132_;
  wire _33133_;
  wire _33134_;
  wire _33135_;
  wire _33136_;
  wire _33137_;
  wire _33138_;
  wire _33139_;
  wire _33140_;
  wire _33141_;
  wire _33142_;
  wire _33143_;
  wire _33144_;
  wire _33145_;
  wire _33146_;
  wire _33147_;
  wire _33148_;
  wire _33149_;
  wire _33150_;
  wire _33151_;
  wire _33152_;
  wire _33153_;
  wire _33154_;
  wire _33155_;
  wire _33156_;
  wire _33157_;
  wire _33158_;
  wire _33159_;
  wire _33160_;
  wire _33161_;
  wire _33162_;
  wire _33163_;
  wire _33164_;
  wire _33165_;
  wire _33166_;
  wire _33167_;
  wire _33168_;
  wire _33169_;
  wire _33170_;
  wire _33171_;
  wire _33172_;
  wire _33173_;
  wire _33174_;
  wire _33175_;
  wire _33176_;
  wire _33177_;
  wire _33178_;
  wire _33179_;
  wire _33180_;
  wire _33181_;
  wire _33182_;
  wire _33183_;
  wire _33184_;
  wire _33185_;
  wire _33186_;
  wire _33187_;
  wire _33188_;
  wire _33189_;
  wire _33190_;
  wire _33191_;
  wire _33192_;
  wire _33193_;
  wire _33194_;
  wire _33195_;
  wire _33196_;
  wire _33197_;
  wire _33198_;
  wire _33199_;
  wire _33200_;
  wire _33201_;
  wire _33202_;
  wire _33203_;
  wire _33204_;
  wire _33205_;
  wire _33206_;
  wire _33207_;
  wire _33208_;
  wire _33209_;
  wire _33210_;
  wire _33211_;
  wire _33212_;
  wire _33213_;
  wire _33214_;
  wire _33215_;
  wire _33216_;
  wire _33217_;
  wire _33218_;
  wire _33219_;
  wire _33220_;
  wire _33221_;
  wire _33222_;
  wire _33223_;
  wire _33224_;
  wire _33225_;
  wire _33226_;
  wire _33227_;
  wire _33228_;
  wire _33229_;
  wire _33230_;
  wire _33231_;
  wire _33232_;
  wire _33233_;
  wire _33234_;
  wire _33235_;
  wire _33236_;
  wire _33237_;
  wire _33238_;
  wire _33239_;
  wire _33240_;
  wire _33241_;
  wire _33242_;
  wire _33243_;
  wire _33244_;
  wire _33245_;
  wire _33246_;
  wire _33247_;
  wire _33248_;
  wire _33249_;
  wire _33250_;
  wire _33251_;
  wire _33252_;
  wire _33253_;
  wire _33254_;
  wire _33255_;
  wire _33256_;
  wire _33257_;
  wire _33258_;
  wire _33259_;
  wire _33260_;
  wire _33261_;
  wire _33262_;
  wire _33263_;
  wire _33264_;
  wire _33265_;
  wire _33266_;
  wire _33267_;
  wire _33268_;
  wire _33269_;
  wire _33270_;
  wire _33271_;
  wire _33272_;
  wire _33273_;
  wire _33274_;
  wire _33275_;
  wire _33276_;
  wire _33277_;
  wire _33278_;
  wire _33279_;
  wire _33280_;
  wire _33281_;
  wire _33282_;
  wire _33283_;
  wire _33284_;
  wire _33285_;
  wire _33286_;
  wire _33287_;
  wire _33288_;
  wire _33289_;
  wire _33290_;
  wire _33291_;
  wire _33292_;
  wire _33293_;
  wire _33294_;
  wire _33295_;
  wire _33296_;
  wire _33297_;
  wire _33298_;
  wire _33299_;
  wire _33300_;
  wire _33301_;
  wire _33302_;
  wire _33303_;
  wire _33304_;
  wire _33305_;
  wire _33306_;
  wire _33307_;
  wire _33308_;
  wire _33309_;
  wire _33310_;
  wire _33311_;
  wire _33312_;
  wire _33313_;
  wire _33314_;
  wire _33315_;
  wire _33316_;
  wire _33317_;
  wire _33318_;
  wire _33319_;
  wire _33320_;
  wire _33321_;
  wire _33322_;
  wire _33323_;
  wire _33324_;
  wire _33325_;
  wire _33326_;
  wire _33327_;
  wire _33328_;
  wire _33329_;
  wire _33330_;
  wire _33331_;
  wire _33332_;
  wire _33333_;
  wire _33334_;
  wire _33335_;
  wire _33336_;
  wire _33337_;
  wire _33338_;
  wire _33339_;
  wire _33340_;
  wire _33341_;
  wire _33342_;
  wire _33343_;
  wire _33344_;
  wire _33345_;
  wire _33346_;
  wire _33347_;
  wire _33348_;
  wire _33349_;
  wire _33350_;
  wire _33351_;
  wire _33352_;
  wire _33353_;
  wire _33354_;
  wire _33355_;
  wire _33356_;
  wire _33357_;
  wire _33358_;
  wire _33359_;
  wire _33360_;
  wire _33361_;
  wire _33362_;
  wire _33363_;
  wire _33364_;
  wire _33365_;
  wire _33366_;
  wire _33367_;
  wire _33368_;
  wire _33369_;
  wire _33370_;
  wire _33371_;
  wire _33372_;
  wire _33373_;
  wire _33374_;
  wire _33375_;
  wire _33376_;
  wire _33377_;
  wire _33378_;
  wire _33379_;
  wire _33380_;
  wire _33381_;
  wire _33382_;
  wire _33383_;
  wire _33384_;
  wire _33385_;
  wire _33386_;
  wire _33387_;
  wire _33388_;
  wire _33389_;
  wire _33390_;
  wire _33391_;
  wire _33392_;
  wire _33393_;
  wire _33394_;
  wire _33395_;
  wire _33396_;
  wire _33397_;
  wire _33398_;
  wire _33399_;
  wire _33400_;
  wire _33401_;
  wire _33402_;
  wire _33403_;
  wire _33404_;
  wire _33405_;
  wire _33406_;
  wire _33407_;
  wire _33408_;
  wire _33409_;
  wire _33410_;
  wire _33411_;
  wire _33412_;
  wire _33413_;
  wire _33414_;
  wire _33415_;
  wire _33416_;
  wire _33417_;
  wire _33418_;
  wire _33419_;
  wire _33420_;
  wire _33421_;
  wire _33422_;
  wire _33423_;
  wire _33424_;
  wire _33425_;
  wire _33426_;
  wire _33427_;
  wire _33428_;
  wire _33429_;
  wire _33430_;
  wire _33431_;
  wire _33432_;
  wire _33433_;
  wire _33434_;
  wire _33435_;
  wire _33436_;
  wire _33437_;
  wire _33438_;
  wire _33439_;
  wire _33440_;
  wire _33441_;
  wire _33442_;
  wire _33443_;
  wire _33444_;
  wire _33445_;
  wire _33446_;
  wire _33447_;
  wire _33448_;
  wire _33449_;
  wire _33450_;
  wire _33451_;
  wire _33452_;
  wire _33453_;
  wire _33454_;
  wire _33455_;
  wire _33456_;
  wire _33457_;
  wire _33458_;
  wire _33459_;
  wire _33460_;
  wire _33461_;
  wire _33462_;
  wire _33463_;
  wire _33464_;
  wire _33465_;
  wire _33466_;
  wire _33467_;
  wire _33468_;
  wire _33469_;
  wire _33470_;
  wire _33471_;
  wire _33472_;
  wire _33473_;
  wire _33474_;
  wire _33475_;
  wire _33476_;
  wire _33477_;
  wire _33478_;
  wire _33479_;
  wire _33480_;
  wire _33481_;
  wire _33482_;
  wire _33483_;
  wire _33484_;
  wire _33485_;
  wire _33486_;
  wire _33487_;
  wire _33488_;
  wire _33489_;
  wire _33490_;
  wire _33491_;
  wire _33492_;
  wire _33493_;
  wire _33494_;
  wire _33495_;
  wire _33496_;
  wire _33497_;
  wire _33498_;
  wire _33499_;
  wire _33500_;
  wire _33501_;
  wire _33502_;
  wire _33503_;
  wire _33504_;
  wire _33505_;
  wire _33506_;
  wire _33507_;
  wire _33508_;
  wire _33509_;
  wire _33510_;
  wire _33511_;
  wire _33512_;
  wire _33513_;
  wire _33514_;
  wire _33515_;
  wire _33516_;
  wire _33517_;
  wire _33518_;
  wire _33519_;
  wire _33520_;
  wire _33521_;
  wire _33522_;
  wire _33523_;
  wire _33524_;
  wire _33525_;
  wire _33526_;
  wire _33527_;
  wire _33528_;
  wire _33529_;
  wire _33530_;
  wire _33531_;
  wire _33532_;
  wire _33533_;
  wire _33534_;
  wire _33535_;
  wire _33536_;
  wire _33537_;
  wire _33538_;
  wire _33539_;
  wire _33540_;
  wire _33541_;
  wire _33542_;
  wire _33543_;
  wire _33544_;
  wire _33545_;
  wire _33546_;
  wire _33547_;
  wire _33548_;
  wire _33549_;
  wire _33550_;
  wire _33551_;
  wire _33552_;
  wire _33553_;
  wire _33554_;
  wire _33555_;
  wire _33556_;
  wire _33557_;
  wire _33558_;
  wire _33559_;
  wire _33560_;
  wire _33561_;
  wire _33562_;
  wire _33563_;
  wire _33564_;
  wire _33565_;
  wire _33566_;
  wire _33567_;
  wire _33568_;
  wire _33569_;
  wire _33570_;
  wire _33571_;
  wire _33572_;
  wire _33573_;
  wire _33574_;
  wire _33575_;
  wire _33576_;
  wire _33577_;
  wire _33578_;
  wire _33579_;
  wire _33580_;
  wire _33581_;
  wire _33582_;
  wire _33583_;
  wire _33584_;
  wire _33585_;
  wire _33586_;
  wire _33587_;
  wire _33588_;
  wire _33589_;
  wire _33590_;
  wire _33591_;
  wire _33592_;
  wire _33593_;
  wire _33594_;
  wire _33595_;
  wire _33596_;
  wire _33597_;
  wire _33598_;
  wire _33599_;
  wire _33600_;
  wire _33601_;
  wire _33602_;
  wire _33603_;
  wire _33604_;
  wire _33605_;
  wire _33606_;
  wire _33607_;
  wire _33608_;
  wire _33609_;
  wire _33610_;
  wire _33611_;
  wire _33612_;
  wire _33613_;
  wire _33614_;
  wire _33615_;
  wire _33616_;
  wire _33617_;
  wire _33618_;
  wire _33619_;
  wire _33620_;
  wire _33621_;
  wire _33622_;
  wire _33623_;
  wire _33624_;
  wire _33625_;
  wire _33626_;
  wire _33627_;
  wire _33628_;
  wire _33629_;
  wire _33630_;
  wire _33631_;
  wire _33632_;
  wire _33633_;
  wire _33634_;
  wire _33635_;
  wire _33636_;
  wire _33637_;
  wire _33638_;
  wire _33639_;
  wire _33640_;
  wire _33641_;
  wire _33642_;
  wire _33643_;
  wire _33644_;
  wire _33645_;
  wire _33646_;
  wire _33647_;
  wire _33648_;
  wire _33649_;
  wire _33650_;
  wire _33651_;
  wire _33652_;
  wire _33653_;
  wire _33654_;
  wire _33655_;
  wire _33656_;
  wire _33657_;
  wire _33658_;
  wire _33659_;
  wire _33660_;
  wire _33661_;
  wire _33662_;
  wire _33663_;
  wire _33664_;
  wire _33665_;
  wire _33666_;
  wire _33667_;
  wire _33668_;
  wire _33669_;
  wire _33670_;
  wire _33671_;
  wire _33672_;
  wire _33673_;
  wire _33674_;
  wire _33675_;
  wire _33676_;
  wire _33677_;
  wire _33678_;
  wire _33679_;
  wire _33680_;
  wire _33681_;
  wire _33682_;
  wire _33683_;
  wire _33684_;
  wire _33685_;
  wire _33686_;
  wire _33687_;
  wire _33688_;
  wire _33689_;
  wire _33690_;
  wire _33691_;
  wire _33692_;
  wire _33693_;
  wire _33694_;
  wire _33695_;
  wire _33696_;
  wire _33697_;
  wire _33698_;
  wire _33699_;
  wire _33700_;
  wire _33701_;
  wire _33702_;
  wire _33703_;
  wire _33704_;
  wire _33705_;
  wire _33706_;
  wire _33707_;
  wire _33708_;
  wire _33709_;
  wire _33710_;
  wire _33711_;
  wire _33712_;
  wire _33713_;
  wire _33714_;
  wire _33715_;
  wire _33716_;
  wire _33717_;
  wire _33718_;
  wire _33719_;
  wire _33720_;
  wire _33721_;
  wire _33722_;
  wire _33723_;
  wire _33724_;
  wire _33725_;
  wire _33726_;
  wire _33727_;
  wire _33728_;
  wire _33729_;
  wire _33730_;
  wire _33731_;
  wire _33732_;
  wire _33733_;
  wire _33734_;
  wire _33735_;
  wire _33736_;
  wire _33737_;
  wire _33738_;
  wire _33739_;
  wire _33740_;
  wire _33741_;
  wire _33742_;
  wire _33743_;
  wire _33744_;
  wire _33745_;
  wire _33746_;
  wire _33747_;
  wire _33748_;
  wire _33749_;
  wire _33750_;
  wire _33751_;
  wire _33752_;
  wire _33753_;
  wire _33754_;
  wire _33755_;
  wire _33756_;
  wire _33757_;
  wire _33758_;
  wire _33759_;
  wire _33760_;
  wire _33761_;
  wire _33762_;
  wire _33763_;
  wire _33764_;
  wire _33765_;
  wire _33766_;
  wire _33767_;
  wire _33768_;
  wire _33769_;
  wire _33770_;
  wire _33771_;
  wire _33772_;
  wire _33773_;
  wire _33774_;
  wire _33775_;
  wire _33776_;
  wire _33777_;
  wire _33778_;
  wire _33779_;
  wire _33780_;
  wire _33781_;
  wire _33782_;
  wire _33783_;
  wire _33784_;
  wire _33785_;
  wire _33786_;
  wire _33787_;
  wire _33788_;
  wire _33789_;
  wire _33790_;
  wire _33791_;
  wire _33792_;
  wire _33793_;
  wire _33794_;
  wire _33795_;
  wire _33796_;
  wire _33797_;
  wire _33798_;
  wire _33799_;
  wire _33800_;
  wire _33801_;
  wire _33802_;
  wire _33803_;
  wire _33804_;
  wire _33805_;
  wire _33806_;
  wire _33807_;
  wire _33808_;
  wire _33809_;
  wire _33810_;
  wire _33811_;
  wire _33812_;
  wire _33813_;
  wire _33814_;
  wire _33815_;
  wire _33816_;
  wire _33817_;
  wire _33818_;
  wire _33819_;
  wire _33820_;
  wire _33821_;
  wire _33822_;
  wire _33823_;
  wire _33824_;
  wire _33825_;
  wire _33826_;
  wire _33827_;
  wire _33828_;
  wire _33829_;
  wire _33830_;
  wire _33831_;
  wire _33832_;
  wire _33833_;
  wire _33834_;
  wire _33835_;
  wire _33836_;
  wire _33837_;
  wire _33838_;
  wire _33839_;
  wire _33840_;
  wire _33841_;
  wire _33842_;
  wire _33843_;
  wire _33844_;
  wire _33845_;
  wire _33846_;
  wire _33847_;
  wire _33848_;
  wire _33849_;
  wire _33850_;
  wire _33851_;
  wire _33852_;
  wire _33853_;
  wire _33854_;
  wire _33855_;
  wire _33856_;
  wire _33857_;
  wire _33858_;
  wire _33859_;
  wire _33860_;
  wire _33861_;
  wire _33862_;
  wire _33863_;
  wire _33864_;
  wire _33865_;
  wire _33866_;
  wire _33867_;
  wire _33868_;
  wire _33869_;
  wire _33870_;
  wire _33871_;
  wire _33872_;
  wire _33873_;
  wire _33874_;
  wire _33875_;
  wire _33876_;
  wire _33877_;
  wire _33878_;
  wire _33879_;
  wire _33880_;
  wire _33881_;
  wire _33882_;
  wire _33883_;
  wire _33884_;
  wire _33885_;
  wire _33886_;
  wire _33887_;
  wire _33888_;
  wire _33889_;
  wire _33890_;
  wire _33891_;
  wire _33892_;
  wire _33893_;
  wire _33894_;
  wire _33895_;
  wire _33896_;
  wire _33897_;
  wire _33898_;
  wire _33899_;
  wire _33900_;
  wire _33901_;
  wire _33902_;
  wire _33903_;
  wire _33904_;
  wire _33905_;
  wire _33906_;
  wire _33907_;
  wire _33908_;
  wire _33909_;
  wire _33910_;
  wire _33911_;
  wire _33912_;
  wire _33913_;
  wire _33914_;
  wire _33915_;
  wire _33916_;
  wire _33917_;
  wire _33918_;
  wire _33919_;
  wire _33920_;
  wire _33921_;
  wire _33922_;
  wire _33923_;
  wire _33924_;
  wire _33925_;
  wire _33926_;
  wire _33927_;
  wire _33928_;
  wire _33929_;
  wire _33930_;
  wire _33931_;
  wire _33932_;
  wire _33933_;
  wire _33934_;
  wire _33935_;
  wire _33936_;
  wire _33937_;
  wire _33938_;
  wire _33939_;
  wire _33940_;
  wire _33941_;
  wire _33942_;
  wire _33943_;
  wire _33944_;
  wire _33945_;
  wire _33946_;
  wire _33947_;
  wire _33948_;
  wire _33949_;
  wire _33950_;
  wire _33951_;
  wire _33952_;
  wire _33953_;
  wire _33954_;
  wire _33955_;
  wire _33956_;
  wire _33957_;
  wire _33958_;
  wire _33959_;
  wire _33960_;
  wire _33961_;
  wire _33962_;
  wire _33963_;
  wire _33964_;
  wire _33965_;
  wire _33966_;
  wire _33967_;
  wire _33968_;
  wire _33969_;
  wire _33970_;
  wire _33971_;
  wire _33972_;
  wire _33973_;
  wire _33974_;
  wire _33975_;
  wire _33976_;
  wire _33977_;
  wire _33978_;
  wire _33979_;
  wire _33980_;
  wire _33981_;
  wire _33982_;
  wire _33983_;
  wire _33984_;
  wire _33985_;
  wire _33986_;
  wire _33987_;
  wire _33988_;
  wire _33989_;
  wire _33990_;
  wire _33991_;
  wire _33992_;
  wire _33993_;
  wire _33994_;
  wire _33995_;
  wire _33996_;
  wire _33997_;
  wire _33998_;
  wire _33999_;
  wire _34000_;
  wire _34001_;
  wire _34002_;
  wire _34003_;
  wire _34004_;
  wire _34005_;
  wire _34006_;
  wire _34007_;
  wire _34008_;
  wire _34009_;
  wire _34010_;
  wire _34011_;
  wire _34012_;
  wire _34013_;
  wire _34014_;
  wire _34015_;
  wire _34016_;
  wire _34017_;
  wire _34018_;
  wire _34019_;
  wire _34020_;
  wire _34021_;
  wire _34022_;
  wire _34023_;
  wire _34024_;
  wire _34025_;
  wire _34026_;
  wire _34027_;
  wire _34028_;
  wire _34029_;
  wire _34030_;
  wire _34031_;
  wire _34032_;
  wire _34033_;
  wire _34034_;
  wire _34035_;
  wire _34036_;
  wire _34037_;
  wire _34038_;
  wire _34039_;
  wire _34040_;
  wire _34041_;
  wire _34042_;
  wire _34043_;
  wire _34044_;
  wire _34045_;
  wire _34046_;
  wire _34047_;
  wire _34048_;
  wire _34049_;
  wire _34050_;
  wire _34051_;
  wire _34052_;
  wire _34053_;
  wire _34054_;
  wire _34055_;
  wire _34056_;
  wire _34057_;
  wire _34058_;
  wire _34059_;
  wire _34060_;
  wire _34061_;
  wire _34062_;
  wire _34063_;
  wire _34064_;
  wire _34065_;
  wire _34066_;
  wire _34067_;
  wire _34068_;
  wire _34069_;
  wire _34070_;
  wire _34071_;
  wire _34072_;
  wire _34073_;
  wire _34074_;
  wire _34075_;
  wire _34076_;
  wire _34077_;
  wire _34078_;
  wire _34079_;
  wire _34080_;
  wire _34081_;
  wire _34082_;
  wire _34083_;
  wire _34084_;
  wire _34085_;
  wire _34086_;
  wire _34087_;
  wire _34088_;
  wire _34089_;
  wire _34090_;
  wire _34091_;
  wire _34092_;
  wire _34093_;
  wire _34094_;
  wire _34095_;
  wire _34096_;
  wire _34097_;
  wire _34098_;
  wire _34099_;
  wire _34100_;
  wire _34101_;
  wire _34102_;
  wire _34103_;
  wire _34104_;
  wire _34105_;
  wire _34106_;
  wire _34107_;
  wire _34108_;
  wire _34109_;
  wire _34110_;
  wire _34111_;
  wire _34112_;
  wire _34113_;
  wire _34114_;
  wire _34115_;
  wire _34116_;
  wire _34117_;
  wire _34118_;
  wire _34119_;
  wire _34120_;
  wire _34121_;
  wire _34122_;
  wire _34123_;
  wire _34124_;
  wire _34125_;
  wire _34126_;
  wire _34127_;
  wire _34128_;
  wire _34129_;
  wire _34130_;
  wire _34131_;
  wire _34132_;
  wire _34133_;
  wire _34134_;
  wire _34135_;
  wire _34136_;
  wire _34137_;
  wire _34138_;
  wire _34139_;
  wire _34140_;
  wire _34141_;
  wire _34142_;
  wire _34143_;
  wire _34144_;
  wire _34145_;
  wire _34146_;
  wire _34147_;
  wire _34148_;
  wire _34149_;
  wire _34150_;
  wire _34151_;
  wire _34152_;
  wire _34153_;
  wire _34154_;
  wire _34155_;
  wire _34156_;
  wire _34157_;
  wire _34158_;
  wire _34159_;
  wire _34160_;
  wire _34161_;
  wire _34162_;
  wire _34163_;
  wire _34164_;
  wire _34165_;
  wire _34166_;
  wire _34167_;
  wire _34168_;
  wire _34169_;
  wire _34170_;
  wire _34171_;
  wire _34172_;
  wire _34173_;
  wire _34174_;
  wire _34175_;
  wire _34176_;
  wire _34177_;
  wire _34178_;
  wire _34179_;
  wire _34180_;
  wire _34181_;
  wire _34182_;
  wire _34183_;
  wire _34184_;
  wire _34185_;
  wire _34186_;
  wire _34187_;
  wire _34188_;
  wire _34189_;
  wire _34190_;
  wire _34191_;
  wire _34192_;
  wire _34193_;
  wire _34194_;
  wire _34195_;
  wire _34196_;
  wire _34197_;
  wire _34198_;
  wire _34199_;
  wire _34200_;
  wire _34201_;
  wire _34202_;
  wire _34203_;
  wire _34204_;
  wire _34205_;
  wire _34206_;
  wire _34207_;
  wire _34208_;
  wire _34209_;
  wire _34210_;
  wire _34211_;
  wire _34212_;
  wire _34213_;
  wire _34214_;
  wire _34215_;
  wire _34216_;
  wire _34217_;
  wire _34218_;
  wire _34219_;
  wire _34220_;
  wire _34221_;
  wire _34222_;
  wire _34223_;
  wire _34224_;
  wire _34225_;
  wire _34226_;
  wire _34227_;
  wire _34228_;
  wire _34229_;
  wire _34230_;
  wire _34231_;
  wire _34232_;
  wire _34233_;
  wire _34234_;
  wire _34235_;
  wire _34236_;
  wire _34237_;
  wire _34238_;
  wire _34239_;
  wire _34240_;
  wire _34241_;
  wire _34242_;
  wire _34243_;
  wire _34244_;
  wire _34245_;
  wire _34246_;
  wire _34247_;
  wire _34248_;
  wire _34249_;
  wire _34250_;
  wire _34251_;
  wire _34252_;
  wire _34253_;
  wire _34254_;
  wire _34255_;
  wire _34256_;
  wire _34257_;
  wire _34258_;
  wire _34259_;
  wire _34260_;
  wire _34261_;
  wire _34262_;
  wire _34263_;
  wire _34264_;
  wire _34265_;
  wire _34266_;
  wire _34267_;
  wire _34268_;
  wire _34269_;
  wire _34270_;
  wire _34271_;
  wire _34272_;
  wire _34273_;
  wire _34274_;
  wire _34275_;
  wire _34276_;
  wire _34277_;
  wire _34278_;
  wire _34279_;
  wire _34280_;
  wire _34281_;
  wire _34282_;
  wire _34283_;
  wire _34284_;
  wire _34285_;
  wire _34286_;
  wire _34287_;
  wire _34288_;
  wire _34289_;
  wire _34290_;
  wire _34291_;
  wire _34292_;
  wire _34293_;
  wire _34294_;
  wire _34295_;
  wire _34296_;
  wire _34297_;
  wire _34298_;
  wire _34299_;
  wire _34300_;
  wire _34301_;
  wire _34302_;
  wire _34303_;
  wire _34304_;
  wire _34305_;
  wire _34306_;
  wire _34307_;
  wire _34308_;
  wire _34309_;
  wire _34310_;
  wire _34311_;
  wire _34312_;
  wire _34313_;
  wire _34314_;
  wire _34315_;
  wire _34316_;
  wire _34317_;
  wire _34318_;
  wire _34319_;
  wire _34320_;
  wire _34321_;
  wire _34322_;
  wire _34323_;
  wire _34324_;
  wire _34325_;
  wire _34326_;
  wire _34327_;
  wire _34328_;
  wire _34329_;
  wire _34330_;
  wire _34331_;
  wire _34332_;
  wire _34333_;
  wire _34334_;
  wire _34335_;
  wire _34336_;
  wire _34337_;
  wire _34338_;
  wire _34339_;
  wire _34340_;
  wire _34341_;
  wire _34342_;
  wire _34343_;
  wire _34344_;
  wire _34345_;
  wire _34346_;
  wire _34347_;
  wire _34348_;
  wire _34349_;
  wire _34350_;
  wire _34351_;
  wire _34352_;
  wire _34353_;
  wire _34354_;
  wire _34355_;
  wire _34356_;
  wire _34357_;
  wire _34358_;
  wire _34359_;
  wire _34360_;
  wire _34361_;
  wire _34362_;
  wire _34363_;
  wire _34364_;
  wire _34365_;
  wire _34366_;
  wire _34367_;
  wire _34368_;
  wire _34369_;
  wire _34370_;
  wire _34371_;
  wire _34372_;
  wire _34373_;
  wire _34374_;
  wire _34375_;
  wire _34376_;
  wire _34377_;
  wire _34378_;
  wire _34379_;
  wire _34380_;
  wire _34381_;
  wire _34382_;
  wire _34383_;
  wire _34384_;
  wire _34385_;
  wire _34386_;
  wire _34387_;
  wire _34388_;
  wire _34389_;
  wire _34390_;
  wire _34391_;
  wire _34392_;
  wire _34393_;
  wire _34394_;
  wire _34395_;
  wire _34396_;
  wire _34397_;
  wire _34398_;
  wire _34399_;
  wire _34400_;
  wire _34401_;
  wire _34402_;
  wire _34403_;
  wire _34404_;
  wire _34405_;
  wire _34406_;
  wire _34407_;
  wire _34408_;
  wire _34409_;
  wire _34410_;
  wire _34411_;
  wire _34412_;
  wire _34413_;
  wire _34414_;
  wire _34415_;
  wire _34416_;
  wire _34417_;
  wire _34418_;
  wire _34419_;
  wire _34420_;
  wire _34421_;
  wire _34422_;
  wire _34423_;
  wire _34424_;
  wire _34425_;
  wire _34426_;
  wire _34427_;
  wire _34428_;
  wire _34429_;
  wire _34430_;
  wire _34431_;
  wire _34432_;
  wire _34433_;
  wire _34434_;
  wire _34435_;
  wire _34436_;
  wire _34437_;
  wire _34438_;
  wire _34439_;
  wire _34440_;
  wire _34441_;
  wire _34442_;
  wire _34443_;
  wire _34444_;
  wire _34445_;
  wire _34446_;
  wire _34447_;
  wire _34448_;
  wire _34449_;
  wire _34450_;
  wire _34451_;
  wire _34452_;
  wire _34453_;
  wire _34454_;
  wire _34455_;
  wire _34456_;
  wire _34457_;
  wire _34458_;
  wire _34459_;
  wire _34460_;
  wire _34461_;
  wire _34462_;
  wire _34463_;
  wire _34464_;
  wire _34465_;
  wire _34466_;
  wire _34467_;
  wire _34468_;
  wire _34469_;
  wire _34470_;
  wire _34471_;
  wire _34472_;
  wire _34473_;
  wire _34474_;
  wire _34475_;
  wire _34476_;
  wire _34477_;
  wire _34478_;
  wire _34479_;
  wire _34480_;
  wire _34481_;
  wire _34482_;
  wire _34483_;
  wire _34484_;
  wire _34485_;
  wire _34486_;
  wire _34487_;
  wire _34488_;
  wire _34489_;
  wire _34490_;
  wire _34491_;
  wire _34492_;
  wire _34493_;
  wire _34494_;
  wire _34495_;
  wire _34496_;
  wire _34497_;
  wire _34498_;
  wire _34499_;
  wire _34500_;
  wire _34501_;
  wire _34502_;
  wire _34503_;
  wire _34504_;
  wire _34505_;
  wire _34506_;
  wire _34507_;
  wire _34508_;
  wire _34509_;
  wire _34510_;
  wire _34511_;
  wire _34512_;
  wire _34513_;
  wire _34514_;
  wire _34515_;
  wire _34516_;
  wire _34517_;
  wire _34518_;
  wire _34519_;
  wire _34520_;
  wire _34521_;
  wire _34522_;
  wire _34523_;
  wire _34524_;
  wire _34525_;
  wire _34526_;
  wire _34527_;
  wire _34528_;
  wire _34529_;
  wire _34530_;
  wire _34531_;
  wire _34532_;
  wire _34533_;
  wire _34534_;
  wire _34535_;
  wire _34536_;
  wire _34537_;
  wire _34538_;
  wire _34539_;
  wire _34540_;
  wire _34541_;
  wire _34542_;
  wire _34543_;
  wire _34544_;
  wire _34545_;
  wire _34546_;
  wire _34547_;
  wire _34548_;
  wire _34549_;
  wire _34550_;
  wire _34551_;
  wire _34552_;
  wire _34553_;
  wire _34554_;
  wire _34555_;
  wire _34556_;
  wire _34557_;
  wire _34558_;
  wire _34559_;
  wire _34560_;
  wire _34561_;
  wire _34562_;
  wire _34563_;
  wire _34564_;
  wire _34565_;
  wire _34566_;
  wire _34567_;
  wire _34568_;
  wire _34569_;
  wire _34570_;
  wire _34571_;
  wire _34572_;
  wire _34573_;
  wire _34574_;
  wire _34575_;
  wire _34576_;
  wire _34577_;
  wire _34578_;
  wire _34579_;
  wire _34580_;
  wire _34581_;
  wire _34582_;
  wire _34583_;
  wire _34584_;
  wire _34585_;
  wire _34586_;
  wire _34587_;
  wire _34588_;
  wire _34589_;
  wire _34590_;
  wire _34591_;
  wire _34592_;
  wire _34593_;
  wire _34594_;
  wire _34595_;
  wire _34596_;
  wire _34597_;
  wire _34598_;
  wire _34599_;
  wire _34600_;
  wire _34601_;
  wire _34602_;
  wire _34603_;
  wire _34604_;
  wire _34605_;
  wire _34606_;
  wire _34607_;
  wire _34608_;
  wire _34609_;
  wire _34610_;
  wire _34611_;
  wire _34612_;
  wire _34613_;
  wire _34614_;
  wire _34615_;
  wire _34616_;
  wire _34617_;
  wire _34618_;
  wire _34619_;
  wire _34620_;
  wire _34621_;
  wire _34622_;
  wire _34623_;
  wire _34624_;
  wire _34625_;
  wire _34626_;
  wire _34627_;
  wire _34628_;
  wire _34629_;
  wire _34630_;
  wire _34631_;
  wire _34632_;
  wire _34633_;
  wire _34634_;
  wire _34635_;
  wire _34636_;
  wire _34637_;
  wire _34638_;
  wire _34639_;
  wire _34640_;
  wire _34641_;
  wire _34642_;
  wire _34643_;
  wire _34644_;
  wire _34645_;
  wire _34646_;
  wire _34647_;
  wire _34648_;
  wire _34649_;
  wire _34650_;
  wire _34651_;
  wire _34652_;
  wire _34653_;
  wire _34654_;
  wire _34655_;
  wire _34656_;
  wire _34657_;
  wire _34658_;
  wire _34659_;
  wire _34660_;
  wire _34661_;
  wire _34662_;
  wire _34663_;
  wire _34664_;
  wire _34665_;
  wire _34666_;
  wire _34667_;
  wire _34668_;
  wire _34669_;
  wire _34670_;
  wire _34671_;
  wire _34672_;
  wire _34673_;
  wire _34674_;
  wire _34675_;
  wire _34676_;
  wire _34677_;
  wire _34678_;
  wire _34679_;
  wire _34680_;
  wire _34681_;
  wire _34682_;
  wire _34683_;
  wire _34684_;
  wire _34685_;
  wire _34686_;
  wire _34687_;
  wire _34688_;
  wire _34689_;
  wire _34690_;
  wire _34691_;
  wire _34692_;
  wire _34693_;
  wire _34694_;
  wire _34695_;
  wire _34696_;
  wire _34697_;
  wire _34698_;
  wire _34699_;
  wire _34700_;
  wire _34701_;
  wire _34702_;
  wire _34703_;
  wire _34704_;
  wire _34705_;
  wire _34706_;
  wire _34707_;
  wire _34708_;
  wire _34709_;
  wire _34710_;
  wire _34711_;
  wire _34712_;
  wire _34713_;
  wire _34714_;
  wire _34715_;
  wire _34716_;
  wire _34717_;
  wire _34718_;
  wire _34719_;
  wire _34720_;
  wire _34721_;
  wire _34722_;
  wire _34723_;
  wire _34724_;
  wire _34725_;
  wire _34726_;
  wire _34727_;
  wire _34728_;
  wire _34729_;
  wire _34730_;
  wire _34731_;
  wire _34732_;
  wire _34733_;
  wire _34734_;
  wire _34735_;
  wire _34736_;
  wire _34737_;
  wire _34738_;
  wire _34739_;
  wire _34740_;
  wire _34741_;
  wire _34742_;
  wire _34743_;
  wire _34744_;
  wire _34745_;
  wire _34746_;
  wire _34747_;
  wire _34748_;
  wire _34749_;
  wire _34750_;
  wire _34751_;
  wire _34752_;
  wire _34753_;
  wire _34754_;
  wire _34755_;
  wire _34756_;
  wire _34757_;
  wire _34758_;
  wire _34759_;
  wire _34760_;
  wire _34761_;
  wire _34762_;
  wire _34763_;
  wire _34764_;
  wire _34765_;
  wire _34766_;
  wire _34767_;
  wire _34768_;
  wire _34769_;
  wire _34770_;
  wire _34771_;
  wire _34772_;
  wire _34773_;
  wire _34774_;
  wire _34775_;
  wire _34776_;
  wire _34777_;
  wire _34778_;
  wire _34779_;
  wire _34780_;
  wire _34781_;
  wire _34782_;
  wire _34783_;
  wire _34784_;
  wire _34785_;
  wire _34786_;
  wire _34787_;
  wire _34788_;
  wire _34789_;
  wire _34790_;
  wire _34791_;
  wire _34792_;
  wire _34793_;
  wire _34794_;
  wire _34795_;
  wire _34796_;
  wire _34797_;
  wire _34798_;
  wire _34799_;
  wire _34800_;
  wire _34801_;
  wire _34802_;
  wire _34803_;
  wire _34804_;
  wire _34805_;
  wire _34806_;
  wire _34807_;
  wire _34808_;
  wire _34809_;
  wire _34810_;
  wire _34811_;
  wire _34812_;
  wire _34813_;
  wire _34814_;
  wire _34815_;
  wire _34816_;
  wire _34817_;
  wire _34818_;
  wire _34819_;
  wire _34820_;
  wire _34821_;
  wire _34822_;
  wire _34823_;
  wire _34824_;
  wire _34825_;
  wire _34826_;
  wire _34827_;
  wire _34828_;
  wire _34829_;
  wire _34830_;
  wire _34831_;
  wire _34832_;
  wire _34833_;
  wire _34834_;
  wire _34835_;
  wire _34836_;
  wire _34837_;
  wire _34838_;
  wire _34839_;
  wire _34840_;
  wire _34841_;
  wire _34842_;
  wire _34843_;
  wire _34844_;
  wire _34845_;
  wire _34846_;
  wire _34847_;
  wire _34848_;
  wire _34849_;
  wire _34850_;
  wire _34851_;
  wire _34852_;
  wire _34853_;
  wire _34854_;
  wire _34855_;
  wire _34856_;
  wire _34857_;
  wire _34858_;
  wire _34859_;
  wire _34860_;
  wire _34861_;
  wire _34862_;
  wire _34863_;
  wire _34864_;
  wire _34865_;
  wire _34866_;
  wire _34867_;
  wire _34868_;
  wire _34869_;
  wire _34870_;
  wire _34871_;
  wire _34872_;
  wire _34873_;
  wire _34874_;
  wire _34875_;
  wire _34876_;
  wire _34877_;
  wire _34878_;
  wire _34879_;
  wire _34880_;
  wire _34881_;
  wire _34882_;
  wire _34883_;
  wire _34884_;
  wire _34885_;
  wire _34886_;
  wire _34887_;
  wire _34888_;
  wire _34889_;
  wire _34890_;
  wire _34891_;
  wire _34892_;
  wire _34893_;
  wire _34894_;
  wire _34895_;
  wire _34896_;
  wire _34897_;
  wire _34898_;
  wire _34899_;
  wire _34900_;
  wire _34901_;
  wire _34902_;
  wire _34903_;
  wire _34904_;
  wire _34905_;
  wire _34906_;
  wire _34907_;
  wire _34908_;
  wire _34909_;
  wire _34910_;
  wire _34911_;
  wire _34912_;
  wire _34913_;
  wire _34914_;
  wire _34915_;
  wire _34916_;
  wire _34917_;
  wire _34918_;
  wire _34919_;
  wire _34920_;
  wire _34921_;
  wire _34922_;
  wire _34923_;
  wire _34924_;
  wire _34925_;
  wire _34926_;
  wire _34927_;
  wire _34928_;
  wire _34929_;
  wire _34930_;
  wire _34931_;
  wire _34932_;
  wire _34933_;
  wire _34934_;
  wire _34935_;
  wire _34936_;
  wire _34937_;
  wire _34938_;
  wire _34939_;
  wire _34940_;
  wire _34941_;
  wire _34942_;
  wire _34943_;
  wire _34944_;
  wire _34945_;
  wire _34946_;
  wire _34947_;
  wire _34948_;
  wire _34949_;
  wire _34950_;
  wire _34951_;
  wire _34952_;
  wire _34953_;
  wire _34954_;
  wire _34955_;
  wire _34956_;
  wire _34957_;
  wire _34958_;
  wire _34959_;
  wire _34960_;
  wire _34961_;
  wire _34962_;
  wire _34963_;
  wire _34964_;
  wire _34965_;
  wire _34966_;
  wire _34967_;
  wire _34968_;
  wire _34969_;
  wire _34970_;
  wire _34971_;
  wire _34972_;
  wire _34973_;
  wire _34974_;
  wire _34975_;
  wire _34976_;
  wire _34977_;
  wire _34978_;
  wire _34979_;
  wire _34980_;
  wire _34981_;
  wire _34982_;
  wire _34983_;
  wire _34984_;
  wire _34985_;
  wire _34986_;
  wire _34987_;
  wire _34988_;
  wire _34989_;
  wire _34990_;
  wire _34991_;
  wire _34992_;
  wire _34993_;
  wire _34994_;
  wire _34995_;
  wire _34996_;
  wire _34997_;
  wire _34998_;
  wire _34999_;
  wire _35000_;
  wire _35001_;
  wire _35002_;
  wire _35003_;
  wire _35004_;
  wire _35005_;
  wire _35006_;
  wire _35007_;
  wire _35008_;
  wire _35009_;
  wire _35010_;
  wire _35011_;
  wire _35012_;
  wire _35013_;
  wire _35014_;
  wire _35015_;
  wire _35016_;
  wire _35017_;
  wire _35018_;
  wire _35019_;
  wire _35020_;
  wire _35021_;
  wire _35022_;
  wire _35023_;
  wire _35024_;
  wire _35025_;
  wire _35026_;
  wire _35027_;
  wire _35028_;
  wire _35029_;
  wire _35030_;
  wire _35031_;
  wire _35032_;
  wire _35033_;
  wire _35034_;
  wire _35035_;
  wire _35036_;
  wire _35037_;
  wire _35038_;
  wire _35039_;
  wire _35040_;
  wire _35041_;
  wire _35042_;
  wire _35043_;
  wire _35044_;
  wire _35045_;
  wire _35046_;
  wire _35047_;
  wire _35048_;
  wire _35049_;
  wire _35050_;
  wire _35051_;
  wire _35052_;
  wire _35053_;
  wire _35054_;
  wire _35055_;
  wire _35056_;
  wire _35057_;
  wire _35058_;
  wire _35059_;
  wire _35060_;
  wire _35061_;
  wire _35062_;
  wire _35063_;
  wire _35064_;
  wire _35065_;
  wire _35066_;
  wire _35067_;
  wire _35068_;
  wire _35069_;
  wire _35070_;
  wire _35071_;
  wire _35072_;
  wire _35073_;
  wire _35074_;
  wire _35075_;
  wire _35076_;
  wire _35077_;
  wire _35078_;
  wire _35079_;
  wire _35080_;
  wire _35081_;
  wire _35082_;
  wire _35083_;
  wire _35084_;
  wire _35085_;
  wire _35086_;
  wire _35087_;
  wire _35088_;
  wire _35089_;
  wire _35090_;
  wire _35091_;
  wire _35092_;
  wire _35093_;
  wire _35094_;
  wire _35095_;
  wire _35096_;
  wire _35097_;
  wire _35098_;
  wire _35099_;
  wire _35100_;
  wire _35101_;
  wire _35102_;
  wire _35103_;
  wire _35104_;
  wire _35105_;
  wire _35106_;
  wire _35107_;
  wire _35108_;
  wire _35109_;
  wire _35110_;
  wire _35111_;
  wire _35112_;
  wire _35113_;
  wire _35114_;
  wire _35115_;
  wire _35116_;
  wire _35117_;
  wire _35118_;
  wire _35119_;
  wire _35120_;
  wire _35121_;
  wire _35122_;
  wire _35123_;
  wire _35124_;
  wire _35125_;
  wire _35126_;
  wire _35127_;
  wire _35128_;
  wire _35129_;
  wire _35130_;
  wire _35131_;
  wire _35132_;
  wire _35133_;
  wire _35134_;
  wire _35135_;
  wire _35136_;
  wire _35137_;
  wire _35138_;
  wire _35139_;
  wire _35140_;
  wire _35141_;
  wire _35142_;
  wire _35143_;
  wire _35144_;
  wire _35145_;
  wire _35146_;
  wire _35147_;
  wire _35148_;
  wire _35149_;
  wire _35150_;
  wire _35151_;
  wire _35152_;
  wire _35153_;
  wire _35154_;
  wire _35155_;
  wire _35156_;
  wire _35157_;
  wire _35158_;
  wire _35159_;
  wire _35160_;
  wire _35161_;
  wire _35162_;
  wire _35163_;
  wire _35164_;
  wire _35165_;
  wire _35166_;
  wire _35167_;
  wire _35168_;
  wire _35169_;
  wire _35170_;
  wire _35171_;
  wire _35172_;
  wire _35173_;
  wire _35174_;
  wire _35175_;
  wire _35176_;
  wire _35177_;
  wire _35178_;
  wire _35179_;
  wire _35180_;
  wire _35181_;
  wire _35182_;
  wire _35183_;
  wire _35184_;
  wire _35185_;
  wire _35186_;
  wire _35187_;
  wire _35188_;
  wire _35189_;
  wire _35190_;
  wire _35191_;
  wire _35192_;
  wire _35193_;
  wire _35194_;
  wire _35195_;
  wire _35196_;
  wire _35197_;
  wire _35198_;
  wire _35199_;
  wire _35200_;
  wire _35201_;
  wire _35202_;
  wire _35203_;
  wire _35204_;
  wire _35205_;
  wire _35206_;
  wire _35207_;
  wire _35208_;
  wire _35209_;
  wire _35210_;
  wire _35211_;
  wire _35212_;
  wire _35213_;
  wire _35214_;
  wire _35215_;
  wire _35216_;
  wire _35217_;
  wire _35218_;
  wire _35219_;
  wire _35220_;
  wire _35221_;
  wire _35222_;
  wire _35223_;
  wire _35224_;
  wire _35225_;
  wire _35226_;
  wire _35227_;
  wire _35228_;
  wire _35229_;
  wire _35230_;
  wire _35231_;
  wire _35232_;
  wire _35233_;
  wire _35234_;
  wire _35235_;
  wire _35236_;
  wire _35237_;
  wire _35238_;
  wire _35239_;
  wire _35240_;
  wire _35241_;
  wire _35242_;
  wire _35243_;
  wire _35244_;
  wire _35245_;
  wire _35246_;
  wire _35247_;
  wire _35248_;
  wire _35249_;
  wire _35250_;
  wire _35251_;
  wire _35252_;
  wire _35253_;
  wire _35254_;
  wire _35255_;
  wire _35256_;
  wire _35257_;
  wire _35258_;
  wire _35259_;
  wire _35260_;
  wire _35261_;
  wire _35262_;
  wire _35263_;
  wire _35264_;
  wire _35265_;
  wire _35266_;
  wire _35267_;
  wire _35268_;
  wire _35269_;
  wire _35270_;
  wire _35271_;
  wire _35272_;
  wire _35273_;
  wire _35274_;
  wire _35275_;
  wire _35276_;
  wire _35277_;
  wire _35278_;
  wire _35279_;
  wire _35280_;
  wire _35281_;
  wire _35282_;
  wire _35283_;
  wire _35284_;
  wire _35285_;
  wire _35286_;
  wire _35287_;
  wire _35288_;
  wire _35289_;
  wire _35290_;
  wire _35291_;
  wire _35292_;
  wire _35293_;
  wire _35294_;
  wire _35295_;
  wire _35296_;
  wire _35297_;
  wire _35298_;
  wire _35299_;
  wire _35300_;
  wire _35301_;
  wire _35302_;
  wire _35303_;
  wire _35304_;
  wire _35305_;
  wire _35306_;
  wire _35307_;
  wire _35308_;
  wire _35309_;
  wire _35310_;
  wire _35311_;
  wire _35312_;
  wire _35313_;
  wire _35314_;
  wire _35315_;
  wire _35316_;
  wire _35317_;
  wire _35318_;
  wire _35319_;
  wire _35320_;
  wire _35321_;
  wire _35322_;
  wire _35323_;
  wire _35324_;
  wire _35325_;
  wire _35326_;
  wire _35327_;
  wire _35328_;
  wire _35329_;
  wire _35330_;
  wire _35331_;
  wire _35332_;
  wire _35333_;
  wire _35334_;
  wire _35335_;
  wire _35336_;
  wire _35337_;
  wire _35338_;
  wire _35339_;
  wire _35340_;
  wire _35341_;
  wire _35342_;
  wire _35343_;
  wire _35344_;
  wire _35345_;
  wire _35346_;
  wire _35347_;
  wire _35348_;
  wire _35349_;
  wire _35350_;
  wire _35351_;
  wire _35352_;
  wire _35353_;
  wire _35354_;
  wire _35355_;
  wire _35356_;
  wire _35357_;
  wire _35358_;
  wire _35359_;
  wire _35360_;
  wire _35361_;
  wire _35362_;
  wire _35363_;
  wire _35364_;
  wire _35365_;
  wire _35366_;
  wire _35367_;
  wire _35368_;
  wire _35369_;
  wire _35370_;
  wire _35371_;
  wire _35372_;
  wire _35373_;
  wire _35374_;
  wire _35375_;
  wire _35376_;
  wire _35377_;
  wire _35378_;
  wire _35379_;
  wire _35380_;
  wire _35381_;
  wire _35382_;
  wire _35383_;
  wire _35384_;
  wire _35385_;
  wire _35386_;
  wire _35387_;
  wire _35388_;
  wire _35389_;
  wire _35390_;
  wire _35391_;
  wire _35392_;
  wire _35393_;
  wire _35394_;
  wire _35395_;
  wire _35396_;
  wire _35397_;
  wire _35398_;
  wire _35399_;
  wire _35400_;
  wire _35401_;
  wire _35402_;
  wire _35403_;
  wire _35404_;
  wire _35405_;
  wire _35406_;
  wire _35407_;
  wire _35408_;
  wire _35409_;
  wire _35410_;
  wire _35411_;
  wire _35412_;
  wire _35413_;
  wire _35414_;
  wire _35415_;
  wire _35416_;
  wire _35417_;
  wire _35418_;
  wire _35419_;
  wire _35420_;
  wire _35421_;
  wire _35422_;
  wire _35423_;
  wire _35424_;
  wire _35425_;
  wire _35426_;
  wire _35427_;
  wire _35428_;
  wire _35429_;
  wire _35430_;
  wire _35431_;
  wire _35432_;
  wire _35433_;
  wire _35434_;
  wire _35435_;
  wire _35436_;
  wire _35437_;
  wire _35438_;
  wire _35439_;
  wire _35440_;
  wire _35441_;
  wire _35442_;
  wire _35443_;
  wire _35444_;
  wire _35445_;
  wire _35446_;
  wire _35447_;
  wire _35448_;
  wire _35449_;
  wire _35450_;
  wire _35451_;
  wire _35452_;
  wire _35453_;
  wire _35454_;
  wire _35455_;
  wire _35456_;
  wire _35457_;
  wire _35458_;
  wire _35459_;
  wire _35460_;
  wire _35461_;
  wire _35462_;
  wire _35463_;
  wire _35464_;
  wire _35465_;
  wire _35466_;
  wire _35467_;
  wire _35468_;
  wire _35469_;
  wire _35470_;
  wire _35471_;
  wire _35472_;
  wire _35473_;
  wire _35474_;
  wire _35475_;
  wire _35476_;
  wire _35477_;
  wire _35478_;
  wire _35479_;
  wire _35480_;
  wire _35481_;
  wire _35482_;
  wire _35483_;
  wire _35484_;
  wire _35485_;
  wire _35486_;
  wire _35487_;
  wire _35488_;
  wire _35489_;
  wire _35490_;
  wire _35491_;
  wire _35492_;
  wire _35493_;
  wire _35494_;
  wire _35495_;
  wire _35496_;
  wire _35497_;
  wire _35498_;
  wire _35499_;
  wire _35500_;
  wire _35501_;
  wire _35502_;
  wire _35503_;
  wire _35504_;
  wire _35505_;
  wire _35506_;
  wire _35507_;
  wire _35508_;
  wire _35509_;
  wire _35510_;
  wire _35511_;
  wire _35512_;
  wire _35513_;
  wire _35514_;
  wire _35515_;
  wire _35516_;
  wire _35517_;
  wire _35518_;
  wire _35519_;
  wire _35520_;
  wire _35521_;
  wire _35522_;
  wire _35523_;
  wire _35524_;
  wire _35525_;
  wire _35526_;
  wire _35527_;
  wire _35528_;
  wire _35529_;
  wire _35530_;
  wire _35531_;
  wire _35532_;
  wire _35533_;
  wire _35534_;
  wire _35535_;
  wire _35536_;
  wire _35537_;
  wire _35538_;
  wire _35539_;
  wire _35540_;
  wire _35541_;
  wire _35542_;
  wire _35543_;
  wire _35544_;
  wire _35545_;
  wire _35546_;
  wire _35547_;
  wire _35548_;
  wire _35549_;
  wire _35550_;
  wire _35551_;
  wire _35552_;
  wire _35553_;
  wire _35554_;
  wire _35555_;
  wire _35556_;
  wire _35557_;
  wire _35558_;
  wire _35559_;
  wire _35560_;
  wire _35561_;
  wire _35562_;
  wire _35563_;
  wire _35564_;
  wire _35565_;
  wire _35566_;
  wire _35567_;
  wire _35568_;
  wire _35569_;
  wire _35570_;
  wire _35571_;
  wire _35572_;
  wire _35573_;
  wire _35574_;
  wire _35575_;
  wire _35576_;
  wire _35577_;
  wire _35578_;
  wire _35579_;
  wire _35580_;
  wire _35581_;
  wire _35582_;
  wire _35583_;
  wire _35584_;
  wire _35585_;
  wire _35586_;
  wire _35587_;
  wire _35588_;
  wire _35589_;
  wire _35590_;
  wire _35591_;
  wire _35592_;
  wire _35593_;
  wire _35594_;
  wire _35595_;
  wire _35596_;
  wire _35597_;
  wire _35598_;
  wire _35599_;
  wire _35600_;
  wire _35601_;
  wire _35602_;
  wire _35603_;
  wire _35604_;
  wire _35605_;
  wire _35606_;
  wire _35607_;
  wire _35608_;
  wire _35609_;
  wire _35610_;
  wire _35611_;
  wire _35612_;
  wire _35613_;
  wire _35614_;
  wire _35615_;
  wire _35616_;
  wire _35617_;
  wire _35618_;
  wire _35619_;
  wire _35620_;
  wire _35621_;
  wire _35622_;
  wire _35623_;
  wire _35624_;
  wire _35625_;
  wire _35626_;
  wire _35627_;
  wire _35628_;
  wire _35629_;
  wire _35630_;
  wire _35631_;
  wire _35632_;
  wire _35633_;
  wire _35634_;
  wire _35635_;
  wire _35636_;
  wire _35637_;
  wire _35638_;
  wire _35639_;
  wire _35640_;
  wire _35641_;
  wire _35642_;
  wire _35643_;
  wire _35644_;
  wire _35645_;
  wire _35646_;
  wire _35647_;
  wire _35648_;
  wire _35649_;
  wire _35650_;
  wire _35651_;
  wire _35652_;
  wire _35653_;
  wire _35654_;
  wire _35655_;
  wire _35656_;
  wire _35657_;
  wire _35658_;
  wire _35659_;
  wire _35660_;
  wire _35661_;
  wire _35662_;
  wire _35663_;
  wire _35664_;
  wire _35665_;
  wire _35666_;
  wire _35667_;
  wire _35668_;
  wire _35669_;
  wire _35670_;
  wire _35671_;
  wire _35672_;
  wire _35673_;
  wire _35674_;
  wire _35675_;
  wire _35676_;
  wire _35677_;
  wire _35678_;
  wire _35679_;
  wire _35680_;
  wire _35681_;
  wire _35682_;
  wire _35683_;
  wire _35684_;
  wire _35685_;
  wire _35686_;
  wire _35687_;
  wire _35688_;
  wire _35689_;
  wire _35690_;
  wire _35691_;
  wire _35692_;
  wire _35693_;
  wire _35694_;
  wire _35695_;
  wire _35696_;
  wire _35697_;
  wire _35698_;
  wire _35699_;
  wire _35700_;
  wire _35701_;
  wire _35702_;
  wire _35703_;
  wire _35704_;
  wire _35705_;
  wire _35706_;
  wire _35707_;
  wire _35708_;
  wire _35709_;
  wire _35710_;
  wire _35711_;
  wire _35712_;
  wire _35713_;
  wire _35714_;
  wire _35715_;
  wire _35716_;
  wire _35717_;
  wire _35718_;
  wire _35719_;
  wire _35720_;
  wire _35721_;
  wire _35722_;
  wire _35723_;
  wire _35724_;
  wire _35725_;
  wire _35726_;
  wire _35727_;
  wire _35728_;
  wire _35729_;
  wire _35730_;
  wire _35731_;
  wire _35732_;
  wire _35733_;
  wire _35734_;
  wire _35735_;
  wire _35736_;
  wire _35737_;
  wire _35738_;
  wire _35739_;
  wire _35740_;
  wire _35741_;
  wire _35742_;
  wire _35743_;
  wire _35744_;
  wire _35745_;
  wire _35746_;
  wire _35747_;
  wire _35748_;
  wire _35749_;
  wire _35750_;
  wire _35751_;
  wire _35752_;
  wire _35753_;
  wire _35754_;
  wire _35755_;
  wire _35756_;
  wire _35757_;
  wire _35758_;
  wire _35759_;
  wire _35760_;
  wire _35761_;
  wire _35762_;
  wire _35763_;
  wire _35764_;
  wire _35765_;
  wire _35766_;
  wire _35767_;
  wire _35768_;
  wire _35769_;
  wire _35770_;
  wire _35771_;
  wire _35772_;
  wire _35773_;
  wire _35774_;
  wire _35775_;
  wire _35776_;
  wire _35777_;
  wire _35778_;
  wire _35779_;
  wire _35780_;
  wire _35781_;
  wire _35782_;
  wire _35783_;
  wire _35784_;
  wire _35785_;
  wire _35786_;
  wire _35787_;
  wire _35788_;
  wire _35789_;
  wire _35790_;
  wire _35791_;
  wire _35792_;
  wire _35793_;
  wire _35794_;
  wire _35795_;
  wire _35796_;
  wire _35797_;
  wire _35798_;
  wire _35799_;
  wire _35800_;
  wire _35801_;
  wire _35802_;
  wire _35803_;
  wire _35804_;
  wire _35805_;
  wire _35806_;
  wire _35807_;
  wire _35808_;
  wire _35809_;
  wire _35810_;
  wire _35811_;
  wire _35812_;
  wire _35813_;
  wire _35814_;
  wire _35815_;
  wire _35816_;
  wire _35817_;
  wire _35818_;
  wire _35819_;
  wire _35820_;
  wire _35821_;
  wire _35822_;
  wire _35823_;
  wire _35824_;
  wire _35825_;
  wire _35826_;
  wire _35827_;
  wire _35828_;
  wire _35829_;
  wire _35830_;
  wire _35831_;
  wire _35832_;
  wire _35833_;
  wire _35834_;
  wire _35835_;
  wire _35836_;
  wire _35837_;
  wire _35838_;
  wire _35839_;
  wire _35840_;
  wire _35841_;
  wire _35842_;
  wire _35843_;
  wire _35844_;
  wire _35845_;
  wire _35846_;
  wire _35847_;
  wire _35848_;
  wire _35849_;
  wire _35850_;
  wire _35851_;
  wire _35852_;
  wire _35853_;
  wire _35854_;
  wire _35855_;
  wire _35856_;
  wire _35857_;
  wire _35858_;
  wire _35859_;
  wire _35860_;
  wire _35861_;
  wire _35862_;
  wire _35863_;
  wire _35864_;
  wire _35865_;
  wire _35866_;
  wire _35867_;
  wire _35868_;
  wire _35869_;
  wire _35870_;
  wire _35871_;
  wire _35872_;
  wire _35873_;
  wire _35874_;
  wire _35875_;
  wire _35876_;
  wire _35877_;
  wire _35878_;
  wire _35879_;
  wire _35880_;
  wire _35881_;
  wire _35882_;
  wire _35883_;
  wire _35884_;
  wire _35885_;
  wire _35886_;
  wire _35887_;
  wire _35888_;
  wire _35889_;
  wire _35890_;
  wire _35891_;
  wire _35892_;
  wire _35893_;
  wire _35894_;
  wire _35895_;
  wire _35896_;
  wire _35897_;
  wire _35898_;
  wire _35899_;
  wire _35900_;
  wire _35901_;
  wire _35902_;
  wire _35903_;
  wire _35904_;
  wire _35905_;
  wire _35906_;
  wire _35907_;
  wire _35908_;
  wire _35909_;
  wire _35910_;
  wire _35911_;
  wire _35912_;
  wire _35913_;
  wire _35914_;
  wire _35915_;
  wire _35916_;
  wire _35917_;
  wire _35918_;
  wire _35919_;
  wire _35920_;
  wire _35921_;
  wire _35922_;
  wire _35923_;
  wire _35924_;
  wire _35925_;
  wire _35926_;
  wire _35927_;
  wire _35928_;
  wire _35929_;
  wire _35930_;
  wire _35931_;
  wire _35932_;
  wire _35933_;
  wire _35934_;
  wire _35935_;
  wire _35936_;
  wire _35937_;
  wire _35938_;
  wire _35939_;
  wire _35940_;
  wire _35941_;
  wire _35942_;
  wire _35943_;
  wire _35944_;
  wire _35945_;
  wire _35946_;
  wire _35947_;
  wire _35948_;
  wire _35949_;
  wire _35950_;
  wire _35951_;
  wire _35952_;
  wire _35953_;
  wire _35954_;
  wire _35955_;
  wire _35956_;
  wire _35957_;
  wire _35958_;
  wire _35959_;
  wire _35960_;
  wire _35961_;
  wire _35962_;
  wire _35963_;
  wire _35964_;
  wire _35965_;
  wire _35966_;
  wire _35967_;
  wire _35968_;
  wire _35969_;
  wire _35970_;
  wire _35971_;
  wire _35972_;
  wire _35973_;
  wire _35974_;
  wire _35975_;
  wire _35976_;
  wire _35977_;
  wire _35978_;
  wire _35979_;
  wire _35980_;
  wire _35981_;
  wire _35982_;
  wire _35983_;
  wire _35984_;
  wire _35985_;
  wire _35986_;
  wire _35987_;
  wire _35988_;
  wire _35989_;
  wire _35990_;
  wire _35991_;
  wire _35992_;
  wire _35993_;
  wire _35994_;
  wire _35995_;
  wire _35996_;
  wire _35997_;
  wire _35998_;
  wire _35999_;
  wire _36000_;
  wire _36001_;
  wire _36002_;
  wire _36003_;
  wire _36004_;
  wire _36005_;
  wire _36006_;
  wire _36007_;
  wire _36008_;
  wire _36009_;
  wire _36010_;
  wire _36011_;
  wire _36012_;
  wire _36013_;
  wire _36014_;
  wire _36015_;
  wire _36016_;
  wire _36017_;
  wire _36018_;
  wire _36019_;
  wire _36020_;
  wire _36021_;
  wire _36022_;
  wire _36023_;
  wire _36024_;
  wire _36025_;
  wire _36026_;
  wire _36027_;
  wire _36028_;
  wire _36029_;
  wire _36030_;
  wire _36031_;
  wire _36032_;
  wire _36033_;
  wire _36034_;
  wire _36035_;
  wire _36036_;
  wire _36037_;
  wire _36038_;
  wire _36039_;
  wire _36040_;
  wire _36041_;
  wire _36042_;
  wire _36043_;
  wire _36044_;
  wire _36045_;
  wire _36046_;
  wire _36047_;
  wire _36048_;
  wire _36049_;
  wire _36050_;
  wire _36051_;
  wire _36052_;
  wire _36053_;
  wire _36054_;
  wire _36055_;
  wire _36056_;
  wire _36057_;
  wire _36058_;
  wire _36059_;
  wire _36060_;
  wire _36061_;
  wire _36062_;
  wire _36063_;
  wire _36064_;
  wire _36065_;
  wire _36066_;
  wire _36067_;
  wire _36068_;
  wire _36069_;
  wire _36070_;
  wire _36071_;
  wire _36072_;
  wire _36073_;
  wire _36074_;
  wire _36075_;
  wire _36076_;
  wire _36077_;
  wire _36078_;
  wire _36079_;
  wire _36080_;
  wire _36081_;
  wire _36082_;
  wire _36083_;
  wire _36084_;
  wire _36085_;
  wire _36086_;
  wire _36087_;
  wire _36088_;
  wire _36089_;
  wire _36090_;
  wire _36091_;
  wire _36092_;
  wire _36093_;
  wire _36094_;
  wire _36095_;
  wire _36096_;
  wire _36097_;
  wire _36098_;
  wire _36099_;
  wire _36100_;
  wire _36101_;
  wire _36102_;
  wire _36103_;
  wire _36104_;
  wire _36105_;
  wire _36106_;
  wire _36107_;
  wire _36108_;
  wire _36109_;
  wire _36110_;
  wire _36111_;
  wire _36112_;
  wire _36113_;
  wire _36114_;
  wire _36115_;
  wire _36116_;
  wire _36117_;
  wire _36118_;
  wire _36119_;
  wire _36120_;
  wire _36121_;
  wire _36122_;
  wire _36123_;
  wire _36124_;
  wire _36125_;
  wire _36126_;
  wire _36127_;
  wire _36128_;
  wire _36129_;
  wire _36130_;
  wire _36131_;
  wire _36132_;
  wire _36133_;
  wire _36134_;
  wire _36135_;
  wire _36136_;
  wire _36137_;
  wire _36138_;
  wire _36139_;
  wire _36140_;
  wire _36141_;
  wire _36142_;
  wire _36143_;
  wire _36144_;
  wire _36145_;
  wire _36146_;
  wire _36147_;
  wire _36148_;
  wire _36149_;
  wire _36150_;
  wire _36151_;
  wire _36152_;
  wire _36153_;
  wire _36154_;
  wire _36155_;
  wire _36156_;
  wire _36157_;
  wire _36158_;
  wire _36159_;
  wire _36160_;
  wire _36161_;
  wire _36162_;
  wire _36163_;
  wire _36164_;
  wire _36165_;
  wire _36166_;
  wire _36167_;
  wire _36168_;
  wire _36169_;
  wire _36170_;
  wire _36171_;
  wire _36172_;
  wire _36173_;
  wire _36174_;
  wire _36175_;
  wire _36176_;
  wire _36177_;
  wire _36178_;
  wire _36179_;
  wire _36180_;
  wire _36181_;
  wire _36182_;
  wire _36183_;
  wire _36184_;
  wire _36185_;
  wire _36186_;
  wire _36187_;
  wire _36188_;
  wire _36189_;
  wire _36190_;
  wire _36191_;
  wire _36192_;
  wire _36193_;
  wire _36194_;
  wire _36195_;
  wire _36196_;
  wire _36197_;
  wire _36198_;
  wire _36199_;
  wire _36200_;
  wire _36201_;
  wire _36202_;
  wire _36203_;
  wire _36204_;
  wire _36205_;
  wire _36206_;
  wire _36207_;
  wire _36208_;
  wire _36209_;
  wire _36210_;
  wire _36211_;
  wire _36212_;
  wire _36213_;
  wire _36214_;
  wire _36215_;
  wire _36216_;
  wire _36217_;
  wire _36218_;
  wire _36219_;
  wire _36220_;
  wire _36221_;
  wire _36222_;
  wire _36223_;
  wire _36224_;
  wire _36225_;
  wire _36226_;
  wire _36227_;
  wire _36228_;
  wire _36229_;
  wire _36230_;
  wire _36231_;
  wire _36232_;
  wire _36233_;
  wire _36234_;
  wire _36235_;
  wire _36236_;
  wire _36237_;
  wire _36238_;
  wire _36239_;
  wire _36240_;
  wire _36241_;
  wire _36242_;
  wire _36243_;
  wire _36244_;
  wire _36245_;
  wire _36246_;
  wire _36247_;
  wire _36248_;
  wire _36249_;
  wire _36250_;
  wire _36251_;
  wire _36252_;
  wire _36253_;
  wire _36254_;
  wire _36255_;
  wire _36256_;
  wire _36257_;
  wire _36258_;
  wire _36259_;
  wire _36260_;
  wire _36261_;
  wire _36262_;
  wire _36263_;
  wire _36264_;
  wire _36265_;
  wire _36266_;
  wire _36267_;
  wire _36268_;
  wire _36269_;
  wire _36270_;
  wire _36271_;
  wire _36272_;
  wire _36273_;
  wire _36274_;
  wire _36275_;
  wire _36276_;
  wire _36277_;
  wire _36278_;
  wire _36279_;
  wire _36280_;
  wire _36281_;
  wire _36282_;
  wire _36283_;
  wire _36284_;
  wire _36285_;
  wire _36286_;
  wire _36287_;
  wire _36288_;
  wire _36289_;
  wire _36290_;
  wire _36291_;
  wire _36292_;
  wire _36293_;
  wire _36294_;
  wire _36295_;
  wire _36296_;
  wire _36297_;
  wire _36298_;
  wire _36299_;
  wire _36300_;
  wire _36301_;
  wire _36302_;
  wire _36303_;
  wire _36304_;
  wire _36305_;
  wire _36306_;
  wire _36307_;
  wire _36308_;
  wire _36309_;
  wire _36310_;
  wire _36311_;
  wire _36312_;
  wire _36313_;
  wire _36314_;
  wire _36315_;
  wire _36316_;
  wire _36317_;
  wire _36318_;
  wire _36319_;
  wire _36320_;
  wire _36321_;
  wire _36322_;
  wire _36323_;
  wire _36324_;
  wire _36325_;
  wire _36326_;
  wire _36327_;
  wire _36328_;
  wire _36329_;
  wire _36330_;
  wire _36331_;
  wire _36332_;
  wire _36333_;
  wire _36334_;
  wire _36335_;
  wire _36336_;
  wire _36337_;
  wire _36338_;
  wire _36339_;
  wire _36340_;
  wire _36341_;
  wire _36342_;
  wire _36343_;
  wire _36344_;
  wire _36345_;
  wire _36346_;
  wire _36347_;
  wire _36348_;
  wire _36349_;
  wire _36350_;
  wire _36351_;
  wire _36352_;
  wire _36353_;
  wire _36354_;
  wire _36355_;
  wire _36356_;
  wire _36357_;
  wire _36358_;
  wire _36359_;
  wire _36360_;
  wire _36361_;
  wire _36362_;
  wire _36363_;
  wire _36364_;
  wire _36365_;
  wire _36366_;
  wire _36367_;
  wire _36368_;
  wire _36369_;
  wire _36370_;
  wire _36371_;
  wire _36372_;
  wire _36373_;
  wire _36374_;
  wire _36375_;
  wire _36376_;
  wire _36377_;
  wire _36378_;
  wire _36379_;
  wire _36380_;
  wire _36381_;
  wire _36382_;
  wire _36383_;
  wire _36384_;
  wire _36385_;
  wire _36386_;
  wire _36387_;
  wire _36388_;
  wire _36389_;
  wire _36390_;
  wire _36391_;
  wire _36392_;
  wire _36393_;
  wire _36394_;
  wire _36395_;
  wire _36396_;
  wire _36397_;
  wire _36398_;
  wire _36399_;
  wire _36400_;
  wire _36401_;
  wire _36402_;
  wire _36403_;
  wire _36404_;
  wire _36405_;
  wire _36406_;
  wire _36407_;
  wire _36408_;
  wire _36409_;
  wire _36410_;
  wire _36411_;
  wire _36412_;
  wire _36413_;
  wire _36414_;
  wire _36415_;
  wire _36416_;
  wire _36417_;
  wire _36418_;
  wire _36419_;
  wire _36420_;
  wire _36421_;
  wire _36422_;
  wire _36423_;
  wire _36424_;
  wire _36425_;
  wire _36426_;
  wire _36427_;
  wire _36428_;
  wire _36429_;
  wire _36430_;
  wire _36431_;
  wire _36432_;
  wire _36433_;
  wire _36434_;
  wire _36435_;
  wire _36436_;
  wire _36437_;
  wire _36438_;
  wire _36439_;
  wire _36440_;
  wire _36441_;
  wire _36442_;
  wire _36443_;
  wire _36444_;
  wire _36445_;
  wire _36446_;
  wire _36447_;
  wire _36448_;
  wire _36449_;
  wire _36450_;
  wire _36451_;
  wire _36452_;
  wire _36453_;
  wire _36454_;
  wire _36455_;
  wire _36456_;
  wire _36457_;
  wire _36458_;
  wire _36459_;
  wire _36460_;
  wire _36461_;
  wire _36462_;
  wire _36463_;
  wire _36464_;
  wire _36465_;
  wire _36466_;
  wire _36467_;
  wire _36468_;
  wire _36469_;
  wire _36470_;
  wire _36471_;
  wire _36472_;
  wire _36473_;
  wire _36474_;
  wire _36475_;
  wire _36476_;
  wire _36477_;
  wire _36478_;
  wire _36479_;
  wire _36480_;
  wire _36481_;
  wire _36482_;
  wire _36483_;
  wire _36484_;
  wire _36485_;
  wire _36486_;
  wire _36487_;
  wire _36488_;
  wire _36489_;
  wire _36490_;
  wire _36491_;
  wire _36492_;
  wire _36493_;
  wire _36494_;
  wire _36495_;
  wire _36496_;
  wire _36497_;
  wire _36498_;
  wire _36499_;
  wire _36500_;
  wire _36501_;
  wire _36502_;
  wire _36503_;
  wire _36504_;
  wire _36505_;
  wire _36506_;
  wire _36507_;
  wire _36508_;
  wire _36509_;
  wire _36510_;
  wire _36511_;
  wire _36512_;
  wire _36513_;
  wire _36514_;
  wire _36515_;
  wire _36516_;
  wire _36517_;
  wire _36518_;
  wire _36519_;
  wire _36520_;
  wire _36521_;
  wire _36522_;
  wire _36523_;
  wire _36524_;
  wire _36525_;
  wire _36526_;
  wire _36527_;
  wire _36528_;
  wire _36529_;
  wire _36530_;
  wire _36531_;
  wire _36532_;
  wire _36533_;
  wire _36534_;
  wire _36535_;
  wire _36536_;
  wire _36537_;
  wire _36538_;
  wire _36539_;
  wire _36540_;
  wire _36541_;
  wire _36542_;
  wire _36543_;
  wire _36544_;
  wire _36545_;
  wire _36546_;
  wire _36547_;
  wire _36548_;
  wire _36549_;
  wire _36550_;
  wire _36551_;
  wire _36552_;
  wire _36553_;
  wire _36554_;
  wire _36555_;
  wire _36556_;
  wire _36557_;
  wire _36558_;
  wire _36559_;
  wire _36560_;
  wire _36561_;
  wire _36562_;
  wire _36563_;
  wire _36564_;
  wire _36565_;
  wire _36566_;
  wire _36567_;
  wire _36568_;
  wire _36569_;
  wire _36570_;
  wire _36571_;
  wire _36572_;
  wire _36573_;
  wire _36574_;
  wire _36575_;
  wire _36576_;
  wire _36577_;
  wire _36578_;
  wire _36579_;
  wire _36580_;
  wire _36581_;
  wire _36582_;
  wire _36583_;
  wire _36584_;
  wire _36585_;
  wire _36586_;
  wire _36587_;
  wire _36588_;
  wire _36589_;
  wire _36590_;
  wire _36591_;
  wire _36592_;
  wire _36593_;
  wire _36594_;
  wire _36595_;
  wire _36596_;
  wire _36597_;
  wire _36598_;
  wire _36599_;
  wire _36600_;
  wire _36601_;
  wire _36602_;
  wire _36603_;
  wire _36604_;
  wire _36605_;
  wire _36606_;
  wire _36607_;
  wire _36608_;
  wire _36609_;
  wire _36610_;
  wire _36611_;
  wire _36612_;
  wire _36613_;
  wire _36614_;
  wire _36615_;
  wire _36616_;
  wire _36617_;
  wire _36618_;
  wire _36619_;
  wire _36620_;
  wire _36621_;
  wire _36622_;
  wire _36623_;
  wire _36624_;
  wire _36625_;
  wire _36626_;
  wire _36627_;
  wire _36628_;
  wire _36629_;
  wire _36630_;
  wire _36631_;
  wire _36632_;
  wire _36633_;
  wire _36634_;
  wire _36635_;
  wire _36636_;
  wire _36637_;
  wire _36638_;
  wire _36639_;
  wire _36640_;
  wire _36641_;
  wire _36642_;
  wire _36643_;
  wire _36644_;
  wire _36645_;
  wire _36646_;
  wire _36647_;
  wire _36648_;
  wire _36649_;
  wire _36650_;
  wire _36651_;
  wire _36652_;
  wire _36653_;
  wire _36654_;
  wire _36655_;
  wire _36656_;
  wire _36657_;
  wire _36658_;
  wire _36659_;
  wire _36660_;
  wire _36661_;
  wire _36662_;
  wire _36663_;
  wire _36664_;
  wire _36665_;
  wire _36666_;
  wire _36667_;
  wire _36668_;
  wire _36669_;
  wire _36670_;
  wire _36671_;
  wire _36672_;
  wire _36673_;
  wire _36674_;
  wire _36675_;
  wire _36676_;
  wire _36677_;
  wire _36678_;
  wire _36679_;
  wire _36680_;
  wire _36681_;
  wire _36682_;
  wire _36683_;
  wire _36684_;
  wire _36685_;
  wire _36686_;
  wire _36687_;
  wire _36688_;
  wire _36689_;
  wire _36690_;
  wire _36691_;
  wire _36692_;
  wire _36693_;
  wire _36694_;
  wire _36695_;
  wire _36696_;
  wire _36697_;
  wire _36698_;
  wire _36699_;
  wire _36700_;
  wire _36701_;
  wire _36702_;
  wire _36703_;
  wire _36704_;
  wire _36705_;
  wire _36706_;
  wire _36707_;
  wire _36708_;
  wire _36709_;
  wire _36710_;
  wire _36711_;
  wire _36712_;
  wire _36713_;
  wire _36714_;
  wire _36715_;
  wire _36716_;
  wire _36717_;
  wire _36718_;
  wire _36719_;
  wire _36720_;
  wire _36721_;
  wire _36722_;
  wire _36723_;
  wire _36724_;
  wire _36725_;
  wire _36726_;
  wire _36727_;
  wire _36728_;
  wire _36729_;
  wire _36730_;
  wire _36731_;
  wire _36732_;
  wire _36733_;
  wire _36734_;
  wire _36735_;
  wire _36736_;
  wire _36737_;
  wire _36738_;
  wire _36739_;
  wire _36740_;
  wire _36741_;
  wire _36742_;
  wire _36743_;
  wire _36744_;
  wire _36745_;
  wire _36746_;
  wire _36747_;
  wire _36748_;
  wire _36749_;
  wire _36750_;
  wire _36751_;
  wire _36752_;
  wire _36753_;
  wire _36754_;
  wire _36755_;
  wire _36756_;
  wire _36757_;
  wire _36758_;
  wire _36759_;
  wire _36760_;
  wire _36761_;
  wire _36762_;
  wire _36763_;
  wire _36764_;
  wire _36765_;
  wire _36766_;
  wire _36767_;
  wire _36768_;
  wire _36769_;
  wire _36770_;
  wire _36771_;
  wire _36772_;
  wire _36773_;
  wire _36774_;
  wire _36775_;
  wire _36776_;
  wire _36777_;
  wire _36778_;
  wire _36779_;
  wire _36780_;
  wire _36781_;
  wire _36782_;
  wire _36783_;
  wire _36784_;
  wire _36785_;
  wire _36786_;
  wire _36787_;
  wire _36788_;
  wire _36789_;
  wire _36790_;
  wire _36791_;
  wire _36792_;
  wire _36793_;
  wire _36794_;
  wire _36795_;
  wire _36796_;
  wire _36797_;
  wire _36798_;
  wire _36799_;
  wire _36800_;
  wire _36801_;
  wire _36802_;
  wire _36803_;
  wire _36804_;
  wire _36805_;
  wire _36806_;
  wire _36807_;
  wire _36808_;
  wire _36809_;
  wire _36810_;
  wire _36811_;
  wire _36812_;
  wire _36813_;
  wire _36814_;
  wire _36815_;
  wire _36816_;
  wire _36817_;
  wire _36818_;
  wire _36819_;
  wire _36820_;
  wire _36821_;
  wire _36822_;
  wire _36823_;
  wire _36824_;
  wire _36825_;
  wire _36826_;
  wire _36827_;
  wire _36828_;
  wire _36829_;
  wire _36830_;
  wire _36831_;
  wire _36832_;
  wire _36833_;
  wire _36834_;
  wire _36835_;
  wire _36836_;
  wire _36837_;
  wire _36838_;
  wire _36839_;
  wire _36840_;
  wire _36841_;
  wire _36842_;
  wire _36843_;
  wire _36844_;
  wire _36845_;
  wire _36846_;
  wire _36847_;
  wire _36848_;
  wire _36849_;
  wire _36850_;
  wire _36851_;
  wire _36852_;
  wire _36853_;
  wire _36854_;
  wire _36855_;
  wire _36856_;
  wire _36857_;
  wire _36858_;
  wire _36859_;
  wire _36860_;
  wire _36861_;
  wire _36862_;
  wire _36863_;
  wire _36864_;
  wire _36865_;
  wire _36866_;
  wire _36867_;
  wire _36868_;
  wire _36869_;
  wire _36870_;
  wire _36871_;
  wire _36872_;
  wire _36873_;
  wire _36874_;
  wire _36875_;
  wire _36876_;
  wire _36877_;
  wire _36878_;
  wire _36879_;
  wire _36880_;
  wire _36881_;
  wire _36882_;
  wire _36883_;
  wire _36884_;
  wire _36885_;
  wire _36886_;
  wire _36887_;
  wire _36888_;
  wire _36889_;
  wire _36890_;
  wire _36891_;
  wire _36892_;
  wire _36893_;
  wire _36894_;
  wire _36895_;
  wire _36896_;
  wire _36897_;
  wire _36898_;
  wire _36899_;
  wire _36900_;
  wire _36901_;
  wire _36902_;
  wire _36903_;
  wire _36904_;
  wire _36905_;
  wire _36906_;
  wire _36907_;
  wire _36908_;
  wire _36909_;
  wire _36910_;
  wire _36911_;
  wire _36912_;
  wire _36913_;
  wire _36914_;
  wire _36915_;
  wire _36916_;
  wire _36917_;
  wire _36918_;
  wire _36919_;
  wire _36920_;
  wire _36921_;
  wire _36922_;
  wire _36923_;
  wire _36924_;
  wire _36925_;
  wire _36926_;
  wire _36927_;
  wire _36928_;
  wire _36929_;
  wire _36930_;
  wire _36931_;
  wire _36932_;
  wire _36933_;
  wire _36934_;
  wire _36935_;
  wire _36936_;
  wire _36937_;
  wire _36938_;
  wire _36939_;
  wire _36940_;
  wire _36941_;
  wire _36942_;
  wire _36943_;
  wire _36944_;
  wire _36945_;
  wire _36946_;
  wire _36947_;
  wire _36948_;
  wire _36949_;
  wire _36950_;
  wire _36951_;
  wire _36952_;
  wire _36953_;
  wire _36954_;
  wire _36955_;
  wire _36956_;
  wire _36957_;
  wire _36958_;
  wire _36959_;
  wire _36960_;
  wire _36961_;
  wire _36962_;
  wire _36963_;
  wire _36964_;
  wire _36965_;
  wire _36966_;
  wire _36967_;
  wire _36968_;
  wire _36969_;
  wire _36970_;
  wire _36971_;
  wire _36972_;
  wire _36973_;
  wire _36974_;
  wire _36975_;
  wire _36976_;
  wire _36977_;
  wire _36978_;
  wire _36979_;
  wire _36980_;
  wire _36981_;
  wire _36982_;
  wire _36983_;
  wire _36984_;
  wire _36985_;
  wire _36986_;
  wire _36987_;
  wire _36988_;
  wire _36989_;
  wire _36990_;
  wire _36991_;
  wire _36992_;
  wire _36993_;
  wire _36994_;
  wire _36995_;
  wire _36996_;
  wire _36997_;
  wire _36998_;
  wire _36999_;
  wire _37000_;
  wire _37001_;
  wire _37002_;
  wire _37003_;
  wire _37004_;
  wire _37005_;
  wire _37006_;
  wire _37007_;
  wire _37008_;
  wire _37009_;
  wire _37010_;
  wire _37011_;
  wire _37012_;
  wire _37013_;
  wire _37014_;
  wire _37015_;
  wire _37016_;
  wire _37017_;
  wire _37018_;
  wire _37019_;
  wire _37020_;
  wire _37021_;
  wire _37022_;
  wire _37023_;
  wire _37024_;
  wire _37025_;
  wire _37026_;
  wire _37027_;
  wire _37028_;
  wire _37029_;
  wire _37030_;
  wire _37031_;
  wire _37032_;
  wire _37033_;
  wire _37034_;
  wire _37035_;
  wire _37036_;
  wire _37037_;
  wire _37038_;
  wire _37039_;
  wire _37040_;
  wire _37041_;
  wire _37042_;
  wire _37043_;
  wire _37044_;
  wire _37045_;
  wire _37046_;
  wire _37047_;
  wire _37048_;
  wire _37049_;
  wire _37050_;
  wire _37051_;
  wire _37052_;
  wire _37053_;
  wire _37054_;
  wire _37055_;
  wire _37056_;
  wire _37057_;
  wire _37058_;
  wire _37059_;
  wire _37060_;
  wire _37061_;
  wire _37062_;
  wire _37063_;
  wire _37064_;
  wire _37065_;
  wire _37066_;
  wire _37067_;
  wire _37068_;
  wire _37069_;
  wire _37070_;
  wire _37071_;
  wire _37072_;
  wire _37073_;
  wire _37074_;
  wire _37075_;
  wire _37076_;
  wire _37077_;
  wire _37078_;
  wire _37079_;
  wire _37080_;
  wire _37081_;
  wire _37082_;
  wire _37083_;
  wire _37084_;
  wire _37085_;
  wire _37086_;
  wire _37087_;
  wire _37088_;
  wire _37089_;
  wire _37090_;
  wire _37091_;
  wire _37092_;
  wire _37093_;
  wire _37094_;
  wire _37095_;
  wire _37096_;
  wire _37097_;
  wire _37098_;
  wire _37099_;
  wire _37100_;
  wire _37101_;
  wire _37102_;
  wire _37103_;
  wire _37104_;
  wire _37105_;
  wire _37106_;
  wire _37107_;
  wire _37108_;
  wire _37109_;
  wire _37110_;
  wire _37111_;
  wire _37112_;
  wire _37113_;
  wire _37114_;
  wire _37115_;
  wire _37116_;
  wire _37117_;
  wire _37118_;
  wire _37119_;
  wire _37120_;
  wire _37121_;
  wire _37122_;
  wire _37123_;
  wire _37124_;
  wire _37125_;
  wire _37126_;
  wire _37127_;
  wire _37128_;
  wire _37129_;
  wire _37130_;
  wire _37131_;
  wire _37132_;
  wire _37133_;
  wire _37134_;
  wire _37135_;
  wire _37136_;
  wire _37137_;
  wire _37138_;
  wire _37139_;
  wire _37140_;
  wire _37141_;
  wire _37142_;
  wire _37143_;
  wire _37144_;
  wire _37145_;
  wire _37146_;
  wire _37147_;
  wire _37148_;
  wire _37149_;
  wire _37150_;
  wire _37151_;
  wire _37152_;
  wire _37153_;
  wire _37154_;
  wire _37155_;
  wire _37156_;
  wire _37157_;
  wire _37158_;
  wire _37159_;
  wire _37160_;
  wire _37161_;
  wire _37162_;
  wire _37163_;
  wire _37164_;
  wire _37165_;
  wire _37166_;
  wire _37167_;
  wire _37168_;
  wire _37169_;
  wire _37170_;
  wire _37171_;
  wire _37172_;
  wire _37173_;
  wire _37174_;
  wire _37175_;
  wire _37176_;
  wire _37177_;
  wire _37178_;
  wire _37179_;
  wire _37180_;
  wire _37181_;
  wire _37182_;
  wire _37183_;
  wire _37184_;
  wire _37185_;
  wire _37186_;
  wire _37187_;
  wire _37188_;
  wire _37189_;
  wire _37190_;
  wire _37191_;
  wire _37192_;
  wire _37193_;
  wire _37194_;
  wire _37195_;
  wire _37196_;
  wire _37197_;
  wire _37198_;
  wire _37199_;
  wire _37200_;
  wire _37201_;
  wire _37202_;
  wire _37203_;
  wire _37204_;
  wire _37205_;
  wire _37206_;
  wire _37207_;
  wire _37208_;
  wire _37209_;
  wire _37210_;
  wire _37211_;
  wire _37212_;
  wire _37213_;
  wire _37214_;
  wire _37215_;
  wire _37216_;
  wire _37217_;
  wire _37218_;
  wire _37219_;
  wire _37220_;
  wire _37221_;
  wire _37222_;
  wire _37223_;
  wire _37224_;
  wire _37225_;
  wire _37226_;
  wire _37227_;
  wire _37228_;
  wire _37229_;
  wire _37230_;
  wire _37231_;
  wire _37232_;
  wire _37233_;
  wire _37234_;
  wire _37235_;
  wire _37236_;
  wire _37237_;
  wire _37238_;
  wire _37239_;
  wire _37240_;
  wire _37241_;
  wire _37242_;
  wire _37243_;
  wire _37244_;
  wire _37245_;
  wire _37246_;
  wire _37247_;
  wire _37248_;
  wire _37249_;
  wire _37250_;
  wire _37251_;
  wire _37252_;
  wire _37253_;
  wire _37254_;
  wire _37255_;
  wire _37256_;
  wire _37257_;
  wire _37258_;
  wire _37259_;
  wire _37260_;
  wire _37261_;
  wire _37262_;
  wire _37263_;
  wire _37264_;
  wire _37265_;
  wire _37266_;
  wire _37267_;
  wire _37268_;
  wire _37269_;
  wire _37270_;
  wire _37271_;
  wire _37272_;
  wire _37273_;
  wire _37274_;
  wire _37275_;
  wire _37276_;
  wire _37277_;
  wire _37278_;
  wire _37279_;
  wire _37280_;
  wire _37281_;
  wire _37282_;
  wire _37283_;
  wire _37284_;
  wire _37285_;
  wire _37286_;
  wire _37287_;
  wire _37288_;
  wire _37289_;
  wire _37290_;
  wire _37291_;
  wire _37292_;
  wire _37293_;
  wire _37294_;
  wire _37295_;
  wire _37296_;
  wire _37297_;
  wire _37298_;
  wire _37299_;
  wire _37300_;
  wire _37301_;
  wire _37302_;
  wire _37303_;
  wire _37304_;
  wire _37305_;
  wire _37306_;
  wire _37307_;
  wire _37308_;
  wire _37309_;
  wire _37310_;
  wire _37311_;
  wire _37312_;
  wire _37313_;
  wire _37314_;
  wire _37315_;
  wire _37316_;
  wire _37317_;
  wire _37318_;
  wire _37319_;
  wire _37320_;
  wire _37321_;
  wire _37322_;
  wire _37323_;
  wire _37324_;
  wire _37325_;
  wire _37326_;
  wire _37327_;
  wire _37328_;
  wire _37329_;
  wire _37330_;
  wire _37331_;
  wire _37332_;
  wire _37333_;
  wire _37334_;
  wire _37335_;
  wire _37336_;
  wire _37337_;
  wire _37338_;
  wire _37339_;
  wire _37340_;
  wire _37341_;
  wire _37342_;
  wire _37343_;
  wire _37344_;
  wire _37345_;
  wire _37346_;
  wire _37347_;
  wire _37348_;
  wire _37349_;
  wire _37350_;
  wire _37351_;
  wire _37352_;
  wire _37353_;
  wire _37354_;
  wire _37355_;
  wire _37356_;
  wire _37357_;
  wire _37358_;
  wire _37359_;
  wire _37360_;
  wire _37361_;
  wire _37362_;
  wire _37363_;
  wire _37364_;
  wire _37365_;
  wire _37366_;
  wire _37367_;
  wire _37368_;
  wire _37369_;
  wire _37370_;
  wire _37371_;
  wire _37372_;
  wire _37373_;
  wire _37374_;
  wire _37375_;
  wire _37376_;
  wire _37377_;
  wire _37378_;
  wire _37379_;
  wire _37380_;
  wire _37381_;
  wire _37382_;
  wire _37383_;
  wire _37384_;
  wire _37385_;
  wire _37386_;
  wire _37387_;
  wire _37388_;
  wire _37389_;
  wire _37390_;
  wire _37391_;
  wire _37392_;
  wire _37393_;
  wire _37394_;
  wire _37395_;
  wire _37396_;
  wire _37397_;
  wire _37398_;
  wire _37399_;
  wire _37400_;
  wire _37401_;
  wire _37402_;
  wire _37403_;
  wire _37404_;
  wire _37405_;
  wire _37406_;
  wire _37407_;
  wire _37408_;
  wire _37409_;
  wire _37410_;
  wire _37411_;
  wire _37412_;
  wire _37413_;
  wire _37414_;
  wire _37415_;
  wire _37416_;
  wire _37417_;
  wire _37418_;
  wire _37419_;
  wire _37420_;
  wire _37421_;
  wire _37422_;
  wire _37423_;
  wire _37424_;
  wire _37425_;
  wire _37426_;
  wire _37427_;
  wire _37428_;
  wire _37429_;
  wire _37430_;
  wire _37431_;
  wire _37432_;
  wire _37433_;
  wire _37434_;
  wire _37435_;
  wire _37436_;
  wire _37437_;
  wire _37438_;
  wire _37439_;
  wire _37440_;
  wire _37441_;
  wire _37442_;
  wire _37443_;
  wire _37444_;
  wire _37445_;
  wire _37446_;
  wire _37447_;
  wire _37448_;
  wire _37449_;
  wire _37450_;
  wire _37451_;
  wire _37452_;
  wire _37453_;
  wire _37454_;
  wire _37455_;
  wire _37456_;
  wire _37457_;
  wire _37458_;
  wire _37459_;
  wire _37460_;
  wire _37461_;
  wire _37462_;
  wire _37463_;
  wire _37464_;
  wire _37465_;
  wire _37466_;
  wire _37467_;
  wire _37468_;
  wire _37469_;
  wire _37470_;
  wire _37471_;
  wire _37472_;
  wire _37473_;
  wire _37474_;
  wire _37475_;
  wire _37476_;
  wire _37477_;
  wire _37478_;
  wire _37479_;
  wire _37480_;
  wire _37481_;
  wire _37482_;
  wire _37483_;
  wire _37484_;
  wire _37485_;
  wire _37486_;
  wire _37487_;
  wire _37488_;
  wire _37489_;
  wire _37490_;
  wire _37491_;
  wire _37492_;
  wire _37493_;
  wire _37494_;
  wire _37495_;
  wire _37496_;
  wire _37497_;
  wire _37498_;
  wire _37499_;
  wire _37500_;
  wire _37501_;
  wire _37502_;
  wire _37503_;
  wire _37504_;
  wire _37505_;
  wire _37506_;
  wire _37507_;
  wire _37508_;
  wire _37509_;
  wire _37510_;
  wire _37511_;
  wire _37512_;
  wire _37513_;
  wire _37514_;
  wire _37515_;
  wire _37516_;
  wire _37517_;
  wire _37518_;
  wire _37519_;
  wire _37520_;
  wire _37521_;
  wire _37522_;
  wire _37523_;
  wire _37524_;
  wire _37525_;
  wire _37526_;
  wire _37527_;
  wire _37528_;
  wire _37529_;
  wire _37530_;
  wire _37531_;
  wire _37532_;
  wire _37533_;
  wire _37534_;
  wire _37535_;
  wire _37536_;
  wire _37537_;
  wire _37538_;
  wire _37539_;
  wire _37540_;
  wire _37541_;
  wire _37542_;
  wire _37543_;
  wire _37544_;
  wire _37545_;
  wire _37546_;
  wire _37547_;
  wire _37548_;
  wire _37549_;
  wire _37550_;
  wire _37551_;
  wire _37552_;
  wire _37553_;
  wire _37554_;
  wire _37555_;
  wire _37556_;
  wire _37557_;
  wire _37558_;
  wire _37559_;
  wire _37560_;
  wire _37561_;
  wire _37562_;
  wire _37563_;
  wire _37564_;
  wire _37565_;
  wire _37566_;
  wire _37567_;
  wire _37568_;
  wire _37569_;
  wire _37570_;
  wire _37571_;
  wire _37572_;
  wire _37573_;
  wire _37574_;
  wire _37575_;
  wire _37576_;
  wire _37577_;
  wire _37578_;
  wire _37579_;
  wire _37580_;
  wire _37581_;
  wire _37582_;
  wire _37583_;
  wire _37584_;
  wire _37585_;
  wire _37586_;
  wire _37587_;
  wire _37588_;
  wire _37589_;
  wire _37590_;
  wire _37591_;
  wire _37592_;
  wire _37593_;
  wire _37594_;
  wire _37595_;
  wire _37596_;
  wire _37597_;
  wire _37598_;
  wire _37599_;
  wire _37600_;
  wire _37601_;
  wire _37602_;
  wire _37603_;
  wire _37604_;
  wire _37605_;
  wire _37606_;
  wire _37607_;
  wire _37608_;
  wire _37609_;
  wire _37610_;
  wire _37611_;
  wire _37612_;
  wire _37613_;
  wire _37614_;
  wire _37615_;
  wire _37616_;
  wire _37617_;
  wire _37618_;
  wire _37619_;
  wire _37620_;
  wire _37621_;
  wire _37622_;
  wire _37623_;
  wire _37624_;
  wire _37625_;
  wire _37626_;
  wire _37627_;
  wire _37628_;
  wire _37629_;
  wire _37630_;
  wire _37631_;
  wire _37632_;
  wire _37633_;
  wire _37634_;
  wire _37635_;
  wire _37636_;
  wire _37637_;
  wire _37638_;
  wire _37639_;
  wire _37640_;
  wire _37641_;
  wire _37642_;
  wire _37643_;
  wire _37644_;
  wire _37645_;
  wire _37646_;
  wire _37647_;
  wire _37648_;
  wire _37649_;
  wire _37650_;
  wire _37651_;
  wire _37652_;
  wire _37653_;
  wire _37654_;
  wire _37655_;
  wire _37656_;
  wire _37657_;
  wire _37658_;
  wire _37659_;
  wire _37660_;
  wire _37661_;
  wire _37662_;
  wire _37663_;
  wire _37664_;
  wire _37665_;
  wire _37666_;
  wire _37667_;
  wire _37668_;
  wire _37669_;
  wire _37670_;
  wire _37671_;
  wire _37672_;
  wire _37673_;
  wire _37674_;
  wire _37675_;
  wire _37676_;
  wire _37677_;
  wire _37678_;
  wire _37679_;
  wire _37680_;
  wire _37681_;
  wire _37682_;
  wire _37683_;
  wire _37684_;
  wire _37685_;
  wire _37686_;
  wire _37687_;
  wire _37688_;
  wire _37689_;
  wire _37690_;
  wire _37691_;
  wire _37692_;
  wire _37693_;
  wire _37694_;
  wire _37695_;
  wire _37696_;
  wire _37697_;
  wire _37698_;
  wire _37699_;
  wire _37700_;
  wire _37701_;
  wire _37702_;
  wire _37703_;
  wire _37704_;
  wire _37705_;
  wire _37706_;
  wire _37707_;
  wire _37708_;
  wire _37709_;
  wire _37710_;
  wire _37711_;
  wire _37712_;
  wire _37713_;
  wire _37714_;
  wire _37715_;
  wire _37716_;
  wire _37717_;
  wire _37718_;
  wire _37719_;
  wire _37720_;
  wire _37721_;
  wire _37722_;
  wire _37723_;
  wire _37724_;
  wire _37725_;
  wire _37726_;
  wire _37727_;
  wire _37728_;
  wire _37729_;
  wire _37730_;
  wire _37731_;
  wire _37732_;
  wire _37733_;
  wire _37734_;
  wire _37735_;
  wire _37736_;
  wire _37737_;
  wire _37738_;
  wire _37739_;
  wire _37740_;
  wire _37741_;
  wire _37742_;
  wire _37743_;
  wire _37744_;
  wire _37745_;
  wire _37746_;
  wire _37747_;
  wire _37748_;
  wire _37749_;
  wire _37750_;
  wire _37751_;
  wire _37752_;
  wire _37753_;
  wire _37754_;
  wire _37755_;
  wire _37756_;
  wire _37757_;
  wire _37758_;
  wire _37759_;
  wire _37760_;
  wire _37761_;
  wire _37762_;
  wire _37763_;
  wire _37764_;
  wire _37765_;
  wire _37766_;
  wire _37767_;
  wire _37768_;
  wire _37769_;
  wire _37770_;
  wire _37771_;
  wire _37772_;
  wire _37773_;
  wire _37774_;
  wire _37775_;
  wire _37776_;
  wire _37777_;
  wire _37778_;
  wire _37779_;
  wire _37780_;
  wire _37781_;
  wire _37782_;
  wire _37783_;
  wire _37784_;
  wire _37785_;
  wire _37786_;
  wire _37787_;
  wire _37788_;
  wire _37789_;
  wire _37790_;
  wire _37791_;
  wire _37792_;
  wire _37793_;
  wire _37794_;
  wire _37795_;
  wire _37796_;
  wire _37797_;
  wire _37798_;
  wire _37799_;
  wire _37800_;
  wire _37801_;
  wire _37802_;
  wire _37803_;
  wire _37804_;
  wire _37805_;
  wire _37806_;
  wire _37807_;
  wire _37808_;
  wire _37809_;
  wire _37810_;
  wire _37811_;
  wire _37812_;
  wire _37813_;
  wire _37814_;
  wire _37815_;
  wire _37816_;
  wire _37817_;
  wire _37818_;
  wire _37819_;
  wire _37820_;
  wire _37821_;
  wire _37822_;
  wire _37823_;
  wire _37824_;
  wire _37825_;
  wire _37826_;
  wire _37827_;
  wire _37828_;
  wire _37829_;
  wire _37830_;
  wire _37831_;
  wire _37832_;
  wire _37833_;
  wire _37834_;
  wire _37835_;
  wire _37836_;
  wire _37837_;
  wire _37838_;
  wire _37839_;
  wire _37840_;
  wire _37841_;
  wire _37842_;
  wire _37843_;
  wire _37844_;
  wire _37845_;
  wire _37846_;
  wire _37847_;
  wire _37848_;
  wire _37849_;
  wire _37850_;
  wire _37851_;
  wire _37852_;
  wire _37853_;
  wire _37854_;
  wire _37855_;
  wire _37856_;
  wire _37857_;
  wire _37858_;
  wire _37859_;
  wire _37860_;
  wire _37861_;
  wire _37862_;
  wire _37863_;
  wire _37864_;
  wire _37865_;
  wire _37866_;
  wire _37867_;
  wire _37868_;
  wire _37869_;
  wire _37870_;
  wire _37871_;
  wire _37872_;
  wire _37873_;
  wire _37874_;
  wire _37875_;
  wire _37876_;
  wire _37877_;
  wire _37878_;
  wire _37879_;
  wire _37880_;
  wire _37881_;
  wire _37882_;
  wire _37883_;
  wire _37884_;
  wire _37885_;
  wire _37886_;
  wire _37887_;
  wire _37888_;
  wire _37889_;
  wire _37890_;
  wire _37891_;
  wire _37892_;
  wire _37893_;
  wire _37894_;
  wire _37895_;
  wire _37896_;
  wire _37897_;
  wire _37898_;
  wire _37899_;
  wire _37900_;
  wire _37901_;
  wire _37902_;
  wire _37903_;
  wire _37904_;
  wire _37905_;
  wire _37906_;
  wire _37907_;
  wire _37908_;
  wire _37909_;
  wire _37910_;
  wire _37911_;
  wire _37912_;
  wire _37913_;
  wire _37914_;
  wire _37915_;
  wire _37916_;
  wire _37917_;
  wire _37918_;
  wire _37919_;
  wire _37920_;
  wire _37921_;
  wire _37922_;
  wire _37923_;
  wire _37924_;
  wire _37925_;
  wire _37926_;
  wire _37927_;
  wire _37928_;
  wire _37929_;
  wire _37930_;
  wire _37931_;
  wire _37932_;
  wire _37933_;
  wire _37934_;
  wire _37935_;
  wire _37936_;
  wire _37937_;
  wire _37938_;
  wire _37939_;
  wire _37940_;
  wire _37941_;
  wire _37942_;
  wire _37943_;
  wire _37944_;
  wire _37945_;
  wire _37946_;
  wire _37947_;
  wire _37948_;
  wire _37949_;
  wire _37950_;
  wire _37951_;
  wire _37952_;
  wire _37953_;
  wire _37954_;
  wire _37955_;
  wire _37956_;
  wire _37957_;
  wire _37958_;
  wire _37959_;
  wire _37960_;
  wire _37961_;
  wire _37962_;
  wire _37963_;
  wire _37964_;
  wire _37965_;
  wire _37966_;
  wire _37967_;
  wire _37968_;
  wire _37969_;
  wire _37970_;
  wire _37971_;
  wire _37972_;
  wire _37973_;
  wire _37974_;
  wire _37975_;
  wire _37976_;
  wire _37977_;
  wire _37978_;
  wire _37979_;
  wire _37980_;
  wire _37981_;
  wire _37982_;
  wire _37983_;
  wire _37984_;
  wire _37985_;
  wire _37986_;
  wire _37987_;
  wire _37988_;
  wire _37989_;
  wire _37990_;
  wire _37991_;
  wire _37992_;
  wire _37993_;
  wire _37994_;
  wire _37995_;
  wire _37996_;
  wire _37997_;
  wire _37998_;
  wire _37999_;
  wire _38000_;
  wire _38001_;
  wire _38002_;
  wire _38003_;
  wire _38004_;
  wire _38005_;
  wire _38006_;
  wire _38007_;
  wire _38008_;
  wire _38009_;
  wire _38010_;
  wire _38011_;
  wire _38012_;
  wire _38013_;
  wire _38014_;
  wire _38015_;
  wire _38016_;
  wire _38017_;
  wire _38018_;
  wire _38019_;
  wire _38020_;
  wire _38021_;
  wire _38022_;
  wire _38023_;
  wire _38024_;
  wire _38025_;
  wire _38026_;
  wire _38027_;
  wire _38028_;
  wire _38029_;
  wire _38030_;
  wire _38031_;
  wire _38032_;
  wire _38033_;
  wire _38034_;
  wire _38035_;
  wire _38036_;
  wire _38037_;
  wire _38038_;
  wire _38039_;
  wire _38040_;
  wire _38041_;
  wire _38042_;
  wire _38043_;
  wire _38044_;
  wire _38045_;
  wire _38046_;
  wire _38047_;
  wire _38048_;
  wire _38049_;
  wire _38050_;
  wire _38051_;
  wire _38052_;
  wire _38053_;
  wire _38054_;
  wire _38055_;
  wire _38056_;
  wire _38057_;
  wire _38058_;
  wire _38059_;
  wire _38060_;
  wire _38061_;
  wire _38062_;
  wire _38063_;
  wire _38064_;
  wire _38065_;
  wire _38066_;
  wire _38067_;
  wire _38068_;
  wire _38069_;
  wire _38070_;
  wire _38071_;
  wire _38072_;
  wire _38073_;
  wire _38074_;
  wire _38075_;
  wire _38076_;
  wire _38077_;
  wire _38078_;
  wire _38079_;
  wire _38080_;
  wire _38081_;
  wire _38082_;
  wire _38083_;
  wire _38084_;
  wire _38085_;
  wire _38086_;
  wire _38087_;
  wire _38088_;
  wire _38089_;
  wire _38090_;
  wire _38091_;
  wire _38092_;
  wire _38093_;
  wire _38094_;
  wire _38095_;
  wire _38096_;
  wire _38097_;
  wire _38098_;
  wire _38099_;
  wire _38100_;
  wire _38101_;
  wire _38102_;
  wire _38103_;
  wire _38104_;
  wire _38105_;
  wire _38106_;
  wire _38107_;
  wire _38108_;
  wire _38109_;
  wire _38110_;
  wire _38111_;
  wire _38112_;
  wire _38113_;
  wire _38114_;
  wire _38115_;
  wire _38116_;
  wire _38117_;
  wire _38118_;
  wire _38119_;
  wire _38120_;
  wire _38121_;
  wire _38122_;
  wire _38123_;
  wire _38124_;
  wire _38125_;
  wire _38126_;
  wire _38127_;
  wire _38128_;
  wire _38129_;
  wire _38130_;
  wire _38131_;
  wire _38132_;
  wire _38133_;
  wire _38134_;
  wire _38135_;
  wire _38136_;
  wire _38137_;
  wire _38138_;
  wire _38139_;
  wire _38140_;
  wire _38141_;
  wire _38142_;
  wire _38143_;
  wire _38144_;
  wire _38145_;
  wire _38146_;
  wire _38147_;
  wire _38148_;
  wire _38149_;
  wire _38150_;
  wire _38151_;
  wire _38152_;
  wire _38153_;
  wire _38154_;
  wire _38155_;
  wire _38156_;
  wire _38157_;
  wire _38158_;
  wire _38159_;
  wire _38160_;
  wire _38161_;
  wire _38162_;
  wire _38163_;
  wire _38164_;
  wire _38165_;
  wire _38166_;
  wire _38167_;
  wire _38168_;
  wire _38169_;
  wire _38170_;
  wire _38171_;
  wire _38172_;
  wire _38173_;
  wire _38174_;
  wire _38175_;
  wire _38176_;
  wire _38177_;
  wire _38178_;
  wire _38179_;
  wire _38180_;
  wire _38181_;
  wire _38182_;
  wire _38183_;
  wire _38184_;
  wire _38185_;
  wire _38186_;
  wire _38187_;
  wire _38188_;
  wire _38189_;
  wire _38190_;
  wire _38191_;
  wire _38192_;
  wire _38193_;
  wire _38194_;
  wire _38195_;
  wire _38196_;
  wire _38197_;
  wire _38198_;
  wire _38199_;
  wire _38200_;
  wire _38201_;
  wire _38202_;
  wire _38203_;
  wire _38204_;
  wire _38205_;
  wire _38206_;
  wire _38207_;
  wire _38208_;
  wire _38209_;
  wire _38210_;
  wire _38211_;
  wire _38212_;
  wire _38213_;
  wire _38214_;
  wire _38215_;
  wire _38216_;
  wire _38217_;
  wire _38218_;
  wire _38219_;
  wire _38220_;
  wire _38221_;
  wire _38222_;
  wire _38223_;
  wire _38224_;
  wire _38225_;
  wire _38226_;
  wire _38227_;
  wire _38228_;
  wire _38229_;
  wire _38230_;
  wire _38231_;
  wire _38232_;
  wire _38233_;
  wire _38234_;
  wire _38235_;
  wire _38236_;
  wire _38237_;
  wire _38238_;
  wire _38239_;
  wire _38240_;
  wire _38241_;
  wire _38242_;
  wire _38243_;
  wire _38244_;
  wire _38245_;
  wire _38246_;
  wire _38247_;
  wire _38248_;
  wire _38249_;
  wire _38250_;
  wire _38251_;
  wire _38252_;
  wire _38253_;
  wire _38254_;
  wire _38255_;
  wire _38256_;
  wire _38257_;
  wire _38258_;
  wire _38259_;
  wire _38260_;
  wire _38261_;
  wire _38262_;
  wire _38263_;
  wire _38264_;
  wire _38265_;
  wire _38266_;
  wire _38267_;
  wire _38268_;
  wire _38269_;
  wire _38270_;
  wire _38271_;
  wire _38272_;
  wire _38273_;
  wire _38274_;
  wire _38275_;
  wire _38276_;
  wire _38277_;
  wire _38278_;
  wire _38279_;
  wire _38280_;
  wire _38281_;
  wire _38282_;
  wire _38283_;
  wire _38284_;
  wire _38285_;
  wire _38286_;
  wire _38287_;
  wire _38288_;
  wire _38289_;
  wire _38290_;
  wire _38291_;
  wire _38292_;
  wire _38293_;
  wire _38294_;
  wire _38295_;
  wire _38296_;
  wire _38297_;
  wire _38298_;
  wire _38299_;
  wire _38300_;
  wire _38301_;
  wire _38302_;
  wire _38303_;
  wire _38304_;
  wire _38305_;
  wire _38306_;
  wire _38307_;
  wire _38308_;
  wire _38309_;
  wire _38310_;
  wire _38311_;
  wire _38312_;
  wire _38313_;
  wire _38314_;
  wire _38315_;
  wire _38316_;
  wire _38317_;
  wire _38318_;
  wire _38319_;
  wire _38320_;
  wire _38321_;
  wire _38322_;
  wire _38323_;
  wire _38324_;
  wire _38325_;
  wire _38326_;
  wire _38327_;
  wire _38328_;
  wire _38329_;
  wire _38330_;
  wire _38331_;
  wire _38332_;
  wire _38333_;
  wire _38334_;
  wire _38335_;
  wire _38336_;
  wire _38337_;
  wire _38338_;
  wire _38339_;
  wire _38340_;
  wire _38341_;
  wire _38342_;
  wire _38343_;
  wire _38344_;
  wire _38345_;
  wire _38346_;
  wire _38347_;
  wire _38348_;
  wire _38349_;
  wire _38350_;
  wire _38351_;
  wire _38352_;
  wire _38353_;
  wire _38354_;
  wire _38355_;
  wire _38356_;
  wire _38357_;
  wire _38358_;
  wire _38359_;
  wire _38360_;
  wire _38361_;
  wire _38362_;
  wire _38363_;
  wire _38364_;
  wire _38365_;
  wire _38366_;
  wire _38367_;
  wire _38368_;
  wire _38369_;
  wire _38370_;
  wire _38371_;
  wire _38372_;
  wire _38373_;
  wire _38374_;
  wire _38375_;
  wire _38376_;
  wire _38377_;
  wire _38378_;
  wire _38379_;
  wire _38380_;
  wire _38381_;
  wire _38382_;
  wire _38383_;
  wire _38384_;
  wire _38385_;
  wire _38386_;
  wire _38387_;
  wire _38388_;
  wire _38389_;
  wire _38390_;
  wire _38391_;
  wire _38392_;
  wire _38393_;
  wire _38394_;
  wire _38395_;
  wire _38396_;
  wire _38397_;
  wire _38398_;
  wire _38399_;
  wire _38400_;
  wire _38401_;
  wire _38402_;
  wire _38403_;
  wire _38404_;
  wire _38405_;
  wire _38406_;
  wire _38407_;
  wire _38408_;
  wire _38409_;
  wire _38410_;
  wire _38411_;
  wire _38412_;
  wire _38413_;
  wire _38414_;
  wire _38415_;
  wire _38416_;
  wire _38417_;
  wire _38418_;
  wire _38419_;
  wire _38420_;
  wire _38421_;
  wire _38422_;
  wire _38423_;
  wire _38424_;
  wire _38425_;
  wire _38426_;
  wire _38427_;
  wire _38428_;
  wire _38429_;
  wire _38430_;
  wire _38431_;
  wire _38432_;
  wire _38433_;
  wire _38434_;
  wire _38435_;
  wire _38436_;
  wire _38437_;
  wire _38438_;
  wire _38439_;
  wire _38440_;
  wire _38441_;
  wire _38442_;
  wire _38443_;
  wire _38444_;
  wire _38445_;
  wire _38446_;
  wire _38447_;
  wire _38448_;
  wire _38449_;
  wire _38450_;
  wire _38451_;
  wire _38452_;
  wire _38453_;
  wire _38454_;
  wire _38455_;
  wire _38456_;
  wire _38457_;
  wire _38458_;
  wire _38459_;
  wire _38460_;
  wire _38461_;
  wire _38462_;
  wire _38463_;
  wire _38464_;
  wire _38465_;
  wire _38466_;
  wire _38467_;
  wire _38468_;
  wire _38469_;
  wire _38470_;
  wire _38471_;
  wire _38472_;
  wire _38473_;
  wire _38474_;
  wire _38475_;
  wire _38476_;
  wire _38477_;
  wire _38478_;
  wire _38479_;
  wire _38480_;
  wire _38481_;
  wire _38482_;
  wire _38483_;
  wire _38484_;
  wire _38485_;
  wire _38486_;
  wire _38487_;
  wire _38488_;
  wire _38489_;
  wire _38490_;
  wire _38491_;
  wire _38492_;
  wire _38493_;
  wire _38494_;
  wire _38495_;
  wire _38496_;
  wire _38497_;
  wire _38498_;
  wire _38499_;
  wire _38500_;
  wire _38501_;
  wire _38502_;
  wire _38503_;
  wire _38504_;
  wire _38505_;
  wire _38506_;
  wire _38507_;
  wire _38508_;
  wire _38509_;
  wire _38510_;
  wire _38511_;
  wire _38512_;
  wire _38513_;
  wire _38514_;
  wire _38515_;
  wire _38516_;
  wire _38517_;
  wire _38518_;
  wire _38519_;
  wire _38520_;
  wire _38521_;
  wire _38522_;
  wire _38523_;
  wire _38524_;
  wire _38525_;
  wire _38526_;
  wire _38527_;
  wire _38528_;
  wire _38529_;
  wire _38530_;
  wire _38531_;
  wire _38532_;
  wire _38533_;
  wire _38534_;
  wire _38535_;
  wire _38536_;
  wire _38537_;
  wire _38538_;
  wire _38539_;
  wire _38540_;
  wire _38541_;
  wire _38542_;
  wire _38543_;
  wire _38544_;
  wire _38545_;
  wire _38546_;
  wire _38547_;
  wire _38548_;
  wire _38549_;
  wire _38550_;
  wire _38551_;
  wire _38552_;
  wire _38553_;
  wire _38554_;
  wire _38555_;
  wire _38556_;
  wire _38557_;
  wire _38558_;
  wire _38559_;
  wire _38560_;
  wire _38561_;
  wire _38562_;
  wire _38563_;
  wire _38564_;
  wire _38565_;
  wire _38566_;
  wire _38567_;
  wire _38568_;
  wire _38569_;
  wire _38570_;
  wire _38571_;
  wire _38572_;
  wire _38573_;
  wire _38574_;
  wire _38575_;
  wire _38576_;
  wire _38577_;
  wire _38578_;
  wire _38579_;
  wire _38580_;
  wire _38581_;
  wire _38582_;
  wire _38583_;
  wire _38584_;
  wire _38585_;
  wire _38586_;
  wire _38587_;
  wire _38588_;
  wire _38589_;
  wire _38590_;
  wire _38591_;
  wire _38592_;
  wire _38593_;
  wire _38594_;
  wire _38595_;
  wire _38596_;
  wire _38597_;
  wire _38598_;
  wire _38599_;
  wire _38600_;
  wire _38601_;
  wire _38602_;
  wire _38603_;
  wire _38604_;
  wire _38605_;
  wire _38606_;
  wire _38607_;
  wire _38608_;
  wire _38609_;
  wire _38610_;
  wire _38611_;
  wire _38612_;
  wire _38613_;
  wire _38614_;
  wire _38615_;
  wire _38616_;
  wire _38617_;
  wire _38618_;
  wire _38619_;
  wire _38620_;
  wire _38621_;
  wire _38622_;
  wire _38623_;
  wire _38624_;
  wire _38625_;
  wire _38626_;
  wire _38627_;
  wire _38628_;
  wire _38629_;
  wire _38630_;
  wire _38631_;
  wire _38632_;
  wire _38633_;
  wire _38634_;
  wire _38635_;
  wire _38636_;
  wire _38637_;
  wire _38638_;
  wire _38639_;
  wire _38640_;
  wire _38641_;
  wire _38642_;
  wire _38643_;
  wire _38644_;
  wire _38645_;
  wire _38646_;
  wire _38647_;
  wire _38648_;
  wire _38649_;
  wire _38650_;
  wire _38651_;
  wire _38652_;
  wire _38653_;
  wire _38654_;
  wire _38655_;
  wire _38656_;
  wire _38657_;
  wire _38658_;
  wire _38659_;
  wire _38660_;
  wire _38661_;
  wire _38662_;
  wire _38663_;
  wire _38664_;
  wire _38665_;
  wire _38666_;
  wire _38667_;
  wire _38668_;
  wire _38669_;
  wire _38670_;
  wire _38671_;
  wire _38672_;
  wire _38673_;
  wire _38674_;
  wire _38675_;
  wire _38676_;
  wire _38677_;
  wire _38678_;
  wire _38679_;
  wire _38680_;
  wire _38681_;
  wire _38682_;
  wire _38683_;
  wire _38684_;
  wire _38685_;
  wire _38686_;
  wire _38687_;
  wire _38688_;
  wire _38689_;
  wire _38690_;
  wire _38691_;
  wire _38692_;
  wire _38693_;
  wire _38694_;
  wire _38695_;
  wire _38696_;
  wire _38697_;
  wire _38698_;
  wire _38699_;
  wire _38700_;
  wire _38701_;
  wire _38702_;
  wire _38703_;
  wire _38704_;
  wire _38705_;
  wire _38706_;
  wire _38707_;
  wire _38708_;
  wire _38709_;
  wire _38710_;
  wire _38711_;
  wire _38712_;
  wire _38713_;
  wire _38714_;
  wire _38715_;
  wire _38716_;
  wire _38717_;
  wire _38718_;
  wire _38719_;
  wire _38720_;
  wire _38721_;
  wire _38722_;
  wire _38723_;
  wire _38724_;
  wire _38725_;
  wire _38726_;
  wire _38727_;
  wire _38728_;
  wire _38729_;
  wire _38730_;
  wire _38731_;
  wire _38732_;
  wire _38733_;
  wire _38734_;
  wire _38735_;
  wire _38736_;
  wire _38737_;
  wire _38738_;
  wire _38739_;
  wire _38740_;
  wire _38741_;
  wire _38742_;
  wire _38743_;
  wire _38744_;
  wire _38745_;
  wire _38746_;
  wire _38747_;
  wire _38748_;
  wire _38749_;
  wire _38750_;
  wire _38751_;
  wire _38752_;
  wire _38753_;
  wire _38754_;
  wire _38755_;
  wire _38756_;
  wire _38757_;
  wire _38758_;
  wire _38759_;
  wire _38760_;
  wire _38761_;
  wire _38762_;
  wire _38763_;
  wire _38764_;
  wire _38765_;
  wire _38766_;
  wire _38767_;
  wire _38768_;
  wire _38769_;
  wire _38770_;
  wire _38771_;
  wire _38772_;
  wire _38773_;
  wire _38774_;
  wire _38775_;
  wire _38776_;
  wire _38777_;
  wire _38778_;
  wire _38779_;
  wire _38780_;
  wire _38781_;
  wire _38782_;
  wire _38783_;
  wire _38784_;
  wire _38785_;
  wire _38786_;
  wire _38787_;
  wire _38788_;
  wire _38789_;
  wire _38790_;
  wire _38791_;
  wire _38792_;
  wire _38793_;
  wire _38794_;
  wire _38795_;
  wire _38796_;
  wire _38797_;
  wire _38798_;
  wire _38799_;
  wire _38800_;
  wire _38801_;
  wire _38802_;
  wire _38803_;
  wire _38804_;
  wire _38805_;
  wire _38806_;
  wire _38807_;
  wire _38808_;
  wire _38809_;
  wire _38810_;
  wire _38811_;
  wire _38812_;
  wire _38813_;
  wire _38814_;
  wire _38815_;
  wire _38816_;
  wire _38817_;
  wire _38818_;
  wire _38819_;
  wire _38820_;
  wire _38821_;
  wire _38822_;
  wire _38823_;
  wire _38824_;
  wire _38825_;
  wire _38826_;
  wire _38827_;
  wire _38828_;
  wire _38829_;
  wire _38830_;
  wire _38831_;
  wire _38832_;
  wire _38833_;
  wire _38834_;
  wire _38835_;
  wire _38836_;
  wire _38837_;
  wire _38838_;
  wire _38839_;
  wire _38840_;
  wire _38841_;
  wire _38842_;
  wire _38843_;
  wire _38844_;
  wire _38845_;
  wire _38846_;
  wire _38847_;
  wire _38848_;
  wire _38849_;
  wire _38850_;
  wire _38851_;
  wire _38852_;
  wire _38853_;
  wire _38854_;
  wire _38855_;
  wire _38856_;
  wire _38857_;
  wire _38858_;
  wire _38859_;
  wire _38860_;
  wire _38861_;
  wire _38862_;
  wire _38863_;
  wire _38864_;
  wire _38865_;
  wire _38866_;
  wire _38867_;
  wire _38868_;
  wire _38869_;
  wire _38870_;
  wire _38871_;
  wire _38872_;
  wire _38873_;
  wire _38874_;
  wire _38875_;
  wire _38876_;
  wire _38877_;
  wire _38878_;
  wire _38879_;
  wire _38880_;
  wire _38881_;
  wire _38882_;
  wire _38883_;
  wire _38884_;
  wire _38885_;
  wire _38886_;
  wire _38887_;
  wire _38888_;
  wire _38889_;
  wire _38890_;
  wire _38891_;
  wire _38892_;
  wire _38893_;
  wire _38894_;
  wire _38895_;
  wire _38896_;
  wire _38897_;
  wire _38898_;
  wire _38899_;
  wire _38900_;
  wire _38901_;
  wire _38902_;
  wire _38903_;
  wire _38904_;
  wire _38905_;
  wire _38906_;
  wire _38907_;
  wire _38908_;
  wire _38909_;
  wire _38910_;
  wire _38911_;
  wire _38912_;
  wire _38913_;
  wire _38914_;
  wire _38915_;
  wire _38916_;
  wire _38917_;
  wire _38918_;
  wire _38919_;
  wire _38920_;
  wire _38921_;
  wire _38922_;
  wire _38923_;
  wire _38924_;
  wire _38925_;
  wire _38926_;
  wire _38927_;
  wire _38928_;
  wire _38929_;
  wire _38930_;
  wire _38931_;
  wire _38932_;
  wire _38933_;
  wire _38934_;
  wire _38935_;
  wire _38936_;
  wire _38937_;
  wire _38938_;
  wire _38939_;
  wire _38940_;
  wire _38941_;
  wire _38942_;
  wire _38943_;
  wire _38944_;
  wire _38945_;
  wire _38946_;
  wire _38947_;
  wire _38948_;
  wire _38949_;
  wire _38950_;
  wire _38951_;
  wire _38952_;
  wire _38953_;
  wire _38954_;
  wire _38955_;
  wire _38956_;
  wire _38957_;
  wire _38958_;
  wire _38959_;
  wire _38960_;
  wire _38961_;
  wire _38962_;
  wire _38963_;
  wire _38964_;
  wire _38965_;
  wire _38966_;
  wire _38967_;
  wire _38968_;
  wire _38969_;
  wire _38970_;
  wire _38971_;
  wire _38972_;
  wire _38973_;
  wire _38974_;
  wire _38975_;
  wire _38976_;
  wire _38977_;
  wire _38978_;
  wire _38979_;
  wire _38980_;
  wire _38981_;
  wire _38982_;
  wire _38983_;
  wire _38984_;
  wire _38985_;
  wire _38986_;
  wire _38987_;
  wire _38988_;
  wire _38989_;
  wire _38990_;
  wire _38991_;
  wire _38992_;
  wire _38993_;
  wire _38994_;
  wire _38995_;
  wire _38996_;
  wire _38997_;
  wire _38998_;
  wire _38999_;
  wire _39000_;
  wire _39001_;
  wire _39002_;
  wire _39003_;
  wire _39004_;
  wire _39005_;
  wire _39006_;
  wire _39007_;
  wire _39008_;
  wire _39009_;
  wire _39010_;
  wire _39011_;
  wire _39012_;
  wire _39013_;
  wire _39014_;
  wire _39015_;
  wire _39016_;
  wire _39017_;
  wire _39018_;
  wire _39019_;
  wire _39020_;
  wire _39021_;
  wire _39022_;
  wire _39023_;
  wire _39024_;
  wire _39025_;
  wire _39026_;
  wire _39027_;
  wire _39028_;
  wire _39029_;
  wire _39030_;
  wire _39031_;
  wire _39032_;
  wire _39033_;
  wire _39034_;
  wire _39035_;
  wire _39036_;
  wire _39037_;
  wire _39038_;
  wire _39039_;
  wire _39040_;
  wire _39041_;
  wire _39042_;
  wire _39043_;
  wire _39044_;
  wire _39045_;
  wire _39046_;
  wire _39047_;
  wire _39048_;
  wire _39049_;
  wire _39050_;
  wire _39051_;
  wire _39052_;
  wire _39053_;
  wire _39054_;
  wire _39055_;
  wire _39056_;
  wire _39057_;
  wire _39058_;
  wire _39059_;
  wire _39060_;
  wire _39061_;
  wire _39062_;
  wire _39063_;
  wire _39064_;
  wire _39065_;
  wire _39066_;
  wire _39067_;
  wire _39068_;
  wire _39069_;
  wire _39070_;
  wire _39071_;
  wire _39072_;
  wire _39073_;
  wire _39074_;
  wire _39075_;
  wire _39076_;
  wire _39077_;
  wire _39078_;
  wire _39079_;
  wire _39080_;
  wire _39081_;
  wire _39082_;
  wire _39083_;
  wire _39084_;
  wire _39085_;
  wire _39086_;
  wire _39087_;
  wire _39088_;
  wire _39089_;
  wire _39090_;
  wire _39091_;
  wire _39092_;
  wire _39093_;
  wire _39094_;
  wire _39095_;
  wire _39096_;
  wire _39097_;
  wire _39098_;
  wire _39099_;
  wire _39100_;
  wire _39101_;
  wire _39102_;
  wire _39103_;
  wire _39104_;
  wire _39105_;
  wire _39106_;
  wire _39107_;
  wire _39108_;
  wire _39109_;
  wire _39110_;
  wire _39111_;
  wire _39112_;
  wire _39113_;
  wire _39114_;
  wire _39115_;
  wire _39116_;
  wire _39117_;
  wire _39118_;
  wire _39119_;
  wire _39120_;
  wire _39121_;
  wire _39122_;
  wire _39123_;
  wire _39124_;
  wire _39125_;
  wire _39126_;
  wire _39127_;
  wire _39128_;
  wire _39129_;
  wire _39130_;
  wire _39131_;
  wire _39132_;
  wire _39133_;
  wire _39134_;
  wire _39135_;
  wire _39136_;
  wire _39137_;
  wire _39138_;
  wire _39139_;
  wire _39140_;
  wire _39141_;
  wire _39142_;
  wire _39143_;
  wire _39144_;
  wire _39145_;
  wire _39146_;
  wire _39147_;
  wire _39148_;
  wire _39149_;
  wire _39150_;
  wire _39151_;
  wire _39152_;
  wire _39153_;
  wire _39154_;
  wire _39155_;
  wire _39156_;
  wire _39157_;
  wire _39158_;
  wire _39159_;
  wire _39160_;
  wire _39161_;
  wire _39162_;
  wire _39163_;
  wire _39164_;
  wire _39165_;
  wire _39166_;
  wire _39167_;
  wire _39168_;
  wire _39169_;
  wire _39170_;
  wire _39171_;
  wire _39172_;
  wire _39173_;
  wire _39174_;
  wire _39175_;
  wire _39176_;
  wire _39177_;
  wire _39178_;
  wire _39179_;
  wire _39180_;
  wire _39181_;
  wire _39182_;
  wire _39183_;
  wire _39184_;
  wire _39185_;
  wire _39186_;
  wire _39187_;
  wire _39188_;
  wire _39189_;
  wire _39190_;
  wire _39191_;
  wire _39192_;
  wire _39193_;
  wire _39194_;
  wire _39195_;
  wire _39196_;
  wire _39197_;
  wire _39198_;
  wire _39199_;
  wire _39200_;
  wire _39201_;
  wire _39202_;
  wire _39203_;
  wire _39204_;
  wire _39205_;
  wire _39206_;
  wire _39207_;
  wire _39208_;
  wire _39209_;
  wire _39210_;
  wire _39211_;
  wire _39212_;
  wire _39213_;
  wire _39214_;
  wire _39215_;
  wire _39216_;
  wire _39217_;
  wire _39218_;
  wire _39219_;
  wire _39220_;
  wire _39221_;
  wire _39222_;
  wire _39223_;
  wire _39224_;
  wire _39225_;
  wire _39226_;
  wire _39227_;
  wire _39228_;
  wire _39229_;
  wire _39230_;
  wire _39231_;
  wire _39232_;
  wire _39233_;
  wire _39234_;
  wire _39235_;
  wire _39236_;
  wire _39237_;
  wire _39238_;
  wire _39239_;
  wire _39240_;
  wire _39241_;
  wire _39242_;
  wire _39243_;
  wire _39244_;
  wire _39245_;
  wire _39246_;
  wire _39247_;
  wire _39248_;
  wire _39249_;
  wire _39250_;
  wire _39251_;
  wire _39252_;
  wire _39253_;
  wire _39254_;
  wire _39255_;
  wire _39256_;
  wire _39257_;
  wire _39258_;
  wire _39259_;
  wire _39260_;
  wire _39261_;
  wire _39262_;
  wire _39263_;
  wire _39264_;
  wire _39265_;
  wire _39266_;
  wire _39267_;
  wire _39268_;
  wire _39269_;
  wire _39270_;
  wire _39271_;
  wire _39272_;
  wire _39273_;
  wire _39274_;
  wire _39275_;
  wire _39276_;
  wire _39277_;
  wire _39278_;
  wire _39279_;
  wire _39280_;
  wire _39281_;
  wire _39282_;
  wire _39283_;
  wire _39284_;
  wire _39285_;
  wire _39286_;
  wire _39287_;
  wire _39288_;
  wire _39289_;
  wire _39290_;
  wire _39291_;
  wire _39292_;
  wire _39293_;
  wire _39294_;
  wire _39295_;
  wire _39296_;
  wire _39297_;
  wire _39298_;
  wire _39299_;
  wire _39300_;
  wire _39301_;
  wire _39302_;
  wire _39303_;
  wire _39304_;
  wire _39305_;
  wire _39306_;
  wire _39307_;
  wire _39308_;
  wire _39309_;
  wire _39310_;
  wire _39311_;
  wire _39312_;
  wire _39313_;
  wire _39314_;
  wire _39315_;
  wire _39316_;
  wire _39317_;
  wire _39318_;
  wire _39319_;
  wire _39320_;
  wire _39321_;
  wire _39322_;
  wire _39323_;
  wire _39324_;
  wire _39325_;
  wire _39326_;
  wire _39327_;
  wire _39328_;
  wire _39329_;
  wire _39330_;
  wire _39331_;
  wire _39332_;
  wire _39333_;
  wire _39334_;
  wire _39335_;
  wire _39336_;
  wire _39337_;
  wire _39338_;
  wire _39339_;
  wire _39340_;
  wire _39341_;
  wire _39342_;
  wire _39343_;
  wire _39344_;
  wire _39345_;
  wire _39346_;
  wire _39347_;
  wire _39348_;
  wire _39349_;
  wire _39350_;
  wire _39351_;
  wire _39352_;
  wire _39353_;
  wire _39354_;
  wire _39355_;
  wire _39356_;
  wire _39357_;
  wire _39358_;
  wire _39359_;
  wire _39360_;
  wire _39361_;
  wire _39362_;
  wire _39363_;
  wire _39364_;
  wire _39365_;
  wire _39366_;
  wire _39367_;
  wire _39368_;
  wire _39369_;
  wire _39370_;
  wire _39371_;
  wire _39372_;
  wire _39373_;
  wire _39374_;
  wire _39375_;
  wire _39376_;
  wire _39377_;
  wire _39378_;
  wire _39379_;
  wire _39380_;
  wire _39381_;
  wire _39382_;
  wire _39383_;
  wire _39384_;
  wire _39385_;
  wire _39386_;
  wire _39387_;
  wire _39388_;
  wire _39389_;
  wire _39390_;
  wire _39391_;
  wire _39392_;
  wire _39393_;
  wire _39394_;
  wire _39395_;
  wire _39396_;
  wire _39397_;
  wire _39398_;
  wire _39399_;
  wire _39400_;
  wire _39401_;
  wire _39402_;
  wire _39403_;
  wire _39404_;
  wire _39405_;
  wire _39406_;
  wire _39407_;
  wire _39408_;
  wire _39409_;
  wire _39410_;
  wire _39411_;
  wire _39412_;
  wire _39413_;
  wire _39414_;
  wire _39415_;
  wire _39416_;
  wire _39417_;
  wire _39418_;
  wire _39419_;
  wire _39420_;
  wire _39421_;
  wire _39422_;
  wire _39423_;
  wire _39424_;
  wire _39425_;
  wire _39426_;
  wire _39427_;
  wire _39428_;
  wire _39429_;
  wire _39430_;
  wire _39431_;
  wire _39432_;
  wire _39433_;
  wire _39434_;
  wire _39435_;
  wire _39436_;
  wire _39437_;
  wire _39438_;
  wire _39439_;
  wire _39440_;
  wire _39441_;
  wire _39442_;
  wire _39443_;
  wire _39444_;
  wire _39445_;
  wire _39446_;
  wire _39447_;
  wire _39448_;
  wire _39449_;
  wire _39450_;
  wire _39451_;
  wire _39452_;
  wire _39453_;
  wire _39454_;
  wire _39455_;
  wire _39456_;
  wire _39457_;
  wire _39458_;
  wire _39459_;
  wire _39460_;
  wire _39461_;
  wire _39462_;
  wire _39463_;
  wire _39464_;
  wire _39465_;
  wire _39466_;
  wire _39467_;
  wire _39468_;
  wire _39469_;
  wire _39470_;
  wire _39471_;
  wire _39472_;
  wire _39473_;
  wire _39474_;
  wire _39475_;
  wire _39476_;
  wire _39477_;
  wire _39478_;
  wire _39479_;
  wire _39480_;
  wire _39481_;
  wire _39482_;
  wire _39483_;
  wire _39484_;
  wire _39485_;
  wire _39486_;
  wire _39487_;
  wire _39488_;
  wire _39489_;
  wire _39490_;
  wire _39491_;
  wire _39492_;
  wire _39493_;
  wire _39494_;
  wire _39495_;
  wire _39496_;
  wire _39497_;
  wire _39498_;
  wire _39499_;
  wire _39500_;
  wire _39501_;
  wire _39502_;
  wire _39503_;
  wire _39504_;
  wire _39505_;
  wire _39506_;
  wire _39507_;
  wire _39508_;
  wire _39509_;
  wire _39510_;
  wire _39511_;
  wire _39512_;
  wire _39513_;
  wire _39514_;
  wire _39515_;
  wire _39516_;
  wire _39517_;
  wire _39518_;
  wire _39519_;
  wire _39520_;
  wire _39521_;
  wire _39522_;
  wire _39523_;
  wire _39524_;
  wire _39525_;
  wire _39526_;
  wire _39527_;
  wire _39528_;
  wire _39529_;
  wire _39530_;
  wire _39531_;
  wire _39532_;
  wire _39533_;
  wire _39534_;
  wire _39535_;
  wire _39536_;
  wire _39537_;
  wire _39538_;
  wire _39539_;
  wire _39540_;
  wire _39541_;
  wire _39542_;
  wire _39543_;
  wire _39544_;
  wire _39545_;
  wire _39546_;
  wire _39547_;
  wire _39548_;
  wire _39549_;
  wire _39550_;
  wire _39551_;
  wire _39552_;
  wire _39553_;
  wire _39554_;
  wire _39555_;
  wire _39556_;
  wire _39557_;
  wire _39558_;
  wire _39559_;
  wire _39560_;
  wire _39561_;
  wire _39562_;
  wire _39563_;
  wire _39564_;
  wire _39565_;
  wire _39566_;
  wire _39567_;
  wire _39568_;
  wire _39569_;
  wire _39570_;
  wire _39571_;
  wire _39572_;
  wire _39573_;
  wire _39574_;
  wire _39575_;
  wire _39576_;
  wire _39577_;
  wire _39578_;
  wire _39579_;
  wire _39580_;
  wire _39581_;
  wire _39582_;
  wire _39583_;
  wire _39584_;
  wire _39585_;
  wire _39586_;
  wire _39587_;
  wire _39588_;
  wire _39589_;
  wire _39590_;
  wire _39591_;
  wire _39592_;
  wire _39593_;
  wire _39594_;
  wire _39595_;
  wire _39596_;
  wire _39597_;
  wire _39598_;
  wire _39599_;
  wire _39600_;
  wire _39601_;
  wire _39602_;
  wire _39603_;
  wire _39604_;
  wire _39605_;
  wire _39606_;
  wire _39607_;
  wire _39608_;
  wire _39609_;
  wire _39610_;
  wire _39611_;
  wire _39612_;
  wire _39613_;
  wire _39614_;
  wire _39615_;
  wire _39616_;
  wire _39617_;
  wire _39618_;
  wire _39619_;
  wire _39620_;
  wire _39621_;
  wire _39622_;
  wire _39623_;
  wire _39624_;
  wire _39625_;
  wire _39626_;
  wire _39627_;
  wire _39628_;
  wire _39629_;
  wire _39630_;
  wire _39631_;
  wire _39632_;
  wire _39633_;
  wire _39634_;
  wire _39635_;
  wire _39636_;
  wire _39637_;
  wire _39638_;
  wire _39639_;
  wire _39640_;
  wire _39641_;
  wire _39642_;
  wire _39643_;
  wire _39644_;
  wire _39645_;
  wire _39646_;
  wire _39647_;
  wire _39648_;
  wire _39649_;
  wire _39650_;
  wire _39651_;
  wire _39652_;
  wire _39653_;
  wire _39654_;
  wire _39655_;
  wire _39656_;
  wire _39657_;
  wire _39658_;
  wire _39659_;
  wire _39660_;
  wire _39661_;
  wire _39662_;
  wire _39663_;
  wire _39664_;
  wire _39665_;
  wire _39666_;
  wire _39667_;
  wire _39668_;
  wire _39669_;
  wire _39670_;
  wire _39671_;
  wire _39672_;
  wire _39673_;
  wire _39674_;
  wire _39675_;
  wire _39676_;
  wire _39677_;
  wire _39678_;
  wire _39679_;
  wire _39680_;
  wire _39681_;
  wire _39682_;
  wire _39683_;
  wire _39684_;
  wire _39685_;
  wire _39686_;
  wire _39687_;
  wire _39688_;
  wire _39689_;
  wire _39690_;
  wire _39691_;
  wire _39692_;
  wire _39693_;
  wire _39694_;
  wire _39695_;
  wire _39696_;
  wire _39697_;
  wire _39698_;
  wire _39699_;
  wire _39700_;
  wire _39701_;
  wire _39702_;
  wire _39703_;
  wire _39704_;
  wire _39705_;
  wire _39706_;
  wire _39707_;
  wire _39708_;
  wire _39709_;
  wire _39710_;
  wire _39711_;
  wire _39712_;
  wire _39713_;
  wire _39714_;
  wire _39715_;
  wire _39716_;
  wire _39717_;
  wire _39718_;
  wire _39719_;
  wire _39720_;
  wire _39721_;
  wire _39722_;
  wire _39723_;
  wire _39724_;
  wire _39725_;
  wire _39726_;
  wire _39727_;
  wire _39728_;
  wire _39729_;
  wire _39730_;
  wire _39731_;
  wire _39732_;
  wire _39733_;
  wire _39734_;
  wire _39735_;
  wire _39736_;
  wire _39737_;
  wire _39738_;
  wire _39739_;
  wire _39740_;
  wire _39741_;
  wire _39742_;
  wire _39743_;
  wire _39744_;
  wire _39745_;
  wire _39746_;
  wire _39747_;
  wire _39748_;
  wire _39749_;
  wire _39750_;
  wire _39751_;
  wire _39752_;
  wire _39753_;
  wire _39754_;
  wire _39755_;
  wire _39756_;
  wire _39757_;
  wire _39758_;
  wire _39759_;
  wire _39760_;
  wire _39761_;
  wire _39762_;
  wire _39763_;
  wire _39764_;
  wire _39765_;
  wire _39766_;
  wire _39767_;
  wire _39768_;
  wire _39769_;
  wire _39770_;
  wire _39771_;
  wire _39772_;
  wire _39773_;
  wire _39774_;
  wire _39775_;
  wire _39776_;
  wire _39777_;
  wire _39778_;
  wire _39779_;
  wire _39780_;
  wire _39781_;
  wire _39782_;
  wire _39783_;
  wire _39784_;
  wire _39785_;
  wire _39786_;
  wire _39787_;
  wire _39788_;
  wire _39789_;
  wire _39790_;
  wire _39791_;
  wire _39792_;
  wire _39793_;
  wire _39794_;
  wire _39795_;
  wire _39796_;
  wire _39797_;
  wire _39798_;
  wire _39799_;
  wire _39800_;
  wire _39801_;
  wire _39802_;
  wire _39803_;
  wire _39804_;
  wire _39805_;
  wire _39806_;
  wire _39807_;
  wire _39808_;
  wire _39809_;
  wire _39810_;
  wire _39811_;
  wire _39812_;
  wire _39813_;
  wire _39814_;
  wire _39815_;
  wire _39816_;
  wire _39817_;
  wire _39818_;
  wire _39819_;
  wire _39820_;
  wire _39821_;
  wire _39822_;
  wire _39823_;
  wire _39824_;
  wire _39825_;
  wire _39826_;
  wire _39827_;
  wire _39828_;
  wire _39829_;
  wire _39830_;
  wire _39831_;
  wire _39832_;
  wire _39833_;
  wire _39834_;
  wire _39835_;
  wire _39836_;
  wire _39837_;
  wire _39838_;
  wire _39839_;
  wire _39840_;
  wire _39841_;
  wire _39842_;
  wire _39843_;
  wire _39844_;
  wire _39845_;
  wire _39846_;
  wire _39847_;
  wire _39848_;
  wire _39849_;
  wire _39850_;
  wire _39851_;
  wire _39852_;
  wire _39853_;
  wire _39854_;
  wire _39855_;
  wire _39856_;
  wire _39857_;
  wire _39858_;
  wire _39859_;
  wire _39860_;
  wire _39861_;
  wire _39862_;
  wire _39863_;
  wire _39864_;
  wire _39865_;
  wire _39866_;
  wire _39867_;
  wire _39868_;
  wire _39869_;
  wire _39870_;
  wire _39871_;
  wire _39872_;
  wire _39873_;
  wire _39874_;
  wire _39875_;
  wire _39876_;
  wire _39877_;
  wire _39878_;
  wire _39879_;
  wire _39880_;
  wire _39881_;
  wire _39882_;
  wire _39883_;
  wire _39884_;
  wire _39885_;
  wire _39886_;
  wire _39887_;
  wire _39888_;
  wire _39889_;
  wire _39890_;
  wire _39891_;
  wire _39892_;
  wire _39893_;
  wire _39894_;
  wire _39895_;
  wire _39896_;
  wire _39897_;
  wire _39898_;
  wire _39899_;
  wire _39900_;
  wire _39901_;
  wire _39902_;
  wire _39903_;
  wire _39904_;
  wire _39905_;
  wire _39906_;
  wire _39907_;
  wire _39908_;
  wire _39909_;
  wire _39910_;
  wire _39911_;
  wire _39912_;
  wire _39913_;
  wire _39914_;
  wire _39915_;
  wire _39916_;
  wire _39917_;
  wire _39918_;
  wire _39919_;
  wire _39920_;
  wire _39921_;
  wire _39922_;
  wire _39923_;
  wire _39924_;
  wire _39925_;
  wire _39926_;
  wire _39927_;
  wire _39928_;
  wire _39929_;
  wire _39930_;
  wire _39931_;
  wire _39932_;
  wire _39933_;
  wire _39934_;
  wire _39935_;
  wire _39936_;
  wire _39937_;
  wire _39938_;
  wire _39939_;
  wire _39940_;
  wire _39941_;
  wire _39942_;
  wire _39943_;
  wire _39944_;
  wire _39945_;
  wire _39946_;
  wire _39947_;
  wire _39948_;
  wire _39949_;
  wire _39950_;
  wire _39951_;
  wire _39952_;
  wire _39953_;
  wire _39954_;
  wire _39955_;
  wire _39956_;
  wire _39957_;
  wire _39958_;
  wire _39959_;
  wire _39960_;
  wire _39961_;
  wire _39962_;
  wire _39963_;
  wire _39964_;
  wire _39965_;
  wire _39966_;
  wire _39967_;
  wire _39968_;
  wire _39969_;
  wire _39970_;
  wire _39971_;
  wire _39972_;
  wire _39973_;
  wire _39974_;
  wire _39975_;
  wire _39976_;
  wire _39977_;
  wire _39978_;
  wire _39979_;
  wire _39980_;
  wire _39981_;
  wire _39982_;
  wire _39983_;
  wire _39984_;
  wire _39985_;
  wire _39986_;
  wire _39987_;
  wire _39988_;
  wire _39989_;
  wire _39990_;
  wire _39991_;
  wire _39992_;
  wire _39993_;
  wire _39994_;
  wire _39995_;
  wire _39996_;
  wire _39997_;
  wire _39998_;
  wire _39999_;
  wire _40000_;
  wire _40001_;
  wire _40002_;
  wire _40003_;
  wire _40004_;
  wire _40005_;
  wire _40006_;
  wire _40007_;
  wire _40008_;
  wire _40009_;
  wire _40010_;
  wire _40011_;
  wire _40012_;
  wire _40013_;
  wire _40014_;
  wire _40015_;
  wire _40016_;
  wire _40017_;
  wire _40018_;
  wire _40019_;
  wire _40020_;
  wire _40021_;
  wire _40022_;
  wire _40023_;
  wire _40024_;
  wire _40025_;
  wire _40026_;
  wire _40027_;
  wire _40028_;
  wire _40029_;
  wire _40030_;
  wire _40031_;
  wire _40032_;
  wire _40033_;
  wire _40034_;
  wire _40035_;
  wire _40036_;
  wire _40037_;
  wire _40038_;
  wire _40039_;
  wire _40040_;
  wire _40041_;
  wire _40042_;
  wire _40043_;
  wire _40044_;
  wire _40045_;
  wire _40046_;
  wire _40047_;
  wire _40048_;
  wire _40049_;
  wire _40050_;
  wire _40051_;
  wire _40052_;
  wire _40053_;
  wire _40054_;
  wire _40055_;
  wire _40056_;
  wire _40057_;
  wire _40058_;
  wire _40059_;
  wire _40060_;
  wire _40061_;
  wire _40062_;
  wire _40063_;
  wire _40064_;
  wire _40065_;
  wire _40066_;
  wire _40067_;
  wire _40068_;
  wire _40069_;
  wire _40070_;
  wire _40071_;
  wire _40072_;
  wire _40073_;
  wire _40074_;
  wire _40075_;
  wire _40076_;
  wire _40077_;
  wire _40078_;
  wire _40079_;
  wire _40080_;
  wire _40081_;
  wire _40082_;
  wire _40083_;
  wire _40084_;
  wire _40085_;
  wire _40086_;
  wire _40087_;
  wire _40088_;
  wire _40089_;
  wire _40090_;
  wire _40091_;
  wire _40092_;
  wire _40093_;
  wire _40094_;
  wire _40095_;
  wire _40096_;
  wire _40097_;
  wire _40098_;
  wire _40099_;
  wire _40100_;
  wire _40101_;
  wire _40102_;
  wire _40103_;
  wire _40104_;
  wire _40105_;
  wire _40106_;
  wire _40107_;
  wire _40108_;
  wire _40109_;
  wire _40110_;
  wire _40111_;
  wire _40112_;
  wire _40113_;
  wire _40114_;
  wire _40115_;
  wire _40116_;
  wire _40117_;
  wire _40118_;
  wire _40119_;
  wire _40120_;
  wire _40121_;
  wire _40122_;
  wire _40123_;
  wire _40124_;
  wire _40125_;
  wire _40126_;
  wire _40127_;
  wire _40128_;
  wire _40129_;
  wire _40130_;
  wire _40131_;
  wire _40132_;
  wire _40133_;
  wire _40134_;
  wire _40135_;
  wire _40136_;
  wire _40137_;
  wire _40138_;
  wire _40139_;
  wire _40140_;
  wire _40141_;
  wire _40142_;
  wire _40143_;
  wire _40144_;
  wire _40145_;
  wire _40146_;
  wire _40147_;
  wire _40148_;
  wire _40149_;
  wire _40150_;
  wire _40151_;
  wire _40152_;
  wire _40153_;
  wire _40154_;
  wire _40155_;
  wire _40156_;
  wire _40157_;
  wire _40158_;
  wire _40159_;
  wire _40160_;
  wire _40161_;
  wire _40162_;
  wire _40163_;
  wire _40164_;
  wire _40165_;
  wire _40166_;
  wire _40167_;
  wire _40168_;
  wire _40169_;
  wire _40170_;
  wire _40171_;
  wire _40172_;
  wire _40173_;
  wire _40174_;
  wire _40175_;
  wire _40176_;
  wire _40177_;
  wire _40178_;
  wire _40179_;
  wire _40180_;
  wire _40181_;
  wire _40182_;
  wire _40183_;
  wire _40184_;
  wire _40185_;
  wire _40186_;
  wire _40187_;
  wire _40188_;
  wire _40189_;
  wire _40190_;
  wire _40191_;
  wire _40192_;
  wire _40193_;
  wire _40194_;
  wire _40195_;
  wire _40196_;
  wire _40197_;
  wire _40198_;
  wire _40199_;
  wire _40200_;
  wire _40201_;
  wire _40202_;
  wire _40203_;
  wire _40204_;
  wire _40205_;
  wire _40206_;
  wire _40207_;
  wire _40208_;
  wire _40209_;
  wire _40210_;
  wire _40211_;
  wire _40212_;
  wire _40213_;
  wire _40214_;
  wire _40215_;
  wire _40216_;
  wire _40217_;
  wire _40218_;
  wire _40219_;
  wire _40220_;
  wire _40221_;
  wire _40222_;
  wire _40223_;
  wire _40224_;
  wire _40225_;
  wire _40226_;
  wire _40227_;
  wire _40228_;
  wire _40229_;
  wire _40230_;
  wire _40231_;
  wire _40232_;
  wire _40233_;
  wire _40234_;
  wire _40235_;
  wire _40236_;
  wire _40237_;
  wire _40238_;
  wire _40239_;
  wire _40240_;
  wire _40241_;
  wire _40242_;
  wire _40243_;
  wire _40244_;
  wire _40245_;
  wire _40246_;
  wire _40247_;
  wire _40248_;
  wire _40249_;
  wire _40250_;
  wire _40251_;
  wire _40252_;
  wire _40253_;
  wire _40254_;
  wire _40255_;
  wire _40256_;
  wire _40257_;
  wire _40258_;
  wire _40259_;
  wire _40260_;
  wire _40261_;
  wire _40262_;
  wire _40263_;
  wire _40264_;
  wire _40265_;
  wire _40266_;
  wire _40267_;
  wire _40268_;
  wire _40269_;
  wire _40270_;
  wire _40271_;
  wire _40272_;
  wire _40273_;
  wire _40274_;
  wire _40275_;
  wire _40276_;
  wire _40277_;
  wire _40278_;
  wire _40279_;
  wire _40280_;
  wire _40281_;
  wire _40282_;
  wire _40283_;
  wire _40284_;
  wire _40285_;
  wire _40286_;
  wire _40287_;
  wire _40288_;
  wire _40289_;
  wire _40290_;
  wire _40291_;
  wire _40292_;
  wire _40293_;
  wire _40294_;
  wire _40295_;
  wire _40296_;
  wire _40297_;
  wire _40298_;
  wire _40299_;
  wire _40300_;
  wire _40301_;
  wire _40302_;
  wire _40303_;
  wire _40304_;
  wire _40305_;
  wire _40306_;
  wire _40307_;
  wire _40308_;
  wire _40309_;
  wire _40310_;
  wire _40311_;
  wire _40312_;
  wire _40313_;
  wire _40314_;
  wire _40315_;
  wire _40316_;
  wire _40317_;
  wire _40318_;
  wire _40319_;
  wire _40320_;
  wire _40321_;
  wire _40322_;
  wire _40323_;
  wire _40324_;
  wire _40325_;
  wire _40326_;
  wire _40327_;
  wire _40328_;
  wire _40329_;
  wire _40330_;
  wire _40331_;
  wire _40332_;
  wire _40333_;
  wire _40334_;
  wire _40335_;
  wire _40336_;
  wire _40337_;
  wire _40338_;
  wire _40339_;
  wire _40340_;
  wire _40341_;
  wire _40342_;
  wire _40343_;
  wire _40344_;
  wire _40345_;
  wire _40346_;
  wire _40347_;
  wire _40348_;
  wire _40349_;
  wire _40350_;
  wire _40351_;
  wire _40352_;
  wire _40353_;
  wire _40354_;
  wire _40355_;
  wire _40356_;
  wire _40357_;
  wire _40358_;
  wire _40359_;
  wire _40360_;
  wire _40361_;
  wire _40362_;
  wire _40363_;
  wire _40364_;
  wire _40365_;
  wire _40366_;
  wire _40367_;
  wire _40368_;
  wire _40369_;
  wire _40370_;
  wire _40371_;
  wire _40372_;
  wire _40373_;
  wire _40374_;
  wire _40375_;
  wire _40376_;
  wire _40377_;
  wire _40378_;
  wire _40379_;
  wire _40380_;
  wire _40381_;
  wire _40382_;
  wire _40383_;
  wire _40384_;
  wire _40385_;
  wire _40386_;
  wire _40387_;
  wire _40388_;
  wire _40389_;
  wire _40390_;
  wire _40391_;
  wire _40392_;
  wire _40393_;
  wire _40394_;
  wire _40395_;
  wire _40396_;
  wire _40397_;
  wire _40398_;
  wire _40399_;
  wire _40400_;
  wire _40401_;
  wire _40402_;
  wire _40403_;
  wire _40404_;
  wire _40405_;
  wire _40406_;
  wire _40407_;
  wire _40408_;
  wire _40409_;
  wire _40410_;
  wire _40411_;
  wire _40412_;
  wire _40413_;
  wire _40414_;
  wire _40415_;
  wire _40416_;
  wire _40417_;
  wire _40418_;
  wire _40419_;
  wire _40420_;
  wire _40421_;
  wire _40422_;
  wire _40423_;
  wire _40424_;
  wire _40425_;
  wire _40426_;
  wire _40427_;
  wire _40428_;
  wire _40429_;
  wire _40430_;
  wire _40431_;
  wire _40432_;
  wire _40433_;
  wire _40434_;
  wire _40435_;
  wire _40436_;
  wire _40437_;
  wire _40438_;
  wire _40439_;
  wire _40440_;
  wire _40441_;
  wire _40442_;
  wire _40443_;
  wire _40444_;
  wire _40445_;
  wire _40446_;
  wire _40447_;
  wire _40448_;
  wire _40449_;
  wire _40450_;
  wire _40451_;
  wire _40452_;
  wire _40453_;
  wire _40454_;
  wire _40455_;
  wire _40456_;
  wire _40457_;
  wire _40458_;
  wire _40459_;
  wire _40460_;
  wire _40461_;
  wire _40462_;
  wire _40463_;
  wire _40464_;
  wire _40465_;
  wire _40466_;
  wire _40467_;
  wire _40468_;
  wire _40469_;
  wire _40470_;
  wire _40471_;
  wire _40472_;
  wire _40473_;
  wire _40474_;
  wire _40475_;
  wire _40476_;
  wire _40477_;
  wire _40478_;
  wire _40479_;
  wire _40480_;
  wire _40481_;
  wire _40482_;
  wire _40483_;
  wire _40484_;
  wire _40485_;
  wire _40486_;
  wire _40487_;
  wire _40488_;
  wire _40489_;
  wire _40490_;
  wire _40491_;
  wire _40492_;
  wire _40493_;
  wire _40494_;
  wire _40495_;
  wire _40496_;
  wire _40497_;
  wire _40498_;
  wire _40499_;
  wire _40500_;
  wire _40501_;
  wire _40502_;
  wire _40503_;
  wire _40504_;
  wire _40505_;
  wire _40506_;
  wire _40507_;
  wire _40508_;
  wire _40509_;
  wire _40510_;
  wire _40511_;
  wire _40512_;
  wire _40513_;
  wire _40514_;
  wire _40515_;
  wire _40516_;
  wire _40517_;
  wire _40518_;
  wire _40519_;
  wire _40520_;
  wire _40521_;
  wire _40522_;
  wire _40523_;
  wire _40524_;
  wire _40525_;
  wire _40526_;
  wire _40527_;
  wire _40528_;
  wire _40529_;
  wire _40530_;
  wire _40531_;
  wire _40532_;
  wire _40533_;
  wire _40534_;
  wire _40535_;
  wire _40536_;
  wire _40537_;
  wire _40538_;
  wire _40539_;
  wire _40540_;
  wire _40541_;
  wire _40542_;
  wire _40543_;
  wire _40544_;
  wire _40545_;
  wire _40546_;
  wire _40547_;
  wire _40548_;
  wire _40549_;
  wire _40550_;
  wire _40551_;
  wire _40552_;
  wire _40553_;
  wire _40554_;
  wire _40555_;
  wire _40556_;
  wire _40557_;
  wire _40558_;
  wire _40559_;
  wire _40560_;
  wire _40561_;
  wire _40562_;
  wire _40563_;
  wire _40564_;
  wire _40565_;
  wire _40566_;
  wire _40567_;
  wire _40568_;
  wire _40569_;
  wire _40570_;
  wire _40571_;
  wire _40572_;
  wire _40573_;
  wire _40574_;
  wire _40575_;
  wire _40576_;
  wire _40577_;
  wire _40578_;
  wire _40579_;
  wire _40580_;
  wire _40581_;
  wire _40582_;
  wire _40583_;
  wire _40584_;
  wire _40585_;
  wire _40586_;
  wire _40587_;
  wire _40588_;
  wire _40589_;
  wire _40590_;
  wire _40591_;
  wire _40592_;
  wire _40593_;
  wire _40594_;
  wire _40595_;
  wire _40596_;
  wire _40597_;
  wire _40598_;
  wire _40599_;
  wire _40600_;
  wire _40601_;
  wire _40602_;
  wire _40603_;
  wire _40604_;
  wire _40605_;
  wire _40606_;
  wire _40607_;
  wire _40608_;
  wire _40609_;
  wire _40610_;
  wire _40611_;
  wire _40612_;
  wire _40613_;
  wire _40614_;
  wire _40615_;
  wire _40616_;
  wire _40617_;
  wire _40618_;
  wire _40619_;
  wire _40620_;
  wire _40621_;
  wire _40622_;
  wire _40623_;
  wire _40624_;
  wire _40625_;
  wire _40626_;
  wire _40627_;
  wire _40628_;
  wire _40629_;
  wire _40630_;
  wire _40631_;
  wire _40632_;
  wire _40633_;
  wire _40634_;
  wire _40635_;
  wire _40636_;
  wire _40637_;
  wire _40638_;
  wire _40639_;
  wire _40640_;
  wire _40641_;
  wire _40642_;
  wire _40643_;
  wire _40644_;
  wire _40645_;
  wire _40646_;
  wire _40647_;
  wire _40648_;
  wire _40649_;
  wire _40650_;
  wire _40651_;
  wire _40652_;
  wire _40653_;
  wire _40654_;
  wire _40655_;
  wire _40656_;
  wire _40657_;
  wire _40658_;
  wire _40659_;
  wire _40660_;
  wire _40661_;
  wire _40662_;
  wire _40663_;
  wire _40664_;
  wire _40665_;
  wire _40666_;
  wire _40667_;
  wire _40668_;
  wire _40669_;
  wire _40670_;
  wire _40671_;
  wire _40672_;
  wire _40673_;
  wire _40674_;
  wire _40675_;
  wire _40676_;
  wire _40677_;
  wire _40678_;
  wire _40679_;
  wire _40680_;
  wire _40681_;
  wire _40682_;
  wire _40683_;
  wire _40684_;
  wire _40685_;
  wire _40686_;
  wire _40687_;
  wire _40688_;
  wire _40689_;
  wire _40690_;
  wire _40691_;
  wire _40692_;
  wire _40693_;
  wire _40694_;
  wire _40695_;
  wire _40696_;
  wire _40697_;
  wire _40698_;
  wire _40699_;
  wire _40700_;
  wire _40701_;
  wire _40702_;
  wire _40703_;
  wire _40704_;
  wire _40705_;
  wire _40706_;
  wire _40707_;
  wire _40708_;
  wire _40709_;
  wire _40710_;
  wire _40711_;
  wire _40712_;
  wire _40713_;
  wire _40714_;
  wire _40715_;
  wire _40716_;
  wire _40717_;
  wire _40718_;
  wire _40719_;
  wire _40720_;
  wire _40721_;
  wire _40722_;
  wire _40723_;
  wire _40724_;
  wire _40725_;
  wire _40726_;
  wire _40727_;
  wire _40728_;
  wire _40729_;
  wire _40730_;
  wire _40731_;
  wire _40732_;
  wire _40733_;
  wire _40734_;
  wire _40735_;
  wire _40736_;
  wire _40737_;
  wire _40738_;
  wire _40739_;
  wire _40740_;
  wire _40741_;
  wire _40742_;
  wire _40743_;
  wire _40744_;
  wire _40745_;
  wire _40746_;
  wire _40747_;
  wire _40748_;
  wire _40749_;
  wire _40750_;
  wire _40751_;
  wire _40752_;
  wire _40753_;
  wire _40754_;
  wire _40755_;
  wire _40756_;
  wire _40757_;
  wire _40758_;
  wire _40759_;
  wire _40760_;
  wire _40761_;
  wire _40762_;
  wire _40763_;
  wire _40764_;
  wire _40765_;
  wire _40766_;
  wire _40767_;
  wire _40768_;
  wire _40769_;
  wire _40770_;
  wire _40771_;
  wire _40772_;
  wire _40773_;
  wire _40774_;
  wire _40775_;
  wire _40776_;
  wire _40777_;
  wire _40778_;
  wire _40779_;
  wire _40780_;
  wire _40781_;
  wire _40782_;
  wire _40783_;
  wire _40784_;
  wire _40785_;
  wire _40786_;
  wire _40787_;
  wire _40788_;
  wire _40789_;
  wire _40790_;
  wire _40791_;
  wire _40792_;
  wire _40793_;
  wire _40794_;
  wire _40795_;
  wire _40796_;
  wire _40797_;
  wire _40798_;
  wire _40799_;
  wire _40800_;
  wire _40801_;
  wire _40802_;
  wire _40803_;
  wire _40804_;
  wire _40805_;
  wire _40806_;
  wire _40807_;
  wire _40808_;
  wire _40809_;
  wire _40810_;
  wire _40811_;
  wire _40812_;
  wire _40813_;
  wire _40814_;
  wire _40815_;
  wire _40816_;
  wire _40817_;
  wire _40818_;
  wire _40819_;
  wire _40820_;
  wire _40821_;
  wire _40822_;
  wire _40823_;
  wire _40824_;
  wire _40825_;
  wire _40826_;
  wire _40827_;
  wire _40828_;
  wire _40829_;
  wire _40830_;
  wire _40831_;
  wire _40832_;
  wire _40833_;
  wire _40834_;
  wire _40835_;
  wire _40836_;
  wire _40837_;
  wire _40838_;
  wire _40839_;
  wire _40840_;
  wire _40841_;
  wire _40842_;
  wire _40843_;
  wire _40844_;
  wire _40845_;
  wire _40846_;
  wire _40847_;
  wire _40848_;
  wire _40849_;
  wire _40850_;
  wire _40851_;
  wire _40852_;
  wire _40853_;
  wire _40854_;
  wire _40855_;
  wire _40856_;
  wire _40857_;
  wire _40858_;
  wire _40859_;
  wire _40860_;
  wire _40861_;
  wire _40862_;
  wire _40863_;
  wire _40864_;
  wire _40865_;
  wire _40866_;
  wire _40867_;
  wire _40868_;
  wire _40869_;
  wire _40870_;
  wire _40871_;
  wire _40872_;
  wire _40873_;
  wire _40874_;
  wire _40875_;
  wire _40876_;
  wire _40877_;
  wire _40878_;
  wire _40879_;
  wire _40880_;
  wire _40881_;
  wire _40882_;
  wire _40883_;
  wire _40884_;
  wire _40885_;
  wire _40886_;
  wire _40887_;
  wire _40888_;
  wire _40889_;
  wire _40890_;
  wire _40891_;
  wire _40892_;
  wire _40893_;
  wire _40894_;
  wire _40895_;
  wire _40896_;
  wire _40897_;
  wire _40898_;
  wire _40899_;
  wire _40900_;
  wire _40901_;
  wire _40902_;
  wire _40903_;
  wire _40904_;
  wire _40905_;
  wire _40906_;
  wire _40907_;
  wire _40908_;
  wire _40909_;
  wire _40910_;
  wire _40911_;
  wire _40912_;
  wire _40913_;
  wire _40914_;
  wire _40915_;
  wire _40916_;
  wire _40917_;
  wire _40918_;
  wire _40919_;
  wire _40920_;
  wire _40921_;
  wire _40922_;
  wire _40923_;
  wire _40924_;
  wire _40925_;
  wire _40926_;
  wire _40927_;
  wire _40928_;
  wire _40929_;
  wire _40930_;
  wire _40931_;
  wire _40932_;
  wire _40933_;
  wire _40934_;
  wire _40935_;
  wire _40936_;
  wire _40937_;
  wire _40938_;
  wire _40939_;
  wire _40940_;
  wire _40941_;
  wire _40942_;
  wire _40943_;
  wire _40944_;
  wire _40945_;
  wire _40946_;
  wire _40947_;
  wire _40948_;
  wire _40949_;
  wire _40950_;
  wire _40951_;
  wire _40952_;
  wire _40953_;
  wire _40954_;
  wire _40955_;
  wire _40956_;
  wire _40957_;
  wire _40958_;
  wire _40959_;
  wire _40960_;
  wire _40961_;
  wire _40962_;
  wire _40963_;
  wire _40964_;
  wire _40965_;
  wire _40966_;
  wire _40967_;
  wire _40968_;
  wire _40969_;
  wire _40970_;
  wire _40971_;
  wire _40972_;
  wire _40973_;
  wire _40974_;
  wire _40975_;
  wire _40976_;
  wire _40977_;
  wire _40978_;
  wire _40979_;
  wire _40980_;
  wire _40981_;
  wire _40982_;
  wire _40983_;
  wire _40984_;
  wire _40985_;
  wire _40986_;
  wire _40987_;
  wire _40988_;
  wire _40989_;
  wire _40990_;
  wire _40991_;
  wire _40992_;
  wire _40993_;
  wire _40994_;
  wire _40995_;
  wire _40996_;
  wire _40997_;
  wire _40998_;
  wire _40999_;
  wire _41000_;
  wire _41001_;
  wire _41002_;
  wire _41003_;
  wire _41004_;
  wire _41005_;
  wire _41006_;
  wire _41007_;
  wire _41008_;
  wire _41009_;
  wire _41010_;
  wire _41011_;
  wire _41012_;
  wire _41013_;
  wire _41014_;
  wire _41015_;
  wire _41016_;
  wire _41017_;
  wire _41018_;
  wire _41019_;
  wire _41020_;
  wire _41021_;
  wire _41022_;
  wire _41023_;
  wire _41024_;
  wire _41025_;
  wire _41026_;
  wire _41027_;
  wire _41028_;
  wire _41029_;
  wire _41030_;
  wire _41031_;
  wire _41032_;
  wire _41033_;
  wire _41034_;
  wire _41035_;
  wire _41036_;
  wire _41037_;
  wire _41038_;
  wire _41039_;
  wire _41040_;
  wire _41041_;
  wire _41042_;
  wire _41043_;
  wire _41044_;
  wire _41045_;
  wire _41046_;
  wire _41047_;
  wire _41048_;
  wire _41049_;
  wire _41050_;
  wire _41051_;
  wire _41052_;
  wire _41053_;
  wire _41054_;
  wire _41055_;
  wire _41056_;
  wire _41057_;
  wire _41058_;
  wire _41059_;
  wire _41060_;
  wire _41061_;
  wire _41062_;
  wire _41063_;
  wire _41064_;
  wire _41065_;
  wire _41066_;
  wire _41067_;
  wire _41068_;
  wire _41069_;
  wire _41070_;
  wire _41071_;
  wire _41072_;
  wire _41073_;
  wire _41074_;
  wire _41075_;
  wire _41076_;
  wire _41077_;
  wire _41078_;
  wire _41079_;
  wire _41080_;
  wire _41081_;
  wire _41082_;
  wire _41083_;
  wire _41084_;
  wire _41085_;
  wire _41086_;
  wire _41087_;
  wire _41088_;
  wire _41089_;
  wire _41090_;
  wire _41091_;
  wire _41092_;
  wire _41093_;
  wire _41094_;
  wire _41095_;
  wire _41096_;
  wire _41097_;
  wire _41098_;
  wire _41099_;
  wire _41100_;
  wire _41101_;
  wire _41102_;
  wire _41103_;
  wire _41104_;
  wire _41105_;
  wire _41106_;
  wire _41107_;
  wire _41108_;
  wire _41109_;
  wire _41110_;
  wire _41111_;
  wire _41112_;
  wire _41113_;
  wire _41114_;
  wire _41115_;
  wire _41116_;
  wire _41117_;
  wire _41118_;
  wire _41119_;
  wire _41120_;
  wire _41121_;
  wire _41122_;
  wire _41123_;
  wire _41124_;
  wire _41125_;
  wire _41126_;
  wire _41127_;
  wire _41128_;
  wire _41129_;
  wire _41130_;
  wire _41131_;
  wire _41132_;
  wire _41133_;
  wire _41134_;
  wire _41135_;
  wire _41136_;
  wire _41137_;
  wire _41138_;
  wire _41139_;
  wire _41140_;
  wire _41141_;
  wire _41142_;
  wire _41143_;
  wire _41144_;
  wire _41145_;
  wire _41146_;
  wire _41147_;
  wire _41148_;
  wire _41149_;
  wire _41150_;
  wire _41151_;
  wire _41152_;
  wire _41153_;
  wire _41154_;
  wire _41155_;
  wire _41156_;
  wire _41157_;
  wire _41158_;
  wire _41159_;
  wire _41160_;
  wire _41161_;
  wire _41162_;
  wire _41163_;
  wire _41164_;
  wire _41165_;
  wire _41166_;
  wire _41167_;
  wire _41168_;
  wire _41169_;
  wire _41170_;
  wire _41171_;
  wire _41172_;
  wire _41173_;
  wire _41174_;
  wire _41175_;
  wire _41176_;
  wire _41177_;
  wire _41178_;
  wire _41179_;
  wire _41180_;
  wire _41181_;
  wire _41182_;
  wire _41183_;
  wire _41184_;
  wire _41185_;
  wire _41186_;
  wire _41187_;
  wire _41188_;
  wire _41189_;
  wire _41190_;
  wire _41191_;
  wire _41192_;
  wire _41193_;
  wire _41194_;
  wire _41195_;
  wire _41196_;
  wire _41197_;
  wire _41198_;
  wire _41199_;
  wire _41200_;
  wire _41201_;
  wire _41202_;
  wire _41203_;
  wire _41204_;
  wire _41205_;
  wire _41206_;
  wire _41207_;
  wire _41208_;
  wire _41209_;
  wire _41210_;
  wire _41211_;
  wire _41212_;
  wire _41213_;
  wire _41214_;
  wire _41215_;
  wire _41216_;
  wire _41217_;
  wire _41218_;
  wire _41219_;
  wire _41220_;
  wire _41221_;
  wire _41222_;
  wire _41223_;
  wire _41224_;
  wire _41225_;
  wire _41226_;
  wire _41227_;
  wire _41228_;
  wire _41229_;
  wire _41230_;
  wire _41231_;
  wire _41232_;
  wire _41233_;
  wire _41234_;
  wire _41235_;
  wire _41236_;
  wire _41237_;
  wire _41238_;
  wire _41239_;
  wire _41240_;
  wire _41241_;
  wire _41242_;
  wire _41243_;
  wire _41244_;
  wire _41245_;
  wire _41246_;
  wire _41247_;
  wire _41248_;
  wire _41249_;
  wire _41250_;
  wire _41251_;
  wire _41252_;
  wire _41253_;
  wire _41254_;
  wire _41255_;
  wire _41256_;
  wire _41257_;
  wire _41258_;
  wire _41259_;
  wire _41260_;
  wire _41261_;
  wire _41262_;
  wire _41263_;
  wire _41264_;
  wire _41265_;
  wire _41266_;
  wire _41267_;
  wire _41268_;
  wire _41269_;
  wire _41270_;
  wire _41271_;
  wire _41272_;
  wire _41273_;
  wire _41274_;
  wire _41275_;
  wire _41276_;
  wire _41277_;
  wire _41278_;
  wire _41279_;
  wire _41280_;
  wire _41281_;
  wire _41282_;
  wire _41283_;
  wire _41284_;
  wire _41285_;
  wire _41286_;
  wire _41287_;
  wire _41288_;
  wire _41289_;
  wire _41290_;
  wire _41291_;
  wire _41292_;
  wire _41293_;
  wire _41294_;
  wire _41295_;
  wire _41296_;
  wire _41297_;
  wire _41298_;
  wire _41299_;
  wire _41300_;
  wire _41301_;
  wire _41302_;
  wire _41303_;
  wire _41304_;
  wire _41305_;
  wire _41306_;
  wire _41307_;
  wire _41308_;
  wire _41309_;
  wire _41310_;
  wire _41311_;
  wire _41312_;
  wire _41313_;
  wire _41314_;
  wire _41315_;
  wire _41316_;
  wire _41317_;
  wire _41318_;
  wire _41319_;
  wire _41320_;
  wire _41321_;
  wire _41322_;
  wire _41323_;
  wire _41324_;
  wire _41325_;
  wire _41326_;
  wire _41327_;
  wire _41328_;
  wire _41329_;
  wire _41330_;
  wire _41331_;
  wire _41332_;
  wire _41333_;
  wire _41334_;
  wire _41335_;
  wire _41336_;
  wire _41337_;
  wire _41338_;
  wire _41339_;
  wire _41340_;
  wire _41341_;
  wire _41342_;
  wire _41343_;
  wire _41344_;
  wire _41345_;
  wire _41346_;
  wire _41347_;
  wire _41348_;
  wire _41349_;
  wire _41350_;
  wire _41351_;
  wire _41352_;
  wire _41353_;
  wire _41354_;
  wire _41355_;
  wire _41356_;
  wire _41357_;
  wire _41358_;
  wire _41359_;
  wire _41360_;
  wire _41361_;
  wire _41362_;
  wire _41363_;
  wire _41364_;
  wire _41365_;
  wire _41366_;
  wire _41367_;
  wire _41368_;
  wire _41369_;
  wire _41370_;
  wire _41371_;
  wire _41372_;
  wire _41373_;
  wire _41374_;
  wire _41375_;
  wire _41376_;
  wire _41377_;
  wire _41378_;
  wire _41379_;
  wire _41380_;
  wire _41381_;
  wire _41382_;
  wire _41383_;
  wire _41384_;
  wire _41385_;
  wire _41386_;
  wire _41387_;
  wire _41388_;
  wire _41389_;
  wire _41390_;
  wire _41391_;
  wire _41392_;
  wire _41393_;
  wire _41394_;
  wire _41395_;
  wire _41396_;
  wire _41397_;
  wire _41398_;
  wire _41399_;
  wire _41400_;
  wire _41401_;
  wire _41402_;
  wire _41403_;
  wire _41404_;
  wire _41405_;
  wire _41406_;
  wire _41407_;
  wire _41408_;
  wire _41409_;
  wire _41410_;
  wire _41411_;
  wire _41412_;
  wire _41413_;
  wire _41414_;
  wire _41415_;
  wire _41416_;
  wire _41417_;
  wire _41418_;
  wire _41419_;
  wire _41420_;
  wire _41421_;
  wire _41422_;
  wire _41423_;
  wire _41424_;
  wire _41425_;
  wire _41426_;
  wire _41427_;
  wire _41428_;
  wire _41429_;
  wire _41430_;
  wire _41431_;
  wire _41432_;
  wire _41433_;
  wire _41434_;
  wire _41435_;
  wire _41436_;
  wire _41437_;
  wire _41438_;
  wire _41439_;
  wire _41440_;
  wire _41441_;
  wire _41442_;
  wire _41443_;
  wire _41444_;
  wire _41445_;
  wire _41446_;
  wire _41447_;
  wire _41448_;
  wire _41449_;
  wire _41450_;
  wire _41451_;
  wire _41452_;
  wire _41453_;
  wire _41454_;
  wire _41455_;
  wire _41456_;
  wire _41457_;
  wire _41458_;
  wire _41459_;
  wire _41460_;
  wire _41461_;
  wire _41462_;
  wire _41463_;
  wire _41464_;
  wire _41465_;
  wire _41466_;
  wire _41467_;
  wire _41468_;
  wire _41469_;
  wire _41470_;
  wire _41471_;
  wire _41472_;
  wire _41473_;
  wire _41474_;
  wire _41475_;
  wire _41476_;
  wire _41477_;
  wire _41478_;
  wire _41479_;
  wire _41480_;
  wire _41481_;
  wire _41482_;
  wire _41483_;
  wire _41484_;
  wire _41485_;
  wire _41486_;
  wire _41487_;
  wire _41488_;
  wire _41489_;
  wire _41490_;
  wire _41491_;
  wire _41492_;
  wire _41493_;
  wire _41494_;
  wire _41495_;
  wire _41496_;
  wire _41497_;
  wire _41498_;
  wire _41499_;
  wire _41500_;
  wire _41501_;
  wire _41502_;
  wire _41503_;
  wire _41504_;
  wire _41505_;
  wire _41506_;
  wire _41507_;
  wire _41508_;
  wire _41509_;
  wire _41510_;
  wire _41511_;
  wire _41512_;
  wire _41513_;
  wire _41514_;
  wire _41515_;
  wire _41516_;
  wire _41517_;
  wire _41518_;
  wire _41519_;
  wire _41520_;
  wire _41521_;
  wire _41522_;
  wire _41523_;
  wire _41524_;
  wire _41525_;
  wire _41526_;
  wire _41527_;
  wire _41528_;
  wire _41529_;
  wire _41530_;
  wire _41531_;
  wire _41532_;
  wire _41533_;
  wire _41534_;
  wire _41535_;
  wire _41536_;
  wire _41537_;
  wire _41538_;
  wire _41539_;
  wire _41540_;
  wire _41541_;
  wire _41542_;
  wire _41543_;
  wire _41544_;
  wire _41545_;
  wire _41546_;
  wire _41547_;
  wire _41548_;
  wire _41549_;
  wire _41550_;
  wire _41551_;
  wire _41552_;
  wire _41553_;
  wire _41554_;
  wire _41555_;
  wire _41556_;
  wire _41557_;
  wire _41558_;
  wire _41559_;
  wire _41560_;
  wire _41561_;
  wire _41562_;
  wire _41563_;
  wire _41564_;
  wire _41565_;
  wire _41566_;
  wire _41567_;
  wire _41568_;
  wire _41569_;
  wire _41570_;
  wire _41571_;
  wire _41572_;
  wire _41573_;
  wire _41574_;
  wire _41575_;
  wire _41576_;
  wire _41577_;
  wire _41578_;
  wire _41579_;
  wire _41580_;
  wire _41581_;
  wire _41582_;
  wire _41583_;
  wire _41584_;
  wire _41585_;
  wire _41586_;
  wire _41587_;
  wire _41588_;
  wire _41589_;
  wire _41590_;
  wire _41591_;
  wire _41592_;
  wire _41593_;
  wire _41594_;
  wire _41595_;
  wire _41596_;
  wire _41597_;
  wire _41598_;
  wire _41599_;
  wire _41600_;
  wire _41601_;
  wire _41602_;
  wire _41603_;
  wire _41604_;
  wire _41605_;
  wire _41606_;
  wire _41607_;
  wire _41608_;
  wire _41609_;
  wire _41610_;
  wire _41611_;
  wire _41612_;
  wire _41613_;
  wire _41614_;
  wire _41615_;
  wire _41616_;
  wire _41617_;
  wire _41618_;
  wire _41619_;
  wire _41620_;
  wire _41621_;
  wire _41622_;
  wire _41623_;
  wire _41624_;
  wire _41625_;
  wire _41626_;
  wire _41627_;
  wire _41628_;
  wire _41629_;
  wire _41630_;
  wire _41631_;
  wire _41632_;
  wire _41633_;
  wire _41634_;
  wire _41635_;
  wire _41636_;
  wire _41637_;
  wire _41638_;
  wire _41639_;
  wire _41640_;
  wire _41641_;
  wire _41642_;
  wire _41643_;
  wire _41644_;
  wire _41645_;
  wire _41646_;
  wire _41647_;
  wire _41648_;
  wire _41649_;
  wire _41650_;
  wire _41651_;
  wire _41652_;
  wire _41653_;
  wire _41654_;
  wire _41655_;
  wire _41656_;
  wire _41657_;
  wire _41658_;
  wire _41659_;
  wire _41660_;
  wire _41661_;
  wire _41662_;
  wire _41663_;
  wire _41664_;
  wire _41665_;
  wire _41666_;
  wire _41667_;
  wire _41668_;
  wire _41669_;
  wire _41670_;
  wire _41671_;
  wire _41672_;
  wire _41673_;
  wire _41674_;
  wire _41675_;
  wire _41676_;
  wire _41677_;
  wire _41678_;
  wire _41679_;
  wire _41680_;
  wire _41681_;
  wire _41682_;
  wire _41683_;
  wire _41684_;
  wire _41685_;
  wire _41686_;
  wire _41687_;
  wire _41688_;
  wire _41689_;
  wire _41690_;
  wire _41691_;
  wire _41692_;
  wire _41693_;
  wire _41694_;
  wire _41695_;
  wire _41696_;
  wire _41697_;
  wire _41698_;
  wire _41699_;
  wire _41700_;
  wire _41701_;
  wire _41702_;
  wire _41703_;
  wire _41704_;
  wire _41705_;
  wire _41706_;
  wire _41707_;
  wire _41708_;
  wire _41709_;
  wire _41710_;
  wire _41711_;
  wire _41712_;
  wire _41713_;
  wire _41714_;
  wire _41715_;
  wire _41716_;
  wire _41717_;
  wire _41718_;
  wire _41719_;
  wire _41720_;
  wire _41721_;
  wire _41722_;
  wire _41723_;
  wire _41724_;
  wire _41725_;
  wire _41726_;
  wire _41727_;
  wire _41728_;
  wire _41729_;
  wire _41730_;
  wire _41731_;
  wire _41732_;
  wire _41733_;
  wire _41734_;
  wire _41735_;
  wire _41736_;
  wire _41737_;
  wire _41738_;
  wire _41739_;
  wire _41740_;
  wire _41741_;
  wire _41742_;
  wire _41743_;
  wire _41744_;
  wire _41745_;
  wire _41746_;
  wire _41747_;
  wire _41748_;
  wire _41749_;
  wire _41750_;
  wire _41751_;
  wire _41752_;
  wire _41753_;
  wire _41754_;
  wire _41755_;
  wire _41756_;
  wire _41757_;
  wire _41758_;
  wire _41759_;
  wire _41760_;
  wire _41761_;
  wire _41762_;
  wire _41763_;
  wire _41764_;
  wire _41765_;
  wire _41766_;
  wire _41767_;
  wire _41768_;
  wire _41769_;
  wire _41770_;
  wire _41771_;
  wire _41772_;
  wire _41773_;
  wire _41774_;
  wire _41775_;
  wire _41776_;
  wire _41777_;
  wire _41778_;
  wire _41779_;
  wire _41780_;
  wire _41781_;
  wire _41782_;
  wire _41783_;
  wire _41784_;
  wire _41785_;
  wire _41786_;
  wire _41787_;
  wire _41788_;
  wire _41789_;
  wire _41790_;
  wire _41791_;
  wire _41792_;
  wire _41793_;
  wire _41794_;
  wire _41795_;
  wire _41796_;
  wire _41797_;
  wire _41798_;
  wire _41799_;
  wire _41800_;
  wire _41801_;
  wire _41802_;
  wire _41803_;
  wire _41804_;
  wire _41805_;
  wire _41806_;
  wire _41807_;
  wire _41808_;
  wire _41809_;
  wire _41810_;
  wire _41811_;
  wire _41812_;
  wire _41813_;
  wire _41814_;
  wire _41815_;
  wire _41816_;
  wire _41817_;
  wire _41818_;
  wire _41819_;
  wire _41820_;
  wire _41821_;
  wire _41822_;
  wire _41823_;
  wire _41824_;
  wire _41825_;
  wire _41826_;
  wire _41827_;
  wire _41828_;
  wire _41829_;
  wire _41830_;
  wire _41831_;
  wire _41832_;
  wire _41833_;
  wire _41834_;
  wire _41835_;
  wire _41836_;
  wire _41837_;
  wire _41838_;
  wire _41839_;
  wire _41840_;
  wire _41841_;
  wire _41842_;
  wire _41843_;
  wire _41844_;
  wire _41845_;
  wire _41846_;
  wire _41847_;
  wire _41848_;
  wire _41849_;
  wire _41850_;
  wire _41851_;
  wire _41852_;
  wire _41853_;
  wire _41854_;
  wire _41855_;
  wire _41856_;
  wire _41857_;
  wire _41858_;
  wire _41859_;
  wire _41860_;
  wire _41861_;
  wire _41862_;
  wire _41863_;
  wire _41864_;
  wire _41865_;
  wire _41866_;
  wire _41867_;
  wire _41868_;
  wire _41869_;
  wire _41870_;
  wire _41871_;
  wire _41872_;
  wire _41873_;
  wire _41874_;
  wire _41875_;
  wire _41876_;
  wire _41877_;
  wire _41878_;
  wire _41879_;
  wire _41880_;
  wire _41881_;
  wire _41882_;
  wire _41883_;
  wire _41884_;
  wire _41885_;
  wire _41886_;
  wire _41887_;
  wire _41888_;
  wire _41889_;
  wire _41890_;
  wire _41891_;
  wire _41892_;
  wire _41893_;
  wire _41894_;
  wire _41895_;
  wire _41896_;
  wire _41897_;
  wire _41898_;
  wire _41899_;
  wire _41900_;
  wire _41901_;
  wire _41902_;
  wire _41903_;
  wire _41904_;
  wire _41905_;
  wire _41906_;
  wire _41907_;
  wire _41908_;
  wire _41909_;
  wire _41910_;
  wire _41911_;
  wire _41912_;
  wire _41913_;
  wire _41914_;
  wire _41915_;
  wire _41916_;
  wire _41917_;
  wire _41918_;
  wire _41919_;
  wire _41920_;
  wire _41921_;
  wire _41922_;
  wire _41923_;
  wire _41924_;
  wire _41925_;
  wire _41926_;
  wire _41927_;
  wire _41928_;
  wire _41929_;
  wire _41930_;
  wire _41931_;
  wire _41932_;
  wire _41933_;
  wire _41934_;
  wire _41935_;
  wire _41936_;
  wire _41937_;
  wire _41938_;
  wire _41939_;
  wire _41940_;
  wire _41941_;
  wire _41942_;
  wire _41943_;
  wire _41944_;
  wire _41945_;
  wire _41946_;
  wire _41947_;
  wire _41948_;
  wire _41949_;
  wire _41950_;
  wire _41951_;
  wire _41952_;
  wire _41953_;
  wire _41954_;
  wire _41955_;
  wire _41956_;
  wire _41957_;
  wire _41958_;
  wire _41959_;
  wire _41960_;
  wire _41961_;
  wire _41962_;
  wire _41963_;
  wire _41964_;
  wire _41965_;
  wire _41966_;
  wire _41967_;
  wire _41968_;
  wire _41969_;
  wire _41970_;
  wire _41971_;
  wire _41972_;
  wire _41973_;
  wire _41974_;
  wire _41975_;
  wire _41976_;
  wire _41977_;
  wire _41978_;
  wire _41979_;
  wire _41980_;
  wire _41981_;
  wire _41982_;
  wire _41983_;
  wire _41984_;
  wire _41985_;
  wire _41986_;
  wire _41987_;
  wire _41988_;
  wire _41989_;
  wire _41990_;
  wire _41991_;
  wire _41992_;
  wire _41993_;
  wire _41994_;
  wire _41995_;
  wire _41996_;
  wire _41997_;
  wire _41998_;
  wire _41999_;
  wire _42000_;
  wire _42001_;
  wire _42002_;
  wire _42003_;
  wire _42004_;
  wire _42005_;
  wire _42006_;
  wire _42007_;
  wire _42008_;
  wire _42009_;
  wire _42010_;
  wire _42011_;
  wire _42012_;
  wire _42013_;
  wire _42014_;
  wire _42015_;
  wire _42016_;
  wire _42017_;
  wire _42018_;
  wire _42019_;
  wire _42020_;
  wire _42021_;
  wire _42022_;
  wire _42023_;
  wire _42024_;
  wire _42025_;
  wire _42026_;
  wire _42027_;
  wire _42028_;
  wire _42029_;
  wire _42030_;
  wire _42031_;
  wire _42032_;
  wire _42033_;
  wire _42034_;
  wire _42035_;
  wire _42036_;
  wire _42037_;
  wire _42038_;
  wire _42039_;
  wire _42040_;
  wire _42041_;
  wire _42042_;
  wire _42043_;
  wire _42044_;
  wire _42045_;
  wire _42046_;
  wire _42047_;
  wire _42048_;
  wire _42049_;
  wire _42050_;
  wire _42051_;
  wire _42052_;
  wire _42053_;
  wire _42054_;
  wire _42055_;
  wire _42056_;
  wire _42057_;
  wire _42058_;
  wire _42059_;
  wire _42060_;
  wire _42061_;
  wire _42062_;
  wire _42063_;
  wire _42064_;
  wire _42065_;
  wire _42066_;
  wire _42067_;
  wire _42068_;
  wire _42069_;
  wire _42070_;
  wire _42071_;
  wire _42072_;
  wire _42073_;
  wire _42074_;
  wire _42075_;
  wire _42076_;
  wire _42077_;
  wire _42078_;
  wire _42079_;
  wire _42080_;
  wire _42081_;
  wire _42082_;
  wire _42083_;
  wire _42084_;
  wire _42085_;
  wire _42086_;
  wire _42087_;
  wire _42088_;
  wire _42089_;
  wire _42090_;
  wire _42091_;
  wire _42092_;
  wire _42093_;
  wire _42094_;
  wire _42095_;
  wire _42096_;
  wire _42097_;
  wire _42098_;
  wire _42099_;
  wire _42100_;
  wire _42101_;
  wire _42102_;
  wire _42103_;
  wire _42104_;
  wire _42105_;
  wire _42106_;
  wire _42107_;
  wire _42108_;
  wire _42109_;
  wire _42110_;
  wire _42111_;
  wire _42112_;
  wire _42113_;
  wire _42114_;
  wire _42115_;
  wire _42116_;
  wire _42117_;
  wire _42118_;
  wire _42119_;
  wire _42120_;
  wire _42121_;
  wire _42122_;
  wire _42123_;
  wire _42124_;
  wire _42125_;
  wire _42126_;
  wire _42127_;
  wire _42128_;
  wire _42129_;
  wire _42130_;
  wire _42131_;
  wire _42132_;
  wire _42133_;
  wire _42134_;
  wire _42135_;
  wire _42136_;
  wire _42137_;
  wire _42138_;
  wire _42139_;
  wire _42140_;
  wire _42141_;
  wire _42142_;
  wire _42143_;
  wire _42144_;
  wire _42145_;
  wire _42146_;
  wire _42147_;
  wire _42148_;
  wire _42149_;
  wire _42150_;
  wire _42151_;
  wire _42152_;
  wire _42153_;
  wire _42154_;
  wire _42155_;
  wire _42156_;
  wire _42157_;
  wire _42158_;
  wire _42159_;
  wire _42160_;
  wire _42161_;
  wire _42162_;
  wire _42163_;
  wire _42164_;
  wire _42165_;
  wire _42166_;
  wire _42167_;
  wire _42168_;
  wire _42169_;
  wire _42170_;
  wire _42171_;
  wire _42172_;
  wire _42173_;
  wire _42174_;
  wire _42175_;
  wire _42176_;
  wire _42177_;
  wire _42178_;
  wire _42179_;
  wire _42180_;
  wire _42181_;
  wire _42182_;
  wire _42183_;
  wire _42184_;
  wire _42185_;
  wire _42186_;
  wire _42187_;
  wire _42188_;
  wire _42189_;
  wire _42190_;
  wire _42191_;
  wire _42192_;
  wire _42193_;
  wire _42194_;
  wire _42195_;
  wire _42196_;
  wire _42197_;
  wire _42198_;
  wire _42199_;
  wire _42200_;
  wire _42201_;
  wire _42202_;
  wire _42203_;
  wire _42204_;
  wire _42205_;
  wire _42206_;
  wire _42207_;
  wire _42208_;
  wire _42209_;
  wire _42210_;
  wire _42211_;
  wire _42212_;
  wire _42213_;
  wire _42214_;
  wire _42215_;
  wire _42216_;
  wire _42217_;
  wire _42218_;
  wire _42219_;
  wire _42220_;
  wire _42221_;
  wire _42222_;
  wire _42223_;
  wire _42224_;
  wire _42225_;
  wire _42226_;
  wire _42227_;
  wire _42228_;
  wire _42229_;
  wire _42230_;
  wire _42231_;
  wire _42232_;
  wire _42233_;
  wire _42234_;
  wire _42235_;
  wire _42236_;
  wire _42237_;
  wire _42238_;
  wire _42239_;
  wire _42240_;
  wire _42241_;
  wire _42242_;
  wire _42243_;
  wire _42244_;
  wire _42245_;
  wire _42246_;
  wire _42247_;
  wire _42248_;
  wire _42249_;
  wire _42250_;
  wire _42251_;
  wire _42252_;
  wire _42253_;
  wire _42254_;
  wire _42255_;
  wire _42256_;
  wire _42257_;
  wire _42258_;
  wire _42259_;
  wire _42260_;
  wire _42261_;
  wire _42262_;
  wire _42263_;
  wire _42264_;
  wire _42265_;
  wire _42266_;
  wire _42267_;
  wire _42268_;
  wire _42269_;
  wire _42270_;
  wire _42271_;
  wire _42272_;
  wire _42273_;
  wire _42274_;
  wire _42275_;
  wire _42276_;
  wire _42277_;
  wire _42278_;
  wire _42279_;
  wire _42280_;
  wire _42281_;
  wire _42282_;
  wire _42283_;
  wire _42284_;
  wire _42285_;
  wire _42286_;
  wire _42287_;
  wire _42288_;
  wire _42289_;
  wire _42290_;
  wire _42291_;
  wire _42292_;
  wire _42293_;
  wire _42294_;
  wire _42295_;
  wire _42296_;
  wire _42297_;
  wire _42298_;
  wire _42299_;
  wire _42300_;
  wire _42301_;
  wire _42302_;
  wire _42303_;
  wire _42304_;
  wire _42305_;
  wire _42306_;
  wire _42307_;
  wire _42308_;
  wire _42309_;
  wire _42310_;
  wire _42311_;
  wire _42312_;
  wire _42313_;
  wire _42314_;
  wire _42315_;
  wire _42316_;
  wire _42317_;
  wire _42318_;
  wire _42319_;
  wire _42320_;
  wire _42321_;
  wire _42322_;
  wire _42323_;
  wire _42324_;
  wire _42325_;
  wire _42326_;
  wire _42327_;
  wire _42328_;
  wire _42329_;
  wire _42330_;
  wire _42331_;
  wire _42332_;
  wire _42333_;
  wire _42334_;
  wire _42335_;
  wire _42336_;
  wire _42337_;
  wire _42338_;
  wire _42339_;
  wire _42340_;
  wire _42341_;
  wire _42342_;
  wire _42343_;
  wire _42344_;
  wire _42345_;
  wire _42346_;
  wire _42347_;
  wire _42348_;
  wire _42349_;
  wire _42350_;
  wire _42351_;
  wire _42352_;
  wire _42353_;
  wire _42354_;
  wire _42355_;
  wire _42356_;
  wire _42357_;
  wire _42358_;
  wire _42359_;
  wire _42360_;
  wire _42361_;
  wire _42362_;
  wire _42363_;
  wire _42364_;
  wire _42365_;
  wire _42366_;
  wire _42367_;
  wire _42368_;
  wire _42369_;
  wire _42370_;
  wire _42371_;
  wire _42372_;
  wire _42373_;
  wire _42374_;
  wire _42375_;
  wire _42376_;
  wire _42377_;
  wire _42378_;
  wire _42379_;
  wire _42380_;
  wire _42381_;
  wire _42382_;
  wire _42383_;
  wire _42384_;
  wire _42385_;
  wire _42386_;
  wire _42387_;
  wire _42388_;
  wire _42389_;
  wire _42390_;
  wire _42391_;
  wire _42392_;
  wire _42393_;
  wire _42394_;
  wire _42395_;
  wire _42396_;
  wire _42397_;
  wire _42398_;
  wire _42399_;
  wire _42400_;
  wire _42401_;
  wire _42402_;
  wire _42403_;
  wire _42404_;
  wire _42405_;
  wire _42406_;
  wire _42407_;
  wire _42408_;
  wire _42409_;
  wire _42410_;
  wire _42411_;
  wire _42412_;
  wire _42413_;
  wire _42414_;
  wire _42415_;
  wire _42416_;
  wire _42417_;
  wire _42418_;
  wire _42419_;
  wire _42420_;
  wire _42421_;
  wire _42422_;
  wire _42423_;
  wire _42424_;
  wire _42425_;
  wire _42426_;
  wire _42427_;
  wire _42428_;
  wire _42429_;
  wire _42430_;
  wire _42431_;
  wire _42432_;
  wire _42433_;
  wire _42434_;
  wire _42435_;
  wire _42436_;
  wire _42437_;
  wire _42438_;
  wire _42439_;
  wire _42440_;
  wire _42441_;
  wire _42442_;
  wire _42443_;
  wire _42444_;
  wire _42445_;
  wire _42446_;
  wire _42447_;
  wire _42448_;
  wire _42449_;
  wire _42450_;
  wire _42451_;
  wire _42452_;
  wire _42453_;
  wire _42454_;
  wire _42455_;
  wire _42456_;
  wire _42457_;
  wire _42458_;
  wire _42459_;
  wire _42460_;
  wire _42461_;
  wire _42462_;
  wire _42463_;
  wire _42464_;
  wire _42465_;
  wire _42466_;
  wire _42467_;
  wire _42468_;
  wire _42469_;
  wire _42470_;
  wire _42471_;
  wire _42472_;
  wire _42473_;
  wire _42474_;
  wire _42475_;
  wire _42476_;
  wire _42477_;
  wire _42478_;
  wire _42479_;
  wire _42480_;
  wire _42481_;
  wire _42482_;
  wire _42483_;
  wire _42484_;
  wire _42485_;
  wire _42486_;
  wire _42487_;
  wire _42488_;
  wire _42489_;
  wire _42490_;
  wire _42491_;
  wire _42492_;
  wire _42493_;
  wire _42494_;
  wire _42495_;
  wire _42496_;
  wire _42497_;
  wire _42498_;
  wire _42499_;
  wire _42500_;
  wire _42501_;
  wire _42502_;
  wire _42503_;
  wire _42504_;
  wire _42505_;
  wire _42506_;
  wire _42507_;
  wire _42508_;
  wire _42509_;
  wire _42510_;
  wire _42511_;
  wire _42512_;
  wire _42513_;
  wire _42514_;
  wire _42515_;
  wire _42516_;
  wire _42517_;
  wire _42518_;
  wire _42519_;
  wire _42520_;
  wire _42521_;
  wire _42522_;
  wire _42523_;
  wire _42524_;
  wire _42525_;
  wire _42526_;
  wire _42527_;
  wire _42528_;
  wire _42529_;
  wire _42530_;
  wire _42531_;
  wire _42532_;
  wire _42533_;
  wire _42534_;
  wire _42535_;
  wire _42536_;
  wire _42537_;
  wire _42538_;
  wire _42539_;
  wire _42540_;
  wire _42541_;
  wire _42542_;
  wire _42543_;
  wire _42544_;
  wire _42545_;
  wire _42546_;
  wire _42547_;
  wire _42548_;
  wire _42549_;
  wire _42550_;
  wire _42551_;
  wire _42552_;
  wire _42553_;
  wire _42554_;
  wire _42555_;
  wire _42556_;
  wire _42557_;
  wire _42558_;
  wire _42559_;
  wire _42560_;
  wire _42561_;
  wire _42562_;
  wire _42563_;
  wire _42564_;
  wire _42565_;
  wire _42566_;
  wire _42567_;
  wire _42568_;
  wire _42569_;
  wire _42570_;
  wire _42571_;
  wire _42572_;
  wire _42573_;
  wire _42574_;
  wire _42575_;
  wire _42576_;
  wire _42577_;
  wire _42578_;
  wire _42579_;
  wire _42580_;
  wire _42581_;
  wire _42582_;
  wire _42583_;
  wire _42584_;
  wire _42585_;
  wire _42586_;
  wire _42587_;
  wire _42588_;
  wire _42589_;
  wire _42590_;
  wire _42591_;
  wire _42592_;
  wire _42593_;
  wire _42594_;
  wire _42595_;
  wire _42596_;
  wire _42597_;
  wire _42598_;
  wire _42599_;
  wire _42600_;
  wire _42601_;
  wire _42602_;
  wire _42603_;
  wire _42604_;
  wire _42605_;
  wire _42606_;
  wire _42607_;
  wire _42608_;
  wire _42609_;
  wire _42610_;
  wire _42611_;
  wire _42612_;
  wire _42613_;
  wire _42614_;
  wire _42615_;
  wire _42616_;
  wire _42617_;
  wire _42618_;
  wire _42619_;
  wire _42620_;
  wire _42621_;
  wire _42622_;
  wire _42623_;
  wire _42624_;
  wire _42625_;
  wire _42626_;
  wire _42627_;
  wire _42628_;
  wire _42629_;
  wire _42630_;
  wire _42631_;
  wire _42632_;
  wire _42633_;
  wire _42634_;
  wire _42635_;
  wire _42636_;
  wire _42637_;
  wire _42638_;
  wire _42639_;
  wire _42640_;
  wire _42641_;
  wire _42642_;
  wire _42643_;
  wire _42644_;
  wire _42645_;
  wire _42646_;
  wire _42647_;
  wire _42648_;
  wire _42649_;
  wire _42650_;
  wire _42651_;
  wire _42652_;
  wire _42653_;
  wire _42654_;
  wire _42655_;
  wire _42656_;
  wire _42657_;
  wire _42658_;
  wire _42659_;
  wire _42660_;
  wire _42661_;
  wire _42662_;
  wire _42663_;
  wire _42664_;
  wire _42665_;
  wire _42666_;
  wire _42667_;
  wire _42668_;
  wire _42669_;
  wire _42670_;
  wire _42671_;
  wire _42672_;
  wire _42673_;
  wire _42674_;
  wire _42675_;
  wire _42676_;
  wire _42677_;
  wire _42678_;
  wire _42679_;
  wire _42680_;
  wire _42681_;
  wire _42682_;
  wire _42683_;
  wire _42684_;
  wire _42685_;
  wire _42686_;
  wire _42687_;
  wire _42688_;
  wire _42689_;
  wire _42690_;
  wire _42691_;
  wire _42692_;
  wire _42693_;
  wire _42694_;
  wire _42695_;
  wire _42696_;
  wire _42697_;
  wire _42698_;
  wire _42699_;
  wire _42700_;
  wire _42701_;
  wire _42702_;
  wire _42703_;
  wire _42704_;
  wire _42705_;
  wire _42706_;
  wire _42707_;
  wire _42708_;
  wire _42709_;
  wire _42710_;
  wire _42711_;
  wire _42712_;
  wire _42713_;
  wire _42714_;
  wire _42715_;
  wire _42716_;
  wire _42717_;
  wire _42718_;
  wire _42719_;
  wire _42720_;
  wire _42721_;
  wire _42722_;
  wire _42723_;
  wire _42724_;
  wire _42725_;
  wire _42726_;
  wire _42727_;
  wire _42728_;
  wire _42729_;
  wire _42730_;
  wire _42731_;
  wire _42732_;
  wire _42733_;
  wire _42734_;
  wire _42735_;
  wire _42736_;
  wire _42737_;
  wire _42738_;
  wire _42739_;
  wire _42740_;
  wire _42741_;
  wire _42742_;
  wire _42743_;
  wire _42744_;
  wire _42745_;
  wire _42746_;
  wire _42747_;
  wire _42748_;
  wire _42749_;
  wire _42750_;
  wire _42751_;
  wire _42752_;
  wire _42753_;
  wire _42754_;
  wire _42755_;
  wire _42756_;
  wire _42757_;
  wire _42758_;
  wire _42759_;
  wire _42760_;
  wire _42761_;
  wire _42762_;
  wire _42763_;
  wire _42764_;
  wire _42765_;
  wire _42766_;
  wire _42767_;
  wire _42768_;
  wire _42769_;
  wire _42770_;
  wire _42771_;
  wire _42772_;
  wire _42773_;
  wire _42774_;
  wire _42775_;
  wire _42776_;
  wire _42777_;
  wire _42778_;
  wire _42779_;
  wire _42780_;
  wire _42781_;
  wire _42782_;
  wire _42783_;
  wire _42784_;
  wire _42785_;
  wire _42786_;
  wire _42787_;
  wire _42788_;
  wire _42789_;
  wire _42790_;
  wire _42791_;
  wire _42792_;
  wire _42793_;
  wire _42794_;
  wire _42795_;
  wire _42796_;
  wire _42797_;
  wire _42798_;
  wire _42799_;
  wire _42800_;
  wire _42801_;
  wire _42802_;
  wire _42803_;
  wire _42804_;
  wire _42805_;
  wire _42806_;
  wire _42807_;
  wire _42808_;
  wire _42809_;
  wire _42810_;
  wire _42811_;
  wire _42812_;
  wire _42813_;
  wire _42814_;
  wire _42815_;
  wire _42816_;
  wire _42817_;
  wire _42818_;
  wire _42819_;
  wire _42820_;
  wire _42821_;
  wire _42822_;
  wire _42823_;
  wire _42824_;
  wire _42825_;
  wire _42826_;
  wire _42827_;
  wire _42828_;
  wire _42829_;
  wire _42830_;
  wire _42831_;
  wire _42832_;
  wire _42833_;
  wire _42834_;
  wire _42835_;
  wire _42836_;
  wire _42837_;
  wire _42838_;
  wire _42839_;
  wire _42840_;
  wire _42841_;
  wire _42842_;
  wire _42843_;
  wire _42844_;
  wire _42845_;
  wire _42846_;
  wire _42847_;
  wire _42848_;
  wire _42849_;
  wire _42850_;
  wire _42851_;
  wire _42852_;
  wire _42853_;
  wire _42854_;
  wire _42855_;
  wire _42856_;
  wire _42857_;
  wire _42858_;
  wire _42859_;
  wire _42860_;
  wire _42861_;
  wire _42862_;
  wire _42863_;
  wire _42864_;
  wire _42865_;
  wire _42866_;
  wire _42867_;
  wire _42868_;
  wire _42869_;
  wire _42870_;
  wire _42871_;
  wire _42872_;
  wire _42873_;
  wire _42874_;
  wire _42875_;
  wire _42876_;
  wire _42877_;
  wire _42878_;
  wire _42879_;
  wire _42880_;
  wire _42881_;
  wire _42882_;
  wire _42883_;
  wire _42884_;
  wire _42885_;
  wire _42886_;
  wire _42887_;
  wire _42888_;
  wire _42889_;
  wire _42890_;
  wire _42891_;
  wire _42892_;
  wire _42893_;
  wire _42894_;
  wire _42895_;
  wire _42896_;
  wire _42897_;
  wire _42898_;
  wire _42899_;
  wire _42900_;
  wire _42901_;
  wire _42902_;
  wire _42903_;
  wire _42904_;
  wire _42905_;
  wire _42906_;
  wire _42907_;
  wire _42908_;
  wire _42909_;
  wire _42910_;
  wire _42911_;
  wire _42912_;
  wire _42913_;
  wire _42914_;
  wire _42915_;
  wire _42916_;
  wire _42917_;
  wire _42918_;
  wire _42919_;
  wire _42920_;
  wire _42921_;
  wire _42922_;
  wire _42923_;
  wire _42924_;
  wire _42925_;
  wire _42926_;
  wire _42927_;
  wire _42928_;
  wire _42929_;
  wire _42930_;
  wire _42931_;
  wire _42932_;
  wire _42933_;
  wire _42934_;
  wire _42935_;
  wire _42936_;
  wire _42937_;
  wire _42938_;
  wire _42939_;
  wire _42940_;
  wire _42941_;
  wire _42942_;
  wire _42943_;
  wire _42944_;
  wire _42945_;
  wire _42946_;
  wire _42947_;
  wire _42948_;
  wire _42949_;
  wire _42950_;
  wire _42951_;
  wire _42952_;
  wire _42953_;
  wire _42954_;
  wire _42955_;
  wire _42956_;
  wire _42957_;
  wire _42958_;
  wire _42959_;
  wire _42960_;
  wire _42961_;
  wire _42962_;
  wire _42963_;
  wire _42964_;
  wire _42965_;
  wire _42966_;
  wire _42967_;
  wire _42968_;
  wire _42969_;
  wire _42970_;
  wire _42971_;
  wire _42972_;
  wire _42973_;
  wire _42974_;
  wire _42975_;
  wire _42976_;
  wire _42977_;
  wire _42978_;
  wire _42979_;
  wire _42980_;
  wire _42981_;
  wire _42982_;
  wire _42983_;
  wire _42984_;
  wire _42985_;
  wire _42986_;
  wire _42987_;
  wire _42988_;
  wire _42989_;
  wire _42990_;
  wire _42991_;
  wire _42992_;
  wire _42993_;
  wire _42994_;
  wire _42995_;
  wire _42996_;
  wire _42997_;
  wire _42998_;
  wire _42999_;
  wire _43000_;
  wire _43001_;
  wire _43002_;
  wire _43003_;
  wire _43004_;
  wire _43005_;
  wire _43006_;
  wire _43007_;
  wire _43008_;
  wire _43009_;
  wire _43010_;
  wire _43011_;
  wire _43012_;
  wire _43013_;
  wire _43014_;
  wire _43015_;
  wire _43016_;
  wire _43017_;
  wire _43018_;
  wire _43019_;
  wire _43020_;
  wire _43021_;
  wire _43022_;
  wire _43023_;
  wire _43024_;
  wire _43025_;
  wire _43026_;
  wire _43027_;
  wire _43028_;
  wire _43029_;
  wire _43030_;
  wire _43031_;
  wire _43032_;
  wire _43033_;
  wire _43034_;
  wire _43035_;
  wire _43036_;
  wire _43037_;
  wire _43038_;
  wire _43039_;
  wire _43040_;
  wire _43041_;
  wire _43042_;
  wire _43043_;
  wire _43044_;
  wire _43045_;
  wire _43046_;
  wire _43047_;
  wire _43048_;
  wire _43049_;
  wire _43050_;
  wire _43051_;
  wire _43052_;
  wire _43053_;
  wire _43054_;
  wire _43055_;
  wire _43056_;
  wire _43057_;
  wire _43058_;
  wire _43059_;
  wire _43060_;
  wire _43061_;
  wire _43062_;
  wire _43063_;
  wire _43064_;
  wire _43065_;
  wire _43066_;
  wire _43067_;
  wire _43068_;
  wire _43069_;
  wire _43070_;
  wire _43071_;
  wire _43072_;
  wire _43073_;
  wire _43074_;
  wire _43075_;
  wire _43076_;
  wire _43077_;
  wire _43078_;
  wire _43079_;
  wire _43080_;
  wire _43081_;
  wire _43082_;
  wire _43083_;
  wire _43084_;
  wire _43085_;
  wire _43086_;
  wire _43087_;
  wire _43088_;
  wire _43089_;
  wire _43090_;
  wire _43091_;
  wire _43092_;
  wire _43093_;
  wire _43094_;
  wire _43095_;
  wire _43096_;
  wire _43097_;
  wire _43098_;
  wire _43099_;
  wire _43100_;
  wire _43101_;
  wire _43102_;
  wire _43103_;
  wire _43104_;
  wire _43105_;
  wire _43106_;
  wire _43107_;
  wire _43108_;
  wire _43109_;
  wire _43110_;
  wire _43111_;
  wire _43112_;
  wire _43113_;
  wire _43114_;
  wire _43115_;
  wire _43116_;
  wire _43117_;
  wire _43118_;
  wire _43119_;
  wire _43120_;
  wire _43121_;
  wire _43122_;
  wire _43123_;
  wire _43124_;
  wire _43125_;
  wire _43126_;
  wire _43127_;
  wire _43128_;
  wire _43129_;
  wire _43130_;
  wire _43131_;
  wire _43132_;
  wire _43133_;
  wire _43134_;
  wire _43135_;
  wire _43136_;
  wire _43137_;
  wire _43138_;
  wire _43139_;
  wire _43140_;
  wire _43141_;
  wire _43142_;
  wire _43143_;
  wire _43144_;
  wire _43145_;
  wire _43146_;
  wire _43147_;
  wire _43148_;
  wire _43149_;
  wire _43150_;
  wire _43151_;
  wire _43152_;
  wire _43153_;
  wire _43154_;
  wire _43155_;
  wire _43156_;
  wire _43157_;
  wire _43158_;
  wire _43159_;
  wire _43160_;
  wire _43161_;
  wire _43162_;
  wire _43163_;
  wire _43164_;
  wire _43165_;
  wire _43166_;
  wire _43167_;
  wire _43168_;
  wire _43169_;
  wire _43170_;
  wire _43171_;
  wire _43172_;
  wire _43173_;
  wire _43174_;
  wire _43175_;
  wire _43176_;
  wire _43177_;
  wire _43178_;
  wire _43179_;
  wire _43180_;
  wire _43181_;
  wire _43182_;
  wire _43183_;
  wire _43184_;
  wire _43185_;
  wire _43186_;
  wire _43187_;
  wire _43188_;
  wire _43189_;
  wire _43190_;
  wire _43191_;
  wire _43192_;
  wire _43193_;
  wire _43194_;
  wire _43195_;
  wire _43196_;
  wire _43197_;
  wire _43198_;
  wire _43199_;
  wire _43200_;
  wire _43201_;
  wire _43202_;
  wire _43203_;
  wire _43204_;
  wire _43205_;
  wire _43206_;
  wire _43207_;
  wire _43208_;
  wire _43209_;
  wire _43210_;
  wire _43211_;
  wire _43212_;
  wire _43213_;
  wire _43214_;
  wire _43215_;
  wire _43216_;
  wire _43217_;
  wire _43218_;
  wire _43219_;
  wire _43220_;
  wire _43221_;
  wire _43222_;
  wire _43223_;
  wire _43224_;
  wire _43225_;
  wire _43226_;
  wire _43227_;
  wire _43228_;
  wire _43229_;
  wire _43230_;
  wire _43231_;
  wire _43232_;
  wire _43233_;
  wire _43234_;
  wire _43235_;
  wire _43236_;
  wire _43237_;
  wire _43238_;
  wire _43239_;
  wire _43240_;
  wire _43241_;
  wire _43242_;
  wire _43243_;
  wire _43244_;
  wire _43245_;
  wire _43246_;
  wire _43247_;
  wire _43248_;
  wire _43249_;
  wire _43250_;
  wire _43251_;
  wire _43252_;
  wire _43253_;
  wire _43254_;
  wire _43255_;
  wire _43256_;
  wire _43257_;
  wire _43258_;
  wire _43259_;
  wire _43260_;
  wire _43261_;
  wire _43262_;
  wire _43263_;
  wire _43264_;
  wire _43265_;
  wire _43266_;
  wire _43267_;
  wire _43268_;
  wire _43269_;
  wire _43270_;
  wire _43271_;
  wire _43272_;
  wire _43273_;
  wire _43274_;
  wire _43275_;
  wire _43276_;
  wire _43277_;
  wire _43278_;
  wire _43279_;
  wire _43280_;
  wire _43281_;
  wire _43282_;
  wire _43283_;
  wire _43284_;
  wire _43285_;
  wire _43286_;
  wire _43287_;
  wire _43288_;
  wire _43289_;
  wire _43290_;
  wire _43291_;
  wire _43292_;
  wire _43293_;
  wire _43294_;
  wire _43295_;
  wire _43296_;
  wire _43297_;
  wire _43298_;
  wire _43299_;
  wire _43300_;
  wire _43301_;
  wire _43302_;
  wire _43303_;
  wire _43304_;
  wire _43305_;
  wire _43306_;
  wire _43307_;
  wire _43308_;
  wire _43309_;
  wire _43310_;
  wire _43311_;
  wire _43312_;
  wire _43313_;
  wire _43314_;
  wire _43315_;
  wire _43316_;
  wire _43317_;
  wire _43318_;
  wire _43319_;
  wire _43320_;
  wire _43321_;
  wire _43322_;
  wire _43323_;
  wire _43324_;
  wire _43325_;
  wire _43326_;
  wire _43327_;
  wire _43328_;
  wire _43329_;
  wire _43330_;
  wire _43331_;
  wire _43332_;
  wire _43333_;
  wire _43334_;
  wire _43335_;
  wire _43336_;
  wire _43337_;
  wire _43338_;
  wire _43339_;
  wire _43340_;
  wire _43341_;
  wire _43342_;
  wire _43343_;
  wire _43344_;
  wire _43345_;
  wire _43346_;
  wire _43347_;
  wire _43348_;
  wire _43349_;
  wire _43350_;
  wire _43351_;
  wire _43352_;
  wire _43353_;
  wire _43354_;
  wire _43355_;
  wire _43356_;
  wire _43357_;
  wire _43358_;
  wire _43359_;
  wire _43360_;
  wire _43361_;
  wire _43362_;
  wire _43363_;
  wire _43364_;
  wire _43365_;
  wire _43366_;
  wire _43367_;
  wire _43368_;
  wire _43369_;
  wire _43370_;
  wire _43371_;
  wire _43372_;
  wire _43373_;
  wire _43374_;
  wire _43375_;
  wire _43376_;
  wire _43377_;
  wire _43378_;
  wire _43379_;
  wire _43380_;
  wire _43381_;
  wire _43382_;
  wire _43383_;
  wire _43384_;
  wire _43385_;
  wire _43386_;
  wire _43387_;
  wire _43388_;
  wire _43389_;
  wire _43390_;
  wire _43391_;
  wire _43392_;
  wire _43393_;
  wire _43394_;
  wire _43395_;
  wire _43396_;
  wire _43397_;
  wire _43398_;
  wire _43399_;
  wire _43400_;
  wire _43401_;
  wire _43402_;
  wire _43403_;
  wire _43404_;
  wire _43405_;
  wire _43406_;
  wire _43407_;
  wire _43408_;
  wire _43409_;
  wire _43410_;
  wire _43411_;
  wire _43412_;
  wire _43413_;
  wire _43414_;
  wire _43415_;
  wire _43416_;
  wire _43417_;
  wire _43418_;
  wire _43419_;
  wire _43420_;
  wire _43421_;
  wire _43422_;
  wire _43423_;
  wire _43424_;
  wire _43425_;
  wire _43426_;
  wire _43427_;
  wire _43428_;
  wire _43429_;
  wire _43430_;
  wire _43431_;
  wire _43432_;
  wire _43433_;
  wire _43434_;
  wire _43435_;
  wire _43436_;
  wire _43437_;
  wire _43438_;
  wire _43439_;
  wire _43440_;
  wire _43441_;
  wire _43442_;
  wire _43443_;
  wire _43444_;
  wire _43445_;
  wire _43446_;
  wire _43447_;
  wire _43448_;
  wire _43449_;
  wire _43450_;
  wire _43451_;
  wire _43452_;
  wire _43453_;
  wire _43454_;
  wire _43455_;
  wire _43456_;
  wire _43457_;
  wire _43458_;
  wire _43459_;
  wire _43460_;
  wire _43461_;
  wire _43462_;
  wire _43463_;
  wire _43464_;
  wire _43465_;
  wire _43466_;
  wire _43467_;
  wire _43468_;
  wire _43469_;
  wire _43470_;
  wire _43471_;
  wire _43472_;
  wire _43473_;
  wire _43474_;
  wire _43475_;
  wire _43476_;
  wire _43477_;
  wire _43478_;
  wire _43479_;
  wire _43480_;
  wire _43481_;
  wire _43482_;
  wire _43483_;
  wire _43484_;
  wire _43485_;
  wire _43486_;
  wire _43487_;
  wire _43488_;
  wire _43489_;
  wire _43490_;
  wire _43491_;
  wire _43492_;
  wire _43493_;
  wire _43494_;
  wire _43495_;
  wire _43496_;
  wire _43497_;
  wire _43498_;
  wire _43499_;
  wire _43500_;
  wire _43501_;
  wire _43502_;
  wire _43503_;
  wire _43504_;
  wire _43505_;
  wire _43506_;
  wire _43507_;
  wire _43508_;
  wire _43509_;
  wire _43510_;
  wire _43511_;
  wire _43512_;
  wire _43513_;
  wire _43514_;
  wire _43515_;
  wire _43516_;
  wire _43517_;
  wire _43518_;
  wire _43519_;
  wire _43520_;
  wire _43521_;
  wire _43522_;
  wire _43523_;
  wire _43524_;
  wire _43525_;
  wire _43526_;
  wire _43527_;
  wire _43528_;
  wire _43529_;
  wire _43530_;
  wire _43531_;
  wire _43532_;
  wire _43533_;
  wire [7:0] ACC_gm;
  wire [7:0] acc;
  input clk;
  wire [31:0] cxrom_data_out;
  wire \oc8051_gm_cxrom_1.cell0.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell0.data ;
  wire \oc8051_gm_cxrom_1.cell0.rst ;
  wire \oc8051_gm_cxrom_1.cell0.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell0.word ;
  wire \oc8051_gm_cxrom_1.cell1.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell1.data ;
  wire \oc8051_gm_cxrom_1.cell1.rst ;
  wire \oc8051_gm_cxrom_1.cell1.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell1.word ;
  wire \oc8051_gm_cxrom_1.cell10.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell10.data ;
  wire \oc8051_gm_cxrom_1.cell10.rst ;
  wire \oc8051_gm_cxrom_1.cell10.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell10.word ;
  wire \oc8051_gm_cxrom_1.cell11.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell11.data ;
  wire \oc8051_gm_cxrom_1.cell11.rst ;
  wire \oc8051_gm_cxrom_1.cell11.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell11.word ;
  wire \oc8051_gm_cxrom_1.cell12.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell12.data ;
  wire \oc8051_gm_cxrom_1.cell12.rst ;
  wire \oc8051_gm_cxrom_1.cell12.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell12.word ;
  wire \oc8051_gm_cxrom_1.cell13.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell13.data ;
  wire \oc8051_gm_cxrom_1.cell13.rst ;
  wire \oc8051_gm_cxrom_1.cell13.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell13.word ;
  wire \oc8051_gm_cxrom_1.cell14.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell14.data ;
  wire \oc8051_gm_cxrom_1.cell14.rst ;
  wire \oc8051_gm_cxrom_1.cell14.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell14.word ;
  wire \oc8051_gm_cxrom_1.cell15.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell15.data ;
  wire \oc8051_gm_cxrom_1.cell15.rst ;
  wire \oc8051_gm_cxrom_1.cell15.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell15.word ;
  wire \oc8051_gm_cxrom_1.cell2.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell2.data ;
  wire \oc8051_gm_cxrom_1.cell2.rst ;
  wire \oc8051_gm_cxrom_1.cell2.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell2.word ;
  wire \oc8051_gm_cxrom_1.cell3.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell3.data ;
  wire \oc8051_gm_cxrom_1.cell3.rst ;
  wire \oc8051_gm_cxrom_1.cell3.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell3.word ;
  wire \oc8051_gm_cxrom_1.cell4.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell4.data ;
  wire \oc8051_gm_cxrom_1.cell4.rst ;
  wire \oc8051_gm_cxrom_1.cell4.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell4.word ;
  wire \oc8051_gm_cxrom_1.cell5.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell5.data ;
  wire \oc8051_gm_cxrom_1.cell5.rst ;
  wire \oc8051_gm_cxrom_1.cell5.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell5.word ;
  wire \oc8051_gm_cxrom_1.cell6.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell6.data ;
  wire \oc8051_gm_cxrom_1.cell6.rst ;
  wire \oc8051_gm_cxrom_1.cell6.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell6.word ;
  wire \oc8051_gm_cxrom_1.cell7.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell7.data ;
  wire \oc8051_gm_cxrom_1.cell7.rst ;
  wire \oc8051_gm_cxrom_1.cell7.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell7.word ;
  wire \oc8051_gm_cxrom_1.cell8.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell8.data ;
  wire \oc8051_gm_cxrom_1.cell8.rst ;
  wire \oc8051_gm_cxrom_1.cell8.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell8.word ;
  wire \oc8051_gm_cxrom_1.cell9.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell9.data ;
  wire \oc8051_gm_cxrom_1.cell9.rst ;
  wire \oc8051_gm_cxrom_1.cell9.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell9.word ;
  wire \oc8051_gm_cxrom_1.clk ;
  wire [31:0] \oc8051_gm_cxrom_1.cxrom_data_out ;
  wire [15:0] \oc8051_gm_cxrom_1.rd_addr_0 ;
  wire \oc8051_gm_cxrom_1.rst ;
  wire [127:0] \oc8051_gm_cxrom_1.word_in ;
  wire [7:0] \oc8051_golden_model_1.ACC ;
  wire [7:0] \oc8051_golden_model_1.ACC_03 ;
  wire [7:0] \oc8051_golden_model_1.ACC_13 ;
  wire [7:0] \oc8051_golden_model_1.ACC_23 ;
  wire [7:0] \oc8051_golden_model_1.ACC_33 ;
  wire [7:0] \oc8051_golden_model_1.ACC_c4 ;
  wire [7:0] \oc8051_golden_model_1.ACC_d6 ;
  wire [7:0] \oc8051_golden_model_1.ACC_d7 ;
  wire [7:0] \oc8051_golden_model_1.ACC_e4 ;
  wire [7:0] \oc8051_golden_model_1.B ;
  wire [7:0] \oc8051_golden_model_1.DPH ;
  wire [7:0] \oc8051_golden_model_1.DPL ;
  wire [7:0] \oc8051_golden_model_1.IE ;
  wire [7:0] \oc8051_golden_model_1.IP ;
  wire [7:0] \oc8051_golden_model_1.IRAM[0] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[10] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[11] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[12] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[13] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[14] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[15] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[1] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[2] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[3] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[4] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[5] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[6] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[7] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[8] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[9] ;
  wire [7:0] \oc8051_golden_model_1.P0 ;
  wire [7:0] \oc8051_golden_model_1.P1 ;
  wire [7:0] \oc8051_golden_model_1.P2 ;
  wire [7:0] \oc8051_golden_model_1.P3 ;
  wire [15:0] \oc8051_golden_model_1.PC ;
  wire [7:0] \oc8051_golden_model_1.PCON ;
  wire [15:0] \oc8051_golden_model_1.PC_22 ;
  wire [15:0] \oc8051_golden_model_1.PC_32 ;
  wire [7:0] \oc8051_golden_model_1.PSW ;
  wire [7:0] \oc8051_golden_model_1.PSW_13 ;
  wire [7:0] \oc8051_golden_model_1.PSW_24 ;
  wire [7:0] \oc8051_golden_model_1.PSW_25 ;
  wire [7:0] \oc8051_golden_model_1.PSW_26 ;
  wire [7:0] \oc8051_golden_model_1.PSW_27 ;
  wire [7:0] \oc8051_golden_model_1.PSW_28 ;
  wire [7:0] \oc8051_golden_model_1.PSW_29 ;
  wire [7:0] \oc8051_golden_model_1.PSW_2a ;
  wire [7:0] \oc8051_golden_model_1.PSW_2b ;
  wire [7:0] \oc8051_golden_model_1.PSW_2c ;
  wire [7:0] \oc8051_golden_model_1.PSW_2d ;
  wire [7:0] \oc8051_golden_model_1.PSW_2e ;
  wire [7:0] \oc8051_golden_model_1.PSW_2f ;
  wire [7:0] \oc8051_golden_model_1.PSW_33 ;
  wire [7:0] \oc8051_golden_model_1.PSW_34 ;
  wire [7:0] \oc8051_golden_model_1.PSW_35 ;
  wire [7:0] \oc8051_golden_model_1.PSW_36 ;
  wire [7:0] \oc8051_golden_model_1.PSW_37 ;
  wire [7:0] \oc8051_golden_model_1.PSW_38 ;
  wire [7:0] \oc8051_golden_model_1.PSW_39 ;
  wire [7:0] \oc8051_golden_model_1.PSW_3a ;
  wire [7:0] \oc8051_golden_model_1.PSW_3b ;
  wire [7:0] \oc8051_golden_model_1.PSW_3c ;
  wire [7:0] \oc8051_golden_model_1.PSW_3d ;
  wire [7:0] \oc8051_golden_model_1.PSW_3e ;
  wire [7:0] \oc8051_golden_model_1.PSW_3f ;
  wire [7:0] \oc8051_golden_model_1.PSW_72 ;
  wire [7:0] \oc8051_golden_model_1.PSW_82 ;
  wire [7:0] \oc8051_golden_model_1.PSW_84 ;
  wire [7:0] \oc8051_golden_model_1.PSW_94 ;
  wire [7:0] \oc8051_golden_model_1.PSW_95 ;
  wire [7:0] \oc8051_golden_model_1.PSW_96 ;
  wire [7:0] \oc8051_golden_model_1.PSW_97 ;
  wire [7:0] \oc8051_golden_model_1.PSW_98 ;
  wire [7:0] \oc8051_golden_model_1.PSW_99 ;
  wire [7:0] \oc8051_golden_model_1.PSW_9a ;
  wire [7:0] \oc8051_golden_model_1.PSW_9b ;
  wire [7:0] \oc8051_golden_model_1.PSW_9c ;
  wire [7:0] \oc8051_golden_model_1.PSW_9d ;
  wire [7:0] \oc8051_golden_model_1.PSW_9e ;
  wire [7:0] \oc8051_golden_model_1.PSW_9f ;
  wire [7:0] \oc8051_golden_model_1.PSW_a0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a2 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_ba ;
  wire [7:0] \oc8051_golden_model_1.PSW_bb ;
  wire [7:0] \oc8051_golden_model_1.PSW_bc ;
  wire [7:0] \oc8051_golden_model_1.PSW_bd ;
  wire [7:0] \oc8051_golden_model_1.PSW_be ;
  wire [7:0] \oc8051_golden_model_1.PSW_bf ;
  wire [7:0] \oc8051_golden_model_1.PSW_c3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d4 ;
  wire [7:0] \oc8051_golden_model_1.RD_IRAM_0 ;
  wire [7:0] \oc8051_golden_model_1.RD_IRAM_1 ;
  wire [3:0] \oc8051_golden_model_1.RD_IRAM_ADDR ;
  wire [15:0] \oc8051_golden_model_1.RD_ROM_0_ADDR ;
  wire [7:0] \oc8051_golden_model_1.SBUF ;
  wire [7:0] \oc8051_golden_model_1.SCON ;
  wire [7:0] \oc8051_golden_model_1.SP ;
  wire [7:0] \oc8051_golden_model_1.TCON ;
  wire [7:0] \oc8051_golden_model_1.TH0 ;
  wire [7:0] \oc8051_golden_model_1.TH1 ;
  wire [7:0] \oc8051_golden_model_1.TL0 ;
  wire [7:0] \oc8051_golden_model_1.TL1 ;
  wire [7:0] \oc8051_golden_model_1.TMOD ;
  wire \oc8051_golden_model_1.clk ;
  wire [1:0] \oc8051_golden_model_1.n0006 ;
  wire [7:0] \oc8051_golden_model_1.n0007 ;
  wire [7:0] \oc8051_golden_model_1.n0011 ;
  wire [7:0] \oc8051_golden_model_1.n0019 ;
  wire [7:0] \oc8051_golden_model_1.n0023 ;
  wire [7:0] \oc8051_golden_model_1.n0027 ;
  wire [7:0] \oc8051_golden_model_1.n0031 ;
  wire [7:0] \oc8051_golden_model_1.n0035 ;
  wire [7:0] \oc8051_golden_model_1.n0039 ;
  wire [7:0] \oc8051_golden_model_1.n0561 ;
  wire [7:0] \oc8051_golden_model_1.n0594 ;
  wire [15:0] \oc8051_golden_model_1.n0701 ;
  wire [15:0] \oc8051_golden_model_1.n0733 ;
  wire [7:0] \oc8051_golden_model_1.n0994 ;
  wire [3:0] \oc8051_golden_model_1.n1071 ;
  wire [3:0] \oc8051_golden_model_1.n1073 ;
  wire [3:0] \oc8051_golden_model_1.n1075 ;
  wire [3:0] \oc8051_golden_model_1.n1076 ;
  wire [3:0] \oc8051_golden_model_1.n1077 ;
  wire [3:0] \oc8051_golden_model_1.n1078 ;
  wire [3:0] \oc8051_golden_model_1.n1079 ;
  wire [3:0] \oc8051_golden_model_1.n1080 ;
  wire [3:0] \oc8051_golden_model_1.n1081 ;
  wire \oc8051_golden_model_1.n1118 ;
  wire \oc8051_golden_model_1.n1146 ;
  wire [8:0] \oc8051_golden_model_1.n1147 ;
  wire [8:0] \oc8051_golden_model_1.n1148 ;
  wire [7:0] \oc8051_golden_model_1.n1149 ;
  wire \oc8051_golden_model_1.n1150 ;
  wire \oc8051_golden_model_1.n1151 ;
  wire [2:0] \oc8051_golden_model_1.n1152 ;
  wire \oc8051_golden_model_1.n1153 ;
  wire [1:0] \oc8051_golden_model_1.n1154 ;
  wire [7:0] \oc8051_golden_model_1.n1155 ;
  wire [15:0] \oc8051_golden_model_1.n1181 ;
  wire [7:0] \oc8051_golden_model_1.n1183 ;
  wire [8:0] \oc8051_golden_model_1.n1185 ;
  wire [8:0] \oc8051_golden_model_1.n1189 ;
  wire \oc8051_golden_model_1.n1190 ;
  wire [3:0] \oc8051_golden_model_1.n1191 ;
  wire [4:0] \oc8051_golden_model_1.n1192 ;
  wire [4:0] \oc8051_golden_model_1.n1196 ;
  wire \oc8051_golden_model_1.n1197 ;
  wire [8:0] \oc8051_golden_model_1.n1198 ;
  wire \oc8051_golden_model_1.n1206 ;
  wire [7:0] \oc8051_golden_model_1.n1207 ;
  wire [8:0] \oc8051_golden_model_1.n1211 ;
  wire \oc8051_golden_model_1.n1212 ;
  wire [4:0] \oc8051_golden_model_1.n1217 ;
  wire \oc8051_golden_model_1.n1218 ;
  wire \oc8051_golden_model_1.n1226 ;
  wire [7:0] \oc8051_golden_model_1.n1227 ;
  wire [8:0] \oc8051_golden_model_1.n1229 ;
  wire [8:0] \oc8051_golden_model_1.n1231 ;
  wire \oc8051_golden_model_1.n1232 ;
  wire [3:0] \oc8051_golden_model_1.n1233 ;
  wire [4:0] \oc8051_golden_model_1.n1234 ;
  wire [4:0] \oc8051_golden_model_1.n1236 ;
  wire \oc8051_golden_model_1.n1237 ;
  wire [8:0] \oc8051_golden_model_1.n1238 ;
  wire \oc8051_golden_model_1.n1245 ;
  wire [7:0] \oc8051_golden_model_1.n1246 ;
  wire [8:0] \oc8051_golden_model_1.n1249 ;
  wire \oc8051_golden_model_1.n1250 ;
  wire \oc8051_golden_model_1.n1257 ;
  wire [7:0] \oc8051_golden_model_1.n1258 ;
  wire [8:0] \oc8051_golden_model_1.n1260 ;
  wire [8:0] \oc8051_golden_model_1.n1262 ;
  wire \oc8051_golden_model_1.n1263 ;
  wire [4:0] \oc8051_golden_model_1.n1264 ;
  wire [4:0] \oc8051_golden_model_1.n1266 ;
  wire \oc8051_golden_model_1.n1267 ;
  wire [8:0] \oc8051_golden_model_1.n1268 ;
  wire \oc8051_golden_model_1.n1275 ;
  wire [7:0] \oc8051_golden_model_1.n1276 ;
  wire [4:0] \oc8051_golden_model_1.n1278 ;
  wire \oc8051_golden_model_1.n1279 ;
  wire [7:0] \oc8051_golden_model_1.n1280 ;
  wire [8:0] \oc8051_golden_model_1.n1282 ;
  wire \oc8051_golden_model_1.n1283 ;
  wire \oc8051_golden_model_1.n1290 ;
  wire [7:0] \oc8051_golden_model_1.n1291 ;
  wire [7:0] \oc8051_golden_model_1.n1292 ;
  wire [8:0] \oc8051_golden_model_1.n1295 ;
  wire [8:0] \oc8051_golden_model_1.n1296 ;
  wire [7:0] \oc8051_golden_model_1.n1297 ;
  wire \oc8051_golden_model_1.n1298 ;
  wire [7:0] \oc8051_golden_model_1.n1299 ;
  wire [7:0] \oc8051_golden_model_1.n1300 ;
  wire [8:0] \oc8051_golden_model_1.n1303 ;
  wire [8:0] \oc8051_golden_model_1.n1305 ;
  wire \oc8051_golden_model_1.n1306 ;
  wire [4:0] \oc8051_golden_model_1.n1307 ;
  wire [4:0] \oc8051_golden_model_1.n1309 ;
  wire \oc8051_golden_model_1.n1310 ;
  wire \oc8051_golden_model_1.n1317 ;
  wire [7:0] \oc8051_golden_model_1.n1318 ;
  wire [8:0] \oc8051_golden_model_1.n1322 ;
  wire \oc8051_golden_model_1.n1323 ;
  wire [4:0] \oc8051_golden_model_1.n1325 ;
  wire \oc8051_golden_model_1.n1326 ;
  wire \oc8051_golden_model_1.n1333 ;
  wire [7:0] \oc8051_golden_model_1.n1334 ;
  wire [8:0] \oc8051_golden_model_1.n1338 ;
  wire \oc8051_golden_model_1.n1339 ;
  wire [4:0] \oc8051_golden_model_1.n1341 ;
  wire \oc8051_golden_model_1.n1342 ;
  wire \oc8051_golden_model_1.n1349 ;
  wire [7:0] \oc8051_golden_model_1.n1350 ;
  wire [8:0] \oc8051_golden_model_1.n1354 ;
  wire \oc8051_golden_model_1.n1355 ;
  wire [4:0] \oc8051_golden_model_1.n1357 ;
  wire \oc8051_golden_model_1.n1358 ;
  wire \oc8051_golden_model_1.n1365 ;
  wire [7:0] \oc8051_golden_model_1.n1366 ;
  wire \oc8051_golden_model_1.n1520 ;
  wire [6:0] \oc8051_golden_model_1.n1521 ;
  wire [7:0] \oc8051_golden_model_1.n1522 ;
  wire \oc8051_golden_model_1.n1545 ;
  wire [7:0] \oc8051_golden_model_1.n1546 ;
  wire [3:0] \oc8051_golden_model_1.n1553 ;
  wire \oc8051_golden_model_1.n1554 ;
  wire [7:0] \oc8051_golden_model_1.n1555 ;
  wire [7:0] \oc8051_golden_model_1.n1680 ;
  wire \oc8051_golden_model_1.n1683 ;
  wire \oc8051_golden_model_1.n1685 ;
  wire \oc8051_golden_model_1.n1691 ;
  wire [7:0] \oc8051_golden_model_1.n1692 ;
  wire \oc8051_golden_model_1.n1696 ;
  wire \oc8051_golden_model_1.n1698 ;
  wire \oc8051_golden_model_1.n1704 ;
  wire [7:0] \oc8051_golden_model_1.n1705 ;
  wire \oc8051_golden_model_1.n1709 ;
  wire \oc8051_golden_model_1.n1711 ;
  wire \oc8051_golden_model_1.n1717 ;
  wire [7:0] \oc8051_golden_model_1.n1718 ;
  wire \oc8051_golden_model_1.n1722 ;
  wire \oc8051_golden_model_1.n1724 ;
  wire \oc8051_golden_model_1.n1730 ;
  wire [7:0] \oc8051_golden_model_1.n1731 ;
  wire \oc8051_golden_model_1.n1733 ;
  wire [7:0] \oc8051_golden_model_1.n1734 ;
  wire [7:0] \oc8051_golden_model_1.n1735 ;
  wire [15:0] \oc8051_golden_model_1.n1739 ;
  wire \oc8051_golden_model_1.n1745 ;
  wire [7:0] \oc8051_golden_model_1.n1746 ;
  wire \oc8051_golden_model_1.n1749 ;
  wire [7:0] \oc8051_golden_model_1.n1750 ;
  wire \oc8051_golden_model_1.n1765 ;
  wire [7:0] \oc8051_golden_model_1.n1766 ;
  wire \oc8051_golden_model_1.n1771 ;
  wire [7:0] \oc8051_golden_model_1.n1772 ;
  wire \oc8051_golden_model_1.n1777 ;
  wire [7:0] \oc8051_golden_model_1.n1778 ;
  wire \oc8051_golden_model_1.n1783 ;
  wire [7:0] \oc8051_golden_model_1.n1784 ;
  wire \oc8051_golden_model_1.n1789 ;
  wire [7:0] \oc8051_golden_model_1.n1790 ;
  wire [7:0] \oc8051_golden_model_1.n1791 ;
  wire [3:0] \oc8051_golden_model_1.n1792 ;
  wire [7:0] \oc8051_golden_model_1.n1793 ;
  wire [7:0] \oc8051_golden_model_1.n1828 ;
  wire \oc8051_golden_model_1.n1847 ;
  wire [7:0] \oc8051_golden_model_1.n1848 ;
  wire [7:0] \oc8051_golden_model_1.n1852 ;
  wire [3:0] \oc8051_golden_model_1.n1853 ;
  wire [7:0] \oc8051_golden_model_1.n1854 ;
  wire \oc8051_golden_model_1.rst ;
  wire [7:0] \oc8051_top_1.acc ;
  wire [31:0] \oc8051_top_1.cxrom_data_out ;
  wire \oc8051_top_1.cy ;
  wire [1:0] \oc8051_top_1.cy_sel ;
  wire [7:0] \oc8051_top_1.dptr_hi ;
  wire [7:0] \oc8051_top_1.dptr_lo ;
  wire \oc8051_top_1.ea_int ;
  wire [31:0] \oc8051_top_1.idat_onchip ;
  wire \oc8051_top_1.int_ack ;
  wire [7:0] \oc8051_top_1.int_src ;
  wire \oc8051_top_1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.mem_act ;
  wire \oc8051_top_1.oc8051_alu1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.divsrc2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.des2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div0 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.div_out ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.rst ;
  wire [5:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.rst ;
  wire [15:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul ;
  wire \oc8051_top_1.oc8051_alu1.rst ;
  wire \oc8051_top_1.oc8051_alu1.srcAc ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.acc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.clk ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.dptr ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op1_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op2_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op3_r ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.pc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_alu_src_sel1.sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_alu_src_sel1.sel2 ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.sel3 ;
  wire [7:0] \oc8051_top_1.oc8051_comp1.acc ;
  wire \oc8051_top_1.oc8051_comp1.cy ;
  wire \oc8051_top_1.oc8051_cy_select1.cy_in ;
  wire [1:0] \oc8051_top_1.oc8051_cy_select1.cy_sel ;
  wire [3:0] \oc8051_top_1.oc8051_decoder1.alu_op ;
  wire \oc8051_top_1.oc8051_decoder1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.cy_sel ;
  wire \oc8051_top_1.oc8051_decoder1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_decoder1.op ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.psw_set ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_wr_sel ;
  wire \oc8051_top_1.oc8051_decoder1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.src_sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.src_sel2 ;
  wire \oc8051_top_1.oc8051_decoder1.src_sel3 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.state ;
  wire \oc8051_top_1.oc8051_decoder1.wait_data ;
  wire \oc8051_top_1.oc8051_decoder1.wr ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.wr_sfr ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[7] ;
  wire \oc8051_top_1.oc8051_indi_addr1.clk ;
  wire \oc8051_top_1.oc8051_indi_addr1.rst ;
  wire \oc8051_top_1.oc8051_indi_addr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.cdata ;
  wire \oc8051_top_1.oc8051_memory_interface1.cdone ;
  wire \oc8051_top_1.oc8051_memory_interface1.clk ;
  wire \oc8051_top_1.oc8051_memory_interface1.dack_ir ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dadr_o ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dadr_ot ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_ir ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.dmem_wait ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dptr ;
  wire \oc8051_top_1.oc8051_memory_interface1.dstb_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.dwe_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.ea_int ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.iadr_t ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_cur ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_old ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_onchip ;
  wire \oc8051_top_1.oc8051_memory_interface1.imem_wait ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm2_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_t ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_v ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_vec_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.istb_t ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op2_buff ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op3_buff ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.op_pos ;
  wire \oc8051_top_1.oc8051_memory_interface1.out_of_rst ;
  wire [3:0] \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_buf ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log_prev ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_addr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_ind ;
  wire \oc8051_top_1.oc8051_memory_interface1.reti ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ri_r ;
  wire [4:0] \oc8051_top_1.oc8051_memory_interface1.rn_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.sfr ;
  wire \oc8051_top_1.oc8051_memory_interface1.sfr_bit ;
  wire \oc8051_top_1.oc8051_ram_top1.bit_addr_r ;
  wire [2:0] \oc8051_top_1.oc8051_ram_top1.bit_select ;
  wire \oc8051_top_1.oc8051_ram_top1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.rd_data_m ;
  wire \oc8051_top_1.oc8051_ram_top1.rd_en_r ;
  wire \oc8051_top_1.oc8051_ram_top1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.wr_data_r ;
  wire \oc8051_top_1.oc8051_rom1.clk ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.cxrom_data_out ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.data_o ;
  wire \oc8051_top_1.oc8051_rom1.ea_int ;
  wire \oc8051_top_1.oc8051_rom1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.b_reg ;
  wire \oc8051_top_1.oc8051_sfr1.bit_out ;
  wire \oc8051_top_1.oc8051_sfr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.cy ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_lo ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.int_ack ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ip ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.p ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ack ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie1_buff ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.set ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_int ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.intr ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd ;
  wire [11:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp ;
  wire [10:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.p ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.pres_ow ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.prescaler ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.psw_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.rxd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.srcAc ;
  wire \oc8051_top_1.oc8051_sfr1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.t2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.tc2_int ;
  wire \oc8051_top_1.oc8051_sfr1.tclk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.tf0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.txd ;
  wire \oc8051_top_1.oc8051_sfr1.uart_int ;
  wire \oc8051_top_1.oc8051_sfr1.wait_data ;
  wire \oc8051_top_1.oc8051_sfr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.p0_i ;
  wire [7:0] \oc8051_top_1.p0_o ;
  wire [7:0] \oc8051_top_1.p1_i ;
  wire [7:0] \oc8051_top_1.p1_o ;
  wire [7:0] \oc8051_top_1.p2_i ;
  wire [7:0] \oc8051_top_1.p2_o ;
  wire [7:0] \oc8051_top_1.p3_i ;
  wire [7:0] \oc8051_top_1.p3_o ;
  wire [15:0] \oc8051_top_1.pc ;
  wire [15:0] \oc8051_top_1.pc_log ;
  wire [15:0] \oc8051_top_1.pc_log_prev ;
  wire [7:0] \oc8051_top_1.psw ;
  wire [1:0] \oc8051_top_1.psw_set ;
  wire \oc8051_top_1.rd_ind ;
  wire \oc8051_top_1.reti ;
  wire \oc8051_top_1.rxd_i ;
  wire \oc8051_top_1.sfr_bit ;
  wire [7:0] \oc8051_top_1.sfr_out ;
  wire \oc8051_top_1.srcAc ;
  wire [2:0] \oc8051_top_1.src_sel1 ;
  wire [1:0] \oc8051_top_1.src_sel2 ;
  wire \oc8051_top_1.src_sel3 ;
  wire \oc8051_top_1.t0_i ;
  wire \oc8051_top_1.t1_i ;
  wire \oc8051_top_1.t2_i ;
  wire \oc8051_top_1.t2ex_i ;
  wire \oc8051_top_1.txd_o ;
  wire \oc8051_top_1.wait_data ;
  wire \oc8051_top_1.wb_clk_i ;
  wire \oc8051_top_1.wb_rst_i ;
  wire [15:0] \oc8051_top_1.wbd_adr_o ;
  wire \oc8051_top_1.wbd_cyc_o ;
  wire [7:0] \oc8051_top_1.wbd_dat_o ;
  wire \oc8051_top_1.wbd_stb_o ;
  wire \oc8051_top_1.wbd_we_o ;
  wire op0_cnst;
  input [7:0] p0_in;
  wire [7:0] p0_out;
  input [7:0] p1_in;
  wire [7:0] p1_out;
  input [7:0] p2_in;
  wire [7:0] p2_out;
  input [7:0] p3_in;
  wire [7:0] p3_out;
  wire [15:0] pc1;
  wire [15:0] pc2;
  output property_invalid_pc;
  wire [7:0] psw;
  wire [3:0] rd_iram_addr;
  wire [15:0] rd_rom_0_addr;
  input rst;
  input rxd_i;
  input t0_i;
  input t1_i;
  input t2_i;
  input t2ex_i;
  wire txd_o;
  wire [15:0] wbd_adr_o;
  wire wbd_cyc_o;
  wire [7:0] wbd_dat_o;
  wire wbd_stb_o;
  wire wbd_we_o;
  input [127:0] word_in;
  not (_42618_, rst);
  not (_18751_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  not (_18772_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_18773_, \oc8051_top_1.oc8051_decoder1.alu_op [1], _18772_);
  and (_18784_, _18773_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_18795_, \oc8051_top_1.oc8051_decoder1.alu_op [2], _18772_);
  and (_18806_, \oc8051_top_1.oc8051_decoder1.alu_op [3], _18772_);
  nor (_18817_, _18806_, _18795_);
  and (_18828_, _18817_, _18784_);
  nor (_18839_, _18828_, _18751_);
  and (_18850_, _18751_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  not (_18861_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  and (_18872_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _18861_);
  nor (_18883_, _18872_, _18850_);
  not (_18894_, _18883_);
  and (_18905_, _18894_, _18828_);
  or (_18916_, _18905_, _18839_);
  and (_22124_, _18916_, _42618_);
  nor (_18937_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  not (_18948_, _18937_);
  and (_18959_, _18948_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12]);
  and (_18970_, _18948_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8]);
  and (_18981_, _18948_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7]);
  not (_18992_, _18981_);
  not (_19003_, _18872_);
  nor (_19014_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  not (_19025_, \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  and (_19036_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _19025_);
  nor (_19047_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  not (_19058_, \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  nor (_19069_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _19058_);
  nor (_19080_, _19069_, _19047_);
  nor (_19091_, _19080_, _19036_);
  not (_19102_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  and (_19112_, _19036_, _19102_);
  nor (_19123_, _19112_, _19091_);
  and (_19134_, _19123_, _19014_);
  not (_19145_, _19134_);
  and (_19156_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and (_19167_, _19156_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  not (_19178_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and (_19189_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], _19178_);
  and (_19200_, _19189_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor (_19211_, _19200_, _19167_);
  and (_19222_, _19211_, _19145_);
  nor (_19233_, _19222_, _19003_);
  not (_19244_, _18850_);
  nor (_19255_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  nor (_19266_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _19058_);
  nor (_19277_, _19266_, _19255_);
  nor (_19288_, _19277_, _19036_);
  not (_19299_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  and (_19310_, _19036_, _19299_);
  nor (_19321_, _19310_, _19288_);
  and (_19332_, _19321_, _19014_);
  not (_19343_, _19332_);
  and (_19354_, _19156_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  and (_19365_, _19189_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_19376_, _19365_, _19354_);
  and (_19387_, _19376_, _19343_);
  nor (_19398_, _19387_, _19244_);
  nor (_19409_, _19398_, _19233_);
  nor (_19420_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  nor (_19430_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _19058_);
  nor (_19441_, _19430_, _19420_);
  nor (_19452_, _19441_, _19036_);
  not (_19463_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  and (_19474_, _19036_, _19463_);
  nor (_19485_, _19474_, _19452_);
  and (_19496_, _19485_, _19014_);
  not (_19507_, _19496_);
  and (_19517_, _19156_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  and (_19528_, _19189_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_19539_, _19528_, _19517_);
  and (_19550_, _19539_, _19507_);
  nor (_19561_, _19550_, _18894_);
  nor (_19572_, _19561_, _18937_);
  and (_19583_, _19572_, _19409_);
  nor (_19594_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  nor (_19604_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _19058_);
  nor (_19615_, _19604_, _19594_);
  nor (_19626_, _19615_, _19036_);
  not (_19637_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  and (_19648_, _19036_, _19637_);
  nor (_19659_, _19648_, _19626_);
  and (_19670_, _19659_, _19014_);
  not (_19681_, _19670_);
  and (_19691_, _19156_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  and (_19702_, _19189_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor (_19713_, _19702_, _19691_);
  and (_19724_, _19713_, _19681_);
  and (_19735_, _19724_, _18937_);
  nor (_19746_, _19735_, _19583_);
  not (_19768_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  and (_19779_, _19768_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and (_19791_, _19779_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_19803_, _19791_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_19815_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and (_19827_, _19815_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_19839_, _19827_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor (_19840_, _19839_, _19803_);
  not (_19851_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_19862_, _19779_, _19851_);
  and (_19872_, _19862_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  nor (_19883_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_19894_, _19883_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  and (_19905_, _19894_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  nor (_19916_, _19905_, _19872_);
  and (_19927_, _19916_, _19840_);
  and (_19938_, _19883_, _19768_);
  and (_19948_, _19938_, _19659_);
  and (_19959_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and (_19970_, _19959_, _19851_);
  and (_19981_, _19970_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_19992_, _19959_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_20003_, _19992_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [6]);
  nor (_20014_, _20003_, _19981_);
  not (_20025_, _20014_);
  nor (_20035_, _20025_, _19948_);
  and (_20046_, _20035_, _19927_);
  not (_20057_, _20046_);
  and (_20068_, _20057_, _19746_);
  not (_20079_, _20068_);
  nor (_20090_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  nor (_20101_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _19058_);
  nor (_20112_, _20101_, _20090_);
  nor (_20122_, _20112_, _19036_);
  not (_20133_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  and (_20144_, _19036_, _20133_);
  nor (_20155_, _20144_, _20122_);
  and (_20166_, _20155_, _19014_);
  not (_20177_, _20166_);
  and (_20188_, _19156_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  and (_20199_, _19189_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor (_20209_, _20199_, _20188_);
  and (_20220_, _20209_, _20177_);
  nor (_20231_, _20220_, _19003_);
  nor (_20242_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  nor (_20253_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _19058_);
  nor (_20264_, _20253_, _20242_);
  nor (_20275_, _20264_, _19036_);
  not (_20285_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  and (_20296_, _19036_, _20285_);
  nor (_20307_, _20296_, _20275_);
  and (_20318_, _20307_, _19014_);
  not (_20329_, _20318_);
  and (_20340_, _19156_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  and (_20351_, _19189_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor (_20362_, _20351_, _20340_);
  and (_20372_, _20362_, _20329_);
  nor (_20383_, _20372_, _19244_);
  nor (_20394_, _20383_, _20231_);
  nor (_20405_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  nor (_20416_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _19058_);
  nor (_20427_, _20416_, _20405_);
  nor (_20438_, _20427_, _19036_);
  not (_20449_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  and (_20459_, _19036_, _20449_);
  nor (_20470_, _20459_, _20438_);
  and (_20481_, _20470_, _19014_);
  not (_20492_, _20481_);
  and (_20503_, _19156_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  and (_20514_, _19189_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor (_20525_, _20514_, _20503_);
  and (_20536_, _20525_, _20492_);
  nor (_20546_, _20536_, _18894_);
  nor (_20557_, _20546_, _18937_);
  and (_20568_, _20557_, _20394_);
  nor (_20579_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  nor (_20590_, _19058_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [7]);
  nor (_20601_, _20590_, _20579_);
  nor (_20612_, _20601_, _19036_);
  not (_20623_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  and (_20633_, _19036_, _20623_);
  nor (_20644_, _20633_, _20612_);
  and (_20655_, _20644_, _19014_);
  not (_20676_, _20655_);
  and (_20687_, _19156_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  and (_20688_, _19189_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor (_20699_, _20688_, _20687_);
  and (_20719_, _20699_, _20676_);
  and (_20730_, _20719_, _18937_);
  nor (_20731_, _20730_, _20568_);
  and (_20752_, _19791_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_20763_, _19827_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor (_20764_, _20763_, _20752_);
  and (_20775_, _19894_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  and (_20786_, _19862_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  nor (_20797_, _20786_, _20775_);
  and (_20817_, _20797_, _20764_);
  and (_20818_, _20644_, _19938_);
  and (_20829_, _19970_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_20840_, _19992_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [7]);
  nor (_20851_, _20840_, _20829_);
  not (_20862_, _20851_);
  nor (_20873_, _20862_, _20818_);
  and (_20884_, _20873_, _20817_);
  not (_20895_, _20884_);
  and (_20905_, _20895_, _20731_);
  and (_20916_, _20905_, _20079_);
  not (_20927_, _20916_);
  and (_20948_, _19791_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_20949_, _19827_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_20960_, _20949_, _20948_);
  and (_20971_, _19894_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  and (_20982_, _19862_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  nor (_20993_, _20982_, _20971_);
  and (_21003_, _20993_, _20960_);
  and (_21014_, _20307_, _19938_);
  and (_21025_, _19992_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [5]);
  and (_21036_, _19970_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor (_21047_, _21036_, _21025_);
  not (_21058_, _21047_);
  nor (_21069_, _21058_, _21014_);
  and (_21080_, _21069_, _21003_);
  not (_21090_, _21080_);
  and (_21101_, _21090_, _20731_);
  and (_21122_, _19791_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_21123_, _19827_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_21134_, _21123_, _21122_);
  and (_21145_, _19894_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  and (_21156_, _19862_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  nor (_21167_, _21156_, _21145_);
  and (_21178_, _21167_, _21134_);
  and (_21188_, _19938_, _19321_);
  and (_21199_, _19970_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_21210_, _19992_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [4]);
  nor (_21221_, _21210_, _21199_);
  not (_21232_, _21221_);
  nor (_21243_, _21232_, _21188_);
  and (_21254_, _21243_, _21178_);
  not (_21265_, _21254_);
  and (_21276_, _21265_, _19746_);
  and (_21286_, _21101_, _21276_);
  nor (_21297_, _21286_, _20068_);
  and (_21318_, _21286_, _20057_);
  nor (_21319_, _21318_, _21297_);
  and (_21330_, _21319_, _21101_);
  and (_21341_, _20905_, _20068_);
  and (_21352_, _20731_, _20057_);
  and (_21363_, _20895_, _19746_);
  nor (_21373_, _21363_, _21352_);
  nor (_21384_, _21373_, _21341_);
  and (_21395_, _21384_, _21330_);
  and (_21406_, _21384_, _21318_);
  nor (_21417_, _21406_, _21395_);
  nor (_21428_, _21417_, _20927_);
  and (_21439_, _21417_, _20927_);
  nor (_21450_, _21439_, _21428_);
  not (_21461_, _21450_);
  and (_21471_, _21265_, _20731_);
  and (_21482_, _19791_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_21493_, _19827_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_21504_, _21493_, _21482_);
  and (_21515_, _19894_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  and (_21526_, _19862_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  nor (_21537_, _21526_, _21515_);
  and (_21548_, _21537_, _21504_);
  and (_21558_, _20155_, _19938_);
  and (_21569_, _19970_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_21580_, _19992_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [3]);
  nor (_21591_, _21580_, _21569_);
  not (_21602_, _21591_);
  nor (_21613_, _21602_, _21558_);
  and (_21624_, _21613_, _21548_);
  not (_21635_, _21624_);
  and (_21646_, _21635_, _19746_);
  and (_21666_, _21646_, _21471_);
  and (_21667_, _21090_, _19746_);
  nor (_21678_, _21667_, _21471_);
  nor (_21689_, _21678_, _21286_);
  and (_21700_, _21689_, _21666_);
  nor (_21711_, _21101_, _20068_);
  nor (_21722_, _21711_, _21330_);
  and (_21733_, _21722_, _21700_);
  nor (_21744_, _21384_, _21330_);
  nor (_21754_, _21744_, _21395_);
  nor (_21775_, _21754_, _21318_);
  nor (_21776_, _21775_, _21406_);
  and (_21787_, _21776_, _21733_);
  nor (_21798_, _21776_, _21733_);
  nor (_21809_, _21798_, _21787_);
  not (_21820_, _21809_);
  and (_21831_, _19791_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_21841_, _19827_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor (_21852_, _21841_, _21831_);
  and (_21863_, _19894_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  and (_21874_, _19862_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  nor (_21885_, _21874_, _21863_);
  and (_21896_, _21885_, _21852_);
  and (_21907_, _20470_, _19938_);
  and (_21918_, _19992_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [1]);
  and (_21929_, _19970_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor (_21939_, _21929_, _21918_);
  not (_21950_, _21939_);
  nor (_21961_, _21950_, _21907_);
  and (_21972_, _21961_, _21896_);
  not (_21983_, _21972_);
  and (_21994_, _21983_, _20731_);
  and (_22005_, _19791_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_22015_, _19827_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  nor (_22026_, _22015_, _22005_);
  and (_22037_, _19894_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  and (_22048_, _19862_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  nor (_22059_, _22048_, _22037_);
  and (_22070_, _22059_, _22026_);
  and (_22081_, _19938_, _19123_);
  and (_22092_, _19970_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_22102_, _19992_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [2]);
  nor (_22113_, _22102_, _22092_);
  not (_22125_, _22113_);
  nor (_22136_, _22125_, _22081_);
  and (_22147_, _22136_, _22070_);
  not (_22158_, _22147_);
  and (_22169_, _22158_, _19746_);
  and (_22180_, _22169_, _21994_);
  and (_22190_, _21983_, _19746_);
  not (_22201_, _22190_);
  and (_22222_, _22158_, _20731_);
  and (_22223_, _22222_, _22201_);
  and (_22234_, _22223_, _21646_);
  nor (_22245_, _22234_, _22180_);
  and (_22256_, _21635_, _20731_);
  nor (_22267_, _22256_, _21276_);
  nor (_22277_, _22267_, _21666_);
  not (_22288_, _22277_);
  nor (_22299_, _22288_, _22245_);
  nor (_22310_, _21689_, _21666_);
  nor (_22321_, _22310_, _21700_);
  and (_22332_, _22321_, _22299_);
  nor (_22343_, _21722_, _21700_);
  nor (_22354_, _22343_, _21733_);
  and (_22364_, _22354_, _22332_);
  and (_22375_, _19791_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_22386_, _19827_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor (_22397_, _22386_, _22375_);
  and (_22408_, _19894_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  and (_22419_, _19862_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  nor (_22430_, _22419_, _22408_);
  and (_22440_, _22430_, _22397_);
  and (_22451_, _19938_, _19485_);
  and (_22462_, _19992_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [0]);
  and (_22473_, _19970_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_22484_, _22473_, _22462_);
  not (_22495_, _22484_);
  nor (_22516_, _22495_, _22451_);
  and (_22517_, _22516_, _22440_);
  not (_22527_, _22517_);
  and (_22538_, _22527_, _20731_);
  and (_22549_, _22538_, _22190_);
  nor (_22560_, _22169_, _21994_);
  nor (_22571_, _22560_, _22180_);
  and (_22582_, _22571_, _22549_);
  nor (_22593_, _22223_, _21646_);
  nor (_22603_, _22593_, _22234_);
  and (_22624_, _22603_, _22582_);
  and (_22625_, _22288_, _22245_);
  nor (_22636_, _22625_, _22299_);
  and (_22647_, _22636_, _22624_);
  nor (_22658_, _22321_, _22299_);
  nor (_22669_, _22658_, _22332_);
  and (_22680_, _22669_, _22647_);
  nor (_22690_, _22354_, _22332_);
  nor (_22701_, _22690_, _22364_);
  and (_22712_, _22701_, _22680_);
  nor (_22723_, _22712_, _22364_);
  nor (_22734_, _22723_, _21820_);
  nor (_22745_, _22734_, _21787_);
  nor (_22756_, _22745_, _21461_);
  or (_22767_, _22756_, _21341_);
  nor (_22777_, _22767_, _21428_);
  nor (_22788_, _22777_, _18992_);
  and (_22799_, _22777_, _18992_);
  nor (_22810_, _22799_, _22788_);
  not (_22821_, _22810_);
  and (_22842_, _18948_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6]);
  and (_22843_, _22745_, _21461_);
  nor (_22854_, _22843_, _22756_);
  and (_22864_, _22854_, _22842_);
  and (_22875_, _18948_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5]);
  and (_22886_, _22723_, _21820_);
  nor (_22897_, _22886_, _22734_);
  and (_22908_, _22897_, _22875_);
  nor (_22919_, _22897_, _22875_);
  nor (_22930_, _22919_, _22908_);
  not (_22941_, _22930_);
  and (_22951_, _18948_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4]);
  nor (_22962_, _22701_, _22680_);
  nor (_22973_, _22962_, _22712_);
  and (_22984_, _22973_, _22951_);
  nor (_22995_, _22973_, _22951_);
  nor (_23006_, _22995_, _22984_);
  and (_23017_, _18948_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3]);
  nor (_23028_, _22669_, _22647_);
  nor (_23038_, _23028_, _22680_);
  and (_23049_, _23038_, _23017_);
  nor (_23060_, _23038_, _23017_);
  nor (_23071_, _23060_, _23049_);
  not (_23082_, _23071_);
  and (_23103_, _18948_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2]);
  nor (_23104_, _22636_, _22624_);
  nor (_23114_, _23104_, _22647_);
  and (_23125_, _23114_, _23103_);
  and (_23136_, _18948_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1]);
  nor (_23147_, _22603_, _22582_);
  nor (_23158_, _23147_, _22624_);
  and (_23169_, _23158_, _23136_);
  and (_23180_, _18948_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0]);
  nor (_23191_, _22571_, _22549_);
  nor (_23202_, _23191_, _22582_);
  and (_23213_, _23202_, _23180_);
  nor (_23223_, _23158_, _23136_);
  nor (_23234_, _23223_, _23169_);
  and (_23245_, _23234_, _23213_);
  nor (_23256_, _23245_, _23169_);
  not (_23267_, _23256_);
  nor (_23278_, _23114_, _23103_);
  nor (_23289_, _23278_, _23125_);
  and (_23300_, _23289_, _23267_);
  nor (_23311_, _23300_, _23125_);
  nor (_23322_, _23311_, _23082_);
  nor (_23332_, _23322_, _23049_);
  not (_23343_, _23332_);
  and (_23354_, _23343_, _23006_);
  nor (_23365_, _23354_, _22984_);
  nor (_23386_, _23365_, _22941_);
  nor (_23387_, _23386_, _22908_);
  nor (_23398_, _22854_, _22842_);
  nor (_23409_, _23398_, _22864_);
  not (_23420_, _23409_);
  nor (_23431_, _23420_, _23387_);
  nor (_23442_, _23431_, _22864_);
  nor (_23452_, _23442_, _22821_);
  nor (_23463_, _23452_, _22788_);
  not (_23474_, _23463_);
  and (_23485_, _23474_, _18970_);
  and (_23496_, _23485_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  and (_23507_, _18948_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10]);
  and (_23518_, _23507_, _23496_);
  and (_23529_, _23518_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  and (_23540_, _23529_, _18959_);
  not (_23551_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  nor (_23561_, _18937_, _23551_);
  or (_23572_, _23561_, _23540_);
  nand (_23583_, _23540_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  and (_23594_, _23583_, _23572_);
  and (_24283_, _23594_, _42618_);
  nor (_23615_, _18828_, _18861_);
  and (_23626_, _18828_, _18861_);
  or (_23637_, _23626_, _23615_);
  and (_02354_, _23637_, _42618_);
  and (_23658_, _22527_, _19746_);
  and (_02542_, _23658_, _42618_);
  nor (_23678_, _22538_, _22190_);
  nor (_23689_, _23678_, _22549_);
  and (_02700_, _23689_, _42618_);
  nor (_23710_, _23202_, _23180_);
  nor (_23721_, _23710_, _23213_);
  and (_02882_, _23721_, _42618_);
  nor (_23742_, _23234_, _23213_);
  nor (_23753_, _23742_, _23245_);
  and (_03125_, _23753_, _42618_);
  nor (_23773_, _23289_, _23267_);
  nor (_23784_, _23773_, _23300_);
  and (_03328_, _23784_, _42618_);
  and (_23815_, _23311_, _23082_);
  nor (_23816_, _23815_, _23322_);
  and (_03527_, _23816_, _42618_);
  nor (_23837_, _23343_, _23006_);
  nor (_23848_, _23837_, _23354_);
  and (_03728_, _23848_, _42618_);
  and (_23869_, _23365_, _22941_);
  nor (_23879_, _23869_, _23386_);
  and (_03927_, _23879_, _42618_);
  and (_23900_, _23420_, _23387_);
  nor (_23911_, _23900_, _23431_);
  and (_04023_, _23911_, _42618_);
  and (_23932_, _23442_, _22821_);
  nor (_23943_, _23932_, _23452_);
  and (_04123_, _23943_, _42618_);
  nor (_23963_, _23474_, _18970_);
  nor (_23974_, _23963_, _23485_);
  and (_04222_, _23974_, _42618_);
  and (_23995_, _18948_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  nor (_24006_, _23995_, _23485_);
  nor (_24017_, _24006_, _23496_);
  and (_04321_, _24017_, _42618_);
  nor (_24038_, _23507_, _23496_);
  nor (_24048_, _24038_, _23518_);
  and (_04414_, _24048_, _42618_);
  and (_24069_, _18948_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  nor (_24080_, _24069_, _23518_);
  nor (_24091_, _24080_, _23529_);
  and (_04512_, _24091_, _42618_);
  nor (_24112_, _23529_, _18959_);
  nor (_24122_, _24112_, _23540_);
  and (_04611_, _24122_, _42618_);
  and (_24143_, \oc8051_top_1.oc8051_decoder1.alu_op [0], _18772_);
  nor (_24154_, _24143_, _18773_);
  not (_24165_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and (_24176_, _18795_, _24165_);
  and (_24187_, _24176_, _24154_);
  and (_24198_, _24187_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand (_24208_, _24198_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_24219_, _24198_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_24230_, _24219_, _24208_);
  and (_00925_, _24230_, _42618_);
  and (_00951_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _42618_);
  not (_24261_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  and (_24272_, _20536_, _24261_);
  and (_24284_, _20220_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_24294_, _24284_, _24272_);
  nor (_24305_, _24294_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_24316_, _20372_, _24261_);
  and (_24327_, _20719_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_24338_, _24327_, _24316_);
  and (_24349_, _24338_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_24360_, _24349_, _24305_);
  nor (_24371_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nor (_24381_, _24371_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7]);
  and (_24392_, _24371_, _20884_);
  nor (_24403_, _24392_, _24381_);
  not (_24414_, _24403_);
  and (_24425_, _19550_, _24261_);
  and (_24436_, _19222_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_24447_, _24436_, _24425_);
  nor (_24458_, _24447_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_24468_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_24479_, _19387_, _24261_);
  and (_24490_, _19724_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_24501_, _24490_, _24479_);
  nor (_24522_, _24501_, _24468_);
  nor (_24523_, _24522_, _24458_);
  nor (_24534_, _24523_, _24414_);
  and (_24544_, _24523_, _24414_);
  nor (_24555_, _24544_, _24534_);
  nor (_24566_, _24371_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6]);
  and (_24577_, _24371_, _20046_);
  nor (_24588_, _24577_, _24566_);
  not (_24599_, _24588_);
  nor (_24610_, _20536_, _24261_);
  nor (_24621_, _24610_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_24631_, _20220_, _24261_);
  and (_24642_, _20372_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_24653_, _24642_, _24631_);
  nor (_24664_, _24653_, _24468_);
  nor (_24675_, _24664_, _24621_);
  nor (_24686_, _24675_, _24599_);
  and (_24697_, _24675_, _24599_);
  nor (_24707_, _24697_, _24686_);
  not (_24718_, _24707_);
  nor (_24729_, _24371_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5]);
  and (_24740_, _24371_, _21080_);
  nor (_24751_, _24740_, _24729_);
  not (_24762_, _24751_);
  nor (_24773_, _19550_, _24261_);
  nor (_24784_, _24773_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_24794_, _19222_, _24261_);
  and (_24805_, _19387_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_24816_, _24805_, _24794_);
  nor (_24827_, _24816_, _24468_);
  nor (_24838_, _24827_, _24784_);
  nor (_24849_, _24838_, _24762_);
  and (_24860_, _24838_, _24762_);
  and (_24871_, _24294_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_24881_, _24871_);
  nor (_24892_, _24371_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4]);
  and (_24903_, _24371_, _21254_);
  nor (_24914_, _24903_, _24892_);
  and (_24925_, _24914_, _24881_);
  and (_24936_, _24447_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_24947_, _24936_);
  and (_24958_, _24371_, _21624_);
  nor (_24968_, _24371_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3]);
  nor (_24979_, _24968_, _24958_);
  and (_24990_, _24979_, _24947_);
  nor (_25001_, _24979_, _24947_);
  nor (_25012_, _25001_, _24990_);
  not (_25023_, _25012_);
  and (_25034_, _24610_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_25045_, _25034_);
  and (_25065_, _24371_, _22147_);
  nor (_25066_, _24371_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2]);
  nor (_25077_, _25066_, _25065_);
  and (_25088_, _25077_, _25045_);
  and (_25099_, _24773_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_25110_, _25099_);
  nor (_25121_, _24371_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1]);
  and (_25132_, _24371_, _21972_);
  nor (_25143_, _25132_, _25121_);
  nor (_25154_, _25143_, _25110_);
  not (_25165_, _25154_);
  nor (_25176_, _25077_, _25045_);
  nor (_25187_, _25176_, _25088_);
  and (_25198_, _25187_, _25165_);
  nor (_25209_, _25198_, _25088_);
  nor (_25220_, _25209_, _25023_);
  nor (_25231_, _25220_, _24990_);
  nor (_25242_, _24914_, _24881_);
  nor (_25253_, _25242_, _24925_);
  not (_25264_, _25253_);
  nor (_25275_, _25264_, _25231_);
  nor (_25286_, _25275_, _24925_);
  nor (_25297_, _25286_, _24860_);
  nor (_25308_, _25297_, _24849_);
  nor (_25328_, _25308_, _24718_);
  nor (_25329_, _25328_, _24686_);
  not (_25340_, _25329_);
  and (_25351_, _25340_, _24555_);
  or (_25362_, _25351_, _24534_);
  and (_25373_, _20719_, _19724_);
  or (_25384_, _25373_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  not (_25395_, _24501_);
  and (_25406_, _24338_, _25395_);
  nor (_25417_, _24816_, _24653_);
  and (_25428_, _25417_, _25406_);
  or (_25439_, _25428_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_25450_, _25439_, _25384_);
  and (_25461_, _25450_, _25362_);
  and (_25472_, _25461_, _24360_);
  nor (_25483_, _25340_, _24555_);
  or (_25494_, _25483_, _25351_);
  and (_25505_, _25494_, _25472_);
  nor (_25516_, _25472_, _24403_);
  nor (_25527_, _25516_, _25505_);
  not (_25538_, _25527_);
  and (_25549_, _25527_, _24360_);
  not (_25560_, _24523_);
  nor (_25571_, _25472_, _24599_);
  and (_25582_, _25308_, _24718_);
  nor (_25593_, _25582_, _25328_);
  and (_25604_, _25593_, _25472_);
  or (_25615_, _25604_, _25571_);
  and (_25636_, _25615_, _25560_);
  nor (_25637_, _25615_, _25560_);
  nor (_25648_, _25637_, _25636_);
  not (_25659_, _25648_);
  not (_25670_, _24675_);
  nor (_25681_, _25472_, _24762_);
  nor (_25692_, _24860_, _24849_);
  nor (_25702_, _25692_, _25286_);
  and (_25713_, _25692_, _25286_);
  or (_25724_, _25713_, _25702_);
  and (_25735_, _25724_, _25472_);
  or (_25746_, _25735_, _25681_);
  and (_25757_, _25746_, _25670_);
  nor (_25768_, _25746_, _25670_);
  not (_25779_, _24838_);
  and (_25790_, _25264_, _25231_);
  or (_25801_, _25790_, _25275_);
  and (_25812_, _25801_, _25472_);
  nor (_25823_, _25472_, _24914_);
  nor (_25834_, _25823_, _25812_);
  and (_25845_, _25834_, _25779_);
  and (_25856_, _25209_, _25023_);
  nor (_25867_, _25856_, _25220_);
  not (_25878_, _25867_);
  and (_25889_, _25878_, _25472_);
  nor (_25900_, _25472_, _24979_);
  nor (_25911_, _25900_, _25889_);
  and (_25922_, _25911_, _24881_);
  nor (_25933_, _25911_, _24881_);
  nor (_25944_, _25933_, _25922_);
  not (_25965_, _25944_);
  nor (_25966_, _25187_, _25165_);
  nor (_25977_, _25966_, _25198_);
  not (_25988_, _25977_);
  and (_25999_, _25988_, _25472_);
  nor (_26010_, _25472_, _25077_);
  nor (_26021_, _26010_, _25999_);
  and (_26032_, _26021_, _24947_);
  and (_26043_, _25472_, _25099_);
  nor (_26054_, _26043_, _25143_);
  and (_26064_, _26043_, _25143_);
  nor (_26075_, _26064_, _26054_);
  and (_26086_, _26075_, _25045_);
  nor (_26097_, _26075_, _25045_);
  nor (_26108_, _26097_, _26086_);
  and (_26119_, _24371_, _22517_);
  nor (_26130_, _24371_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0]);
  nor (_26141_, _26130_, _26119_);
  nor (_26152_, _26141_, _25110_);
  not (_26163_, _26152_);
  and (_26174_, _26163_, _26108_);
  nor (_26185_, _26174_, _26086_);
  nor (_26196_, _26021_, _24947_);
  nor (_26207_, _26196_, _26032_);
  not (_26218_, _26207_);
  nor (_26229_, _26218_, _26185_);
  nor (_26240_, _26229_, _26032_);
  nor (_26251_, _26240_, _25965_);
  nor (_26262_, _26251_, _25922_);
  nor (_26273_, _25834_, _25779_);
  nor (_26284_, _26273_, _25845_);
  not (_26295_, _26284_);
  nor (_26306_, _26295_, _26262_);
  nor (_26317_, _26306_, _25845_);
  nor (_26328_, _26317_, _25768_);
  nor (_26339_, _26328_, _25757_);
  nor (_26350_, _26339_, _25659_);
  or (_26361_, _26350_, _25636_);
  or (_26372_, _26361_, _25549_);
  and (_26383_, _26372_, _25450_);
  nor (_26394_, _26383_, _25538_);
  and (_26405_, _25549_, _25450_);
  and (_26415_, _26405_, _26361_);
  or (_26426_, _26415_, _26394_);
  and (_00971_, _26426_, _42618_);
  or (_26447_, _25527_, _24360_);
  and (_26458_, _26447_, _26383_);
  and (_02836_, _26458_, _42618_);
  and (_02848_, _25472_, _42618_);
  and (_02870_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _42618_);
  and (_02894_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _42618_);
  and (_02916_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _42618_);
  or (_26519_, _24187_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_26530_, _24198_, rst);
  and (_02927_, _26530_, _26519_);
  and (_26551_, _26458_, _25099_);
  or (_26562_, _26551_, _26141_);
  nand (_26573_, _26551_, _26141_);
  and (_26584_, _26573_, _26562_);
  and (_02940_, _26584_, _42618_);
  nor (_26605_, _26163_, _26108_);
  or (_26616_, _26605_, _26174_);
  nand (_26627_, _26616_, _26458_);
  or (_26638_, _26458_, _26075_);
  and (_26649_, _26638_, _26627_);
  and (_02954_, _26649_, _42618_);
  and (_26670_, _26218_, _26185_);
  or (_26681_, _26670_, _26229_);
  nand (_26692_, _26681_, _26458_);
  or (_26703_, _26458_, _26021_);
  and (_26714_, _26703_, _26692_);
  and (_02967_, _26714_, _42618_);
  and (_26735_, _26240_, _25965_);
  or (_26746_, _26735_, _26251_);
  nand (_26756_, _26746_, _26458_);
  or (_26767_, _26458_, _25911_);
  and (_26778_, _26767_, _26756_);
  and (_02981_, _26778_, _42618_);
  and (_26799_, _26295_, _26262_);
  or (_26810_, _26799_, _26306_);
  nand (_26821_, _26810_, _26458_);
  or (_26832_, _26458_, _25834_);
  and (_26843_, _26832_, _26821_);
  and (_02995_, _26843_, _42618_);
  or (_26864_, _25768_, _25757_);
  and (_26875_, _26864_, _26317_);
  nor (_26886_, _26864_, _26317_);
  or (_26897_, _26886_, _26875_);
  nand (_26908_, _26897_, _26458_);
  or (_26919_, _26458_, _25746_);
  and (_26930_, _26919_, _26908_);
  and (_03008_, _26930_, _42618_);
  and (_26951_, _26339_, _25659_);
  or (_26962_, _26951_, _26350_);
  nand (_26973_, _26962_, _26458_);
  or (_26984_, _26458_, _25615_);
  and (_26995_, _26984_, _26973_);
  and (_03022_, _26995_, _42618_);
  and (_27016_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and (_27027_, _27016_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  and (_27038_, _27027_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  and (_27049_, _27038_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  and (_27060_, _27049_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  not (_27071_, _27060_);
  not (_27082_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_27093_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _18772_);
  and (_27103_, _27093_, _27082_);
  and (_27114_, _27103_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  not (_27125_, _27114_);
  nor (_27136_, _27049_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor (_27147_, _27136_, _27125_);
  and (_27158_, _27147_, _27071_);
  not (_27169_, _27158_);
  and (_27180_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_27191_, _27180_, _27093_);
  not (_27202_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  and (_27213_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _18772_);
  and (_27224_, _27213_, _27202_);
  and (_27245_, _27224_, _27082_);
  and (_27246_, _27245_, \oc8051_top_1.oc8051_memory_interface1.imm_r [5]);
  nor (_27257_, _27246_, _27191_);
  not (_27268_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  and (_27279_, _27103_, _27268_);
  and (_27290_, _27279_, \oc8051_top_1.oc8051_memory_interface1.ri_r [5]);
  and (_27301_, _27224_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_27312_, _27301_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [5]);
  nor (_27323_, _27312_, _27290_);
  and (_27334_, _27323_, _27257_);
  and (_27345_, _27334_, _27169_);
  and (_27356_, _27301_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [4]);
  not (_27367_, _27356_);
  and (_27378_, _27279_, \oc8051_top_1.oc8051_memory_interface1.ri_r [4]);
  nor (_27389_, _27378_, _27191_);
  and (_27400_, _27389_, _27367_);
  nor (_27411_, _27038_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  not (_27422_, _27411_);
  nor (_27433_, _27125_, _27049_);
  and (_27444_, _27433_, _27422_);
  or (_27454_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_27465_, _27454_, _18772_);
  nor (_27476_, _27465_, _27213_);
  and (_27487_, _27476_, \oc8051_top_1.oc8051_memory_interface1.rn_r [4]);
  and (_27498_, _27245_, \oc8051_top_1.oc8051_memory_interface1.imm_r [4]);
  nor (_27509_, _27498_, _27487_);
  not (_27520_, _27509_);
  nor (_27531_, _27520_, _27444_);
  and (_27542_, _27531_, _27400_);
  nor (_27553_, _27542_, _27345_);
  nor (_27564_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  nor (_27575_, _27564_, _27016_);
  and (_27586_, _27575_, _27114_);
  and (_27597_, _27279_, \oc8051_top_1.oc8051_memory_interface1.ri_r [1]);
  nor (_27608_, _27597_, _27586_);
  and (_27619_, _27301_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [1]);
  and (_27630_, _27245_, \oc8051_top_1.oc8051_memory_interface1.imm_r [1]);
  and (_27641_, _27476_, \oc8051_top_1.oc8051_memory_interface1.rn_r [1]);
  or (_27652_, _27641_, _27630_);
  nor (_27663_, _27652_, _27619_);
  and (_27674_, _27663_, _27608_);
  and (_27685_, _27301_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [0]);
  and (_27696_, _27245_, \oc8051_top_1.oc8051_memory_interface1.imm_r [0]);
  nor (_27707_, _27696_, _27685_);
  and (_27718_, _27279_, \oc8051_top_1.oc8051_memory_interface1.ri_r [0]);
  not (_27729_, _27718_);
  not (_27740_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and (_27751_, _27114_, _27740_);
  and (_27762_, _27476_, \oc8051_top_1.oc8051_memory_interface1.rn_r [0]);
  nor (_27773_, _27762_, _27751_);
  and (_27784_, _27773_, _27729_);
  and (_27795_, _27784_, _27707_);
  and (_27806_, _27795_, _27674_);
  not (_27816_, _27038_);
  nor (_27827_, _27027_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor (_27838_, _27827_, _27125_);
  and (_27849_, _27838_, _27816_);
  not (_27860_, _27849_);
  and (_27881_, _27476_, \oc8051_top_1.oc8051_memory_interface1.rn_r [3]);
  and (_27882_, _27279_, \oc8051_top_1.oc8051_memory_interface1.ri_r [3]);
  nor (_27893_, _27882_, _27881_);
  and (_27904_, _27301_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [3]);
  and (_27915_, _27245_, \oc8051_top_1.oc8051_memory_interface1.imm_r [3]);
  nor (_27926_, _27915_, _27904_);
  and (_27937_, _27926_, _27893_);
  and (_27948_, _27937_, _27860_);
  nor (_27959_, _27016_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_27970_, _27959_, _27027_);
  and (_27981_, _27970_, _27114_);
  and (_27992_, _27279_, \oc8051_top_1.oc8051_memory_interface1.ri_r [2]);
  nor (_28003_, _27992_, _27981_);
  and (_28014_, _27301_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [2]);
  and (_28025_, _27245_, \oc8051_top_1.oc8051_memory_interface1.imm_r [2]);
  and (_28036_, _27476_, \oc8051_top_1.oc8051_memory_interface1.rn_r [2]);
  or (_28047_, _28036_, _28025_);
  nor (_28058_, _28047_, _28014_);
  and (_28069_, _28058_, _28003_);
  and (_28080_, _28069_, _27948_);
  and (_28091_, _28080_, _27806_);
  not (_28102_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  and (_28113_, _27060_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor (_28124_, _28113_, _28102_);
  and (_28135_, _28113_, _28102_);
  nor (_28145_, _28135_, _28124_);
  nor (_28156_, _28145_, _27125_);
  not (_28167_, _28156_);
  and (_28188_, _27279_, \oc8051_top_1.oc8051_memory_interface1.ri_r [7]);
  nor (_28189_, _28188_, _27191_);
  and (_28200_, _27301_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [7]);
  and (_28211_, _27245_, \oc8051_top_1.oc8051_memory_interface1.imm_r [7]);
  nor (_28222_, _28211_, _28200_);
  and (_28233_, _28222_, _28189_);
  and (_28244_, _28233_, _28167_);
  not (_28255_, _28113_);
  nor (_28266_, _27060_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor (_28277_, _28266_, _27125_);
  and (_28288_, _28277_, _28255_);
  not (_28299_, _28288_);
  and (_28310_, _27245_, \oc8051_top_1.oc8051_memory_interface1.imm_r [6]);
  nor (_28321_, _28310_, _27191_);
  and (_28332_, _27279_, \oc8051_top_1.oc8051_memory_interface1.ri_r [6]);
  and (_28343_, _27301_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [6]);
  nor (_28354_, _28343_, _28332_);
  and (_28365_, _28354_, _28321_);
  and (_28376_, _28365_, _28299_);
  nor (_28387_, _28376_, _28244_);
  and (_28398_, _28387_, _28091_);
  nand (_28409_, _28398_, _27553_);
  and (_28420_, _26426_, _24187_);
  not (_28431_, _28420_);
  and (_28442_, _23594_, _18828_);
  not (_28453_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  and (_28463_, _24143_, _28453_);
  and (_28474_, _28463_, _18817_);
  nor (_28485_, _20046_, _19724_);
  and (_28496_, _20046_, _19724_);
  nor (_28507_, _28496_, _28485_);
  not (_28518_, _28507_);
  nor (_28539_, _21080_, _20372_);
  nor (_28540_, _21254_, _19387_);
  and (_28551_, _21080_, _20372_);
  nor (_28562_, _28551_, _28539_);
  and (_28573_, _28562_, _28540_);
  nor (_28584_, _28573_, _28539_);
  nor (_28595_, _28584_, _28518_);
  and (_28606_, _21254_, _19387_);
  nor (_28617_, _28606_, _28540_);
  nor (_28628_, _21624_, _20220_);
  and (_28639_, _21624_, _20220_);
  nor (_28650_, _28639_, _28628_);
  nor (_28661_, _22147_, _19222_);
  and (_28672_, _22147_, _19222_);
  nor (_28683_, _28672_, _28661_);
  not (_28694_, _28683_);
  nor (_28705_, _21972_, _20536_);
  nor (_28716_, _22517_, _19550_);
  and (_28727_, _21972_, _20536_);
  nor (_28738_, _28727_, _28705_);
  and (_28749_, _28738_, _28716_);
  nor (_28760_, _28749_, _28705_);
  nor (_28770_, _28760_, _28694_);
  nor (_28781_, _28770_, _28661_);
  nor (_28792_, _28781_, _28650_);
  and (_28803_, _28781_, _28650_);
  nor (_28814_, _28803_, _28792_);
  not (_28825_, \oc8051_top_1.oc8051_sfr1.bit_out );
  and (_28836_, _19036_, _28825_);
  not (_28847_, \oc8051_top_1.oc8051_ram_top1.bit_select [0]);
  and (_28858_, _28847_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_28869_, _28858_, _19080_);
  nor (_28880_, _28869_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  not (_28891_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_28912_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], _28891_);
  and (_28913_, _28912_, _20427_);
  not (_28924_, _28913_);
  and (_28935_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_28946_, _28935_, _20112_);
  nor (_28957_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_28968_, _28957_, _19441_);
  nor (_28979_, _28968_, _28946_);
  and (_28990_, _28979_, _28924_);
  and (_29001_, _28990_, _28880_);
  not (_29012_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_29023_, _28858_, _19615_);
  nor (_29034_, _29023_, _29012_);
  and (_29045_, _28957_, _19277_);
  not (_29056_, _29045_);
  and (_29067_, _28935_, _20601_);
  and (_29077_, _28912_, _20264_);
  nor (_29088_, _29077_, _29067_);
  and (_29099_, _29088_, _29056_);
  and (_29110_, _29099_, _29034_);
  nor (_29121_, _29110_, _29001_);
  nor (_29132_, _29121_, _19036_);
  nor (_29143_, _29132_, _28836_);
  and (_29154_, \oc8051_top_1.oc8051_decoder1.cy_sel [0], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_29165_, _29154_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  not (_29176_, _29165_);
  and (_29187_, _29176_, _29143_);
  and (_29198_, _29176_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  nor (_29209_, _29198_, _29187_);
  and (_29220_, _22517_, _19550_);
  nor (_29231_, _29220_, _28716_);
  not (_29242_, _29231_);
  nor (_29253_, _29242_, _29209_);
  and (_29264_, _29253_, _28738_);
  and (_29275_, _28760_, _28694_);
  nor (_29286_, _29275_, _28770_);
  and (_29297_, _29286_, _29264_);
  not (_29308_, _29297_);
  nor (_29319_, _29308_, _28814_);
  nor (_29330_, _28781_, _28639_);
  or (_29341_, _29330_, _28628_);
  or (_29352_, _29341_, _29319_);
  and (_29363_, _29352_, _28617_);
  nor (_29373_, _28562_, _28540_);
  nor (_29384_, _29373_, _28573_);
  and (_29395_, _29384_, _29363_);
  and (_29406_, _28584_, _28518_);
  nor (_29417_, _29406_, _28595_);
  and (_29438_, _29417_, _29395_);
  or (_29439_, _29438_, _28595_);
  nor (_29450_, _29439_, _28485_);
  nor (_29461_, _20884_, _20719_);
  and (_29472_, _20884_, _20719_);
  nor (_29483_, _29472_, _29461_);
  not (_29494_, _29483_);
  nor (_29505_, _29494_, _29450_);
  and (_29516_, _29494_, _29450_);
  nor (_29527_, _29516_, _29505_);
  and (_29538_, _29527_, _28474_);
  not (_29549_, _29538_);
  not (_29560_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_29571_, _18773_, _29560_);
  and (_29582_, _29571_, _18817_);
  not (_29593_, _29582_);
  not (_29604_, _19724_);
  nor (_29615_, _20046_, _29604_);
  and (_29626_, _21090_, _20372_);
  not (_29637_, _19387_);
  and (_29648_, _21254_, _29637_);
  nor (_29659_, _29648_, _28562_);
  nor (_29670_, _29659_, _29626_);
  nor (_29680_, _29670_, _28507_);
  nor (_29691_, _29680_, _29615_);
  and (_29712_, _29670_, _28507_);
  nor (_29713_, _29712_, _29680_);
  not (_29724_, _29713_);
  and (_29735_, _29648_, _28562_);
  nor (_29746_, _29735_, _29659_);
  not (_29757_, _29746_);
  not (_29768_, _28617_);
  not (_29779_, _28650_);
  not (_29790_, _19550_);
  and (_29801_, _22517_, _29790_);
  nor (_29812_, _29801_, _28738_);
  not (_29823_, _20536_);
  nor (_29834_, _21972_, _29823_);
  nor (_29845_, _29834_, _29812_);
  nor (_29856_, _29845_, _28683_);
  not (_29867_, _19222_);
  nor (_29878_, _22147_, _29867_);
  nor (_29889_, _29878_, _29856_);
  nor (_29900_, _29889_, _29779_);
  and (_29911_, _29889_, _29779_);
  nor (_29922_, _29911_, _29900_);
  and (_29933_, _29845_, _28683_);
  nor (_29944_, _29933_, _29856_);
  not (_29955_, _29944_);
  and (_29966_, _29801_, _28738_);
  nor (_29976_, _29966_, _29812_);
  not (_29987_, _29976_);
  nor (_29998_, _29231_, _29209_);
  and (_30009_, _29998_, _29987_);
  and (_30020_, _30009_, _29955_);
  and (_30031_, _30020_, _29922_);
  not (_30042_, _20220_);
  or (_30053_, _21624_, _30042_);
  and (_30064_, _21624_, _30042_);
  or (_30075_, _29889_, _30064_);
  and (_30085_, _30075_, _30053_);
  or (_30096_, _30085_, _30031_);
  and (_30107_, _30096_, _29768_);
  and (_30118_, _30107_, _29757_);
  and (_30129_, _30118_, _29724_);
  nor (_30140_, _30129_, _29691_);
  nor (_30151_, _30140_, _29483_);
  and (_30162_, _30140_, _29483_);
  nor (_30173_, _30162_, _30151_);
  nor (_30184_, _30173_, _29593_);
  and (_30194_, _18806_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and (_30205_, _30194_, _29571_);
  nor (_30216_, _22517_, _21972_);
  and (_30227_, _30216_, _22158_);
  and (_30238_, _30227_, _21635_);
  and (_30249_, _30238_, _21265_);
  and (_30260_, _30249_, _21090_);
  and (_30271_, _30260_, _20057_);
  and (_30282_, _30271_, _29209_);
  not (_30293_, _29209_);
  and (_30303_, _21080_, _20046_);
  and (_30314_, _22517_, _21972_);
  and (_30335_, _30314_, _22147_);
  and (_30336_, _30335_, _21624_);
  and (_30347_, _30336_, _21254_);
  and (_30358_, _30347_, _30303_);
  and (_30369_, _30358_, _30293_);
  nor (_30380_, _30369_, _30282_);
  and (_30391_, _30380_, _20884_);
  nor (_30402_, _30380_, _20884_);
  nor (_30412_, _30402_, _30391_);
  and (_30423_, _30412_, _30205_);
  not (_30434_, _20719_);
  nor (_30445_, _29209_, _30434_);
  not (_30456_, _30445_);
  and (_30467_, _29209_, _20884_);
  and (_30478_, _30194_, _18784_);
  not (_30489_, _30478_);
  nor (_30500_, _30489_, _30467_);
  and (_30511_, _30500_, _30456_);
  nor (_30522_, _30511_, _30423_);
  and (_30532_, _28463_, _24176_);
  not (_30543_, _30532_);
  and (_30554_, _22147_, _21972_);
  nor (_30565_, _30554_, _21624_);
  and (_30576_, _30565_, _30532_);
  and (_30587_, _30576_, _21265_);
  nor (_30598_, _30587_, _21090_);
  and (_30609_, _30598_, _20046_);
  nor (_30620_, _30303_, _20884_);
  nor (_30631_, _30620_, _30576_);
  and (_30641_, _30631_, _29209_);
  nor (_30652_, _30641_, _30609_);
  and (_30663_, _30652_, _20884_);
  nor (_30674_, _30652_, _20884_);
  nor (_30685_, _30674_, _30663_);
  nor (_30696_, _30685_, _30543_);
  not (_30707_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and (_30718_, _18806_, _30707_);
  and (_30729_, _30718_, _28463_);
  not (_30740_, _30729_);
  nor (_30750_, _30740_, _29472_);
  and (_30761_, _30718_, _24154_);
  and (_30772_, _30761_, _29483_);
  nor (_30783_, _30772_, _30750_);
  and (_30794_, _30194_, _24154_);
  not (_30805_, _30794_);
  nor (_30816_, _30805_, _22517_);
  and (_30827_, _30718_, _18773_);
  not (_30838_, _30827_);
  nor (_30849_, _30838_, _20046_);
  nor (_30859_, _30849_, _30816_);
  and (_30870_, _30194_, _28463_);
  not (_30881_, _30870_);
  nor (_30892_, _30881_, _29209_);
  and (_30903_, _24176_, _18784_);
  and (_30914_, _30903_, _29461_);
  and (_30925_, _29571_, _24176_);
  and (_30936_, _30925_, _20884_);
  nor (_30947_, _30936_, _30914_);
  and (_30958_, _24154_, _18817_);
  not (_30968_, _30958_);
  nor (_30979_, _30968_, _20884_);
  not (_30990_, _30979_);
  nand (_31001_, _30990_, _30947_);
  nor (_31012_, _31001_, _30892_);
  and (_31023_, _31012_, _30859_);
  and (_31045_, _31023_, _30783_);
  not (_31046_, _31045_);
  nor (_31068_, _31046_, _30696_);
  and (_31069_, _31068_, _30522_);
  not (_31090_, _31069_);
  nor (_31091_, _31090_, _30184_);
  and (_31113_, _31091_, _29549_);
  not (_31114_, _31113_);
  nor (_31125_, _31114_, _28442_);
  and (_31136_, _31125_, _28431_);
  not (_31147_, _31136_);
  or (_31168_, _31147_, _28409_);
  not (_31169_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_31189_, \oc8051_top_1.oc8051_decoder1.wr , _18772_);
  not (_31190_, _31189_);
  nor (_31211_, _31190_, _27103_);
  and (_31212_, _31211_, _31169_);
  not (_31233_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  nand (_31234_, _28409_, _31233_);
  and (_31255_, _31234_, _31212_);
  and (_31256_, _31255_, _31168_);
  nor (_31277_, _31211_, _31233_);
  not (_31278_, _28474_);
  nor (_31299_, _29505_, _29461_);
  nor (_31300_, _31299_, _31278_);
  not (_31320_, _31300_);
  and (_31321_, _20884_, _30434_);
  nor (_31342_, _31321_, _30151_);
  nor (_31343_, _31342_, _29593_);
  and (_31364_, _29209_, _20046_);
  and (_31365_, _31364_, _30598_);
  nor (_31386_, _31365_, _30467_);
  nor (_31387_, _29209_, _20884_);
  not (_31408_, _31387_);
  nor (_31409_, _31408_, _30609_);
  nor (_31429_, _31409_, _30543_);
  and (_31430_, _31429_, _31386_);
  nor (_31451_, _30925_, _30293_);
  and (_31452_, _30805_, _29198_);
  nor (_31473_, _31452_, _29187_);
  not (_31474_, _31473_);
  nor (_31495_, _31474_, _31451_);
  nor (_31496_, _29198_, _29143_);
  not (_31517_, _30761_);
  nor (_31518_, _31517_, _29187_);
  nor (_31538_, _31518_, _30729_);
  nor (_31539_, _31538_, _31496_);
  and (_31560_, _29165_, _29143_);
  and (_31561_, _30718_, _29571_);
  and (_31582_, _30903_, _29143_);
  nor (_31583_, _31582_, _31561_);
  nor (_31604_, _31583_, _31560_);
  nor (_31605_, _30968_, _29209_);
  and (_31626_, _30718_, _18784_);
  not (_31627_, _31626_);
  nor (_31647_, _31627_, _20884_);
  nor (_31648_, _30881_, _22517_);
  or (_31669_, _31648_, _30576_);
  or (_31670_, _31669_, _31647_);
  or (_31691_, _31670_, _31605_);
  or (_31692_, _31691_, _31604_);
  or (_31713_, _31692_, _31539_);
  or (_31714_, _31713_, _31495_);
  nor (_31735_, _31714_, _31430_);
  not (_31736_, _31735_);
  nor (_31756_, _31736_, _31343_);
  and (_31757_, _31756_, _31320_);
  nor (_31768_, _28376_, _27345_);
  not (_31779_, _28244_);
  not (_31790_, _27948_);
  nor (_31801_, _31790_, _27542_);
  and (_31812_, _31801_, _31779_);
  and (_31823_, _31812_, _31768_);
  not (_31834_, _28069_);
  nor (_31845_, _27795_, _27674_);
  and (_31855_, _31845_, _31834_);
  and (_31866_, _31855_, _31823_);
  nand (_31877_, _31866_, _31757_);
  or (_31888_, _31866_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_31899_, _31211_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_31910_, _31899_, _31888_);
  and (_31921_, _31910_, _31877_);
  or (_31932_, _31921_, _31277_);
  or (_31943_, _31932_, _31256_);
  and (_06626_, _31943_, _42618_);
  and (_31963_, _26584_, _24187_);
  not (_31974_, _31963_);
  and (_31985_, _29242_, _29209_);
  nor (_31996_, _31985_, _29253_);
  nand (_32007_, _31996_, _28474_);
  and (_32018_, _30903_, _28716_);
  and (_32029_, _30925_, _22517_);
  nor (_32040_, _32029_, _32018_);
  nor (_32051_, _31517_, _28716_);
  nor (_32062_, _32051_, _30729_);
  or (_32073_, _32062_, _29220_);
  and (_32083_, _30194_, _28453_);
  not (_32094_, _32083_);
  nor (_32105_, _32094_, _21972_);
  and (_32116_, _31561_, _20895_);
  nor (_32127_, _32116_, _32105_);
  and (_32138_, _32127_, _32073_);
  and (_32149_, _32138_, _32040_);
  and (_32160_, _23911_, _18828_);
  and (_32171_, _31996_, _29582_);
  nor (_32182_, _31627_, _29209_);
  nor (_32192_, _30489_, _19550_);
  and (_32203_, _30205_, _22517_);
  nor (_32214_, _32203_, _32192_);
  nor (_32225_, _30958_, _30532_);
  nor (_32236_, _32225_, _22517_);
  not (_32247_, _32236_);
  nand (_32258_, _32247_, _32214_);
  or (_32269_, _32258_, _32182_);
  or (_32280_, _32269_, _32171_);
  nor (_32291_, _32280_, _32160_);
  and (_32301_, _32291_, _32149_);
  and (_32312_, _32301_, _32007_);
  and (_32323_, _32312_, _31974_);
  not (_32334_, _32323_);
  or (_32345_, _32334_, _28409_);
  not (_32356_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nand (_32367_, _28409_, _32356_);
  and (_32378_, _32367_, _31212_);
  and (_32389_, _32378_, _32345_);
  nor (_32399_, _31211_, _32356_);
  not (_32410_, _31757_);
  or (_32421_, _32410_, _28409_);
  and (_32432_, _32367_, _31899_);
  and (_32443_, _32432_, _32421_);
  or (_32454_, _32443_, _32399_);
  or (_32465_, _32454_, _32389_);
  and (_08867_, _32465_, _42618_);
  and (_32486_, _23943_, _18828_);
  not (_32497_, _32486_);
  and (_32508_, _26649_, _24187_);
  nor (_32518_, _28738_, _28716_);
  or (_32529_, _32518_, _28749_);
  and (_32540_, _32529_, _29253_);
  nor (_32551_, _32529_, _29253_);
  or (_32562_, _32551_, _32540_);
  and (_32573_, _32562_, _28474_);
  not (_32584_, _32573_);
  nor (_32595_, _30565_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_32606_, _32595_, _21983_);
  nor (_32617_, _32595_, _21983_);
  nor (_32627_, _32617_, _32606_);
  nor (_32638_, _32627_, _30543_);
  not (_32649_, _32638_);
  and (_32660_, _30761_, _28738_);
  nor (_32671_, _30740_, _28727_);
  not (_32682_, _32671_);
  and (_32693_, _30903_, _28705_);
  and (_32704_, _30925_, _21972_);
  nor (_32715_, _32704_, _32693_);
  nand (_32726_, _32715_, _32682_);
  nor (_32736_, _32726_, _32660_);
  nor (_32747_, _32094_, _22147_);
  not (_32758_, _32747_);
  nor (_32769_, _30968_, _21972_);
  nor (_32780_, _30838_, _22517_);
  nor (_32791_, _32780_, _32769_);
  and (_32802_, _32791_, _32758_);
  and (_32813_, _32802_, _32736_);
  and (_32824_, _32813_, _32649_);
  and (_32835_, _32824_, _32584_);
  nor (_32845_, _30489_, _20536_);
  nor (_32856_, _30314_, _30216_);
  not (_32867_, _32856_);
  nor (_32878_, _32867_, _29209_);
  and (_32889_, _32867_, _29209_);
  nor (_32900_, _32889_, _32878_);
  and (_32911_, _32900_, _30205_);
  nor (_32922_, _32911_, _32845_);
  not (_32933_, _32922_);
  nor (_32944_, _29998_, _29987_);
  nor (_32955_, _32944_, _30009_);
  nor (_32965_, _32955_, _29593_);
  nor (_32976_, _32965_, _32933_);
  and (_32987_, _32976_, _32835_);
  not (_32998_, _32987_);
  nor (_33009_, _32998_, _32508_);
  and (_33020_, _33009_, _32497_);
  not (_33031_, _33020_);
  or (_33042_, _33031_, _28409_);
  not (_33053_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  nand (_33064_, _28409_, _33053_);
  and (_33074_, _33064_, _31212_);
  and (_33085_, _33074_, _33042_);
  nor (_33096_, _31211_, _33053_);
  not (_33107_, _27674_);
  nor (_33118_, _27795_, _33107_);
  and (_33129_, _33118_, _28069_);
  and (_33140_, _33129_, _31823_);
  nand (_33151_, _33140_, _31757_);
  or (_33162_, _33140_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_33172_, _33162_, _31899_);
  and (_33183_, _33172_, _33151_);
  or (_33194_, _33183_, _33096_);
  or (_33205_, _33194_, _33085_);
  and (_08878_, _33205_, _42618_);
  and (_33226_, _26714_, _24187_);
  not (_33237_, _33226_);
  and (_33248_, _23974_, _18828_);
  nor (_33259_, _30489_, _19222_);
  and (_33270_, _30314_, _30293_);
  and (_33281_, _30216_, _29209_);
  nor (_33291_, _33281_, _33270_);
  nor (_33302_, _33291_, _22147_);
  not (_33313_, _30205_);
  and (_33324_, _33291_, _22147_);
  or (_33335_, _33324_, _33313_);
  nor (_33346_, _33335_, _33302_);
  nor (_33357_, _33346_, _33259_);
  nor (_33368_, _30009_, _29955_);
  nor (_33379_, _33368_, _30020_);
  nor (_33390_, _33379_, _29593_);
  and (_33400_, _30761_, _28683_);
  nor (_33411_, _30740_, _28672_);
  not (_33422_, _33411_);
  and (_33433_, _30903_, _28661_);
  and (_33444_, _30925_, _22147_);
  nor (_33455_, _33444_, _33433_);
  nand (_33466_, _33455_, _33422_);
  nor (_33477_, _33466_, _33400_);
  nor (_33488_, _30838_, _21972_);
  not (_33499_, _33488_);
  nor (_33509_, _30968_, _22147_);
  nor (_33520_, _32094_, _21624_);
  nor (_33531_, _33520_, _33509_);
  and (_33542_, _33531_, _33499_);
  and (_33553_, _33542_, _33477_);
  not (_33564_, _33553_);
  nor (_33575_, _33564_, _33390_);
  nor (_33586_, _29286_, _29264_);
  nor (_33597_, _33586_, _31278_);
  and (_33608_, _33597_, _29308_);
  nor (_33618_, _32617_, _22147_);
  and (_33629_, _30554_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_33640_, _33629_, _33618_);
  nor (_33651_, _33640_, _30543_);
  nor (_33662_, _33651_, _33608_);
  and (_33673_, _33662_, _33575_);
  and (_33684_, _33673_, _33357_);
  not (_33695_, _33684_);
  nor (_33706_, _33695_, _33248_);
  and (_33717_, _33706_, _33237_);
  not (_33728_, _33717_);
  or (_33738_, _33728_, _28409_);
  not (_33749_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  nand (_33760_, _28409_, _33749_);
  and (_33771_, _33760_, _31212_);
  and (_33782_, _33771_, _33738_);
  nor (_33793_, _31211_, _33749_);
  nand (_33804_, _31823_, _28069_);
  or (_33815_, _31845_, _33804_);
  and (_33826_, _33815_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_33837_, _28069_, _27795_);
  and (_33847_, _33837_, _33107_);
  not (_33858_, _33847_);
  nor (_33869_, _33858_, _31757_);
  and (_33880_, _28069_, _27674_);
  and (_33891_, _33880_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or (_33902_, _33891_, _33869_);
  and (_33913_, _33902_, _31823_);
  or (_33924_, _33913_, _33826_);
  and (_33935_, _33924_, _31899_);
  or (_33945_, _33935_, _33793_);
  or (_33956_, _33945_, _33782_);
  and (_08889_, _33956_, _42618_);
  and (_33977_, _24017_, _18828_);
  not (_33988_, _33977_);
  and (_33999_, _26778_, _24187_);
  and (_34010_, _29308_, _28814_);
  or (_34021_, _34010_, _31278_);
  nor (_34032_, _34021_, _29319_);
  not (_34043_, _34032_);
  nor (_34054_, _30020_, _29922_);
  nor (_34064_, _34054_, _30031_);
  nor (_34075_, _34064_, _29593_);
  not (_34086_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_34097_, _30554_, _34086_);
  nor (_34108_, _34097_, _21635_);
  or (_34119_, _34108_, _30543_);
  nor (_34130_, _34119_, _30565_);
  nor (_34141_, _34130_, _34075_);
  nor (_34152_, _30489_, _20220_);
  nor (_34163_, _30335_, _29209_);
  nor (_34173_, _30227_, _30293_);
  nor (_34186_, _34173_, _34163_);
  and (_34205_, _34186_, _21635_);
  not (_34216_, _34205_);
  nor (_34227_, _34186_, _21635_);
  nor (_34238_, _34227_, _33313_);
  and (_34249_, _34238_, _34216_);
  nor (_34260_, _34249_, _34152_);
  and (_34271_, _30903_, _28628_);
  and (_34282_, _30925_, _21624_);
  nor (_34292_, _34282_, _34271_);
  nor (_34303_, _32094_, _21254_);
  not (_34314_, _34303_);
  and (_34325_, _34314_, _34292_);
  nor (_34336_, _30740_, _28639_);
  and (_34347_, _30761_, _28650_);
  nor (_34358_, _34347_, _34336_);
  nor (_34369_, _30968_, _21624_);
  nor (_34380_, _30838_, _22147_);
  nor (_34391_, _34380_, _34369_);
  and (_34401_, _34391_, _34358_);
  and (_34412_, _34401_, _34325_);
  and (_34423_, _34412_, _34260_);
  and (_34434_, _34423_, _34141_);
  and (_34445_, _34434_, _34043_);
  not (_34456_, _34445_);
  nor (_34467_, _34456_, _33999_);
  and (_34478_, _34467_, _33988_);
  not (_34489_, _34478_);
  or (_34500_, _34489_, _28409_);
  not (_34510_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nand (_34521_, _28409_, _34510_);
  and (_34532_, _34521_, _31212_);
  and (_34543_, _34532_, _34500_);
  nor (_34554_, _31211_, _34510_);
  and (_34565_, _33804_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_34576_, _31845_, _28069_);
  not (_34587_, _34576_);
  nor (_34598_, _34587_, _31757_);
  nor (_34609_, _33880_, _33837_);
  nor (_34620_, _34609_, _34510_);
  or (_34630_, _34620_, _34598_);
  and (_34641_, _34630_, _31823_);
  or (_34652_, _34641_, _34565_);
  and (_34663_, _34652_, _31899_);
  or (_34674_, _34663_, _34554_);
  or (_34685_, _34674_, _34543_);
  and (_08900_, _34685_, _42618_);
  and (_34706_, _26843_, _24187_);
  not (_34717_, _34706_);
  and (_34727_, _24048_, _18828_);
  nor (_34738_, _30096_, _28617_);
  and (_34749_, _30096_, _28617_);
  nor (_34760_, _34749_, _34738_);
  and (_34771_, _34760_, _29582_);
  not (_34782_, _34771_);
  nor (_34793_, _29352_, _28617_);
  nor (_34804_, _34793_, _29363_);
  and (_34815_, _34804_, _28474_);
  and (_34826_, _29209_, _21265_);
  nor (_34837_, _29209_, _19387_);
  or (_34847_, _34837_, _34826_);
  and (_34858_, _34847_, _30478_);
  and (_34869_, _30238_, _29209_);
  and (_34880_, _30336_, _30293_);
  nor (_34891_, _34880_, _34869_);
  nor (_34902_, _34891_, _21254_);
  not (_34913_, _34902_);
  and (_34924_, _34891_, _21254_);
  nor (_34935_, _34924_, _33313_);
  and (_34946_, _34935_, _34913_);
  nor (_34956_, _34946_, _34858_);
  nor (_34967_, _30576_, _21265_);
  not (_34978_, _34967_);
  nor (_34989_, _30587_, _30543_);
  and (_35000_, _34989_, _34978_);
  not (_35011_, _35000_);
  and (_35022_, _30761_, _28617_);
  and (_35033_, _30903_, _28540_);
  nor (_35044_, _30740_, _28606_);
  and (_35055_, _30925_, _21254_);
  or (_35065_, _35055_, _35044_);
  or (_35076_, _35065_, _35033_);
  nor (_35087_, _35076_, _35022_);
  nor (_35098_, _30968_, _21254_);
  nor (_35109_, _32094_, _21080_);
  nor (_35120_, _30838_, _21624_);
  or (_35131_, _35120_, _35109_);
  nor (_35142_, _35131_, _35098_);
  and (_35153_, _35142_, _35087_);
  and (_35164_, _35153_, _35011_);
  and (_35174_, _35164_, _34956_);
  not (_35185_, _35174_);
  nor (_35196_, _35185_, _34815_);
  and (_35207_, _35196_, _34782_);
  not (_35218_, _35207_);
  nor (_35229_, _35218_, _34727_);
  and (_35240_, _35229_, _34717_);
  not (_35251_, _35240_);
  or (_35262_, _35251_, _28409_);
  not (_35273_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nand (_35283_, _28409_, _35273_);
  and (_35294_, _35283_, _31212_);
  and (_35305_, _35294_, _35262_);
  nor (_35316_, _31211_, _35273_);
  not (_35327_, _31823_);
  and (_35338_, _27806_, _31834_);
  nor (_35349_, _27806_, _31834_);
  nor (_35360_, _35349_, _35338_);
  or (_35371_, _35360_, _35327_);
  and (_35382_, _35371_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_35393_, _35338_, _32410_);
  and (_35403_, _35349_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  or (_35414_, _35403_, _35393_);
  and (_35425_, _35414_, _31823_);
  or (_35436_, _35425_, _35382_);
  and (_35447_, _35436_, _31899_);
  or (_35458_, _35447_, _35316_);
  or (_35469_, _35458_, _35305_);
  and (_08911_, _35469_, _42618_);
  and (_35489_, _26930_, _24187_);
  not (_35500_, _35489_);
  and (_35511_, _24091_, _18828_);
  nor (_35522_, _29384_, _29363_);
  nor (_35533_, _35522_, _29395_);
  and (_35544_, _35533_, _28474_);
  not (_35555_, _35544_);
  nor (_35566_, _30107_, _29757_);
  nor (_35577_, _35566_, _30118_);
  nor (_35588_, _35577_, _29593_);
  nor (_35598_, _29209_, _20372_);
  and (_35609_, _29209_, _21090_);
  nor (_35620_, _35609_, _35598_);
  nor (_35631_, _35620_, _30489_);
  nor (_35642_, _30249_, _30293_);
  nor (_35653_, _30347_, _29209_);
  nor (_35664_, _35653_, _35642_);
  and (_35675_, _35664_, _21090_);
  nor (_35686_, _35664_, _21090_);
  or (_35697_, _35686_, _33313_);
  nor (_35707_, _35697_, _35675_);
  nor (_35718_, _35707_, _35631_);
  not (_35729_, _30641_);
  and (_35740_, _35729_, _30598_);
  nor (_35751_, _30641_, _30587_);
  nor (_35762_, _35751_, _21080_);
  nor (_35773_, _35762_, _35740_);
  nor (_35784_, _35773_, _30543_);
  and (_35795_, _30761_, _28562_);
  nor (_35806_, _30740_, _28551_);
  not (_35817_, _35806_);
  and (_35827_, _30903_, _28539_);
  and (_35838_, _30925_, _21080_);
  nor (_35849_, _35838_, _35827_);
  nand (_35860_, _35849_, _35817_);
  nor (_35871_, _35860_, _35795_);
  nor (_35882_, _32094_, _20046_);
  not (_35893_, _35882_);
  nor (_35904_, _30968_, _21080_);
  nor (_35915_, _30838_, _21254_);
  nor (_35926_, _35915_, _35904_);
  and (_35937_, _35926_, _35893_);
  and (_35948_, _35937_, _35871_);
  not (_35958_, _35948_);
  nor (_35969_, _35958_, _35784_);
  and (_35980_, _35969_, _35718_);
  not (_35991_, _35980_);
  nor (_36002_, _35991_, _35588_);
  and (_36013_, _36002_, _35555_);
  not (_36024_, _36013_);
  nor (_36035_, _36024_, _35511_);
  and (_36046_, _36035_, _35500_);
  not (_36057_, _36046_);
  or (_36068_, _36057_, _28409_);
  not (_36078_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nand (_36089_, _28409_, _36078_);
  and (_36100_, _36089_, _31212_);
  and (_36111_, _36100_, _36068_);
  nor (_36122_, _31211_, _36078_);
  and (_36133_, _33118_, _31834_);
  and (_36144_, _36133_, _31823_);
  nand (_36155_, _36144_, _31757_);
  or (_36166_, _36144_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_36177_, _36166_, _31899_);
  and (_36188_, _36177_, _36155_);
  or (_36199_, _36188_, _36122_);
  or (_36209_, _36199_, _36111_);
  and (_08922_, _36209_, _42618_);
  and (_36230_, _26995_, _24187_);
  and (_36241_, _24122_, _18828_);
  or (_36252_, _29417_, _29395_);
  nor (_36263_, _31278_, _29438_);
  and (_36274_, _36263_, _36252_);
  nor (_36284_, _30118_, _29724_);
  nor (_36295_, _36284_, _30129_);
  nor (_36306_, _36295_, _29593_);
  nor (_36317_, _29209_, _29604_);
  or (_36328_, _36317_, _30489_);
  nor (_36339_, _36328_, _31364_);
  nor (_36350_, _29209_, _21090_);
  nand (_36361_, _36350_, _30347_);
  nand (_36371_, _30260_, _29209_);
  and (_36382_, _36371_, _36361_);
  and (_36393_, _36382_, _20046_);
  nor (_36404_, _36382_, _20046_);
  or (_36415_, _36404_, _33313_);
  nor (_36426_, _36415_, _36393_);
  nor (_36437_, _36426_, _36339_);
  nor (_36448_, _35740_, _20046_);
  and (_36458_, _35740_, _20046_);
  or (_36469_, _36458_, _36448_);
  and (_36480_, _36469_, _30532_);
  and (_36491_, _30761_, _28507_);
  nor (_36502_, _30740_, _28496_);
  not (_36513_, _36502_);
  and (_36524_, _30903_, _28485_);
  and (_36535_, _30925_, _20046_);
  nor (_36545_, _36535_, _36524_);
  nand (_36556_, _36545_, _36513_);
  nor (_36567_, _36556_, _36491_);
  nor (_36578_, _32094_, _20884_);
  nor (_36589_, _30968_, _20046_);
  nor (_36600_, _30838_, _21080_);
  or (_36611_, _36600_, _36589_);
  nor (_36621_, _36611_, _36578_);
  nand (_36632_, _36621_, _36567_);
  nor (_36643_, _36632_, _36480_);
  nand (_36654_, _36643_, _36437_);
  or (_36665_, _36654_, _36306_);
  or (_36676_, _36665_, _36274_);
  or (_36687_, _36676_, _36241_);
  or (_36698_, _36687_, _36230_);
  or (_36708_, _36698_, _28409_);
  not (_36719_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  nand (_36730_, _28409_, _36719_);
  and (_36741_, _36730_, _31212_);
  and (_36752_, _36741_, _36708_);
  nor (_36763_, _31211_, _36719_);
  nor (_36774_, _28069_, _27674_);
  and (_36785_, _36774_, _27795_);
  and (_36795_, _36785_, _31823_);
  nand (_36806_, _36795_, _31757_);
  or (_36817_, _36795_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_36828_, _36817_, _31899_);
  and (_36839_, _36828_, _36806_);
  or (_36850_, _36839_, _36763_);
  or (_36861_, _36850_, _36752_);
  and (_08933_, _36861_, _42618_);
  and (_36882_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_36893_, \oc8051_top_1.oc8051_decoder1.state [0], \oc8051_top_1.oc8051_decoder1.state [1]);
  or (_36903_, _36893_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_36914_, _36903_);
  not (_36925_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  nor (_36936_, \oc8051_top_1.oc8051_memory_interface1.imem_wait , \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and (_36947_, _36936_, _36925_);
  and (_36958_, _36893_, _18772_);
  and (_36969_, _36958_, _36947_);
  and (_36980_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_36991_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], \oc8051_top_1.oc8051_memory_interface1.cdone );
  not (_37002_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_37012_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  not (_37023_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_37034_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_37045_, _37034_, _37023_);
  and (_37056_, _37045_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  and (_37067_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_37078_, _37067_, _37023_);
  and (_37089_, _37078_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_37100_, _37089_, _37056_);
  not (_37111_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_37122_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], _37111_);
  and (_37133_, _37122_, _37023_);
  and (_37144_, _37133_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  not (_37155_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_37166_, _37155_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_37177_, _37166_, _37023_);
  and (_37188_, _37177_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor (_37199_, _37188_, _37144_);
  nor (_37210_, _37034_, _37023_);
  and (_37221_, _37210_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_37232_, _37034_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_37243_, _37232_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor (_37253_, _37243_, _37221_);
  and (_37264_, _37253_, _37199_);
  and (_37275_, _37264_, _37100_);
  nor (_37286_, _37275_, _37012_);
  and (_37297_, _37286_, _37002_);
  nor (_37308_, _37297_, _36991_);
  nor (_37319_, _37308_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_37330_, _37319_, _36980_);
  and (_37341_, _37330_, _36969_);
  not (_37352_, _37341_);
  not (_37363_, _36947_);
  nor (_37373_, _36958_, \oc8051_top_1.oc8051_decoder1.op [3]);
  nor (_37384_, _37373_, _37363_);
  and (_37395_, _37384_, _37352_);
  not (_37406_, _37395_);
  and (_37417_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_37428_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_37439_, _37078_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  and (_37450_, _37177_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor (_37461_, _37450_, _37439_);
  and (_37472_, _37210_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_37482_, _37232_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor (_37493_, _37482_, _37472_);
  and (_37504_, _37045_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  and (_37515_, _37133_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_37526_, _37515_, _37504_);
  and (_37537_, _37526_, _37493_);
  and (_37548_, _37537_, _37461_);
  nor (_37559_, _37548_, _37012_);
  and (_37570_, _37559_, _37002_);
  nor (_37581_, _37570_, _37428_);
  nor (_37591_, _37581_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_37602_, _37591_, _37417_);
  and (_37613_, _37602_, _36969_);
  not (_37624_, _37613_);
  nor (_37635_, _36958_, \oc8051_top_1.oc8051_decoder1.op [0]);
  nor (_37646_, _37635_, _37363_);
  and (_37657_, _37646_, _37624_);
  and (_37668_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  not (_37679_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_37690_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], \oc8051_top_1.oc8051_memory_interface1.cdone );
  or (_37701_, _37012_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_37712_, _37177_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  and (_37723_, _37133_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_37734_, _37723_, _37712_);
  and (_37745_, _37210_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_37756_, _37232_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor (_37765_, _37756_, _37745_);
  and (_37776_, _37045_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  and (_37787_, _37078_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_37798_, _37787_, _37776_);
  and (_37809_, _37798_, _37765_);
  and (_37820_, _37809_, _37734_);
  nor (_37829_, _37820_, _37701_);
  or (_37830_, _37829_, _37690_);
  and (_37831_, _37830_, _37679_);
  nor (_37832_, _37831_, _37668_);
  and (_37833_, _37832_, _36969_);
  not (_37834_, _37833_);
  nor (_37835_, _36958_, \oc8051_top_1.oc8051_decoder1.op [2]);
  nor (_37836_, _37835_, _37363_);
  and (_37837_, _37836_, _37834_);
  not (_37838_, _37837_);
  not (_37839_, _36969_);
  and (_37840_, _37078_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  and (_37841_, _37232_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nor (_37842_, _37841_, _37840_);
  and (_37843_, _37133_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_37844_, _37843_, _37012_);
  and (_37845_, _37844_, _37842_);
  and (_37846_, _37177_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  not (_37847_, _37846_);
  and (_37848_, _37045_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  and (_37849_, _37210_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor (_37850_, _37849_, _37848_);
  and (_37851_, _37850_, _37847_);
  and (_37852_, _37851_, _37845_);
  and (_37853_, _37852_, _37002_);
  nor (_37854_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], _37002_);
  or (_37855_, _37854_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_37856_, _37855_, _37853_);
  and (_37857_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  or (_37858_, _37857_, _37856_);
  nor (_37859_, _37858_, _37839_);
  not (_37860_, _37859_);
  nor (_37861_, _36958_, \oc8051_top_1.oc8051_decoder1.op [1]);
  nor (_37862_, _37861_, _37363_);
  and (_37863_, _37862_, _37860_);
  and (_37864_, _37863_, _37838_);
  and (_37865_, _37864_, _37657_);
  and (_37866_, _37865_, _37406_);
  and (_37867_, _37232_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_37868_, _37045_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  and (_37869_, _37078_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  or (_37870_, _37869_, _37868_);
  or (_37871_, _37870_, _37867_);
  and (_37872_, _37133_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_37873_, _37872_, _37012_);
  and (_37874_, _37210_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_37875_, _37177_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  nor (_37876_, _37875_, _37874_);
  nand (_37877_, _37876_, _37873_);
  nor (_37878_, _37877_, _37871_);
  and (_37879_, _37878_, _37002_);
  nor (_37880_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], _37002_);
  or (_37881_, _37880_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_37882_, _37881_, _37879_);
  and (_37883_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  or (_37884_, _37883_, _37882_);
  nor (_37885_, _37884_, _37839_);
  not (_37886_, _37885_);
  nor (_37887_, _36958_, \oc8051_top_1.oc8051_decoder1.op [4]);
  nor (_37888_, _37887_, _37363_);
  and (_37889_, _37888_, _37886_);
  not (_37890_, _37889_);
  and (_37891_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_37892_, \oc8051_top_1.oc8051_memory_interface1.cdata [5], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_37893_, _37133_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  and (_37894_, _37177_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor (_37895_, _37894_, _37893_);
  and (_37896_, _37210_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_37897_, _37232_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor (_37898_, _37897_, _37896_);
  and (_37899_, _37045_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  and (_37900_, _37078_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_37901_, _37900_, _37899_);
  and (_37902_, _37901_, _37898_);
  and (_37903_, _37902_, _37895_);
  nor (_37904_, _37903_, _37012_);
  and (_37905_, _37904_, _37002_);
  nor (_37906_, _37905_, _37892_);
  nor (_37907_, _37906_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_37908_, _37907_, _37891_);
  and (_37909_, _37908_, _36969_);
  not (_37910_, _37909_);
  nor (_37911_, _36958_, \oc8051_top_1.oc8051_decoder1.op [5]);
  nor (_37912_, _37911_, _37363_);
  and (_37913_, _37912_, _37910_);
  and (_37914_, \oc8051_top_1.oc8051_memory_interface1.dack_ir , \oc8051_top_1.oc8051_memory_interface1.ddat_ir [7]);
  and (_37915_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  and (_37916_, _37045_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  and (_37917_, _37078_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor (_37918_, _37917_, _37916_);
  and (_37919_, _37133_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  and (_37920_, _37177_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  nor (_37921_, _37920_, _37919_);
  and (_37922_, _37210_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_37923_, _37232_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor (_37924_, _37923_, _37922_);
  and (_37925_, _37924_, _37921_);
  and (_37926_, _37925_, _37918_);
  nor (_37927_, _37926_, _37012_);
  and (_37928_, _37927_, _37002_);
  or (_37929_, _37928_, _37915_);
  and (_37930_, _37929_, _37679_);
  nor (_37931_, _37930_, _37914_);
  and (_37932_, _37931_, _36969_);
  not (_37933_, _37932_);
  nor (_37934_, _36958_, \oc8051_top_1.oc8051_decoder1.op [7]);
  nor (_37935_, _37934_, _37363_);
  and (_37936_, _37935_, _37933_);
  not (_37937_, _37936_);
  and (_37938_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_37939_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_37940_, _37210_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_37941_, _37177_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor (_37942_, _37941_, _37940_);
  and (_37943_, _37078_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  and (_37944_, _37133_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_37945_, _37944_, _37943_);
  and (_37946_, _37045_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  and (_37947_, _37232_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor (_37948_, _37947_, _37946_);
  and (_37949_, _37948_, _37945_);
  and (_37950_, _37949_, _37942_);
  nor (_37951_, _37701_, _37950_);
  nor (_37952_, _37951_, _37939_);
  nor (_37953_, _37952_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_37954_, _37953_, _37938_);
  and (_37955_, _37954_, _36969_);
  not (_37956_, _37955_);
  nor (_37957_, _36958_, \oc8051_top_1.oc8051_decoder1.op [6]);
  nor (_37958_, _37957_, _37363_);
  and (_37959_, _37958_, _37956_);
  nor (_37960_, _37959_, _37937_);
  and (_37961_, _37960_, _37913_);
  and (_37962_, _37961_, _37890_);
  and (_37963_, _37962_, _37866_);
  not (_37964_, _37963_);
  and (_37965_, _37959_, _37913_);
  and (_37966_, _37965_, _37937_);
  and (_37967_, _37966_, _37889_);
  and (_37968_, _37866_, _37967_);
  not (_37969_, _37913_);
  and (_37970_, _37960_, _37969_);
  and (_37971_, _37970_, _37889_);
  and (_37972_, _37971_, _37866_);
  nor (_37973_, _37972_, _37968_);
  and (_37974_, _37973_, _37964_);
  and (_37975_, _37970_, _37890_);
  nor (_37976_, _37863_, _37657_);
  nor (_37977_, _37838_, _37395_);
  and (_37978_, _37977_, _37976_);
  and (_37979_, _37978_, _37975_);
  and (_37980_, _37978_, _37962_);
  nor (_37981_, _37980_, _37979_);
  and (_37982_, _37981_, _37974_);
  nor (_37983_, _37982_, _36914_);
  not (_37984_, _37983_);
  and (_37985_, _37959_, _37937_);
  nor (_37986_, _37837_, _37395_);
  and (_37987_, _37976_, _37986_);
  not (_37988_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and (_37989_, _18772_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_37990_, _37989_, _37988_);
  and (_37991_, _37990_, _37987_);
  and (_37992_, _37991_, _37985_);
  not (_37993_, _36893_);
  nor (_37994_, _37981_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_37995_, _37994_, _37993_);
  nor (_37996_, _37995_, _37992_);
  and (_37997_, _37996_, _37984_);
  nor (_37998_, _37997_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_37999_, _37998_, _36882_);
  and (_38000_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_38001_, _37959_, _37969_);
  and (_38002_, _38001_, _37936_);
  and (_38003_, _38002_, _37890_);
  not (_38004_, _37657_);
  and (_38005_, _37864_, _37406_);
  and (_38006_, _38005_, _38004_);
  and (_38007_, _38006_, _38003_);
  and (_38008_, _37961_, _37889_);
  and (_38009_, _38008_, _38005_);
  and (_38010_, _38009_, _38004_);
  nor (_38011_, _38010_, _38007_);
  and (_38012_, _37987_, _37961_);
  not (_38013_, _37863_);
  and (_38014_, _38013_, _37657_);
  and (_38015_, _38014_, _37977_);
  and (_38016_, _38001_, _37937_);
  and (_38017_, _38016_, _37890_);
  and (_38018_, _38017_, _38015_);
  nor (_38019_, _38018_, _38012_);
  and (_38020_, _38002_, _37889_);
  and (_38021_, _38020_, _38015_);
  nor (_38022_, _37959_, _37936_);
  and (_38023_, _38022_, _37969_);
  and (_38024_, _38023_, _37889_);
  and (_38025_, _38024_, _38015_);
  nor (_38026_, _38025_, _38021_);
  and (_38027_, _37967_, _38006_);
  and (_38028_, _38017_, _38005_);
  nor (_38029_, _38028_, _38027_);
  and (_38030_, _38029_, _38026_);
  and (_38031_, _38030_, _38019_);
  and (_38032_, _38031_, _38011_);
  and (_38033_, _37962_, _38006_);
  and (_38034_, _38020_, _38005_);
  and (_38035_, _38034_, _38004_);
  nor (_38036_, _38035_, _38033_);
  and (_38037_, _38022_, _37913_);
  and (_38038_, _38037_, _37889_);
  and (_38039_, _38038_, _37987_);
  not (_38040_, _38039_);
  and (_38041_, _38037_, _37890_);
  and (_38042_, _38041_, _37987_);
  and (_38043_, _38024_, _37987_);
  nor (_38044_, _38043_, _38042_);
  and (_38045_, _38044_, _38040_);
  and (_38046_, _38023_, _37890_);
  and (_38047_, _38046_, _38015_);
  and (_38048_, _37965_, _37936_);
  and (_38049_, _38048_, _37890_);
  and (_38050_, _38049_, _38015_);
  and (_38051_, _37863_, _37837_);
  and (_38052_, _38051_, _37406_);
  and (_38053_, _38052_, _37890_);
  and (_38054_, _38053_, _37961_);
  or (_38055_, _38054_, _38050_);
  nor (_38056_, _38055_, _38047_);
  and (_38057_, _38056_, _38045_);
  and (_38058_, _38057_, _38036_);
  not (_38059_, _38015_);
  and (_38060_, _38016_, _37889_);
  nor (_38061_, _38060_, _38037_);
  nor (_38062_, _38061_, _38059_);
  not (_38063_, _38062_);
  and (_38064_, _37966_, _37890_);
  and (_38065_, _38064_, _38015_);
  and (_38066_, _38015_, _38003_);
  nor (_38067_, _38066_, _38065_);
  and (_38068_, _37987_, _38002_);
  and (_38069_, _38064_, _38005_);
  nor (_38070_, _38069_, _38068_);
  and (_38071_, _38070_, _38067_);
  and (_38072_, _38071_, _38063_);
  and (_38073_, _37975_, _38006_);
  and (_38074_, _38060_, _38005_);
  nor (_38075_, _38074_, _38073_);
  and (_38076_, _38037_, _38006_);
  and (_38077_, _37962_, _37395_);
  nor (_38078_, _38077_, _38076_);
  and (_38079_, _38078_, _38075_);
  and (_38080_, _37971_, _38006_);
  and (_38081_, _37975_, _38015_);
  nor (_38082_, _38081_, _38080_);
  not (_38083_, _38082_);
  nor (_38084_, _37971_, _38008_);
  nor (_38085_, _38084_, _38059_);
  nor (_38086_, _38085_, _38083_);
  and (_38087_, _38086_, _38079_);
  and (_38088_, _38087_, _38072_);
  and (_38089_, _38088_, _38058_);
  and (_38090_, _38089_, _38032_);
  nor (_38091_, _38090_, _36914_);
  and (_38092_, \oc8051_top_1.oc8051_decoder1.state [0], _18772_);
  and (_38093_, _38092_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_38094_, _38093_, _38076_);
  nor (_38095_, _37992_, _38094_);
  not (_38096_, _38095_);
  nor (_38097_, _38096_, _38091_);
  nor (_38098_, _38097_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_38099_, _38098_, _38000_);
  and (_38100_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_38101_, _37395_, _37890_);
  and (_38102_, _38101_, _38051_);
  and (_38103_, _38102_, _37961_);
  and (_38104_, _38052_, _38023_);
  nor (_38105_, _38104_, _38103_);
  and (_38106_, _37975_, _38052_);
  nor (_38107_, _38106_, _38076_);
  and (_38108_, _38107_, _38105_);
  and (_38109_, _38102_, _38016_);
  and (_38110_, _38052_, _38037_);
  or (_38111_, _38110_, _38109_);
  and (_38112_, _38052_, _38002_);
  and (_38113_, _38102_, _37970_);
  nor (_38114_, _38113_, _38112_);
  not (_38115_, _38114_);
  nor (_38116_, _38115_, _38111_);
  and (_38117_, _38116_, _38108_);
  and (_38118_, _38064_, _38052_);
  not (_38119_, _38118_);
  and (_38120_, _38020_, _37987_);
  not (_38121_, _38053_);
  nor (_38122_, _38048_, _38016_);
  nor (_38123_, _38122_, _38121_);
  nor (_38124_, _38123_, _38120_);
  and (_38125_, _38124_, _38119_);
  and (_38126_, _38125_, _37974_);
  and (_38127_, _38126_, _38117_);
  nor (_38128_, _38127_, _36914_);
  and (_38129_, _37992_, _37913_);
  or (_38130_, _38129_, _38094_);
  nor (_38131_, _38130_, _38128_);
  nor (_38132_, _38131_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_38133_, _38132_, _38100_);
  nor (_38134_, _38133_, _38099_);
  and (_38135_, _38134_, _37999_);
  and (_09484_, _38135_, _42618_);
  and (_38136_, _31212_, _27948_);
  and (_38137_, _27542_, _27345_);
  not (_38138_, _28376_);
  nor (_38139_, _38138_, _28244_);
  and (_38140_, _38139_, _38137_);
  and (_38141_, _38140_, _33118_);
  and (_38142_, _38141_, _28069_);
  and (_38143_, _38142_, _38136_);
  not (_38144_, _38143_);
  and (_38145_, _38144_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor (_38146_, _24187_, _18828_);
  and (_38147_, _28463_, _24165_);
  nor (_38148_, _30958_, _38147_);
  and (_38149_, _38148_, _38146_);
  nor (_38150_, _30827_, _32083_);
  and (_38151_, _38150_, _38149_);
  nor (_38152_, _38151_, _20046_);
  not (_38153_, _38152_);
  and (_38154_, _38153_, _36567_);
  and (_38155_, _38154_, _36437_);
  nor (_38156_, _38155_, _38144_);
  nor (_38157_, _38156_, _38145_);
  and (_38158_, _38144_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor (_38159_, _38151_, _21080_);
  not (_38160_, _38159_);
  and (_38161_, _38160_, _35871_);
  and (_38162_, _38161_, _35718_);
  nor (_38163_, _38162_, _38144_);
  nor (_38164_, _38163_, _38158_);
  and (_38165_, _38144_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  nor (_38166_, _38151_, _21254_);
  not (_38167_, _38166_);
  and (_38168_, _38167_, _35087_);
  and (_38169_, _38168_, _34956_);
  nor (_38170_, _38169_, _38144_);
  nor (_38171_, _38170_, _38165_);
  and (_38172_, _38144_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor (_38173_, _38151_, _21624_);
  not (_38174_, _38173_);
  and (_38175_, _38174_, _34292_);
  and (_38176_, _38175_, _34358_);
  and (_38177_, _38176_, _34260_);
  nor (_38178_, _38177_, _38144_);
  nor (_38179_, _38178_, _38172_);
  and (_38180_, _38144_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_38181_, _38151_, _22147_);
  not (_38182_, _38181_);
  and (_38183_, _38182_, _33477_);
  and (_38184_, _38183_, _33357_);
  nor (_38185_, _38184_, _38144_);
  nor (_38186_, _38185_, _38180_);
  and (_38187_, _38144_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  nor (_38188_, _38151_, _21972_);
  not (_38189_, _38188_);
  and (_38190_, _38189_, _32736_);
  and (_38191_, _38190_, _32922_);
  nor (_38192_, _38191_, _38144_);
  nor (_38193_, _38192_, _38187_);
  and (_38194_, _38136_, _28069_);
  and (_38195_, _38194_, _38141_);
  nor (_38196_, _38195_, _27740_);
  nor (_38197_, _31648_, _30816_);
  nor (_38198_, _38149_, _22517_);
  nor (_38199_, _38198_, _32780_);
  and (_38200_, _38199_, _38197_);
  and (_38201_, _38200_, _32214_);
  and (_38202_, _38201_, _32040_);
  and (_38203_, _38202_, _32073_);
  not (_38204_, _38203_);
  and (_38205_, _38204_, _38143_);
  nor (_38206_, _38205_, _38196_);
  and (_38207_, _38206_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and (_38208_, _38207_, _38193_);
  and (_38209_, _38208_, _38186_);
  and (_38210_, _38209_, _38179_);
  and (_38211_, _38210_, _38171_);
  and (_38212_, _38211_, _38164_);
  and (_38213_, _38212_, _38157_);
  nor (_38214_, _38195_, _28102_);
  nand (_38215_, _38214_, _38213_);
  or (_38216_, _38214_, _38213_);
  and (_38217_, _38216_, _27125_);
  and (_38218_, _38217_, _38215_);
  or (_38219_, _38195_, _28156_);
  or (_38220_, _38219_, _38218_);
  nor (_38221_, _38151_, _20884_);
  not (_38222_, _38221_);
  and (_38223_, _38222_, _30947_);
  and (_38224_, _38223_, _30783_);
  and (_38225_, _38224_, _30522_);
  nand (_38226_, _38225_, _38195_);
  and (_38227_, _38226_, _38220_);
  and (_09504_, _38227_, _42618_);
  not (_38228_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and (_38229_, _38206_, _38228_);
  nor (_38230_, _38206_, _38228_);
  nor (_38231_, _38230_, _38229_);
  and (_38232_, _38231_, _27125_);
  nor (_38233_, _38232_, _27751_);
  nor (_38234_, _38233_, _38143_);
  nor (_38235_, _38234_, _38205_);
  nand (_10660_, _38235_, _42618_);
  nor (_38236_, _38207_, _38193_);
  nor (_38237_, _38236_, _38208_);
  nor (_38238_, _38237_, _27114_);
  nor (_38239_, _38238_, _27586_);
  nor (_38240_, _38239_, _38143_);
  nor (_38241_, _38240_, _38192_);
  nand (_10671_, _38241_, _42618_);
  nor (_38242_, _38208_, _38186_);
  nor (_38243_, _38242_, _38209_);
  nor (_38244_, _38243_, _27114_);
  nor (_38245_, _38244_, _27981_);
  nor (_38246_, _38245_, _38143_);
  nor (_38247_, _38246_, _38185_);
  nand (_10682_, _38247_, _42618_);
  nor (_38248_, _38209_, _38179_);
  nor (_38249_, _38248_, _38210_);
  nor (_38250_, _38249_, _27114_);
  nor (_38251_, _38250_, _27849_);
  nor (_38252_, _38251_, _38143_);
  nor (_38253_, _38252_, _38178_);
  nor (_10693_, _38253_, rst);
  nor (_38254_, _38210_, _38171_);
  nor (_38255_, _38254_, _38211_);
  nor (_38256_, _38255_, _27114_);
  nor (_38257_, _38256_, _27444_);
  nor (_38258_, _38257_, _38143_);
  nor (_38259_, _38258_, _38170_);
  nor (_10704_, _38259_, rst);
  nor (_38260_, _38211_, _38164_);
  nor (_38261_, _38260_, _38212_);
  nor (_38262_, _38261_, _27114_);
  nor (_38263_, _38262_, _27158_);
  nor (_38264_, _38263_, _38143_);
  nor (_38265_, _38264_, _38163_);
  nor (_10715_, _38265_, rst);
  nor (_38266_, _38212_, _38157_);
  nor (_38267_, _38266_, _38213_);
  nor (_38268_, _38267_, _27114_);
  nor (_38269_, _38268_, _28288_);
  nor (_38270_, _38269_, _38143_);
  nor (_38271_, _38270_, _38156_);
  nor (_10726_, _38271_, rst);
  and (_38272_, _38140_, _34576_);
  nand (_38273_, _38272_, _38136_);
  nor (_38274_, _38273_, _31136_);
  and (_38275_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], _18772_);
  and (_38276_, _38275_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_38277_, _38273_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_38278_, _38277_, _38276_);
  or (_38279_, _38278_, _38274_);
  nor (_38280_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  not (_38281_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_38282_, _38281_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38283_, _38282_, _38280_);
  nor (_38284_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  not (_38285_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_38286_, _38285_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38287_, _38286_, _38284_);
  not (_38288_, _38287_);
  nor (_38289_, _38288_, _31299_);
  nor (_38290_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  not (_38291_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_38292_, _38291_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38293_, _38292_, _38290_);
  and (_38294_, _38293_, _38289_);
  nor (_38295_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  not (_38296_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_38297_, _38296_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38298_, _38297_, _38295_);
  and (_38299_, _38298_, _38294_);
  and (_38300_, _38299_, _38283_);
  nor (_38301_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  not (_38302_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_38303_, _38302_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38304_, _38303_, _38301_);
  and (_38305_, _38304_, _38300_);
  nor (_38306_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  not (_38307_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_38308_, _38307_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38309_, _38308_, _38306_);
  and (_38310_, _38309_, _38305_);
  nor (_38311_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  not (_38312_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_38313_, _38312_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38314_, _38313_, _38311_);
  and (_38315_, _38314_, _38310_);
  nor (_38316_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  not (_38317_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_38318_, _38317_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38319_, _38318_, _38316_);
  nand (_38320_, _38319_, _38315_);
  or (_38321_, _38319_, _38315_);
  and (_38322_, _38321_, _28474_);
  and (_38323_, _38322_, _38320_);
  not (_38324_, _38323_);
  and (_38325_, _23879_, _18828_);
  and (_38326_, _29209_, _20372_);
  not (_38327_, _38326_);
  and (_38328_, _30271_, _20895_);
  and (_38329_, _38328_, _29790_);
  and (_38330_, _38329_, _29823_);
  and (_38331_, _38330_, _29867_);
  and (_38332_, _38331_, _30042_);
  nor (_38333_, _38332_, _30293_);
  and (_38334_, _29209_, _19387_);
  nor (_38335_, _38334_, _38333_);
  and (_38336_, _38335_, _38327_);
  and (_38337_, _30358_, _20884_);
  and (_38338_, _20220_, _19222_);
  and (_38339_, _20536_, _19550_);
  and (_38340_, _38339_, _38338_);
  and (_38341_, _38340_, _38337_);
  and (_38342_, _20372_, _19387_);
  and (_38343_, _38342_, _38341_);
  nor (_38344_, _38343_, _29209_);
  not (_38345_, _38344_);
  and (_38346_, _38345_, _38336_);
  nor (_38347_, _29209_, _19724_);
  and (_38348_, _29209_, _19724_);
  nor (_38349_, _38348_, _38347_);
  and (_38350_, _38349_, _38346_);
  and (_38351_, _38350_, _30434_);
  nor (_38352_, _38350_, _30434_);
  nor (_38353_, _38352_, _38351_);
  and (_38354_, _38353_, _30205_);
  and (_38355_, _24187_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  and (_38356_, _29209_, _30434_);
  nor (_38357_, _38356_, _31387_);
  nor (_38358_, _38357_, _30489_);
  nor (_38359_, _31627_, _21624_);
  nor (_38360_, _30968_, _20719_);
  or (_38361_, _38360_, _38359_);
  or (_38362_, _38361_, _38358_);
  nor (_38363_, _38362_, _38355_);
  not (_38364_, _38363_);
  nor (_38365_, _38364_, _38354_);
  not (_38366_, _38365_);
  nor (_38367_, _38366_, _38325_);
  and (_38368_, _38367_, _38324_);
  nand (_38369_, _38368_, _38276_);
  and (_38370_, _38369_, _42618_);
  and (_12677_, _38370_, _38279_);
  and (_38371_, _38140_, _33847_);
  and (_38372_, _38371_, _38136_);
  nor (_38373_, _38372_, _38276_);
  not (_38374_, _38373_);
  nand (_38375_, _38374_, _31136_);
  or (_38376_, _38374_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_38377_, _38376_, _42618_);
  and (_12698_, _38377_, _38375_);
  nor (_38378_, _38273_, _32323_);
  and (_38379_, _38273_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or (_38380_, _38379_, _38276_);
  or (_38381_, _38380_, _38378_);
  and (_38382_, _26458_, _24187_);
  not (_38383_, _38382_);
  and (_38384_, _38288_, _31299_);
  nor (_38385_, _38384_, _38289_);
  and (_38386_, _38385_, _28474_);
  nor (_38387_, _31387_, _30467_);
  not (_38388_, _38387_);
  nor (_38389_, _38388_, _30380_);
  nor (_38390_, _38389_, _29790_);
  and (_38391_, _38389_, _29790_);
  or (_38392_, _38391_, _33313_);
  nor (_38393_, _38392_, _38390_);
  nor (_38394_, _30968_, _19550_);
  and (_38395_, _23658_, _18828_);
  nor (_38396_, _31627_, _21254_);
  nor (_38397_, _30489_, _22517_);
  or (_38398_, _38397_, _38396_);
  or (_38399_, _38398_, _38395_);
  nor (_38400_, _38399_, _38394_);
  not (_38401_, _38400_);
  nor (_38402_, _38401_, _38393_);
  not (_38403_, _38402_);
  nor (_38404_, _38403_, _38386_);
  and (_38405_, _38404_, _38383_);
  nand (_38406_, _38405_, _38276_);
  and (_38407_, _38406_, _42618_);
  and (_13613_, _38407_, _38381_);
  nor (_38408_, _38273_, _33020_);
  and (_38409_, _38273_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_38410_, _38409_, _38276_);
  or (_38411_, _38410_, _38408_);
  nor (_38412_, _38293_, _38289_);
  nor (_38413_, _38412_, _38294_);
  and (_38414_, _38413_, _28474_);
  not (_38415_, _38414_);
  and (_38416_, _25472_, _24187_);
  nor (_38417_, _38329_, _30293_);
  and (_38418_, _38337_, _19550_);
  nor (_38419_, _38418_, _29209_);
  or (_38420_, _38419_, _38417_);
  nor (_38421_, _38420_, _29823_);
  and (_38422_, _38420_, _29823_);
  or (_38423_, _38422_, _38421_);
  and (_38424_, _38423_, _30205_);
  nor (_38425_, _30968_, _20536_);
  and (_38426_, _23689_, _18828_);
  nor (_38427_, _31627_, _21080_);
  nor (_38428_, _30489_, _21972_);
  or (_38429_, _38428_, _38427_);
  or (_38430_, _38429_, _38426_);
  nor (_38431_, _38430_, _38425_);
  not (_38432_, _38431_);
  nor (_38433_, _38432_, _38424_);
  not (_38434_, _38433_);
  nor (_38435_, _38434_, _38416_);
  and (_38436_, _38435_, _38415_);
  nand (_38437_, _38436_, _38276_);
  and (_38438_, _38437_, _42618_);
  and (_13624_, _38438_, _38411_);
  nor (_38439_, _38273_, _33717_);
  and (_38440_, _38273_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_38441_, _38440_, _38276_);
  or (_38442_, _38441_, _38439_);
  nor (_38443_, _38298_, _38294_);
  nor (_38444_, _38443_, _38299_);
  and (_38445_, _38444_, _28474_);
  not (_38446_, _38445_);
  and (_38447_, _38418_, _20536_);
  and (_38448_, _38447_, _30293_);
  and (_38449_, _38330_, _29209_);
  nor (_38450_, _38449_, _38448_);
  and (_38451_, _38450_, _19222_);
  nor (_38452_, _38450_, _19222_);
  nor (_38453_, _38452_, _38451_);
  and (_38454_, _38453_, _30205_);
  not (_38455_, _38454_);
  nor (_38456_, _30489_, _22147_);
  and (_38457_, _24187_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  nor (_38458_, _38457_, _38456_);
  and (_38459_, _23721_, _18828_);
  nor (_38460_, _31627_, _20046_);
  nor (_38461_, _30968_, _19222_);
  or (_38462_, _38461_, _38460_);
  nor (_38463_, _38462_, _38459_);
  and (_38464_, _38463_, _38458_);
  and (_38465_, _38464_, _38455_);
  and (_38466_, _38465_, _38446_);
  nand (_38467_, _38466_, _38276_);
  and (_38468_, _38467_, _42618_);
  and (_13635_, _38468_, _38442_);
  nor (_38469_, _38273_, _34478_);
  and (_38470_, _38273_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_38471_, _38470_, _38276_);
  or (_38472_, _38471_, _38469_);
  nor (_38473_, _38299_, _38283_);
  nor (_38474_, _38473_, _38300_);
  and (_38475_, _38474_, _28474_);
  not (_38476_, _38475_);
  and (_38477_, _23753_, _18828_);
  not (_38478_, _38477_);
  nor (_38479_, _38331_, _30042_);
  not (_38480_, _38479_);
  and (_38481_, _38480_, _38333_);
  and (_38482_, _38447_, _19222_);
  nor (_38483_, _38482_, _20220_);
  nor (_38484_, _38483_, _38341_);
  nor (_38485_, _38484_, _29209_);
  nor (_38486_, _38485_, _38481_);
  nor (_38487_, _38486_, _33313_);
  nor (_38488_, _30968_, _20220_);
  nor (_38489_, _30489_, _21624_);
  and (_38490_, _24187_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  or (_38491_, _38490_, _38489_);
  or (_38492_, _38491_, _31647_);
  nor (_38493_, _38492_, _38488_);
  not (_38494_, _38493_);
  nor (_38495_, _38494_, _38487_);
  and (_38496_, _38495_, _38478_);
  and (_38497_, _38496_, _38476_);
  nand (_38498_, _38497_, _38276_);
  and (_38499_, _38498_, _42618_);
  and (_13646_, _38499_, _38472_);
  nor (_38500_, _38273_, _35240_);
  and (_38501_, _38273_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or (_38502_, _38501_, _38276_);
  or (_38503_, _38502_, _38500_);
  nor (_38504_, _38304_, _38300_);
  nor (_38505_, _38504_, _38305_);
  and (_38506_, _38505_, _28474_);
  not (_38507_, _38506_);
  and (_38508_, _23784_, _18828_);
  nor (_38509_, _38341_, _29209_);
  nor (_38510_, _38509_, _38333_);
  nor (_38511_, _38510_, _29637_);
  and (_38512_, _38510_, _29637_);
  nor (_38513_, _38512_, _38511_);
  and (_38514_, _38513_, _30205_);
  and (_38515_, _24187_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  nor (_38516_, _29209_, _21265_);
  or (_38517_, _38516_, _30489_);
  nor (_38518_, _38517_, _38334_);
  nor (_38519_, _31627_, _22517_);
  nor (_38520_, _30968_, _19387_);
  or (_38521_, _38520_, _38519_);
  or (_38522_, _38521_, _38518_);
  nor (_38523_, _38522_, _38515_);
  not (_38524_, _38523_);
  nor (_38525_, _38524_, _38514_);
  not (_38526_, _38525_);
  nor (_38527_, _38526_, _38508_);
  and (_38528_, _38527_, _38507_);
  nand (_38529_, _38528_, _38276_);
  and (_38530_, _38529_, _42618_);
  and (_13657_, _38530_, _38503_);
  nor (_38531_, _38273_, _36046_);
  and (_38532_, _38273_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or (_38533_, _38532_, _38276_);
  or (_38534_, _38533_, _38531_);
  nor (_38535_, _38309_, _38305_);
  not (_38536_, _38535_);
  nor (_38537_, _38310_, _31278_);
  and (_38538_, _38537_, _38536_);
  not (_38539_, _38538_);
  and (_38540_, _23816_, _18828_);
  and (_38541_, _38341_, _19387_);
  nor (_38542_, _38541_, _29209_);
  not (_38543_, _38542_);
  and (_38544_, _38543_, _38335_);
  and (_38545_, _38544_, _20372_);
  nor (_38546_, _38544_, _20372_);
  nor (_38547_, _38546_, _38545_);
  nor (_38548_, _38547_, _33313_);
  and (_38549_, _24187_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  nor (_38550_, _36350_, _30489_);
  and (_38551_, _38550_, _38327_);
  nor (_38552_, _31627_, _21972_);
  nor (_38553_, _30968_, _20372_);
  or (_38554_, _38553_, _38552_);
  or (_38555_, _38554_, _38551_);
  nor (_38556_, _38555_, _38549_);
  not (_38557_, _38556_);
  nor (_38558_, _38557_, _38548_);
  not (_38559_, _38558_);
  nor (_38560_, _38559_, _38540_);
  and (_38561_, _38560_, _38539_);
  nand (_38562_, _38561_, _38276_);
  and (_38563_, _38562_, _42618_);
  and (_13668_, _38563_, _38534_);
  or (_38564_, _38273_, _36698_);
  not (_38565_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  nand (_38566_, _38273_, _38565_);
  and (_38567_, _38566_, _38564_);
  or (_38568_, _38567_, _38276_);
  not (_38569_, _38276_);
  nor (_38570_, _38314_, _38310_);
  nor (_38571_, _38570_, _38315_);
  and (_38572_, _38571_, _28474_);
  and (_38573_, _23848_, _18828_);
  and (_38574_, _38346_, _19724_);
  nor (_38575_, _38346_, _19724_);
  or (_38576_, _38575_, _38574_);
  and (_38577_, _38576_, _30205_);
  or (_38578_, _29209_, _20057_);
  nor (_38579_, _38348_, _30489_);
  and (_38580_, _38579_, _38578_);
  nor (_38581_, _31627_, _22147_);
  nor (_38582_, _30968_, _19724_);
  and (_38583_, _24187_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  or (_38584_, _38583_, _38582_);
  or (_38585_, _38584_, _38581_);
  or (_38586_, _38585_, _38580_);
  or (_38587_, _38586_, _38577_);
  or (_38588_, _38587_, _38573_);
  or (_38589_, _38588_, _38572_);
  or (_38590_, _38589_, _38569_);
  and (_38591_, _38590_, _42618_);
  and (_13679_, _38591_, _38568_);
  nand (_38592_, _38374_, _32323_);
  or (_38593_, _38374_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_38594_, _38593_, _42618_);
  and (_13690_, _38594_, _38592_);
  nand (_38595_, _38374_, _33020_);
  or (_38596_, _38374_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_38597_, _38596_, _42618_);
  and (_13701_, _38597_, _38595_);
  nand (_38598_, _38374_, _33717_);
  or (_38599_, _38374_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_38600_, _38599_, _42618_);
  and (_13711_, _38600_, _38598_);
  nand (_38601_, _38374_, _34478_);
  or (_38602_, _38374_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_38603_, _38602_, _42618_);
  and (_13722_, _38603_, _38601_);
  nand (_38604_, _38374_, _35240_);
  or (_38605_, _38374_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_38606_, _38605_, _42618_);
  and (_13733_, _38606_, _38604_);
  nand (_38607_, _38374_, _36046_);
  or (_38608_, _38374_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_38609_, _38608_, _42618_);
  and (_13744_, _38609_, _38607_);
  or (_38610_, _38373_, _36698_);
  or (_38611_, _38374_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_38612_, _38611_, _42618_);
  and (_13755_, _38612_, _38610_);
  not (_38613_, _27345_);
  nor (_38614_, _28376_, _38613_);
  and (_38615_, _38614_, _31899_);
  and (_38616_, _38615_, _31812_);
  not (_38617_, _31855_);
  nor (_38618_, _38617_, _31757_);
  not (_38619_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_38620_, _31855_, _38619_);
  or (_38621_, _38620_, _38618_);
  and (_38622_, _38621_, _38616_);
  nor (_38623_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  not (_38624_, _38623_);
  nand (_38625_, _38624_, _31757_);
  and (_38626_, _38623_, _38619_);
  nor (_38627_, _38626_, _38616_);
  and (_38628_, _38627_, _38625_);
  nor (_38629_, _27542_, _38613_);
  and (_38630_, _31212_, _28398_);
  and (_38631_, _38630_, _38629_);
  or (_38632_, _38631_, _38628_);
  or (_38633_, _38632_, _38622_);
  nand (_38634_, _38631_, _38225_);
  and (_38635_, _38634_, _42618_);
  and (_15158_, _38635_, _38633_);
  and (_38636_, _38616_, _33129_);
  nand (_38637_, _38636_, _31757_);
  not (_38638_, _38631_);
  or (_38639_, _38636_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_38640_, _38639_, _38638_);
  and (_38641_, _38640_, _38637_);
  nor (_38642_, _38638_, _38191_);
  or (_38645_, _38642_, _38641_);
  and (_17339_, _38645_, _42618_);
  or (_38647_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_38648_, _23943_, _23911_);
  or (_38649_, _38648_, _23974_);
  or (_38650_, _38649_, _24017_);
  or (_38651_, _38650_, _24048_);
  or (_38652_, _38651_, _24091_);
  or (_38653_, _38652_, _24122_);
  or (_38654_, _38653_, _23594_);
  and (_38655_, _38654_, _18828_);
  or (_38657_, _31342_, _30140_);
  not (_38666_, _31321_);
  nand (_38672_, _38666_, _30140_);
  and (_38678_, _38672_, _29582_);
  and (_38681_, _38678_, _38657_);
  not (_38682_, _29461_);
  nand (_38683_, _29450_, _38682_);
  or (_38684_, _29472_, _29450_);
  and (_38685_, _28474_, _38684_);
  and (_38686_, _38685_, _38683_);
  and (_38687_, _38342_, _25373_);
  and (_38688_, _38340_, _24187_);
  nand (_38689_, _38688_, _38687_);
  nand (_38690_, _38689_, \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or (_38691_, _38690_, _38686_);
  or (_38692_, _38691_, _38681_);
  or (_38693_, _38692_, _38655_);
  and (_38694_, _38693_, _38647_);
  or (_38695_, _38694_, _38616_);
  not (_38696_, _38616_);
  and (_38697_, _33858_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_38698_, _38697_, _33869_);
  or (_38699_, _38698_, _38696_);
  and (_38700_, _38699_, _38695_);
  or (_38701_, _38700_, _38631_);
  nand (_38702_, _38631_, _38184_);
  and (_38703_, _38702_, _42618_);
  and (_17350_, _38703_, _38701_);
  and (_38704_, _38616_, _34576_);
  nand (_38707_, _38704_, _31757_);
  or (_38708_, _38704_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_38709_, _38708_, _38638_);
  and (_38710_, _38709_, _38707_);
  nor (_38711_, _38638_, _38177_);
  or (_38712_, _38711_, _38710_);
  and (_17361_, _38712_, _42618_);
  or (_38713_, _38696_, _35360_);
  nor (_38714_, _38638_, _38169_);
  and (_38715_, _38638_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  nor (_38716_, _38715_, _38714_);
  nor (_38743_, _38716_, rst);
  and (_38717_, _38743_, _38713_);
  and (_38718_, _35349_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  or (_38719_, _38718_, _35393_);
  and (_38720_, _38616_, _42618_);
  and (_38721_, _38720_, _38719_);
  or (_17372_, _38721_, _38717_);
  and (_38722_, _38616_, _36133_);
  nand (_38723_, _38722_, _31757_);
  or (_38724_, _38722_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_38725_, _38724_, _38638_);
  and (_38726_, _38725_, _38723_);
  nor (_38727_, _38638_, _38162_);
  or (_38728_, _38727_, _38726_);
  and (_17383_, _38728_, _42618_);
  and (_38729_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or (_38730_, _38729_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_38731_, _30096_, _29582_);
  and (_38732_, _28474_, _29352_);
  nand (_38733_, _30958_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nand (_38734_, _38733_, _38729_);
  or (_38735_, _38734_, _38732_);
  or (_38736_, _38735_, _38731_);
  and (_38737_, _38736_, _38730_);
  or (_38738_, _38737_, _38616_);
  not (_38739_, _36785_);
  nor (_38740_, _38739_, _31757_);
  or (_38742_, _36785_, _34086_);
  nand (_38746_, _38742_, _38616_);
  or (_38752_, _38746_, _38740_);
  and (_38757_, _38752_, _38738_);
  or (_38764_, _38757_, _38631_);
  nand (_38772_, _38631_, _38155_);
  and (_38780_, _38772_, _42618_);
  and (_17394_, _38780_, _38764_);
  not (_38781_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_38782_, _38275_, _38781_);
  and (_38783_, _38782_, _38368_);
  nor (_38784_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_38785_, _38784_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_38786_, _27542_, _38613_);
  and (_38787_, _38786_, _28387_);
  and (_38788_, _38787_, _28091_);
  and (_38789_, _38788_, _31212_);
  nor (_38790_, _38789_, _38785_);
  nor (_38791_, _38790_, _31136_);
  and (_38792_, _27948_, _27542_);
  and (_38793_, _38792_, _31768_);
  not (_38794_, _31899_);
  nor (_38795_, _38794_, _28244_);
  and (_38796_, _38795_, _38793_);
  and (_38797_, _38796_, _31855_);
  and (_38798_, _38797_, _31757_);
  nor (_38799_, _38797_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  not (_38800_, _38799_);
  not (_38801_, _38782_);
  and (_38802_, _38790_, _38801_);
  and (_38803_, _38802_, _38800_);
  not (_38804_, _38803_);
  nor (_38805_, _38804_, _38798_);
  nor (_38806_, _38805_, _38782_);
  not (_38807_, _38806_);
  nor (_38808_, _38807_, _38791_);
  nor (_38809_, _38808_, _38783_);
  and (_17963_, _38809_, _42618_);
  nor (_38810_, _38801_, _38405_);
  not (_38811_, _38790_);
  and (_38812_, _38811_, _32323_);
  and (_38813_, _27806_, _28069_);
  and (_38814_, _32410_, _38813_);
  not (_38815_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_38821_, _38813_, _38815_);
  nor (_38832_, _38821_, _38814_);
  and (_38833_, _38796_, _38801_);
  not (_38834_, _38833_);
  nor (_38835_, _38834_, _38832_);
  nor (_38846_, _38796_, _38815_);
  nor (_38852_, _38846_, _38811_);
  nor (_38853_, _38852_, _38782_);
  or (_38854_, _38853_, _38835_);
  not (_38855_, _38854_);
  nor (_38856_, _38855_, _38812_);
  nor (_38857_, _38856_, _38810_);
  nor (_19757_, _38857_, rst);
  nor (_38858_, _38801_, _38436_);
  and (_38859_, _38811_, _33020_);
  not (_38860_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor (_38861_, _38796_, _38860_);
  nor (_38862_, _38861_, _38811_);
  not (_38863_, _33129_);
  nor (_38864_, _38863_, _31757_);
  nor (_38865_, _33129_, _38860_);
  nor (_38866_, _38865_, _38864_);
  nand (_38867_, _38802_, _38796_);
  or (_38868_, _38867_, _38866_);
  and (_38869_, _38868_, _38862_);
  or (_38870_, _38869_, _38782_);
  nor (_38871_, _38870_, _38859_);
  nor (_38872_, _38871_, _38858_);
  nor (_19769_, _38872_, rst);
  nor (_38873_, _38801_, _38466_);
  and (_38874_, _38811_, _33717_);
  not (_38875_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor (_38876_, _38796_, _38875_);
  nor (_38877_, _38876_, _38811_);
  not (_38878_, _38877_);
  not (_38879_, _38796_);
  nor (_38880_, _33847_, _38875_);
  nor (_38881_, _38880_, _33869_);
  nor (_38882_, _38881_, _38879_);
  nor (_38883_, _38882_, _38878_);
  nor (_38884_, _38883_, _38782_);
  not (_38885_, _38884_);
  nor (_38886_, _38885_, _38874_);
  nor (_38887_, _38886_, _38873_);
  nor (_19780_, _38887_, rst);
  nor (_38888_, _38790_, _34478_);
  and (_38889_, _38802_, _38879_);
  and (_38890_, _38889_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor (_38891_, _38890_, _38888_);
  and (_38892_, _34587_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor (_38893_, _38892_, _34598_);
  nor (_38894_, _38893_, _38834_);
  and (_38895_, _38894_, _38790_);
  nor (_38896_, _38895_, _38782_);
  and (_38897_, _38896_, _38891_);
  and (_38898_, _38782_, _38497_);
  or (_38899_, _38898_, _38897_);
  nor (_19792_, _38899_, rst);
  nor (_38900_, _38790_, _35240_);
  and (_38901_, _38796_, _35338_);
  and (_38902_, _38901_, _31757_);
  nor (_38903_, _38901_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  not (_38904_, _38903_);
  and (_38905_, _38904_, _38802_);
  not (_38906_, _38905_);
  nor (_38907_, _38906_, _38902_);
  or (_38908_, _38907_, _38900_);
  and (_38909_, _38908_, _38801_);
  nor (_38910_, _38801_, _38528_);
  or (_38911_, _38910_, _38909_);
  and (_19804_, _38911_, _42618_);
  nor (_38912_, _38790_, _36046_);
  and (_38913_, _38796_, _36133_);
  nor (_38914_, _38913_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  not (_38915_, _38914_);
  not (_38916_, _38802_);
  and (_38917_, _38913_, _31757_);
  nor (_38918_, _38917_, _38916_);
  and (_38919_, _38918_, _38915_);
  or (_38920_, _38919_, _38912_);
  and (_38921_, _38920_, _38801_);
  nor (_38922_, _38801_, _38561_);
  or (_38923_, _38922_, _38921_);
  and (_19816_, _38923_, _42618_);
  or (_38924_, _38801_, _38589_);
  and (_38925_, _38811_, _36698_);
  and (_38926_, _38796_, _36785_);
  or (_38927_, _38926_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nand (_38928_, _38926_, _31757_);
  and (_38929_, _38928_, _38802_);
  and (_38930_, _38929_, _38927_);
  or (_38931_, _38930_, _38782_);
  or (_38932_, _38931_, _38925_);
  and (_38933_, _38932_, _38924_);
  and (_19828_, _38933_, _42618_);
  and (_38934_, _28376_, _27345_);
  and (_38935_, _38792_, _31779_);
  and (_38936_, _38935_, _38934_);
  and (_38937_, _38936_, _31855_);
  nand (_38938_, _38937_, _31757_);
  or (_38939_, _38937_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_38940_, _38939_, _31899_);
  and (_38941_, _38940_, _38938_);
  and (_38942_, _38140_, _28091_);
  nand (_38943_, _38942_, _38225_);
  or (_38944_, _38942_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_38945_, _38944_, _31212_);
  and (_38946_, _38945_, _38943_);
  not (_38947_, _31211_);
  and (_38948_, _38947_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  or (_38949_, _38948_, rst);
  or (_38950_, _38949_, _38946_);
  or (_31034_, _38950_, _38941_);
  and (_38951_, _38934_, _31812_);
  and (_38952_, _38951_, _31855_);
  nand (_38953_, _38952_, _31757_);
  or (_38954_, _38952_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_38955_, _38954_, _31899_);
  and (_38956_, _38955_, _38953_);
  and (_38957_, _38629_, _38139_);
  and (_38958_, _38957_, _28091_);
  nand (_38959_, _38958_, _38225_);
  or (_38960_, _38958_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_38961_, _38960_, _31212_);
  and (_38962_, _38961_, _38959_);
  and (_38963_, _38947_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  or (_38964_, _38963_, rst);
  or (_38965_, _38964_, _38962_);
  or (_31057_, _38965_, _38956_);
  and (_38966_, _28376_, _38613_);
  and (_38967_, _38966_, _38935_);
  and (_38968_, _38967_, _31855_);
  nand (_38969_, _38968_, _31757_);
  or (_38970_, _38968_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_38971_, _38970_, _31899_);
  and (_38972_, _38971_, _38969_);
  and (_38973_, _38786_, _38139_);
  and (_38974_, _38973_, _28091_);
  not (_38975_, _38974_);
  nor (_38976_, _38975_, _38225_);
  and (_38977_, _38975_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or (_38978_, _38977_, _38976_);
  and (_38979_, _38978_, _31212_);
  and (_38980_, _38947_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or (_38981_, _38980_, rst);
  or (_38982_, _38981_, _38979_);
  or (_31079_, _38982_, _38972_);
  and (_38983_, _38966_, _31812_);
  and (_38984_, _38983_, _31855_);
  nand (_38985_, _38984_, _31757_);
  or (_38986_, _38984_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and (_38987_, _38986_, _31899_);
  and (_38988_, _38987_, _38985_);
  and (_38989_, _38139_, _27553_);
  and (_38990_, _38989_, _28091_);
  not (_38991_, _38990_);
  nor (_38992_, _38991_, _38225_);
  and (_38993_, _38991_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or (_38994_, _38993_, _38992_);
  and (_38995_, _38994_, _31212_);
  and (_38996_, _38947_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or (_38997_, _38996_, rst);
  or (_38998_, _38997_, _38995_);
  or (_31102_, _38998_, _38988_);
  or (_38999_, _38942_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  and (_39000_, _38999_, _31899_);
  and (_39001_, _38936_, _38813_);
  nand (_39002_, _39001_, _31757_);
  and (_39003_, _39002_, _39000_);
  nand (_39004_, _38942_, _38203_);
  and (_39005_, _39004_, _31212_);
  and (_39006_, _39005_, _38999_);
  not (_39007_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  nor (_39008_, _31211_, _39007_);
  or (_39009_, _39008_, rst);
  or (_39010_, _39009_, _39006_);
  or (_40308_, _39010_, _39003_);
  and (_39011_, _33118_, _28080_);
  and (_39012_, _39011_, _38140_);
  nand (_39013_, _39012_, _31757_);
  or (_39014_, _39012_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_39015_, _39014_, _31899_);
  and (_39016_, _39015_, _39013_);
  nand (_39017_, _38942_, _38191_);
  or (_39018_, _38942_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_39019_, _39018_, _31212_);
  and (_39020_, _39019_, _39017_);
  and (_39021_, _38947_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  or (_39022_, _39021_, rst);
  or (_39023_, _39022_, _39020_);
  or (_40310_, _39023_, _39016_);
  not (_39024_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  not (_39025_, _34609_);
  and (_39026_, _38936_, _39025_);
  nor (_39035_, _39026_, _39024_);
  and (_39046_, _33880_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or (_39057_, _39046_, _33869_);
  and (_39066_, _39057_, _38936_);
  or (_39072_, _39066_, _39035_);
  and (_39083_, _39072_, _31899_);
  nand (_39094_, _38942_, _38184_);
  or (_39105_, _38942_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_39116_, _39105_, _31212_);
  and (_39127_, _39116_, _39094_);
  nor (_39138_, _31211_, _39024_);
  or (_39149_, _39138_, rst);
  or (_39160_, _39149_, _39127_);
  or (_40312_, _39160_, _39083_);
  and (_39181_, _38936_, _34576_);
  nand (_39192_, _39181_, _31757_);
  or (_39203_, _39181_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_39214_, _39203_, _31899_);
  and (_39225_, _39214_, _39192_);
  nand (_39236_, _38942_, _38177_);
  or (_39240_, _38942_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_39241_, _39240_, _31212_);
  and (_39242_, _39241_, _39236_);
  and (_39243_, _38947_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or (_39244_, _39243_, rst);
  or (_39245_, _39244_, _39242_);
  or (_40314_, _39245_, _39225_);
  not (_39246_, _38936_);
  or (_39247_, _39246_, _35360_);
  and (_39248_, _39247_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_39249_, _35349_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or (_39250_, _39249_, _35393_);
  and (_39251_, _39250_, _38936_);
  or (_39252_, _39251_, _39248_);
  and (_39253_, _39252_, _31899_);
  nand (_39254_, _38942_, _38169_);
  or (_39255_, _38942_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_39256_, _39255_, _31212_);
  and (_39257_, _39256_, _39254_);
  not (_39258_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  nor (_39259_, _31211_, _39258_);
  or (_39260_, _39259_, rst);
  or (_39261_, _39260_, _39257_);
  or (_40316_, _39261_, _39253_);
  and (_39262_, _38936_, _36133_);
  nand (_39263_, _39262_, _31757_);
  or (_39264_, _39262_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_39265_, _39264_, _31899_);
  and (_39266_, _39265_, _39263_);
  nand (_39267_, _38942_, _38162_);
  or (_39268_, _38942_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_39269_, _39268_, _31212_);
  and (_39270_, _39269_, _39267_);
  and (_39271_, _38947_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  or (_39272_, _39271_, rst);
  or (_39273_, _39272_, _39270_);
  or (_40318_, _39273_, _39266_);
  and (_39274_, _38936_, _36785_);
  nand (_39275_, _39274_, _31757_);
  or (_39276_, _39274_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_39277_, _39276_, _31899_);
  and (_39278_, _39277_, _39275_);
  nand (_39279_, _38942_, _38155_);
  or (_39280_, _38942_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_39281_, _39280_, _31212_);
  and (_39282_, _39281_, _39279_);
  and (_39283_, _38947_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  or (_39284_, _39283_, rst);
  or (_39285_, _39284_, _39282_);
  or (_40320_, _39285_, _39278_);
  and (_39286_, _38951_, _38813_);
  nand (_39287_, _39286_, _31757_);
  or (_39288_, _38958_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and (_39289_, _39288_, _31899_);
  and (_39290_, _39289_, _39287_);
  nand (_39291_, _38958_, _38203_);
  and (_39292_, _39291_, _31212_);
  and (_39293_, _39292_, _39288_);
  not (_39294_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  nor (_39295_, _31211_, _39294_);
  or (_39296_, _39295_, rst);
  or (_39297_, _39296_, _39293_);
  or (_40322_, _39297_, _39290_);
  and (_39298_, _38951_, _33129_);
  nand (_39299_, _39298_, _31757_);
  or (_39300_, _39298_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_39301_, _39300_, _31899_);
  and (_39302_, _39301_, _39299_);
  nand (_39303_, _38958_, _38191_);
  or (_39304_, _38958_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_39305_, _39304_, _31212_);
  and (_39306_, _39305_, _39303_);
  and (_39307_, _38947_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  or (_39308_, _39307_, rst);
  or (_39309_, _39308_, _39306_);
  or (_40324_, _39309_, _39302_);
  and (_39310_, _38951_, _33847_);
  nand (_39311_, _39310_, _31757_);
  or (_39312_, _39310_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_39313_, _39312_, _31899_);
  and (_39314_, _39313_, _39311_);
  nand (_39315_, _38958_, _38184_);
  or (_39316_, _38958_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_39317_, _39316_, _31212_);
  and (_39318_, _39317_, _39315_);
  and (_39319_, _38947_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  or (_39320_, _39319_, rst);
  or (_39321_, _39320_, _39318_);
  or (_40326_, _39321_, _39314_);
  and (_39322_, _38951_, _34576_);
  nand (_39323_, _39322_, _31757_);
  or (_39324_, _39322_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_39325_, _39324_, _31899_);
  and (_39326_, _39325_, _39323_);
  nand (_39327_, _38958_, _38177_);
  or (_39328_, _38958_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_39329_, _39328_, _31212_);
  and (_39330_, _39329_, _39327_);
  and (_39331_, _38947_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or (_39332_, _39331_, rst);
  or (_39333_, _39332_, _39330_);
  or (_40327_, _39333_, _39326_);
  and (_39334_, _38951_, _35338_);
  nand (_39335_, _39334_, _31757_);
  or (_39336_, _39334_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_39337_, _39336_, _31899_);
  and (_39338_, _39337_, _39335_);
  nand (_39339_, _38958_, _38169_);
  or (_39340_, _38958_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_39341_, _39340_, _31212_);
  and (_39342_, _39341_, _39339_);
  not (_39343_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  nor (_39344_, _31211_, _39343_);
  or (_39345_, _39344_, rst);
  or (_39346_, _39345_, _39342_);
  or (_40329_, _39346_, _39338_);
  and (_39347_, _38951_, _36133_);
  nand (_39348_, _39347_, _31757_);
  or (_39349_, _39347_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_39350_, _39349_, _31899_);
  and (_39351_, _39350_, _39348_);
  nand (_39352_, _38958_, _38162_);
  or (_39353_, _38958_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_39354_, _39353_, _31212_);
  and (_39355_, _39354_, _39352_);
  and (_39356_, _38947_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  or (_39357_, _39356_, rst);
  or (_39358_, _39357_, _39355_);
  or (_40331_, _39358_, _39351_);
  and (_39359_, _38951_, _36785_);
  nand (_39360_, _39359_, _31757_);
  or (_39361_, _39359_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_39362_, _39361_, _31899_);
  and (_39363_, _39362_, _39360_);
  nand (_39364_, _38958_, _38155_);
  or (_39365_, _38958_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_39366_, _39365_, _31212_);
  and (_39367_, _39366_, _39364_);
  and (_39368_, _38947_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  or (_39369_, _39368_, rst);
  or (_39370_, _39369_, _39367_);
  or (_40333_, _39370_, _39363_);
  nand (_39371_, _38974_, _31757_);
  or (_39372_, _38974_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and (_39373_, _39372_, _31899_);
  and (_39374_, _39373_, _39371_);
  nor (_39375_, _38975_, _38203_);
  not (_39376_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  nor (_39377_, _38974_, _39376_);
  or (_39378_, _39377_, _39375_);
  and (_39379_, _39378_, _31212_);
  nor (_39380_, _31211_, _39376_);
  or (_39381_, _39380_, rst);
  or (_39382_, _39381_, _39379_);
  or (_40335_, _39382_, _39374_);
  and (_39383_, _38967_, _33129_);
  nand (_39384_, _39383_, _31757_);
  or (_39385_, _39383_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_39386_, _39385_, _31899_);
  and (_39387_, _39386_, _39384_);
  nor (_39388_, _38975_, _38191_);
  and (_39389_, _38975_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or (_39390_, _39389_, _39388_);
  and (_39391_, _39390_, _31212_);
  and (_39392_, _38947_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or (_39393_, _39392_, rst);
  or (_39394_, _39393_, _39391_);
  or (_40337_, _39394_, _39387_);
  and (_39395_, _38967_, _33847_);
  nand (_39396_, _39395_, _31757_);
  or (_39397_, _39395_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_39398_, _39397_, _31899_);
  and (_39399_, _39398_, _39396_);
  nor (_39400_, _38975_, _38184_);
  and (_39401_, _38975_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or (_39402_, _39401_, _39400_);
  and (_39403_, _39402_, _31212_);
  and (_39404_, _38947_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or (_39405_, _39404_, rst);
  or (_39406_, _39405_, _39403_);
  or (_40339_, _39406_, _39399_);
  and (_39407_, _38967_, _34576_);
  nand (_39408_, _39407_, _31757_);
  or (_39409_, _39407_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_39410_, _39409_, _31899_);
  and (_39411_, _39410_, _39408_);
  nor (_39412_, _38975_, _38177_);
  and (_39413_, _38975_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_39414_, _39413_, _39412_);
  and (_39415_, _39414_, _31212_);
  and (_39416_, _38947_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_39417_, _39416_, rst);
  or (_39418_, _39417_, _39415_);
  or (_40341_, _39418_, _39411_);
  and (_39419_, _38967_, _35338_);
  nand (_39420_, _39419_, _31757_);
  or (_39421_, _39419_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_39422_, _39421_, _31899_);
  and (_39423_, _39422_, _39420_);
  nor (_39424_, _38975_, _38169_);
  not (_39425_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  nor (_39426_, _38974_, _39425_);
  or (_39427_, _39426_, _39424_);
  and (_39428_, _39427_, _31212_);
  nor (_39429_, _31211_, _39425_);
  or (_39430_, _39429_, rst);
  or (_39431_, _39430_, _39428_);
  or (_40343_, _39431_, _39423_);
  and (_39432_, _38967_, _36133_);
  nand (_39433_, _39432_, _31757_);
  or (_39434_, _39432_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_39435_, _39434_, _31899_);
  and (_39436_, _39435_, _39433_);
  nor (_39437_, _38975_, _38162_);
  and (_39438_, _38975_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or (_39439_, _39438_, _39437_);
  and (_39440_, _39439_, _31212_);
  and (_39441_, _38947_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or (_39442_, _39441_, rst);
  or (_39443_, _39442_, _39440_);
  or (_40345_, _39443_, _39436_);
  and (_39444_, _38967_, _36785_);
  nand (_39445_, _39444_, _31757_);
  or (_39446_, _39444_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_39447_, _39446_, _31899_);
  and (_39448_, _39447_, _39445_);
  nor (_39449_, _38975_, _38155_);
  and (_39450_, _38975_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or (_39451_, _39450_, _39449_);
  and (_39452_, _39451_, _31212_);
  and (_39453_, _38947_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or (_39454_, _39453_, rst);
  or (_39455_, _39454_, _39452_);
  or (_40347_, _39455_, _39448_);
  and (_39456_, _38983_, _38813_);
  nand (_39461_, _39456_, _31757_);
  or (_39467_, _39456_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and (_39468_, _39467_, _31899_);
  and (_39469_, _39468_, _39461_);
  nor (_39470_, _38991_, _38203_);
  not (_39471_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  nor (_39472_, _38990_, _39471_);
  or (_39473_, _39472_, _39470_);
  and (_39474_, _39473_, _31212_);
  nor (_39475_, _31211_, _39471_);
  or (_39476_, _39475_, rst);
  or (_39477_, _39476_, _39474_);
  or (_40349_, _39477_, _39469_);
  and (_39478_, _38983_, _33129_);
  nand (_39479_, _39478_, _31757_);
  or (_39480_, _39478_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_39481_, _39480_, _31899_);
  and (_39482_, _39481_, _39479_);
  nor (_39483_, _38991_, _38191_);
  and (_39484_, _38991_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or (_39485_, _39484_, _39483_);
  and (_39486_, _39485_, _31212_);
  and (_39487_, _38947_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or (_39488_, _39487_, rst);
  or (_39489_, _39488_, _39486_);
  or (_40351_, _39489_, _39482_);
  and (_39490_, _38983_, _33847_);
  nand (_39491_, _39490_, _31757_);
  or (_39492_, _39490_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_39493_, _39492_, _31899_);
  and (_39494_, _39493_, _39491_);
  nor (_39495_, _38991_, _38184_);
  and (_39496_, _38991_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or (_39497_, _39496_, _39495_);
  and (_39498_, _39497_, _31212_);
  and (_39499_, _38947_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or (_39500_, _39499_, rst);
  or (_39501_, _39500_, _39498_);
  or (_40353_, _39501_, _39494_);
  and (_39502_, _38983_, _34576_);
  nand (_39503_, _39502_, _31757_);
  or (_39504_, _39502_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_39505_, _39504_, _31899_);
  and (_39506_, _39505_, _39503_);
  nor (_39507_, _38991_, _38177_);
  and (_39508_, _38991_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_39509_, _39508_, _39507_);
  and (_39510_, _39509_, _31212_);
  and (_39511_, _38947_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_39512_, _39511_, rst);
  or (_39513_, _39512_, _39510_);
  or (_40355_, _39513_, _39506_);
  and (_39514_, _38983_, _35338_);
  nand (_39515_, _39514_, _31757_);
  or (_39516_, _39514_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_39517_, _39516_, _31899_);
  and (_39518_, _39517_, _39515_);
  nor (_39519_, _38991_, _38169_);
  not (_39520_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  nor (_39521_, _38990_, _39520_);
  or (_39522_, _39521_, _39519_);
  and (_39523_, _39522_, _31212_);
  nor (_39524_, _31211_, _39520_);
  or (_39525_, _39524_, rst);
  or (_39526_, _39525_, _39523_);
  or (_40356_, _39526_, _39518_);
  and (_39527_, _38983_, _36133_);
  nand (_39528_, _39527_, _31757_);
  or (_39529_, _39527_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_39530_, _39529_, _31899_);
  and (_39531_, _39530_, _39528_);
  nor (_39532_, _38991_, _38162_);
  and (_39533_, _38991_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or (_39534_, _39533_, _39532_);
  and (_39535_, _39534_, _31212_);
  and (_39536_, _38947_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or (_39537_, _39536_, rst);
  or (_39538_, _39537_, _39535_);
  or (_40358_, _39538_, _39531_);
  and (_39539_, _38983_, _36785_);
  nand (_39540_, _39539_, _31757_);
  or (_39541_, _39539_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and (_39542_, _39541_, _31899_);
  and (_39543_, _39542_, _39540_);
  nor (_39544_, _38991_, _38155_);
  and (_39545_, _38991_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or (_39546_, _39545_, _39544_);
  and (_39547_, _39546_, _31212_);
  and (_39548_, _38947_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or (_39549_, _39548_, rst);
  or (_39550_, _39549_, _39547_);
  or (_40360_, _39550_, _39543_);
  and (_40810_, t0_i, _42618_);
  and (_40813_, t1_i, _42618_);
  not (_39551_, _31212_);
  nor (_39552_, _39551_, _27948_);
  and (_39553_, _39552_, _34576_);
  and (_39554_, _39553_, _38140_);
  nand (_39565_, _39554_, _38225_);
  nor (_39576_, _28069_, _27948_);
  and (_39587_, _39576_, _38141_);
  and (_39598_, _39587_, _31212_);
  not (_39609_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and (_39616_, _39609_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  not (_39617_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_39618_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _39617_);
  nor (_39619_, _39618_, _39616_);
  or (_39620_, _39619_, _39598_);
  and (_39621_, _39620_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  not (_39622_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  not (_39623_, t1_i);
  and (_39624_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff , _39623_);
  nor (_39625_, _39624_, _39622_);
  not (_39626_, _39625_);
  not (_39627_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and (_39628_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], _39627_);
  nor (_39629_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6], \oc8051_top_1.oc8051_sfr1.pres_ow );
  not (_39630_, _39629_);
  and (_39631_, _39630_, _39628_);
  and (_39632_, _39631_, _39626_);
  not (_39633_, _39632_);
  nand (_39634_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nand (_39635_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  or (_39636_, _39635_, _39634_);
  nor (_39637_, _39636_, _39633_);
  and (_39638_, _39637_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and (_39639_, _39638_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and (_39640_, _39639_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  or (_39641_, _39640_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  not (_39642_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  nor (_39643_, _39636_, _39642_);
  and (_39644_, _39643_, _39632_);
  and (_39645_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and (_39646_, _39645_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and (_39647_, _39646_, _39644_);
  nor (_39648_, _39647_, _39619_);
  and (_39649_, _39648_, _39641_);
  and (_39650_, _39647_, _39616_);
  and (_39651_, _39650_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor (_39652_, _39651_, _39649_);
  nor (_39653_, _39652_, _39598_);
  or (_39654_, _39653_, _39621_);
  or (_39655_, _39554_, _39654_);
  and (_39656_, _39655_, _42618_);
  and (_40816_, _39656_, _39565_);
  and (_39657_, _39552_, _38272_);
  and (_39658_, _39657_, _42618_);
  and (_39659_, _39658_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor (_39660_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  not (_39661_, _39660_);
  and (_39662_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and (_39663_, _39662_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_39664_, _39663_, _39644_);
  and (_39665_, _39664_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and (_39666_, _39665_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and (_39667_, _39666_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and (_39668_, _39667_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and (_39669_, _39668_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor (_39670_, _39669_, _39661_);
  and (_39671_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  not (_39672_, _39618_);
  and (_39673_, _39669_, _39646_);
  nor (_39674_, _39673_, _39672_);
  or (_39675_, _39674_, _39671_);
  or (_39676_, _39646_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and (_39677_, _39676_, _39675_);
  or (_39678_, _39677_, _39670_);
  nor (_39680_, _39668_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor (_39686_, _39680_, _39598_);
  and (_39687_, _39686_, _39678_);
  not (_39688_, _39598_);
  nor (_39689_, _39688_, _38225_);
  or (_39690_, _39689_, _39687_);
  nor (_39691_, _39554_, rst);
  and (_39692_, _39691_, _39690_);
  or (_40819_, _39692_, _39659_);
  and (_39693_, _39633_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  or (_39694_, _39693_, _39673_);
  and (_39695_, _39694_, _39618_);
  or (_39696_, _39693_, _39669_);
  and (_39697_, _39696_, _39660_);
  nand (_39698_, _39632_, _39609_);
  and (_39699_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  and (_39700_, _39699_, _39698_);
  or (_39701_, _39700_, _39650_);
  or (_39702_, _39701_, _39697_);
  nor (_39703_, _39702_, _39695_);
  nor (_39704_, _39703_, _39598_);
  and (_40822_, _39704_, _39691_);
  and (_39705_, _39552_, _35338_);
  and (_39706_, _39705_, _38140_);
  nor (_39707_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  not (_39708_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  not (_39709_, t0_i);
  and (_39710_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , _39709_);
  nor (_39711_, _39710_, _39708_);
  not (_39712_, _39711_);
  not (_39713_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  nor (_39714_, \oc8051_top_1.oc8051_sfr1.pres_ow , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  nor (_39715_, _39714_, _39713_);
  and (_39716_, _39715_, _39712_);
  not (_39717_, _39716_);
  and (_39718_, _39717_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  and (_39719_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_39720_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and (_39721_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and (_39722_, _39721_, _39720_);
  and (_39723_, _39722_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and (_39724_, _39723_, _39716_);
  and (_39725_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_39726_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and (_39727_, _39726_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_39728_, _39727_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_39729_, _39728_, _39725_);
  and (_39730_, _39729_, _39724_);
  and (_39731_, _39730_, _39719_);
  or (_39732_, _39731_, _39718_);
  and (_39733_, _39732_, _39707_);
  and (_39734_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and (_39735_, _39734_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and (_39736_, _39735_, _39723_);
  and (_39737_, _39736_, _39716_);
  or (_39738_, _39737_, _39718_);
  not (_39739_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_39740_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _39739_);
  and (_39741_, _39729_, _39719_);
  or (_39742_, _39741_, _39718_);
  and (_39743_, _39742_, _39740_);
  or (_39744_, _39743_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_39745_, _39744_, _39738_);
  or (_39746_, _39745_, _39733_);
  nand (_39747_, _39746_, _42618_);
  nor (_39748_, _39747_, _39706_);
  and (_39749_, _39552_, _33847_);
  and (_39750_, _39749_, _38140_);
  not (_39751_, _39750_);
  and (_40825_, _39751_, _39748_);
  and (_39752_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and (_39753_, _39752_, _39724_);
  or (_39754_, _39753_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and (_39755_, _39707_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  not (_39756_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_39757_, _39756_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  or (_39758_, _39757_, _39740_);
  and (_39759_, _39735_, _39724_);
  not (_39760_, _39759_);
  and (_39761_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_39762_, _39761_, _39760_);
  or (_39763_, _39762_, _39758_);
  nand (_39767_, _39757_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand (_39775_, _39767_, _39759_);
  and (_39776_, _39775_, _39763_);
  or (_39777_, _39776_, _39755_);
  and (_39778_, _39777_, _39754_);
  or (_39779_, _39778_, _39706_);
  and (_39780_, _39552_, _38371_);
  not (_39781_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and (_39782_, _39706_, _39781_);
  nor (_39783_, _39782_, _39780_);
  and (_39784_, _39783_, _39779_);
  nor (_39785_, _39751_, _38225_);
  or (_39786_, _39785_, _39784_);
  and (_40828_, _39786_, _42618_);
  not (_39787_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and (_39788_, _39716_, _39739_);
  and (_39789_, _39788_, _39736_);
  and (_39790_, _39789_, _39729_);
  and (_39791_, _39790_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nor (_39792_, _39791_, _39787_);
  and (_39793_, _39791_, _39787_);
  or (_39794_, _39793_, _39792_);
  and (_39795_, _39794_, _39758_);
  and (_39796_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], \oc8051_top_1.oc8051_sfr1.pres_ow );
  and (_39797_, _39796_, _39728_);
  and (_39798_, _39797_, _39725_);
  and (_39799_, _39798_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or (_39800_, _39799_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand (_39801_, _39796_, _39741_);
  and (_39802_, _39801_, _39800_);
  and (_39803_, _39802_, _39761_);
  and (_39804_, _39730_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or (_39805_, _39804_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  not (_39806_, _39707_);
  nor (_39807_, _39731_, _39806_);
  and (_39808_, _39807_, _39805_);
  or (_39809_, _39808_, _39803_);
  or (_39810_, _39809_, _39795_);
  or (_39811_, _39810_, _39706_);
  nand (_39812_, _39706_, _38225_);
  and (_39813_, _39812_, _39811_);
  or (_39814_, _39813_, _39750_);
  nand (_39815_, _39750_, _39787_);
  and (_39816_, _39815_, _42618_);
  and (_40831_, _39816_, _39814_);
  not (_39817_, _39796_);
  or (_39818_, _39817_, _39741_);
  or (_39819_, _39796_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 );
  and (_39820_, _39761_, _42618_);
  and (_39821_, _39820_, _39819_);
  nand (_39822_, _39821_, _39818_);
  nor (_39823_, _39822_, _39706_);
  and (_40834_, _39823_, _39751_);
  and (_39824_, _39552_, _38142_);
  or (_39825_, _39824_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and (_39826_, _39825_, _42618_);
  nand (_39827_, _39824_, _38225_);
  and (_40837_, _39827_, _39826_);
  not (_39828_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and (_39829_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  nor (_39830_, _39829_, _39598_);
  and (_39831_, _39830_, _39632_);
  nor (_39832_, _39831_, _39828_);
  and (_39833_, _39831_, _39828_);
  or (_39834_, _39833_, _39832_);
  and (_39835_, _39646_, _39643_);
  and (_39836_, _39835_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  nand (_39837_, _39836_, _39616_);
  nor (_39838_, _39837_, _39598_);
  or (_39839_, _39838_, _39554_);
  or (_39840_, _39839_, _39834_);
  nand (_39841_, _39554_, _38203_);
  and (_39842_, _39841_, _42618_);
  and (_41323_, _39842_, _39840_);
  not (_39847_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nor (_39848_, _39830_, _39847_);
  not (_39849_, _39829_);
  and (_39850_, _39632_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and (_39851_, _39850_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nor (_39852_, _39850_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nor (_39853_, _39852_, _39851_);
  and (_39854_, _39853_, _39849_);
  and (_39855_, _39640_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and (_39856_, _39855_, _39616_);
  and (_39857_, _39856_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nor (_39858_, _39857_, _39854_);
  nor (_39859_, _39858_, _39598_);
  or (_39860_, _39859_, _39554_);
  or (_39861_, _39860_, _39848_);
  nand (_39862_, _39554_, _38191_);
  and (_39863_, _39862_, _42618_);
  and (_41325_, _39863_, _39861_);
  not (_39873_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  nor (_39874_, _39830_, _39873_);
  nor (_39875_, _39851_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  and (_39876_, _39851_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  nor (_39877_, _39876_, _39875_);
  and (_39878_, _39877_, _39849_);
  and (_39879_, _39650_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nor (_39880_, _39879_, _39878_);
  nor (_39881_, _39880_, _39598_);
  or (_39882_, _39881_, _39874_);
  and (_39883_, _39882_, _39691_);
  not (_39884_, _38184_);
  and (_39885_, _39658_, _39884_);
  or (_41327_, _39885_, _39883_);
  not (_39886_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nor (_39887_, _39830_, _39886_);
  or (_39888_, _39876_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nor (_39889_, _39829_, _39637_);
  and (_39890_, _39889_, _39888_);
  and (_39891_, _39650_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nor (_39892_, _39891_, _39890_);
  nor (_39893_, _39892_, _39598_);
  or (_39894_, _39893_, _39887_);
  and (_39895_, _39894_, _39691_);
  not (_39896_, _38177_);
  and (_39897_, _39658_, _39896_);
  or (_41328_, _39897_, _39895_);
  nor (_39898_, _39830_, _39642_);
  and (_39899_, _39856_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nor (_39900_, _39637_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  nor (_39901_, _39900_, _39644_);
  and (_39902_, _39901_, _39849_);
  nor (_39903_, _39902_, _39899_);
  nor (_39904_, _39903_, _39598_);
  or (_39905_, _39904_, _39898_);
  and (_39906_, _39905_, _39691_);
  not (_39907_, _38169_);
  and (_39908_, _39658_, _39907_);
  or (_41330_, _39908_, _39906_);
  and (_39909_, _39620_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and (_39910_, _39856_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  not (_39911_, _39619_);
  and (_39912_, _39644_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  nor (_39913_, _39644_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  nor (_39914_, _39913_, _39912_);
  and (_39915_, _39914_, _39911_);
  nor (_39916_, _39915_, _39910_);
  nor (_39917_, _39916_, _39598_);
  or (_39918_, _39917_, _39909_);
  and (_39919_, _39918_, _39691_);
  not (_39920_, _38162_);
  and (_39921_, _39658_, _39920_);
  or (_41332_, _39921_, _39919_);
  and (_39922_, _39620_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and (_39923_, _39616_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and (_39924_, _39923_, _39632_);
  and (_39925_, _39924_, _39835_);
  or (_39926_, _39912_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nand (_39927_, _39926_, _39911_);
  nor (_39928_, _39927_, _39640_);
  nor (_39929_, _39928_, _39925_);
  nor (_39930_, _39929_, _39598_);
  or (_39931_, _39930_, _39922_);
  and (_39932_, _39931_, _39691_);
  not (_39933_, _38155_);
  and (_39934_, _39658_, _39933_);
  or (_41334_, _39934_, _39932_);
  and (_39935_, _39644_, _39617_);
  nor (_39936_, _39646_, _39609_);
  not (_39937_, _39936_);
  and (_39938_, _39937_, _39935_);
  nand (_39939_, _39938_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  or (_39940_, _39938_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and (_39941_, _39940_, _39939_);
  or (_39942_, _39941_, _39598_);
  nand (_39943_, _39598_, _38203_);
  and (_39944_, _39943_, _39691_);
  and (_39945_, _39944_, _39942_);
  and (_39946_, _39658_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  or (_41336_, _39946_, _39945_);
  nand (_39947_, _39598_, _38191_);
  nor (_39948_, _39647_, _39672_);
  not (_39949_, _39948_);
  not (_39950_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  nor (_39951_, _39935_, _39618_);
  nor (_39952_, _39951_, _39950_);
  and (_39953_, _39952_, _39949_);
  or (_39954_, _39953_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nand (_39955_, _39953_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and (_39956_, _39955_, _39954_);
  or (_39957_, _39956_, _39598_);
  and (_39958_, _39957_, _39691_);
  and (_39959_, _39958_, _39947_);
  and (_39960_, _39658_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  or (_41338_, _39960_, _39959_);
  nand (_39961_, _39598_, _38184_);
  or (_39962_, _39936_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  not (_39963_, _39962_);
  and (_39964_, _39662_, _39644_);
  and (_39965_, _39964_, _39963_);
  or (_39966_, _39965_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nand (_39967_, _39664_, _39617_);
  nand (_39968_, _39937_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  or (_39969_, _39968_, _39967_);
  and (_39970_, _39969_, _39966_);
  or (_39971_, _39970_, _39598_);
  and (_39972_, _39971_, _39691_);
  and (_39973_, _39972_, _39961_);
  and (_39974_, _39658_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  or (_41340_, _39974_, _39973_);
  nand (_39975_, _39598_, _38177_);
  and (_39976_, _39665_, _39646_);
  and (_39977_, _39664_, _39646_);
  or (_39978_, _39977_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nand (_39979_, _39978_, _39618_);
  nor (_39980_, _39979_, _39976_);
  and (_39981_, _39967_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nor (_39982_, _39967_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or (_39983_, _39982_, _39981_);
  and (_39984_, _39983_, _39672_);
  or (_39985_, _39984_, _39980_);
  or (_39986_, _39985_, _39598_);
  and (_39987_, _39986_, _39691_);
  and (_39988_, _39987_, _39975_);
  and (_39989_, _39658_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or (_41342_, _39989_, _39988_);
  nand (_39990_, _39598_, _38169_);
  or (_39991_, _39976_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nand (_39992_, _39991_, _39618_);
  and (_39993_, _39976_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nor (_39994_, _39993_, _39992_);
  and (_39995_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and (_39996_, _39662_, _39643_);
  and (_39997_, _39996_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_39998_, _39997_, _39632_);
  and (_39999_, _39998_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or (_40000_, _39999_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nand (_40001_, _39999_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and (_40002_, _40001_, _40000_);
  and (_40003_, _40002_, _39660_);
  or (_40004_, _40003_, _39995_);
  or (_40005_, _40004_, _39994_);
  or (_40006_, _40005_, _39598_);
  and (_40007_, _40006_, _39691_);
  and (_40008_, _40007_, _39990_);
  and (_40009_, _39658_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  or (_41344_, _40009_, _40008_);
  nand (_40010_, _39598_, _38162_);
  not (_40011_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and (_40012_, _39666_, _39660_);
  and (_40013_, _39993_, _39618_);
  nor (_40014_, _40013_, _40012_);
  nand (_40015_, _40014_, _40011_);
  or (_40016_, _40014_, _40011_);
  and (_40017_, _40016_, _40015_);
  or (_40018_, _40017_, _39598_);
  and (_40019_, _40018_, _39691_);
  and (_40020_, _40019_, _40010_);
  and (_40021_, _39658_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  or (_41345_, _40021_, _40020_);
  nand (_40022_, _39598_, _38155_);
  and (_40023_, _39963_, _39667_);
  or (_40024_, _40023_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nand (_40025_, _40023_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and (_40026_, _40025_, _40024_);
  or (_40027_, _40026_, _39598_);
  and (_40028_, _40027_, _39691_);
  and (_40029_, _40028_, _40022_);
  and (_40030_, _39658_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  or (_41347_, _40030_, _40029_);
  nor (_40031_, _39717_, _39706_);
  or (_40032_, _40031_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and (_40033_, _39716_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and (_40034_, _39757_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand (_40035_, _40034_, _39736_);
  nand (_40036_, _40035_, _40033_);
  or (_40037_, _40036_, _39706_);
  and (_40038_, _40037_, _40032_);
  or (_40039_, _40038_, _39750_);
  nand (_40040_, _39750_, _38203_);
  and (_40041_, _40040_, _42618_);
  and (_41349_, _40041_, _40039_);
  nor (_40042_, _40033_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and (_40043_, _40033_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  nor (_40044_, _40043_, _40042_);
  and (_40045_, _39757_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and (_40046_, _40045_, _39759_);
  nor (_40047_, _40046_, _40044_);
  nor (_40048_, _40047_, _39706_);
  and (_40049_, _39706_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  or (_40050_, _40049_, _40048_);
  and (_40051_, _40050_, _39751_);
  nor (_40052_, _39751_, _38191_);
  or (_40053_, _40052_, _40051_);
  and (_41351_, _40053_, _42618_);
  nand (_40054_, _39780_, _38184_);
  and (_40055_, _39706_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  nor (_40056_, _40043_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  and (_40057_, _40033_, _39720_);
  nor (_40058_, _40057_, _40056_);
  and (_40059_, _39757_, _39759_);
  and (_40060_, _40059_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nor (_40061_, _40060_, _40058_);
  nor (_40062_, _40061_, _39706_);
  or (_40063_, _40062_, _40055_);
  or (_40064_, _40063_, _39780_);
  and (_40065_, _40064_, _42618_);
  and (_41353_, _40065_, _40054_);
  nand (_40066_, _39780_, _38177_);
  and (_40067_, _39706_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  and (_40068_, _39722_, _39716_);
  nor (_40069_, _40057_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  nor (_40070_, _40069_, _40068_);
  and (_40071_, _40059_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  nor (_40072_, _40071_, _40070_);
  nor (_40073_, _40072_, _39706_);
  or (_40074_, _40073_, _40067_);
  or (_40075_, _40074_, _39780_);
  and (_40076_, _40075_, _42618_);
  and (_41355_, _40076_, _40066_);
  nand (_40077_, _39780_, _38169_);
  and (_40078_, _39706_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  nor (_40079_, _40068_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  nor (_40080_, _40079_, _39724_);
  and (_40081_, _40059_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nor (_40082_, _40081_, _40080_);
  nor (_40083_, _40082_, _39706_);
  or (_40084_, _40083_, _40078_);
  or (_40085_, _40084_, _39780_);
  and (_40086_, _40085_, _42618_);
  and (_41357_, _40086_, _40077_);
  and (_40087_, _39724_, _39806_);
  and (_40088_, _40087_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  nor (_40089_, _40087_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  nor (_40090_, _40089_, _40088_);
  and (_40091_, _40059_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nor (_40092_, _40091_, _40090_);
  nor (_40093_, _40092_, _39706_);
  and (_40094_, _39706_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  or (_40095_, _40094_, _40093_);
  and (_40096_, _40095_, _39751_);
  nor (_40097_, _39751_, _38162_);
  or (_40098_, _40097_, _40096_);
  and (_41359_, _40098_, _42618_);
  not (_40099_, _40088_);
  nor (_40100_, _40099_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and (_40101_, _39757_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_40102_, _40101_, _39716_);
  and (_40103_, _40102_, _39736_);
  nor (_40104_, _40103_, _40100_);
  nor (_40105_, _40104_, _39706_);
  or (_40106_, _40099_, _39706_);
  and (_40107_, _40106_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  or (_40108_, _40107_, _40105_);
  and (_40109_, _40108_, _39751_);
  nor (_40110_, _39751_, _38155_);
  or (_40111_, _40110_, _40109_);
  and (_41361_, _40111_, _42618_);
  or (_40112_, _39789_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand (_40113_, _40112_, _39758_);
  and (_40114_, _39789_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nor (_40115_, _40114_, _40113_);
  and (_40116_, _39796_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or (_40117_, _39796_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand (_40118_, _40117_, _39761_);
  nor (_40119_, _40118_, _40116_);
  and (_40120_, _39724_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or (_40121_, _39724_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand (_40122_, _40121_, _39707_);
  nor (_40123_, _40122_, _40120_);
  or (_40124_, _40123_, _40119_);
  or (_40125_, _40124_, _40115_);
  or (_40126_, _40125_, _39706_);
  nand (_40127_, _39706_, _38203_);
  and (_40128_, _40127_, _40126_);
  or (_40129_, _40128_, _39750_);
  or (_40130_, _39751_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and (_40131_, _40130_, _42618_);
  and (_41362_, _40131_, _40129_);
  nand (_40132_, _39706_, _38191_);
  or (_40133_, _40114_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and (_40134_, _39737_, _39726_);
  not (_40135_, _40134_);
  or (_40136_, _40135_, _39757_);
  and (_40137_, _40136_, _39758_);
  and (_40138_, _40137_, _40133_);
  not (_40139_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nor (_40140_, _40116_, _40139_);
  and (_40141_, _40116_, _40139_);
  or (_40142_, _40141_, _40140_);
  and (_40143_, _40142_, _39761_);
  or (_40144_, _40120_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and (_40145_, _40120_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nor (_40146_, _40145_, _39806_);
  and (_40147_, _40146_, _40144_);
  or (_40148_, _40147_, _40143_);
  or (_40149_, _40148_, _40138_);
  or (_40150_, _40149_, _39706_);
  and (_40151_, _40150_, _40132_);
  or (_40152_, _40151_, _39750_);
  nand (_40153_, _39750_, _40139_);
  and (_40154_, _40153_, _42618_);
  and (_41364_, _40154_, _40152_);
  nand (_40155_, _39706_, _38184_);
  and (_40156_, _39726_, _39716_);
  and (_40157_, _40156_, _39723_);
  or (_40158_, _40157_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_40159_, _39727_, _39724_);
  nor (_40160_, _40159_, _39806_);
  and (_40161_, _40160_, _40158_);
  or (_40162_, _40134_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_40163_, _39737_, _39727_);
  not (_40164_, _40163_);
  and (_40165_, _40164_, _39740_);
  and (_40166_, _40165_, _40162_);
  and (_40167_, _39726_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_40168_, _40167_, _39796_);
  or (_40169_, _40168_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_40170_, _39796_, _39727_);
  nand (_40171_, _40170_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_40172_, _40171_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_40173_, _40172_, _40169_);
  or (_40174_, _40173_, _40166_);
  or (_40175_, _40174_, _40161_);
  or (_40176_, _40175_, _39706_);
  and (_40177_, _40176_, _40155_);
  or (_40178_, _40177_, _39750_);
  or (_40179_, _39751_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_40180_, _40179_, _42618_);
  and (_41366_, _40180_, _40178_);
  nand (_40181_, _39706_, _38177_);
  not (_40182_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_40183_, _40163_, _39739_);
  nor (_40184_, _40183_, _40182_);
  and (_40185_, _40183_, _40182_);
  or (_40186_, _40185_, _40184_);
  and (_40187_, _40186_, _39758_);
  or (_40188_, _40170_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  not (_40189_, _39797_);
  and (_40190_, _40189_, _39761_);
  and (_40191_, _40190_, _40188_);
  or (_40192_, _40159_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_40193_, _39728_, _39724_);
  nor (_40194_, _40193_, _39806_);
  and (_40195_, _40194_, _40192_);
  or (_40196_, _40195_, _40191_);
  or (_40197_, _40196_, _40187_);
  or (_40198_, _40197_, _39706_);
  and (_40199_, _40198_, _40181_);
  or (_40200_, _40199_, _39750_);
  nand (_40201_, _39750_, _40182_);
  and (_40202_, _40201_, _42618_);
  and (_41368_, _40202_, _40200_);
  nand (_40203_, _39706_, _38169_);
  or (_40204_, _40193_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_40205_, _40157_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_40206_, _40205_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_40207_, _40206_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nor (_40208_, _40207_, _39806_);
  and (_40209_, _40208_, _40204_);
  and (_40210_, _39737_, _39728_);
  nand (_40211_, _40210_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or (_40212_, _40210_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_40213_, _40212_, _39740_);
  and (_40214_, _40213_, _40211_);
  and (_40215_, _39797_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or (_40216_, _40215_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_40217_, _40216_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_40218_, _39797_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nand (_40219_, _40218_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_40220_, _40219_, _40217_);
  or (_40221_, _40220_, _40214_);
  or (_40222_, _40221_, _40209_);
  or (_40223_, _40222_, _39706_);
  and (_40224_, _40223_, _40203_);
  or (_40225_, _40224_, _39750_);
  or (_40226_, _39751_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_40227_, _40226_, _42618_);
  and (_41370_, _40227_, _40225_);
  nand (_40228_, _39706_, _38162_);
  not (_40229_, _40207_);
  nor (_40230_, _40229_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_40231_, _40229_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  or (_40232_, _40231_, _40230_);
  and (_40233_, _40232_, _39707_);
  nor (_40234_, _40211_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  or (_40235_, _40234_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nand (_40236_, _40234_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_40237_, _40236_, _39758_);
  and (_40238_, _40237_, _40235_);
  not (_40239_, _39798_);
  and (_40240_, _40239_, _39761_);
  or (_40241_, _40218_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_40242_, _40241_, _40240_);
  or (_40243_, _40242_, _40238_);
  or (_40244_, _40243_, _40233_);
  nor (_40245_, _40244_, _39706_);
  nor (_40246_, _40245_, _39780_);
  and (_40247_, _40246_, _40228_);
  and (_40248_, _39750_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  or (_40249_, _40248_, _40247_);
  and (_41372_, _40249_, _42618_);
  or (_40250_, _39790_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nand (_40251_, _40250_, _39758_);
  nor (_40252_, _40251_, _39791_);
  or (_40253_, _39798_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  not (_40254_, _39799_);
  and (_40255_, _40254_, _39761_);
  and (_40256_, _40255_, _40253_);
  or (_40257_, _39730_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nor (_40258_, _39804_, _39806_);
  and (_40259_, _40258_, _40257_);
  or (_40260_, _40259_, _40256_);
  nor (_40261_, _40260_, _40252_);
  nor (_40262_, _40261_, _39706_);
  and (_40263_, _39706_, _39933_);
  or (_40264_, _40263_, _40262_);
  and (_40265_, _40264_, _39751_);
  and (_40266_, _39750_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or (_40267_, _40266_, _40265_);
  and (_41374_, _40267_, _42618_);
  nor (_40268_, _39824_, _39756_);
  and (_40269_, _39824_, _38204_);
  or (_40270_, _40269_, _40268_);
  and (_41376_, _40270_, _42618_);
  or (_40271_, _39824_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_40272_, _40271_, _42618_);
  nand (_40273_, _39824_, _38191_);
  and (_41378_, _40273_, _40272_);
  or (_40274_, _39824_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and (_40275_, _40274_, _42618_);
  nand (_40276_, _39824_, _38184_);
  and (_41379_, _40276_, _40275_);
  or (_40277_, _39824_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  and (_40278_, _40277_, _42618_);
  nand (_40279_, _39824_, _38177_);
  and (_41381_, _40279_, _40278_);
  or (_40280_, _39824_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and (_40281_, _40280_, _42618_);
  nand (_40282_, _39824_, _38169_);
  and (_41383_, _40282_, _40281_);
  or (_40283_, _39824_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_40284_, _40283_, _42618_);
  nand (_40285_, _39824_, _38162_);
  and (_41385_, _40285_, _40284_);
  or (_40286_, _39824_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and (_40287_, _40286_, _42618_);
  nand (_40288_, _39824_, _38155_);
  and (_41387_, _40288_, _40287_);
  not (_40289_, _27542_);
  nor (_40290_, _38794_, _27948_);
  nand (_40291_, _40290_, _40289_);
  nor (_40292_, _40291_, _28244_);
  and (_40293_, _40292_, _38966_);
  and (_40294_, _40293_, _31855_);
  nand (_40295_, _40294_, _31757_);
  and (_40296_, _38136_, _31855_);
  and (_40297_, _40296_, _38989_);
  not (_40298_, _40297_);
  or (_40299_, _40294_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and (_40300_, _40299_, _40298_);
  and (_40301_, _40300_, _40295_);
  nor (_40302_, _40298_, _38225_);
  or (_40303_, _40302_, _40301_);
  and (_42556_, _40303_, _42618_);
  and (_40304_, _39552_, _38813_);
  and (_40305_, _40304_, _38973_);
  not (_40306_, _40305_);
  and (_40307_, _31790_, _27542_);
  and (_40309_, _40307_, _38795_);
  and (_40311_, _40309_, _38966_);
  and (_40313_, _40311_, _31855_);
  or (_40315_, _40313_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_40317_, _40315_, _40306_);
  nand (_40319_, _40313_, _31757_);
  and (_40321_, _40319_, _40317_);
  nor (_40323_, _40306_, _38225_);
  or (_40325_, _40323_, _40321_);
  and (_42559_, _40325_, _42618_);
  and (_40328_, _40304_, _38140_);
  and (_40330_, _40290_, _27542_);
  and (_40332_, _40330_, _31779_);
  and (_40334_, _40332_, _38934_);
  nand (_40336_, _40334_, _27795_);
  and (_40338_, _40336_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or (_40340_, _40338_, _40328_);
  or (_40342_, _27806_, _33837_);
  and (_40344_, _40342_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or (_40346_, _40344_, _38740_);
  and (_40348_, _40346_, _40334_);
  or (_40350_, _40348_, _40340_);
  nand (_40352_, _40328_, _38155_);
  and (_40354_, _40352_, _42618_);
  and (_42561_, _40354_, _40350_);
  not (_40357_, _40328_);
  nor (_40359_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 );
  nor (_40361_, _40359_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff );
  not (_40362_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  not (_40363_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  not (_40364_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_40365_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _40364_);
  and (_40366_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_40367_, _40366_, _40365_);
  nor (_40368_, _40367_, _40363_);
  or (_40369_, _40368_, _40362_);
  and (_40370_, _40364_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  and (_40371_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  nor (_40372_, _40371_, _40370_);
  nor (_40373_, _40372_, _40363_);
  and (_40374_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _40364_);
  and (_40375_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_40376_, _40375_, _40374_);
  nand (_40377_, _40376_, _40373_);
  or (_40378_, _40377_, _40369_);
  and (_40379_, _40378_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or (_40380_, _40379_, _40361_);
  and (_40381_, _38140_, _31855_);
  and (_40382_, _40381_, _40290_);
  or (_40383_, _40382_, _40380_);
  and (_40384_, _40383_, _40357_);
  nand (_40385_, _40382_, _31757_);
  and (_40386_, _40385_, _40384_);
  nor (_40387_, _40357_, _38225_);
  or (_40388_, _40387_, _40386_);
  and (_42564_, _40388_, _42618_);
  and (_40389_, _39587_, _31899_);
  nand (_40390_, _40389_, _31757_);
  not (_40391_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff );
  and (_40392_, _40391_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  nor (_40393_, _40376_, _40363_);
  not (_40394_, _40393_);
  or (_40395_, _40394_, _40373_);
  or (_40396_, _40395_, _40369_);
  and (_40397_, _40396_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or (_40398_, _40397_, _40392_);
  or (_40399_, _40398_, _40389_);
  and (_40400_, _40399_, _40357_);
  and (_40401_, _40400_, _40390_);
  nor (_40402_, _40357_, _38162_);
  or (_40403_, _40402_, _40401_);
  and (_42566_, _40403_, _42618_);
  not (_40404_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  or (_40405_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff , _40404_);
  nand (_40406_, _40368_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  or (_40407_, _40393_, _40373_);
  or (_40408_, _40407_, _40406_);
  and (_40409_, _40408_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or (_40410_, _40409_, _40405_);
  and (_40411_, _40290_, _38142_);
  or (_40412_, _40411_, _40410_);
  and (_40413_, _40412_, _40357_);
  nand (_40414_, _40411_, _31757_);
  and (_40415_, _40414_, _40413_);
  nor (_40416_, _40357_, _38191_);
  or (_40417_, _40416_, _40415_);
  and (_42568_, _40417_, _42618_);
  and (_40418_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or (_40419_, _40406_, _40395_);
  and (_40420_, _40419_, _40418_);
  and (_40421_, _40290_, _38272_);
  or (_40422_, _40421_, _40420_);
  and (_40423_, _40422_, _40357_);
  nand (_40424_, _40421_, _31757_);
  and (_40425_, _40424_, _40423_);
  nor (_40426_, _40357_, _38177_);
  or (_40427_, _40426_, _40425_);
  and (_42570_, _40427_, _42618_);
  nand (_40428_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nand (_40429_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _40364_);
  and (_40430_, _40429_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_40431_, _40430_, _40428_);
  or (_40432_, _40431_, _40363_);
  and (_40433_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_40434_, _40433_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  not (_40435_, _40434_);
  and (_40436_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_40437_, _40436_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  not (_40438_, _40437_);
  and (_40439_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_40440_, _40439_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_40441_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and (_40442_, _40441_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  nor (_40443_, _40442_, _40440_);
  and (_40444_, _40443_, _40438_);
  and (_40445_, _40444_, _40435_);
  not (_40446_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  nor (_40447_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  nor (_40448_, _40447_, _40446_);
  nand (_40449_, _40448_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  not (_40450_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  nor (_40451_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  nor (_40452_, _40451_, _40450_);
  and (_40453_, _40452_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  not (_40454_, _40453_);
  and (_40455_, _40454_, _40449_);
  nand (_40456_, _40455_, _40445_);
  and (_40457_, _40456_, _40432_);
  and (_40458_, \oc8051_top_1.oc8051_memory_interface1.reti , \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  nor (_40459_, _40458_, _40364_);
  and (_40460_, _40459_, _40457_);
  not (_40461_, _40460_);
  not (_40462_, _40459_);
  and (_40463_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _40363_);
  not (_40464_, _40463_);
  not (_40465_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_40466_, _40448_, _40465_);
  not (_40467_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_40468_, _40452_, _40467_);
  nor (_40469_, _40468_, _40466_);
  not (_40470_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_40471_, _40433_, _40470_);
  not (_40472_, _40471_);
  and (_40473_, _40472_, _40469_);
  nor (_40474_, _40473_, _40464_);
  not (_40475_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_40476_, _40436_, _40475_);
  not (_40477_, _40476_);
  not (_40478_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_40479_, _40439_, _40478_);
  not (_40480_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and (_40481_, _40441_, _40480_);
  nor (_40482_, _40481_, _40479_);
  and (_40483_, _40482_, _40477_);
  nor (_40484_, _40483_, _40464_);
  nor (_40485_, _40484_, _40474_);
  or (_40486_, _40485_, _40462_);
  and (_40487_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [1], _42618_);
  and (_40488_, _40487_, _40486_);
  and (_42605_, _40488_, _40461_);
  nor (_40489_, _40458_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  not (_40490_, _40489_);
  not (_40491_, _40457_);
  and (_40492_, _40485_, _40491_);
  nor (_40493_, _40492_, _40490_);
  nand (_40494_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [1], _42618_);
  nor (_42607_, _40494_, _40493_);
  and (_40495_, _40455_, _40435_);
  nand (_40496_, _40495_, _40457_);
  or (_40497_, _40474_, _40457_);
  and (_40498_, _40497_, _40459_);
  and (_40499_, _40498_, _40496_);
  or (_40500_, _40499_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  nor (_40501_, _40462_, _40457_);
  nand (_40502_, _40501_, _40484_);
  or (_40503_, _40461_, _40444_);
  and (_40504_, _40503_, _42618_);
  and (_40505_, _40504_, _40502_);
  and (_42609_, _40505_, _40500_);
  and (_40506_, _40496_, _40489_);
  or (_40507_, _40506_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  and (_40508_, _40489_, _40457_);
  not (_40509_, _40508_);
  or (_40510_, _40509_, _40444_);
  or (_40511_, _40474_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  nand (_40512_, _40489_, _40484_);
  and (_40513_, _40512_, _40511_);
  or (_40514_, _40513_, _40457_);
  and (_40515_, _40514_, _42618_);
  and (_40516_, _40515_, _40510_);
  and (_42611_, _40516_, _40507_);
  nand (_40517_, _40492_, _40363_);
  nor (_40518_, _40364_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  nand (_40519_, _40518_, _40458_);
  and (_40520_, _40519_, _42618_);
  and (_42613_, _40520_, _40517_);
  and (_40521_, _40492_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  and (_40522_, _40364_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  nor (_40523_, _40522_, _40518_);
  nor (_40524_, _40523_, _40491_);
  or (_40525_, _40524_, _40458_);
  or (_40526_, _40525_, _40521_);
  not (_40527_, _40458_);
  or (_40528_, _40523_, _40527_);
  and (_40529_, _40528_, _42618_);
  and (_42615_, _40529_, _40526_);
  and (_40530_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _42618_);
  and (_42616_, _40530_, _40458_);
  nor (_42621_, _40359_, rst);
  and (_42623_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _42618_);
  nor (_40531_, _40492_, _40458_);
  and (_40532_, _40458_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  or (_40533_, _40532_, _40531_);
  and (_00130_, _40533_, _42618_);
  and (_40534_, _40458_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  or (_40535_, _40534_, _40531_);
  and (_00132_, _40535_, _42618_);
  and (_40536_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _42618_);
  and (_00134_, _40536_, _40458_);
  not (_40537_, _40481_);
  nor (_40538_, _40468_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nor (_40539_, _40538_, _40466_);
  or (_40540_, _40539_, _40471_);
  and (_40541_, _40540_, _40537_);
  or (_40542_, _40541_, _40479_);
  nor (_40543_, _40485_, _40457_);
  and (_40544_, _40543_, _40477_);
  and (_40545_, _40544_, _40542_);
  not (_40546_, _40442_);
  or (_40547_, _40453_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_40548_, _40547_, _40449_);
  or (_40549_, _40548_, _40434_);
  and (_40550_, _40549_, _40546_);
  or (_40551_, _40550_, _40440_);
  and (_40552_, _40457_, _40438_);
  and (_40553_, _40552_, _40551_);
  or (_40554_, _40553_, _40458_);
  or (_40555_, _40554_, _40545_);
  or (_40556_, _40527_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_40557_, _40556_, _42618_);
  and (_00136_, _40557_, _40555_);
  not (_40558_, _40440_);
  or (_40559_, _40442_, _40434_);
  and (_40560_, _40455_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or (_40561_, _40560_, _40559_);
  and (_40562_, _40561_, _40558_);
  and (_40563_, _40562_, _40552_);
  nor (_40564_, _40479_, _40476_);
  or (_40565_, _40481_, _40471_);
  and (_40566_, _40469_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or (_40567_, _40566_, _40565_);
  and (_40568_, _40567_, _40564_);
  and (_40569_, _40568_, _40543_);
  or (_40570_, _40569_, _40458_);
  or (_40571_, _40570_, _40563_);
  or (_40578_, _40527_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and (_40579_, _40578_, _42618_);
  and (_00138_, _40579_, _40571_);
  or (_40590_, _40471_, _40464_);
  nor (_40596_, _40590_, _40469_);
  nand (_40599_, _40596_, _40483_);
  nor (_40600_, _40599_, _40457_);
  not (_40601_, _40455_);
  and (_40602_, _40601_, _40445_);
  and (_40603_, _40602_, _40432_);
  or (_40604_, _40603_, _40458_);
  or (_40605_, _40604_, _40600_);
  or (_40606_, _40527_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  and (_40607_, _40606_, _42618_);
  and (_00139_, _40607_, _40605_);
  and (_40608_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _42618_);
  and (_00141_, _40608_, _40458_);
  and (_40609_, _40458_, _40364_);
  or (_40610_, _40609_, _40493_);
  or (_40611_, _40610_, _40501_);
  and (_00143_, _40611_, _42618_);
  not (_40617_, _40531_);
  and (_40621_, _40617_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  not (_40622_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  and (_40624_, _40453_, _40364_);
  or (_40625_, _40624_, _40622_);
  nor (_40631_, _40449_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_40634_, _40631_, _40434_);
  nand (_40635_, _40634_, _40625_);
  or (_40636_, _40435_, _40366_);
  and (_40639_, _40636_, _40635_);
  or (_40645_, _40639_, _40442_);
  or (_40647_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _40364_);
  or (_40648_, _40647_, _40546_);
  and (_40650_, _40648_, _40558_);
  and (_40656_, _40650_, _40645_);
  and (_40659_, _40440_, _40366_);
  or (_40660_, _40659_, _40437_);
  or (_40661_, _40660_, _40656_);
  or (_40664_, _40647_, _40438_);
  and (_40670_, _40664_, _40457_);
  and (_40672_, _40670_, _40661_);
  and (_40675_, _40468_, _40364_);
  or (_40676_, _40675_, _40622_);
  and (_40682_, _40466_, _40364_);
  nor (_40684_, _40682_, _40471_);
  nand (_40686_, _40684_, _40676_);
  or (_40687_, _40472_, _40366_);
  and (_40693_, _40687_, _40686_);
  or (_40696_, _40693_, _40481_);
  not (_40697_, _40479_);
  or (_40699_, _40647_, _40537_);
  and (_40705_, _40699_, _40697_);
  and (_40708_, _40705_, _40696_);
  and (_40709_, _40479_, _40366_);
  or (_40710_, _40709_, _40476_);
  or (_40713_, _40710_, _40708_);
  and (_40719_, _40647_, _40543_);
  or (_40721_, _40719_, _40544_);
  and (_40722_, _40721_, _40713_);
  or (_40725_, _40722_, _40672_);
  and (_40731_, _40725_, _40527_);
  or (_40733_, _40731_, _40621_);
  and (_00145_, _40733_, _42618_);
  and (_40735_, _40617_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  or (_40741_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _40364_);
  and (_40744_, _40741_, _40438_);
  or (_40745_, _40744_, _40444_);
  or (_40747_, _40624_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_40753_, _40747_, _40634_);
  nand (_40756_, _40434_, _40375_);
  nand (_40757_, _40756_, _40443_);
  or (_40758_, _40757_, _40753_);
  and (_40763_, _40758_, _40745_);
  and (_40768_, _40437_, _40375_);
  or (_40769_, _40768_, _40763_);
  and (_40770_, _40769_, _40457_);
  and (_40775_, _40482_, _40471_);
  or (_40780_, _40775_, _40476_);
  and (_40781_, _40780_, _40375_);
  or (_40782_, _40675_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_40786_, _40684_, _40482_);
  and (_40792_, _40786_, _40782_);
  not (_40793_, _40482_);
  and (_40794_, _40741_, _40793_);
  or (_40798_, _40794_, _40792_);
  and (_40803_, _40798_, _40477_);
  or (_40804_, _40803_, _40781_);
  and (_40805_, _40804_, _40543_);
  or (_40806_, _40805_, _40770_);
  and (_40807_, _40806_, _40527_);
  or (_40808_, _40807_, _40735_);
  and (_00147_, _40808_, _42618_);
  and (_40809_, _40617_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  not (_40811_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  and (_40812_, _40453_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_40814_, _40812_, _40811_);
  nor (_40815_, _40449_, _40364_);
  nor (_40817_, _40815_, _40434_);
  nand (_40818_, _40817_, _40814_);
  or (_40820_, _40435_, _40365_);
  and (_40821_, _40820_, _40818_);
  or (_40823_, _40821_, _40442_);
  or (_40824_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_40826_, _40824_, _40546_);
  and (_40827_, _40826_, _40558_);
  and (_40829_, _40827_, _40823_);
  and (_40830_, _40440_, _40365_);
  or (_40832_, _40830_, _40437_);
  or (_40833_, _40832_, _40829_);
  or (_40835_, _40824_, _40438_);
  and (_40836_, _40835_, _40457_);
  and (_40838_, _40836_, _40833_);
  and (_40839_, _40468_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_40840_, _40839_, _40811_);
  and (_40841_, _40466_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_40842_, _40841_, _40471_);
  nand (_40843_, _40842_, _40840_);
  or (_40844_, _40472_, _40365_);
  and (_40845_, _40844_, _40843_);
  or (_40846_, _40845_, _40481_);
  or (_40847_, _40824_, _40537_);
  and (_40848_, _40847_, _40697_);
  and (_40849_, _40848_, _40846_);
  and (_40850_, _40479_, _40365_);
  or (_40851_, _40850_, _40476_);
  or (_40852_, _40851_, _40849_);
  and (_40853_, _40824_, _40543_);
  or (_40854_, _40853_, _40544_);
  and (_40855_, _40854_, _40852_);
  or (_40856_, _40855_, _40838_);
  and (_40857_, _40856_, _40527_);
  or (_40858_, _40857_, _40809_);
  and (_00149_, _40858_, _42618_);
  and (_40859_, _40617_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  or (_40860_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_40861_, _40860_, _40438_);
  or (_40862_, _40861_, _40444_);
  or (_40863_, _40812_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_40864_, _40863_, _40817_);
  nand (_40865_, _40434_, _40374_);
  nand (_40866_, _40865_, _40443_);
  or (_40867_, _40866_, _40864_);
  and (_40868_, _40867_, _40862_);
  and (_40869_, _40437_, _40374_);
  or (_40870_, _40869_, _40868_);
  and (_40871_, _40870_, _40457_);
  and (_40872_, _40780_, _40374_);
  or (_40873_, _40839_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_40874_, _40842_, _40482_);
  and (_40875_, _40874_, _40873_);
  and (_40876_, _40860_, _40793_);
  or (_40877_, _40876_, _40875_);
  and (_40878_, _40877_, _40477_);
  or (_40879_, _40878_, _40872_);
  and (_40880_, _40879_, _40543_);
  or (_40881_, _40880_, _40871_);
  and (_40882_, _40881_, _40527_);
  or (_40883_, _40882_, _40859_);
  and (_00150_, _40883_, _42618_);
  or (_40884_, _40490_, _40485_);
  and (_40885_, _40884_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0]);
  or (_40886_, _40885_, _40508_);
  and (_00152_, _40886_, _42618_);
  and (_40887_, _40486_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0]);
  or (_40888_, _40887_, _40460_);
  and (_00154_, _40888_, _42618_);
  and (_40889_, _40334_, _38813_);
  or (_40890_, _40889_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and (_40891_, _40890_, _40357_);
  nand (_40892_, _40889_, _31757_);
  and (_40893_, _40892_, _40891_);
  nor (_40894_, _40357_, _38203_);
  or (_40895_, _40894_, _40893_);
  and (_00156_, _40895_, _42618_);
  not (_40896_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  nand (_40897_, _40334_, _33847_);
  nand (_40898_, _40897_, _40896_);
  and (_40899_, _40898_, _40357_);
  or (_40900_, _40897_, _32410_);
  and (_40901_, _40900_, _40899_);
  nor (_40902_, _40357_, _38184_);
  or (_40903_, _40902_, _40901_);
  and (_00158_, _40903_, _42618_);
  nand (_40904_, _40334_, _35338_);
  nor (_40905_, _40904_, _31757_);
  and (_40906_, _40904_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  or (_40907_, _40906_, _40328_);
  or (_40908_, _40907_, _40905_);
  nand (_40909_, _40328_, _38169_);
  and (_40910_, _40909_, _42618_);
  and (_00160_, _40910_, _40908_);
  and (_40911_, _40311_, _38813_);
  or (_40912_, _40911_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_40913_, _40912_, _40306_);
  nand (_40914_, _40911_, _31757_);
  and (_40915_, _40914_, _40913_);
  nor (_40916_, _40306_, _38203_);
  or (_40917_, _40916_, _40915_);
  and (_00161_, _40917_, _42618_);
  and (_40918_, _40311_, _33129_);
  or (_40919_, _40918_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_40920_, _40919_, _40306_);
  nand (_40921_, _40918_, _31757_);
  and (_40922_, _40921_, _40920_);
  nor (_40923_, _40306_, _38191_);
  or (_40924_, _40923_, _40922_);
  and (_00163_, _40924_, _42618_);
  nand (_40925_, _40311_, _39025_);
  and (_40926_, _40925_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_40927_, _40926_, _40305_);
  and (_40928_, _33880_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_40929_, _40928_, _33869_);
  and (_40930_, _40929_, _40311_);
  or (_40931_, _40930_, _40927_);
  nand (_40932_, _40305_, _38184_);
  and (_40933_, _40932_, _42618_);
  and (_00165_, _40933_, _40931_);
  and (_40934_, _40311_, _34576_);
  or (_40935_, _40934_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_40936_, _40935_, _40306_);
  nand (_40937_, _40934_, _31757_);
  and (_40938_, _40937_, _40936_);
  nor (_40939_, _40306_, _38177_);
  or (_40940_, _40939_, _40938_);
  and (_00167_, _40940_, _42618_);
  and (_40941_, _40311_, _35338_);
  or (_40942_, _40941_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  and (_40943_, _40942_, _40306_);
  nand (_40944_, _40941_, _31757_);
  and (_40945_, _40944_, _40943_);
  nor (_40946_, _40306_, _38169_);
  or (_40947_, _40946_, _40945_);
  and (_00169_, _40947_, _42618_);
  and (_40948_, _40311_, _36133_);
  or (_40949_, _40948_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and (_40950_, _40949_, _40306_);
  nand (_40951_, _40948_, _31757_);
  and (_40952_, _40951_, _40950_);
  nor (_40953_, _40306_, _38162_);
  or (_40954_, _40953_, _40952_);
  and (_00171_, _40954_, _42618_);
  and (_40955_, _40311_, _36785_);
  or (_40956_, _40955_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_40957_, _40956_, _40306_);
  nand (_40958_, _40955_, _31757_);
  and (_40959_, _40958_, _40957_);
  nor (_40960_, _40306_, _38155_);
  or (_40961_, _40960_, _40959_);
  and (_00173_, _40961_, _42618_);
  and (_40962_, _40293_, _38813_);
  nand (_40963_, _40962_, _31757_);
  or (_40964_, _40962_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_40965_, _40964_, _40298_);
  and (_40966_, _40965_, _40963_);
  nor (_40967_, _40298_, _38203_);
  or (_40968_, _40967_, _40966_);
  and (_00174_, _40968_, _42618_);
  and (_40969_, _40293_, _33129_);
  nand (_40970_, _40969_, _31757_);
  or (_40971_, _40969_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_40972_, _40971_, _40298_);
  and (_40973_, _40972_, _40970_);
  nor (_40974_, _40298_, _38191_);
  or (_40975_, _40974_, _40973_);
  and (_00176_, _40975_, _42618_);
  and (_40976_, _33880_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_40977_, _40976_, _33869_);
  and (_40978_, _40977_, _40293_);
  nand (_40979_, _40293_, _39025_);
  and (_40980_, _40979_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_40981_, _40980_, _40297_);
  or (_40982_, _40981_, _40978_);
  nand (_40983_, _40297_, _38184_);
  and (_40984_, _40983_, _42618_);
  and (_00178_, _40984_, _40982_);
  and (_40985_, _40293_, _34576_);
  nand (_40986_, _40985_, _31757_);
  or (_40987_, _40985_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_40988_, _40987_, _40986_);
  or (_40989_, _40988_, _40297_);
  nand (_40990_, _40297_, _38177_);
  and (_40991_, _40990_, _42618_);
  and (_00180_, _40991_, _40989_);
  and (_40992_, _40293_, _35338_);
  nand (_40993_, _40992_, _31757_);
  or (_40994_, _40992_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_40995_, _40994_, _40298_);
  and (_40996_, _40995_, _40993_);
  nor (_40997_, _40298_, _38169_);
  or (_40998_, _40997_, _40996_);
  and (_00182_, _40998_, _42618_);
  and (_40999_, _40293_, _36133_);
  nand (_41000_, _40999_, _31757_);
  or (_41001_, _40999_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_41002_, _41001_, _41000_);
  or (_41003_, _41002_, _40297_);
  nand (_41004_, _40297_, _38162_);
  and (_41005_, _41004_, _42618_);
  and (_00184_, _41005_, _41003_);
  and (_41006_, _40293_, _36785_);
  nand (_41007_, _41006_, _31757_);
  or (_41008_, _41006_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and (_41009_, _41008_, _41007_);
  or (_41010_, _41009_, _40297_);
  nand (_41011_, _40297_, _38155_);
  and (_41012_, _41011_, _42618_);
  and (_00185_, _41012_, _41010_);
  and (_41013_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  not (_41014_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  nor (_41015_, _40359_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf );
  and (_41016_, _41015_, _41014_);
  not (_41017_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  nor (_41018_, _41017_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  or (_41019_, _41018_, _41016_);
  nor (_41020_, _41019_, _41013_);
  or (_41021_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  nand (_41022_, _41021_, _42618_);
  nor (_00545_, _41022_, _41020_);
  nor (_41023_, _41020_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or (_41024_, _41023_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  nand (_41025_, _41023_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  and (_41026_, _41025_, _42618_);
  and (_00548_, _41026_, _41024_);
  not (_41027_, rxd_i);
  and (_41028_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r , _41027_);
  nor (_41029_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  not (_41030_, _41029_);
  and (_41031_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re );
  and (_41032_, _41031_, _41030_);
  and (_41033_, _41032_, _41028_);
  not (_41034_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  and (_41035_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], _41034_);
  and (_41036_, _41035_, _41029_);
  or (_41037_, _41036_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  or (_41038_, _41037_, _41033_);
  and (_41039_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _42618_);
  and (_00551_, _41039_, _41038_);
  and (_41040_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  and (_41041_, _41040_, _41030_);
  not (_41042_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  nor (_41043_, _41029_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and (_41044_, _41043_, _41042_);
  nor (_41045_, _41044_, _41041_);
  not (_41046_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  nor (_41047_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _41046_);
  not (_41048_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  nor (_41049_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], _41048_);
  and (_41050_, _41049_, _41047_);
  not (_41051_, _41050_);
  or (_41052_, _41051_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  and (_41053_, _41050_, _41041_);
  and (_41054_, _41041_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_41055_, _41054_, _41053_);
  and (_41056_, _41055_, _41052_);
  or (_41057_, _41056_, _41045_);
  not (_41058_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  nand (_41059_, _41029_, \oc8051_top_1.oc8051_sfr1.pres_ow );
  nor (_41060_, _41059_, _41058_);
  not (_41061_, _41060_);
  or (_41062_, _41061_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  nand (_41063_, _41062_, _41057_);
  nand (_00554_, _41063_, _41039_);
  not (_41064_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r );
  not (_41065_, _41041_);
  nor (_41066_, _41042_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re );
  not (_41067_, _41066_);
  not (_41068_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor (_41069_, _41029_, _41068_);
  and (_41070_, _41069_, _41067_);
  and (_41071_, _41070_, _41065_);
  nor (_41072_, _41071_, _41064_);
  and (_41073_, _41071_, rxd_i);
  or (_41074_, _41073_, rst);
  or (_00556_, _41074_, _41072_);
  nor (_41075_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and (_41076_, _41075_, _41047_);
  and (_41077_, _41076_, _41054_);
  nand (_41078_, _41077_, _41027_);
  or (_41079_, _41077_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  and (_41080_, _41079_, _42618_);
  and (_00559_, _41080_, _41078_);
  and (_41081_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and (_41082_, _41081_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and (_41083_, _41082_, _41046_);
  and (_41084_, _41083_, _41054_);
  and (_41085_, _41032_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor (_41086_, _41085_, _41054_);
  nor (_41087_, _41082_, _41065_);
  or (_41088_, _41087_, _41086_);
  and (_41089_, _41088_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  or (_41090_, _41089_, _41084_);
  and (_00562_, _41090_, _42618_);
  and (_41091_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], _42618_);
  nand (_41092_, _41091_, _41068_);
  nand (_41093_, _41039_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  nand (_00564_, _41093_, _41092_);
  and (_41094_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _41068_);
  not (_41095_, _41032_);
  nand (_41096_, _41036_, _41058_);
  and (_41097_, _41096_, _41095_);
  and (_41098_, _41097_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  or (_41099_, _41098_, _41041_);
  or (_41100_, _41050_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  nor (_41101_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  nand (_41102_, _41101_, _41053_);
  and (_41103_, _41102_, _41100_);
  and (_41104_, _41103_, _41099_);
  or (_41105_, _41104_, _41060_);
  nand (_41106_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  nand (_41107_, _41106_, _41041_);
  or (_41108_, _41107_, _41051_);
  and (_41109_, _41108_, _41061_);
  or (_41110_, _41109_, rxd_i);
  and (_41111_, _41110_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and (_41112_, _41111_, _41105_);
  or (_41113_, _41112_, _41094_);
  and (_00567_, _41113_, _42618_);
  and (_41114_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  not (_41115_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and (_41116_, _41015_, _41115_);
  or (_41117_, _41116_, _41018_);
  nor (_41118_, _41117_, _41114_);
  or (_41119_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nand (_41120_, _41119_, _42618_);
  nor (_00570_, _41120_, _41118_);
  nor (_41121_, _41118_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or (_41122_, _41121_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nand (_41123_, _41121_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  and (_41124_, _41123_, _42618_);
  and (_00572_, _41124_, _41122_);
  not (_41125_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  nor (_41126_, _31834_, _27948_);
  and (_41127_, _41126_, _33118_);
  and (_41128_, _41127_, _31212_);
  and (_41129_, _41128_, _38957_);
  and (_41130_, _41129_, _42618_);
  nand (_41131_, _41130_, _41125_);
  nor (_41132_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  not (_41133_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  nor (_41134_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  and (_41135_, _41134_, _41133_);
  and (_41136_, _41135_, _41132_);
  not (_41137_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  nor (_41138_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  nor (_41139_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  and (_41140_, _41139_, _41138_);
  and (_41141_, _41140_, _41137_);
  and (_41142_, _41141_, _41136_);
  not (_41143_, _41142_);
  or (_41144_, _41143_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  or (_41145_, _41142_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  not (_41146_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  nor (_41147_, _41059_, _41146_);
  and (_41148_, _41147_, _41145_);
  and (_41149_, _41148_, _41144_);
  nor (_41150_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  nor (_41151_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  and (_41152_, _41151_, _41150_);
  and (_41153_, _41030_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr );
  and (_41154_, _41153_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  and (_41155_, _41154_, _41152_);
  not (_41156_, _41155_);
  or (_41157_, _41156_, _41145_);
  and (_41158_, _41152_, _41153_);
  or (_41159_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd , _41146_);
  nor (_41160_, _41159_, _41158_);
  nor (_41161_, _41160_, _41147_);
  and (_41162_, _41161_, _41157_);
  nor (_41163_, _41162_, _41149_);
  nor (_41164_, _41129_, rst);
  nand (_41165_, _41164_, _41163_);
  and (_00575_, _41165_, _41131_);
  nor (_41166_, _41143_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  nand (_41167_, _41158_, _41166_);
  and (_41168_, _41147_, _41142_);
  or (_41169_, _41146_, rst);
  nor (_41170_, _41169_, _41168_);
  and (_41171_, _41170_, _41167_);
  or (_00578_, _41171_, _41130_);
  or (_41172_, _41156_, _41166_);
  or (_41173_, _41158_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  and (_41174_, _41059_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  and (_41175_, _41174_, _41173_);
  and (_41176_, _41175_, _41172_);
  or (_41177_, _41176_, _41168_);
  and (_00580_, _41177_, _41164_);
  and (_41178_, _41154_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  and (_41179_, _41178_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  and (_41180_, _41179_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  nand (_41181_, _41180_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  or (_41182_, _41180_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  and (_41183_, _41182_, _41181_);
  and (_00583_, _41183_, _41164_);
  nor (_41184_, _41155_, _41147_);
  and (_41185_, _41184_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  and (_41186_, _41185_, _41164_);
  and (_41187_, _41130_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  or (_00586_, _41187_, _41186_);
  and (_41188_, _40296_, _38140_);
  or (_41189_, _41188_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  and (_41190_, _41189_, _42618_);
  nand (_41191_, _41188_, _38225_);
  and (_00588_, _41191_, _41190_);
  and (_41192_, _40292_, _38934_);
  and (_41193_, _41192_, _31855_);
  nand (_41194_, _41193_, _31757_);
  and (_41195_, _40304_, _38957_);
  not (_41196_, _41195_);
  or (_41197_, _41193_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  and (_41198_, _41197_, _41196_);
  and (_41199_, _41198_, _41194_);
  nor (_41200_, _41196_, _38225_);
  or (_41201_, _41200_, _41199_);
  and (_00591_, _41201_, _42618_);
  nor (_41202_, _41060_, _41053_);
  not (_41203_, _41202_);
  nor (_41204_, _41097_, _41041_);
  nor (_41205_, _41204_, _41203_);
  nor (_41206_, _41205_, _41068_);
  or (_41207_, _41206_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  or (_41208_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1], _41068_);
  or (_41209_, _41208_, _41202_);
  and (_41210_, _41209_, _42618_);
  and (_01206_, _41210_, _41207_);
  or (_41211_, _41206_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1]);
  or (_41212_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2], _41068_);
  or (_41213_, _41212_, _41202_);
  and (_41214_, _41213_, _42618_);
  and (_01208_, _41214_, _41211_);
  or (_41215_, _41206_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2]);
  or (_41216_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _41068_);
  or (_41217_, _41216_, _41202_);
  and (_41218_, _41217_, _42618_);
  and (_01210_, _41218_, _41215_);
  or (_41219_, _41206_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  or (_41220_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _41068_);
  or (_41221_, _41220_, _41202_);
  and (_41222_, _41221_, _42618_);
  and (_01212_, _41222_, _41219_);
  or (_41223_, _41206_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  or (_41224_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _41068_);
  or (_41225_, _41224_, _41202_);
  and (_41226_, _41225_, _42618_);
  and (_01214_, _41226_, _41223_);
  or (_41227_, _41206_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  or (_41228_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _41068_);
  or (_41229_, _41228_, _41202_);
  and (_41230_, _41229_, _42618_);
  and (_01216_, _41230_, _41227_);
  or (_41231_, _41206_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  or (_41232_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _41068_);
  or (_41233_, _41232_, _41202_);
  and (_41234_, _41233_, _42618_);
  and (_01218_, _41234_, _41231_);
  or (_41235_, _41206_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  or (_41236_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8], _41068_);
  or (_41237_, _41236_, _41202_);
  and (_41238_, _41237_, _42618_);
  and (_01220_, _41238_, _41235_);
  nor (_41239_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , rst);
  and (_41240_, _41239_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  or (_41241_, _41051_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  or (_41242_, _41050_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  and (_41243_, _41242_, _41041_);
  and (_41244_, _41243_, _41241_);
  or (_41245_, _41032_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  and (_41246_, _41245_, _41096_);
  and (_41247_, _41246_, _41065_);
  or (_41248_, _41247_, _41244_);
  or (_41249_, _41248_, _41060_);
  or (_41250_, _41061_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  and (_41251_, _41250_, _41039_);
  and (_41252_, _41251_, _41249_);
  or (_01221_, _41252_, _41240_);
  and (_41253_, _41050_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  and (_41254_, _41253_, _41097_);
  or (_41255_, _41254_, _41205_);
  and (_41256_, _41255_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  and (_41257_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9], _41068_);
  nand (_41258_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor (_41259_, _41258_, _41202_);
  or (_41260_, _41259_, _41257_);
  or (_41261_, _41260_, _41256_);
  and (_01223_, _41261_, _42618_);
  not (_41262_, _41206_);
  and (_41263_, _41262_, _41091_);
  or (_41264_, _41254_, _41203_);
  and (_41265_, _41039_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  and (_41266_, _41265_, _41264_);
  or (_01225_, _41266_, _41263_);
  or (_41267_, _41084_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0]);
  nand (_41268_, _41084_, _41027_);
  and (_41269_, _41268_, _42618_);
  and (_01227_, _41269_, _41267_);
  or (_41270_, _41086_, _41048_);
  or (_41271_, _41054_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and (_41272_, _41271_, _42618_);
  and (_01229_, _41272_, _41270_);
  and (_41273_, _41086_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  nor (_41274_, _41075_, _41081_);
  and (_41275_, _41274_, _41054_);
  or (_41276_, _41275_, _41273_);
  and (_01231_, _41276_, _42618_);
  and (_41277_, _41088_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and (_41278_, _41081_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and (_41279_, _41278_, _41087_);
  or (_41280_, _41279_, _41277_);
  and (_01233_, _41280_, _42618_);
  and (_41281_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _41068_);
  and (_41282_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_41283_, _41282_, _41281_);
  and (_01235_, _41283_, _42618_);
  and (_41284_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _41068_);
  and (_41285_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_41286_, _41285_, _41284_);
  and (_01237_, _41286_, _42618_);
  and (_41287_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _41068_);
  and (_41288_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_41289_, _41288_, _41287_);
  and (_01239_, _41289_, _42618_);
  and (_41290_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _41068_);
  and (_41291_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_41292_, _41291_, _41290_);
  and (_01241_, _41292_, _42618_);
  and (_41293_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _41068_);
  and (_41294_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_41295_, _41294_, _41293_);
  and (_01243_, _41295_, _42618_);
  and (_41296_, _41039_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  or (_01245_, _41296_, _41240_);
  and (_41297_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_41298_, _41297_, _41257_);
  and (_01247_, _41298_, _42618_);
  nor (_41299_, _41154_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  nor (_41300_, _41299_, _41178_);
  and (_01249_, _41300_, _41164_);
  nor (_41301_, _41178_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  nor (_41302_, _41301_, _41179_);
  and (_01251_, _41302_, _41164_);
  nor (_41303_, _41179_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  nor (_41304_, _41303_, _41180_);
  and (_01253_, _41304_, _41164_);
  and (_41305_, _41142_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  or (_41306_, _41305_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  and (_41307_, _41306_, _41147_);
  or (_41308_, _41155_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  or (_41309_, _41184_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  and (_41310_, _41309_, _41308_);
  nor (_41311_, _41310_, _41307_);
  nor (_41312_, _41311_, _41129_);
  nor (_41313_, _41030_, _38203_);
  and (_41314_, _41313_, _41129_);
  or (_41315_, _41314_, _41312_);
  and (_01255_, _41315_, _42618_);
  not (_41316_, _41184_);
  and (_41317_, _41316_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  and (_41318_, _41184_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  or (_41319_, _41318_, _41317_);
  and (_41320_, _41319_, _41164_);
  nand (_41321_, _41029_, _38191_);
  nand (_41322_, _41030_, _38203_);
  and (_41324_, _41322_, _41130_);
  and (_41326_, _41324_, _41321_);
  or (_01256_, _41326_, _41320_);
  nor (_41329_, _41184_, _41137_);
  and (_41331_, _41184_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  or (_41333_, _41331_, _41329_);
  and (_41335_, _41333_, _41164_);
  nand (_41337_, _41029_, _38184_);
  nand (_41339_, _41030_, _38191_);
  and (_41341_, _41339_, _41130_);
  and (_41343_, _41341_, _41337_);
  or (_01258_, _41343_, _41335_);
  nand (_41346_, _41184_, _41137_);
  or (_41348_, _41184_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  and (_41350_, _41348_, _41346_);
  and (_41352_, _41350_, _41164_);
  nand (_41354_, _41030_, _38184_);
  nand (_41356_, _41029_, _38177_);
  and (_41358_, _41356_, _41130_);
  and (_41360_, _41358_, _41354_);
  or (_01260_, _41360_, _41352_);
  nand (_41363_, _41184_, _41133_);
  or (_41365_, _41184_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  and (_41367_, _41365_, _41363_);
  and (_41369_, _41367_, _41164_);
  nand (_41371_, _41030_, _38177_);
  nand (_41373_, _41029_, _38169_);
  and (_41375_, _41373_, _41130_);
  and (_41377_, _41375_, _41371_);
  or (_01262_, _41377_, _41369_);
  or (_41380_, _41316_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  or (_41382_, _41184_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  and (_41384_, _41382_, _41380_);
  and (_41386_, _41384_, _41164_);
  nand (_41388_, _41029_, _38162_);
  nand (_41389_, _41030_, _38169_);
  and (_41390_, _41389_, _41130_);
  and (_41391_, _41390_, _41388_);
  or (_01264_, _41391_, _41386_);
  or (_41392_, _41316_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  or (_41393_, _41184_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  and (_41394_, _41393_, _41392_);
  and (_41395_, _41394_, _41164_);
  nand (_41396_, _41029_, _38155_);
  nand (_41397_, _41030_, _38162_);
  and (_41398_, _41397_, _41130_);
  and (_41399_, _41398_, _41396_);
  or (_01266_, _41399_, _41395_);
  or (_41400_, _41316_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  or (_41401_, _41184_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  and (_41402_, _41401_, _41400_);
  and (_41403_, _41402_, _41164_);
  nand (_41404_, _41029_, _38225_);
  nand (_41405_, _41030_, _38155_);
  and (_41406_, _41405_, _41130_);
  and (_41407_, _41406_, _41404_);
  or (_01268_, _41407_, _41403_);
  and (_41408_, _41129_, _41030_);
  nand (_41409_, _41408_, _38225_);
  and (_41410_, _41184_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  and (_41411_, _41316_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  or (_41412_, _41411_, _41410_);
  or (_41413_, _41412_, _41129_);
  and (_41414_, _41413_, _42618_);
  and (_01270_, _41414_, _41409_);
  or (_41415_, _41316_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  or (_41416_, _41184_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  and (_41417_, _41416_, _41415_);
  and (_41418_, _41417_, _41164_);
  or (_41419_, _41017_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  and (_41420_, _41419_, _41030_);
  and (_41421_, _41420_, _41130_);
  or (_01272_, _41421_, _41418_);
  nand (_41422_, _41188_, _38203_);
  or (_41423_, _41188_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  and (_41424_, _41423_, _42618_);
  and (_01274_, _41424_, _41422_);
  or (_41425_, _41188_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  and (_41426_, _41425_, _42618_);
  nand (_41427_, _41188_, _38191_);
  and (_01276_, _41427_, _41426_);
  or (_41428_, _41188_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  and (_41429_, _41428_, _42618_);
  nand (_41430_, _41188_, _38184_);
  and (_01278_, _41430_, _41429_);
  or (_41431_, _41188_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  and (_41432_, _41431_, _42618_);
  nand (_41433_, _41188_, _38177_);
  and (_01280_, _41433_, _41432_);
  or (_41434_, _41188_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  and (_41435_, _41434_, _42618_);
  nand (_41436_, _41188_, _38169_);
  and (_01282_, _41436_, _41435_);
  or (_41437_, _41188_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  and (_41438_, _41437_, _42618_);
  nand (_41439_, _41188_, _38162_);
  and (_01284_, _41439_, _41438_);
  or (_41440_, _41188_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  and (_41441_, _41440_, _42618_);
  nand (_41442_, _41188_, _38155_);
  and (_01286_, _41442_, _41441_);
  not (_41443_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  or (_41444_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _41443_);
  or (_41445_, _41444_, _41029_);
  nor (_41446_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and (_41447_, _41446_, _41445_);
  or (_41448_, _41447_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or (_41449_, _41448_, _41192_);
  or (_41450_, _38813_, _41034_);
  nand (_41451_, _41450_, _41192_);
  or (_41452_, _41451_, _38814_);
  and (_41453_, _41452_, _41449_);
  or (_41454_, _41453_, _41195_);
  nand (_41455_, _41195_, _38203_);
  and (_41456_, _41455_, _42618_);
  and (_01288_, _41456_, _41454_);
  or (_41457_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  or (_41458_, _41457_, _41192_);
  nand (_41459_, _38863_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  nand (_41460_, _41459_, _41192_);
  or (_41461_, _41460_, _38864_);
  and (_41462_, _41461_, _41458_);
  or (_41463_, _41462_, _41195_);
  nand (_41464_, _41195_, _38191_);
  and (_41465_, _41464_, _42618_);
  and (_01290_, _41465_, _41463_);
  not (_41466_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  and (_41467_, _41043_, _41466_);
  and (_41468_, _41467_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  not (_41469_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  nor (_41470_, _41467_, _41469_);
  or (_41471_, _41470_, _41468_);
  or (_41472_, _41471_, _41192_);
  or (_41473_, _33847_, _41469_);
  nand (_41474_, _41473_, _41192_);
  or (_41475_, _41474_, _33869_);
  and (_41476_, _41475_, _41472_);
  or (_41477_, _41476_, _41195_);
  nand (_41478_, _41195_, _38184_);
  and (_41479_, _41478_, _42618_);
  and (_01291_, _41479_, _41477_);
  and (_41480_, _41192_, _34576_);
  nand (_41481_, _41480_, _31757_);
  or (_41482_, _41480_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  and (_41483_, _41482_, _41196_);
  and (_41484_, _41483_, _41481_);
  nor (_41485_, _41196_, _38177_);
  or (_41486_, _41485_, _41484_);
  and (_01293_, _41486_, _42618_);
  and (_41487_, _41192_, _35338_);
  nand (_41488_, _41487_, _31757_);
  or (_41489_, _41487_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and (_41490_, _41489_, _41196_);
  and (_41491_, _41490_, _41488_);
  nor (_41492_, _41196_, _38169_);
  or (_41493_, _41492_, _41491_);
  and (_01295_, _41493_, _42618_);
  and (_41494_, _41192_, _36133_);
  nand (_41495_, _41494_, _31757_);
  or (_41496_, _41494_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  and (_41497_, _41496_, _41196_);
  and (_41498_, _41497_, _41495_);
  nor (_41499_, _41196_, _38162_);
  or (_41500_, _41499_, _41498_);
  and (_01297_, _41500_, _42618_);
  and (_41501_, _41192_, _36785_);
  nand (_41502_, _41501_, _31757_);
  or (_41503_, _41501_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  and (_41504_, _41503_, _41196_);
  and (_41505_, _41504_, _41502_);
  nor (_41506_, _41196_, _38155_);
  or (_41507_, _41506_, _41505_);
  and (_01299_, _41507_, _42618_);
  and (_01626_, t2_i, _42618_);
  nor (_41508_, t2_i, rst);
  and (_01628_, _41508_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r );
  nand (_41509_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r , _42618_);
  nor (_01631_, _41509_, t2ex_i);
  and (_01634_, t2ex_i, _42618_);
  and (_41510_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  nor (_41511_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and (_41512_, _41511_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and (_41513_, _41512_, _41510_);
  not (_41514_, _41513_);
  and (_41515_, _41514_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and (_41516_, _41513_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  nor (_41517_, _41516_, _41515_);
  and (_41518_, _38137_, _28387_);
  and (_41519_, _41518_, _39749_);
  nor (_41520_, _41519_, _41517_);
  and (_41521_, _27795_, _33107_);
  and (_41522_, _41126_, _41521_);
  and (_41523_, _41518_, _41522_);
  and (_41524_, _41523_, _31212_);
  not (_41525_, _41524_);
  nor (_41526_, _41525_, _38225_);
  or (_41527_, _41526_, _41520_);
  and (_41528_, _41518_, _39553_);
  not (_41529_, _41528_);
  and (_41530_, _41529_, _41527_);
  and (_41531_, _41528_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  or (_41532_, _41531_, _41530_);
  and (_01637_, _41532_, _42618_);
  nand (_41533_, _41528_, _38225_);
  nor (_41534_, _41519_, _41514_);
  or (_41535_, _41534_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  not (_41536_, _41534_);
  or (_41537_, _41536_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  and (_41538_, _41537_, _41535_);
  or (_41539_, _41538_, _41528_);
  and (_41540_, _41539_, _42618_);
  and (_01640_, _41540_, _41533_);
  and (_41541_, _41518_, _39705_);
  and (_41542_, _39552_, _36133_);
  and (_41543_, _41542_, _41518_);
  nor (_41544_, _41543_, _41541_);
  not (_41545_, _41511_);
  or (_41546_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1], \oc8051_top_1.oc8051_sfr1.pres_ow );
  not (_41547_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or (_41548_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _41547_);
  and (_41549_, _41548_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and (_41550_, _41549_, _41546_);
  and (_41551_, _41550_, _41545_);
  and (_41552_, _41551_, _41544_);
  and (_41553_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and (_41554_, _41553_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and (_41555_, _41554_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and (_41556_, _41555_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and (_41557_, _41556_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and (_41558_, _41557_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and (_41559_, _41558_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and (_41560_, _41559_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and (_41561_, _41560_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and (_41562_, _41561_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and (_41563_, _41562_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and (_41564_, _41563_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and (_41565_, _41564_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  and (_41566_, _41565_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  and (_41567_, _41566_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  not (_41568_, _41567_);
  nand (_41569_, _41568_, _41552_);
  or (_41570_, _41552_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  and (_41571_, _41570_, _42618_);
  and (_01643_, _41571_, _41569_);
  nand (_41572_, _41541_, _38225_);
  and (_41573_, _41518_, _36133_);
  and (_41574_, _41573_, _39552_);
  not (_41575_, _41574_);
  not (_41576_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and (_41577_, _41510_, _41576_);
  and (_41578_, _41577_, _41511_);
  and (_41579_, _41578_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  not (_41580_, _41578_);
  not (_41581_, _41512_);
  and (_41582_, _41581_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and (_41583_, _41567_, _41550_);
  and (_41584_, _41583_, _41582_);
  and (_41585_, _41558_, _41550_);
  or (_41586_, _41585_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  nand (_41587_, _41585_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and (_41588_, _41587_, _41586_);
  or (_41589_, _41588_, _41584_);
  and (_41590_, _41589_, _41580_);
  or (_41591_, _41590_, _41579_);
  or (_41592_, _41591_, _41541_);
  and (_41593_, _41592_, _41575_);
  and (_41594_, _41593_, _41572_);
  and (_41595_, _41574_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or (_41596_, _41595_, _41594_);
  and (_01646_, _41596_, _42618_);
  and (_41597_, _41566_, _41550_);
  or (_41598_, _41597_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  nand (_41599_, _41581_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  nand (_41600_, _41599_, _41583_);
  and (_41601_, _41600_, _41598_);
  or (_41602_, _41601_, _41578_);
  or (_41603_, _41580_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  and (_41604_, _41603_, _41544_);
  and (_41605_, _41604_, _41602_);
  and (_41606_, _41541_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  or (_41607_, _41606_, _41605_);
  not (_41608_, _38225_);
  and (_41609_, _41543_, _41608_);
  or (_41610_, _41609_, _41607_);
  and (_01649_, _41610_, _42618_);
  and (_41611_, _41580_, _41550_);
  and (_41612_, _41611_, _41511_);
  nand (_41613_, _41612_, _41567_);
  nand (_41614_, _41613_, _41544_);
  or (_41615_, _41544_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and (_41616_, _41615_, _42618_);
  and (_01652_, _41616_, _41614_);
  or (_41617_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and (_41618_, _40309_, _38614_);
  or (_41619_, _41618_, _41617_);
  nand (_41620_, _38617_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  nand (_41621_, _41620_, _41618_);
  or (_41622_, _41621_, _38618_);
  and (_41623_, _41622_, _41619_);
  and (_41624_, _41518_, _40304_);
  or (_41625_, _41624_, _41623_);
  nand (_41626_, _41624_, _38225_);
  and (_41627_, _41626_, _42618_);
  and (_01655_, _41627_, _41625_);
  or (_41628_, _41513_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  not (_41629_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  nand (_41630_, _41513_, _41629_);
  and (_41631_, _41630_, _41628_);
  or (_41632_, _41631_, _41519_);
  nand (_41633_, _41519_, _38203_);
  and (_41634_, _41633_, _41632_);
  or (_41635_, _41634_, _41528_);
  not (_41636_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  nand (_41637_, _41528_, _41636_);
  and (_41638_, _41637_, _42618_);
  and (_02111_, _41638_, _41635_);
  nand (_41639_, _41519_, _38191_);
  and (_41640_, _41514_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and (_41641_, _41513_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  or (_41642_, _41641_, _41640_);
  or (_41643_, _41642_, _41519_);
  and (_41644_, _41643_, _41639_);
  or (_41645_, _41644_, _41528_);
  or (_41646_, _41529_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and (_41647_, _41646_, _42618_);
  and (_02113_, _41647_, _41645_);
  nand (_41648_, _41519_, _38184_);
  and (_41649_, _41514_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and (_41650_, _41513_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or (_41651_, _41650_, _41649_);
  or (_41652_, _41651_, _41519_);
  and (_41653_, _41652_, _41648_);
  or (_41654_, _41653_, _41528_);
  or (_41655_, _41529_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and (_41656_, _41655_, _42618_);
  and (_02115_, _41656_, _41654_);
  nand (_41657_, _41519_, _38177_);
  and (_41658_, _41514_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and (_41659_, _41513_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or (_41660_, _41659_, _41658_);
  or (_41661_, _41660_, _41519_);
  and (_41662_, _41661_, _41657_);
  or (_41663_, _41662_, _41528_);
  or (_41664_, _41529_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and (_41665_, _41664_, _42618_);
  and (_02117_, _41665_, _41663_);
  nand (_41666_, _41519_, _38169_);
  not (_41667_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  nor (_41668_, _41513_, _41667_);
  and (_41669_, _41513_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or (_41670_, _41669_, _41668_);
  or (_41671_, _41670_, _41519_);
  and (_41672_, _41671_, _41666_);
  or (_41673_, _41672_, _41528_);
  nand (_41674_, _41528_, _41667_);
  and (_41675_, _41674_, _42618_);
  and (_02118_, _41675_, _41673_);
  and (_41676_, _41514_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and (_41677_, _41513_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  nor (_41678_, _41677_, _41676_);
  nor (_41679_, _41678_, _41519_);
  nor (_41680_, _41525_, _38162_);
  or (_41681_, _41680_, _41679_);
  and (_41682_, _41681_, _41529_);
  and (_41683_, _41528_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  or (_41684_, _41683_, _41682_);
  and (_02120_, _41684_, _42618_);
  and (_41685_, _41514_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and (_41686_, _41513_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  nor (_41687_, _41686_, _41685_);
  nor (_41688_, _41687_, _41519_);
  nor (_41689_, _41525_, _38155_);
  or (_41690_, _41689_, _41688_);
  and (_41691_, _41690_, _41529_);
  and (_41692_, _41528_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  or (_41693_, _41692_, _41691_);
  and (_02122_, _41693_, _42618_);
  or (_41694_, _41534_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  not (_41695_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nand (_41696_, _41534_, _41695_);
  and (_41697_, _41696_, _41694_);
  or (_41698_, _41697_, _41528_);
  nand (_41699_, _41528_, _38203_);
  and (_41700_, _41699_, _42618_);
  and (_02124_, _41700_, _41698_);
  and (_41701_, _41536_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  and (_41702_, _41534_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  or (_41703_, _41702_, _41701_);
  or (_41704_, _41703_, _41528_);
  nand (_41705_, _41528_, _38191_);
  and (_41706_, _41705_, _42618_);
  and (_02125_, _41706_, _41704_);
  nand (_41707_, _41528_, _38184_);
  and (_41708_, _41536_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and (_41709_, _41534_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or (_41710_, _41709_, _41708_);
  or (_41711_, _41710_, _41528_);
  and (_41712_, _41711_, _42618_);
  and (_02127_, _41712_, _41707_);
  nand (_41713_, _41528_, _38177_);
  and (_41714_, _41536_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and (_41715_, _41534_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or (_41716_, _41715_, _41714_);
  or (_41717_, _41716_, _41528_);
  and (_41718_, _41717_, _42618_);
  and (_02129_, _41718_, _41713_);
  nand (_41719_, _41528_, _38169_);
  not (_41720_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  nor (_41721_, _41534_, _41720_);
  and (_41722_, _41534_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or (_41723_, _41722_, _41721_);
  or (_41724_, _41723_, _41528_);
  and (_41725_, _41724_, _42618_);
  and (_02131_, _41725_, _41719_);
  nand (_41726_, _41528_, _38162_);
  and (_41727_, _41536_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and (_41728_, _41534_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or (_41729_, _41728_, _41727_);
  or (_41730_, _41729_, _41528_);
  and (_41731_, _41730_, _42618_);
  and (_02132_, _41731_, _41726_);
  nand (_41732_, _41528_, _38155_);
  and (_41733_, _41536_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and (_41734_, _41534_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or (_41735_, _41734_, _41733_);
  or (_41736_, _41735_, _41528_);
  and (_41737_, _41736_, _42618_);
  and (_02134_, _41737_, _41732_);
  or (_41738_, _41550_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and (_41739_, _41550_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  nor (_41740_, _41512_, _41636_);
  nand (_41741_, _41740_, _41567_);
  nand (_41742_, _41741_, _41739_);
  and (_41743_, _41742_, _41738_);
  or (_41744_, _41743_, _41578_);
  and (_41745_, _41578_, _41636_);
  nor (_41746_, _41745_, _41541_);
  and (_41747_, _41746_, _41744_);
  not (_41748_, _41541_);
  nor (_41749_, _41748_, _38203_);
  or (_41750_, _41749_, _41574_);
  or (_41751_, _41750_, _41747_);
  nand (_41752_, _41543_, _41629_);
  and (_41753_, _41752_, _42618_);
  and (_02136_, _41753_, _41751_);
  and (_41754_, _41581_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and (_41755_, _41754_, _41611_);
  and (_41756_, _41755_, _41567_);
  and (_41757_, _41578_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  or (_41758_, _41739_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  nand (_41759_, _41553_, _41550_);
  and (_41760_, _41759_, _41580_);
  and (_41761_, _41760_, _41758_);
  nor (_41762_, _41761_, _41757_);
  nand (_41763_, _41762_, _41544_);
  or (_41764_, _41763_, _41756_);
  nand (_41765_, _41541_, _38191_);
  or (_41766_, _41575_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and (_41767_, _41766_, _42618_);
  and (_41768_, _41767_, _41765_);
  and (_02138_, _41768_, _41764_);
  and (_41769_, _41581_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and (_41770_, _41769_, _41583_);
  and (_41771_, _41759_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  nor (_41772_, _41759_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or (_41773_, _41772_, _41578_);
  or (_41774_, _41773_, _41771_);
  or (_41775_, _41774_, _41770_);
  nor (_41776_, _41580_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  nor (_41777_, _41776_, _41541_);
  and (_41778_, _41777_, _41775_);
  nor (_41779_, _41748_, _38184_);
  or (_41780_, _41779_, _41778_);
  or (_41781_, _41780_, _41574_);
  or (_41782_, _41575_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and (_41783_, _41782_, _42618_);
  and (_02139_, _41783_, _41781_);
  and (_41784_, _41581_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and (_41785_, _41784_, _41583_);
  nand (_41786_, _41554_, _41550_);
  and (_41787_, _41786_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  nor (_41788_, _41786_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or (_41789_, _41788_, _41578_);
  or (_41790_, _41789_, _41787_);
  or (_41791_, _41790_, _41785_);
  nor (_41792_, _41580_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  nor (_41793_, _41792_, _41541_);
  and (_41794_, _41793_, _41791_);
  nor (_41795_, _41748_, _38177_);
  or (_41796_, _41795_, _41794_);
  or (_41797_, _41796_, _41574_);
  or (_41798_, _41575_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and (_41799_, _41798_, _42618_);
  and (_02141_, _41799_, _41797_);
  nor (_41800_, _41512_, _41667_);
  and (_41801_, _41800_, _41583_);
  not (_41802_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and (_41803_, _41555_, _41550_);
  nor (_41804_, _41803_, _41802_);
  and (_41805_, _41803_, _41802_);
  or (_41806_, _41805_, _41578_);
  or (_41807_, _41806_, _41804_);
  or (_41808_, _41807_, _41801_);
  and (_41809_, _41578_, _41667_);
  nor (_41810_, _41809_, _41541_);
  and (_41811_, _41810_, _41808_);
  nor (_41812_, _41748_, _38169_);
  or (_41813_, _41812_, _41811_);
  or (_41814_, _41813_, _41574_);
  nand (_41815_, _41543_, _41802_);
  and (_41816_, _41815_, _42618_);
  and (_02143_, _41816_, _41814_);
  and (_41817_, _41581_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and (_41818_, _41817_, _41583_);
  nand (_41819_, _41556_, _41550_);
  and (_41820_, _41819_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  nor (_41821_, _41819_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or (_41822_, _41821_, _41578_);
  or (_41823_, _41822_, _41820_);
  or (_41824_, _41823_, _41818_);
  nor (_41825_, _41580_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  nor (_41826_, _41825_, _41541_);
  and (_41827_, _41826_, _41824_);
  nor (_41828_, _41748_, _38162_);
  or (_41829_, _41828_, _41827_);
  or (_41830_, _41829_, _41574_);
  or (_41831_, _41575_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and (_41832_, _41831_, _42618_);
  and (_02145_, _41832_, _41830_);
  nor (_41833_, _41748_, _38155_);
  and (_41834_, _41581_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and (_41835_, _41834_, _41583_);
  and (_41836_, _41557_, _41550_);
  nor (_41837_, _41836_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  nor (_41838_, _41837_, _41585_);
  or (_41839_, _41838_, _41578_);
  or (_41840_, _41839_, _41835_);
  nor (_41841_, _41580_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  nor (_41842_, _41841_, _41541_);
  and (_41843_, _41842_, _41840_);
  or (_41844_, _41843_, _41574_);
  or (_41845_, _41844_, _41833_);
  or (_41846_, _41575_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and (_41847_, _41846_, _42618_);
  and (_02146_, _41847_, _41845_);
  not (_41848_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  nor (_41849_, _41512_, _41848_);
  and (_41850_, _41849_, _41583_);
  and (_41851_, _41559_, _41550_);
  or (_41852_, _41851_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nand (_41853_, _41851_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and (_41854_, _41853_, _41852_);
  or (_41855_, _41854_, _41578_);
  or (_41856_, _41855_, _41850_);
  and (_41857_, _41578_, _41848_);
  nor (_41858_, _41857_, _41541_);
  and (_41859_, _41858_, _41856_);
  and (_41860_, _41541_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  or (_41861_, _41860_, _41574_);
  or (_41862_, _41861_, _41859_);
  nand (_41863_, _41543_, _38203_);
  and (_41864_, _41863_, _42618_);
  and (_02148_, _41864_, _41862_);
  and (_41865_, _41581_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  and (_41866_, _41865_, _41583_);
  and (_41867_, _41560_, _41550_);
  or (_41868_, _41867_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  nand (_41869_, _41867_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and (_41870_, _41869_, _41868_);
  or (_41871_, _41870_, _41578_);
  or (_41872_, _41871_, _41866_);
  nor (_41873_, _41580_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  nor (_41874_, _41873_, _41541_);
  and (_41875_, _41874_, _41872_);
  and (_41876_, _41541_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  or (_41877_, _41876_, _41574_);
  or (_41878_, _41877_, _41875_);
  nand (_41879_, _41574_, _38191_);
  and (_41880_, _41879_, _42618_);
  and (_02150_, _41880_, _41878_);
  and (_41881_, _41581_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and (_41882_, _41881_, _41583_);
  nand (_41883_, _41561_, _41550_);
  and (_41884_, _41883_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  nor (_41885_, _41883_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or (_41886_, _41885_, _41578_);
  or (_41887_, _41886_, _41884_);
  or (_41888_, _41887_, _41882_);
  nor (_41889_, _41580_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  nor (_41890_, _41889_, _41541_);
  and (_41891_, _41890_, _41888_);
  and (_41892_, _41541_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or (_41893_, _41892_, _41574_);
  or (_41894_, _41893_, _41891_);
  nand (_41895_, _41574_, _38184_);
  and (_41896_, _41895_, _42618_);
  and (_02152_, _41896_, _41894_);
  and (_41897_, _41581_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and (_41898_, _41897_, _41583_);
  nand (_41899_, _41562_, _41550_);
  and (_41900_, _41899_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  nor (_41901_, _41899_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or (_41902_, _41901_, _41578_);
  or (_41903_, _41902_, _41900_);
  or (_41904_, _41903_, _41898_);
  nor (_41905_, _41580_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  nor (_41906_, _41905_, _41541_);
  and (_41907_, _41906_, _41904_);
  and (_41908_, _41541_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or (_41909_, _41908_, _41574_);
  or (_41910_, _41909_, _41907_);
  nand (_41911_, _41574_, _38177_);
  and (_41912_, _41911_, _42618_);
  and (_02153_, _41912_, _41910_);
  nor (_41913_, _41512_, _41720_);
  and (_41914_, _41913_, _41583_);
  not (_41915_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and (_41916_, _41563_, _41550_);
  nor (_41917_, _41916_, _41915_);
  and (_41918_, _41916_, _41915_);
  or (_41919_, _41918_, _41578_);
  or (_41920_, _41919_, _41917_);
  or (_41921_, _41920_, _41914_);
  and (_41922_, _41578_, _41720_);
  nor (_41923_, _41922_, _41541_);
  and (_41924_, _41923_, _41921_);
  and (_41925_, _41541_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or (_41926_, _41925_, _41574_);
  or (_41927_, _41926_, _41924_);
  nand (_41928_, _41574_, _38169_);
  and (_41929_, _41928_, _42618_);
  and (_02155_, _41929_, _41927_);
  and (_41930_, _41581_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and (_41931_, _41930_, _41583_);
  nand (_41932_, _41564_, _41550_);
  and (_41933_, _41932_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  nor (_41934_, _41932_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or (_41935_, _41934_, _41578_);
  or (_41936_, _41935_, _41933_);
  or (_41937_, _41936_, _41931_);
  nor (_41938_, _41580_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  nor (_41939_, _41938_, _41541_);
  and (_41940_, _41939_, _41937_);
  and (_41941_, _41541_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or (_41942_, _41941_, _41574_);
  or (_41943_, _41942_, _41940_);
  nand (_41944_, _41574_, _38162_);
  and (_41945_, _41944_, _42618_);
  and (_02157_, _41945_, _41943_);
  and (_41946_, _41581_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and (_41947_, _41946_, _41583_);
  and (_41948_, _41565_, _41550_);
  nor (_41949_, _41948_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  nor (_41950_, _41949_, _41597_);
  or (_41951_, _41950_, _41578_);
  or (_41952_, _41951_, _41947_);
  nor (_41953_, _41580_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  nor (_41954_, _41953_, _41541_);
  and (_41955_, _41954_, _41952_);
  and (_41956_, _41541_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or (_41957_, _41956_, _41574_);
  or (_41958_, _41957_, _41955_);
  nand (_41959_, _41574_, _38155_);
  and (_41960_, _41959_, _42618_);
  and (_02159_, _41960_, _41958_);
  not (_41961_, _41624_);
  and (_41962_, _41618_, _38813_);
  or (_41963_, _41962_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and (_41964_, _41963_, _41961_);
  nand (_41965_, _41962_, _31757_);
  and (_41966_, _41965_, _41964_);
  nor (_41967_, _41961_, _38203_);
  or (_41968_, _41967_, _41966_);
  and (_02160_, _41968_, _42618_);
  and (_41969_, _41618_, _33129_);
  or (_41970_, _41969_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  and (_41971_, _41970_, _41961_);
  nand (_41972_, _41969_, _31757_);
  and (_41973_, _41972_, _41971_);
  nor (_41974_, _41961_, _38191_);
  or (_41975_, _41974_, _41973_);
  and (_02162_, _41975_, _42618_);
  nand (_41976_, _41618_, _39025_);
  and (_41977_, _41976_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or (_41978_, _41977_, _41624_);
  and (_41979_, _33880_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or (_41980_, _41979_, _33869_);
  and (_41981_, _41980_, _41618_);
  or (_41982_, _41981_, _41978_);
  nand (_41983_, _41624_, _38184_);
  and (_41984_, _41983_, _42618_);
  and (_02164_, _41984_, _41982_);
  and (_41985_, _41618_, _34576_);
  or (_41986_, _41985_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and (_41987_, _41986_, _41961_);
  nand (_41988_, _41985_, _31757_);
  and (_41989_, _41988_, _41987_);
  nor (_41990_, _41961_, _38177_);
  or (_41991_, _41990_, _41989_);
  and (_02166_, _41991_, _42618_);
  and (_41992_, _41618_, _35338_);
  or (_41993_, _41992_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and (_41994_, _41993_, _41961_);
  nand (_41995_, _41992_, _31757_);
  and (_41996_, _41995_, _41994_);
  nor (_41997_, _41961_, _38169_);
  or (_41998_, _41997_, _41996_);
  and (_02167_, _41998_, _42618_);
  and (_41999_, _41618_, _36133_);
  or (_42000_, _41999_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and (_42001_, _42000_, _41961_);
  nand (_42002_, _41999_, _31757_);
  and (_42003_, _42002_, _42001_);
  nor (_42004_, _41961_, _38162_);
  or (_42005_, _42004_, _42003_);
  and (_02169_, _42005_, _42618_);
  not (_42006_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and (_42007_, _41510_, _42006_);
  or (_42008_, _42007_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or (_42009_, _42008_, _41618_);
  nand (_42010_, _38739_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  nand (_42011_, _42010_, _41618_);
  or (_42012_, _42011_, _38740_);
  and (_42013_, _42012_, _42009_);
  or (_42014_, _42013_, _41624_);
  nand (_42015_, _41624_, _38155_);
  and (_42016_, _42015_, _42618_);
  and (_02171_, _42016_, _42014_);
  and (_42017_, _38227_, _38135_);
  not (_42018_, _42017_);
  not (_42019_, _38133_);
  and (_42020_, _42019_, _38099_);
  and (_42021_, _38638_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  nor (_42022_, _42021_, _38711_);
  nor (_42023_, _42022_, _31790_);
  and (_42024_, _42022_, _31790_);
  or (_42025_, _42024_, _42023_);
  not (_42026_, _42025_);
  and (_42027_, _37657_, _27795_);
  nor (_42028_, _37657_, _27795_);
  nor (_42029_, _42028_, _42027_);
  and (_42030_, _28376_, _28244_);
  not (_42031_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and (_42032_, _31189_, _42031_);
  and (_42033_, _42032_, _33880_);
  and (_42034_, _42033_, _42030_);
  and (_42035_, _42034_, _42029_);
  and (_42036_, _42035_, _27345_);
  and (_42037_, _38716_, _40289_);
  nor (_42038_, _38716_, _40289_);
  nor (_42039_, _42038_, _42037_);
  and (_42040_, _42039_, _42036_);
  and (_42041_, _42040_, _42026_);
  not (_42042_, _38716_);
  nor (_42043_, _42022_, _38004_);
  and (_42044_, _42043_, _42042_);
  and (_42045_, _42044_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  nor (_42046_, _42022_, _37657_);
  and (_42047_, _42046_, _42042_);
  and (_42048_, _42047_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  nor (_42049_, _42048_, _42045_);
  and (_42050_, _42022_, _37657_);
  and (_42051_, _42050_, _42042_);
  and (_42052_, _42051_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  and (_42053_, _42022_, _38004_);
  and (_42054_, _42053_, _38716_);
  and (_42055_, _42054_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  nor (_42056_, _42055_, _42052_);
  and (_42057_, _42056_, _42049_);
  and (_42058_, _42050_, _38716_);
  and (_42059_, _42058_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  and (_42060_, _42043_, _38716_);
  and (_42061_, _42060_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  nor (_42062_, _42061_, _42059_);
  and (_42063_, _42046_, _38716_);
  and (_42064_, _42063_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  and (_42065_, _42053_, _42042_);
  and (_42066_, _42065_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  nor (_42067_, _42066_, _42064_);
  and (_42068_, _42067_, _42062_);
  and (_42069_, _42068_, _42057_);
  nor (_42070_, _42069_, _42041_);
  and (_42071_, _42041_, _41608_);
  nor (_42072_, _42071_, _42070_);
  not (_42073_, _42072_);
  and (_42074_, _42073_, _42020_);
  not (_42075_, _42074_);
  not (_42076_, _37999_);
  nor (_42077_, _42019_, _38099_);
  and (_42078_, _42077_, _37999_);
  not (_42079_, _36958_);
  and (_42080_, _42079_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [7]);
  and (_42081_, _37210_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_42082_, _37232_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nor (_42083_, _42082_, _42081_);
  and (_42084_, _37045_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  and (_42085_, _37133_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor (_42086_, _42085_, _42084_);
  and (_42087_, _37078_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_42088_, _37177_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_42089_, _42088_, _42087_);
  and (_42090_, _42089_, _42086_);
  and (_42091_, _42090_, _42083_);
  nor (_42092_, _37012_, _42079_);
  not (_42093_, _42092_);
  nor (_42094_, _42093_, _42091_);
  nor (_42095_, _42094_, _42080_);
  not (_42096_, _42095_);
  and (_42097_, _42096_, _42078_);
  nor (_42098_, _42097_, _42076_);
  and (_42099_, _42098_, _42075_);
  and (_42100_, _42099_, _42018_);
  and (_42101_, _37987_, _38008_);
  nor (_42102_, _42101_, _38073_);
  and (_42103_, _37962_, _37987_);
  nor (_42104_, _42103_, _38027_);
  not (_42105_, _42104_);
  nor (_42106_, _42105_, _38080_);
  and (_42107_, _42106_, _42102_);
  and (_42108_, _38045_, _38011_);
  and (_42109_, _42108_, _38036_);
  and (_42110_, _42109_, _42107_);
  nor (_42111_, _42110_, _36914_);
  nor (_42112_, _38043_, _38039_);
  not (_42113_, _37990_);
  nor (_42114_, _42113_, _42112_);
  nor (_42115_, _42114_, _42111_);
  not (_42116_, _42115_);
  and (_42117_, _42116_, _42100_);
  and (_42118_, _42079_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [5]);
  and (_42119_, _37078_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_42120_, _37133_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_42121_, _42120_, _42119_);
  and (_42122_, _37210_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_42123_, _37045_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor (_42124_, _42123_, _42122_);
  and (_42125_, _37232_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_42126_, _37177_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_42127_, _42126_, _42125_);
  and (_42128_, _42127_, _42124_);
  and (_42129_, _42128_, _42121_);
  nor (_42130_, _42129_, _42093_);
  nor (_42131_, _42130_, _42118_);
  not (_42132_, _42131_);
  and (_42133_, _42132_, _42078_);
  not (_42134_, _42133_);
  and (_42135_, _42076_, _38133_);
  and (_42136_, _42135_, _38099_);
  not (_42137_, _38265_);
  and (_42138_, _42137_, _38135_);
  nor (_42139_, _42138_, _42136_);
  and (_42140_, _42139_, _42134_);
  and (_42141_, _38134_, _42076_);
  and (_42142_, _42020_, _37999_);
  and (_42143_, _42063_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  and (_42144_, _42054_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  nor (_42145_, _42144_, _42143_);
  and (_42146_, _42065_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  and (_42147_, _42044_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  nor (_42148_, _42147_, _42146_);
  and (_42149_, _42148_, _42145_);
  and (_42150_, _42047_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  and (_42151_, _42051_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  nor (_42152_, _42151_, _42150_);
  and (_42153_, _42060_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  and (_42154_, _42058_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  nor (_42155_, _42154_, _42153_);
  and (_42156_, _42155_, _42152_);
  and (_42157_, _42156_, _42149_);
  nor (_42158_, _42157_, _42041_);
  and (_42159_, _42041_, _39920_);
  nor (_42160_, _42159_, _42158_);
  not (_42161_, _42160_);
  and (_42162_, _42161_, _42142_);
  nor (_42163_, _42162_, _42141_);
  and (_42164_, _42163_, _42140_);
  not (_42165_, _42164_);
  and (_42166_, _42165_, _42117_);
  and (_42167_, _42060_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  and (_42168_, _42058_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  nor (_42169_, _42168_, _42167_);
  and (_42170_, _42044_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  and (_42171_, _42065_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  nor (_42172_, _42171_, _42170_);
  and (_42173_, _42172_, _42169_);
  and (_42174_, _42054_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  and (_42175_, _42047_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  nor (_42176_, _42175_, _42174_);
  and (_42177_, _42063_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  and (_42178_, _42051_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  nor (_42179_, _42178_, _42177_);
  and (_42180_, _42179_, _42176_);
  and (_42181_, _42180_, _42173_);
  nor (_42182_, _42181_, _42041_);
  and (_42183_, _42041_, _39884_);
  nor (_42184_, _42183_, _42182_);
  not (_42185_, _42184_);
  and (_42186_, _42185_, _42142_);
  not (_42187_, _42186_);
  and (_42188_, _37999_, _38133_);
  and (_42189_, _42188_, _38099_);
  and (_42190_, _42189_, _37837_);
  not (_42191_, _42190_);
  not (_42192_, _38247_);
  and (_42193_, _42192_, _38135_);
  and (_42194_, _42079_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [2]);
  and (_42195_, _37078_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_42196_, _37133_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_42197_, _42196_, _42195_);
  and (_42198_, _37210_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_42199_, _37177_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_42200_, _42199_, _42198_);
  and (_42201_, _37045_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  and (_42202_, _37232_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nor (_42203_, _42202_, _42201_);
  and (_42204_, _42203_, _42200_);
  and (_42205_, _42204_, _42197_);
  nor (_42206_, _42205_, _42093_);
  nor (_42207_, _42206_, _42194_);
  not (_42208_, _42207_);
  and (_42209_, _42208_, _42078_);
  nor (_42210_, _42209_, _42193_);
  and (_42211_, _42210_, _42191_);
  and (_42212_, _42211_, _42187_);
  nor (_42213_, _42212_, _42116_);
  nor (_42214_, _42213_, _42166_);
  not (_42215_, _42214_);
  and (_42216_, _42060_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  and (_42217_, _42063_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  nor (_42218_, _42217_, _42216_);
  and (_42219_, _42058_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  and (_42220_, _42051_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  nor (_42221_, _42220_, _42219_);
  and (_42222_, _42221_, _42218_);
  and (_42223_, _42044_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  and (_42224_, _42054_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  nor (_42225_, _42224_, _42223_);
  and (_42226_, _42047_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  and (_42227_, _42065_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  nor (_42228_, _42227_, _42226_);
  and (_42229_, _42228_, _42225_);
  and (_42230_, _42229_, _42222_);
  nor (_42231_, _42230_, _42041_);
  and (_42232_, _42041_, _39907_);
  nor (_42233_, _42232_, _42231_);
  not (_42234_, _42233_);
  and (_42235_, _42234_, _42142_);
  not (_42236_, _42235_);
  not (_42237_, _38259_);
  and (_42238_, _42237_, _38135_);
  nor (_42239_, _42238_, _42135_);
  and (_42240_, _42079_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [4]);
  and (_42241_, _37078_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_42242_, _37133_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_42243_, _42242_, _42241_);
  and (_42244_, _37210_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_42245_, _37177_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_42246_, _42245_, _42244_);
  and (_42247_, _37045_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  and (_42248_, _37232_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nor (_42249_, _42248_, _42247_);
  and (_42250_, _42249_, _42246_);
  and (_42251_, _42250_, _42243_);
  nor (_42252_, _42251_, _42093_);
  nor (_42253_, _42252_, _42240_);
  not (_42254_, _42253_);
  and (_42255_, _42254_, _42078_);
  and (_42256_, _42189_, _42042_);
  nor (_42257_, _42256_, _42255_);
  and (_42258_, _42257_, _42239_);
  and (_42259_, _42258_, _42236_);
  not (_42260_, _42259_);
  and (_42261_, _42260_, _42117_);
  and (_42262_, _42060_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  and (_42263_, _42054_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  nor (_42264_, _42263_, _42262_);
  and (_42265_, _42044_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  and (_42266_, _42065_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  nor (_42267_, _42266_, _42265_);
  and (_42268_, _42267_, _42264_);
  and (_42269_, _42058_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  and (_42270_, _42047_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  nor (_42271_, _42270_, _42269_);
  and (_42272_, _42063_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  and (_42273_, _42051_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  nor (_42274_, _42273_, _42272_);
  and (_42275_, _42274_, _42271_);
  and (_42276_, _42275_, _42268_);
  nor (_42277_, _42276_, _42041_);
  not (_42278_, _38191_);
  and (_42279_, _42041_, _42278_);
  nor (_42280_, _42279_, _42277_);
  not (_42281_, _42280_);
  and (_42282_, _42281_, _42142_);
  not (_42283_, _42282_);
  and (_42284_, _42020_, _42076_);
  and (_42285_, _42079_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [1]);
  and (_42286_, _37210_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_42287_, _37232_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor (_42288_, _42287_, _42286_);
  and (_42289_, _37078_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_42290_, _37177_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_42291_, _42290_, _42289_);
  and (_42292_, _37045_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  and (_42293_, _37133_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_42294_, _42293_, _42292_);
  and (_42295_, _42294_, _42291_);
  and (_42296_, _42295_, _42288_);
  nor (_42297_, _42296_, _42093_);
  nor (_42298_, _42297_, _42285_);
  not (_42299_, _42298_);
  and (_42300_, _42299_, _42078_);
  nor (_42301_, _42300_, _42284_);
  not (_42302_, _38241_);
  and (_42303_, _42302_, _38135_);
  and (_42304_, _42189_, _37863_);
  nor (_42305_, _42304_, _42303_);
  and (_42306_, _42305_, _42301_);
  and (_42307_, _42306_, _42283_);
  nor (_42308_, _42307_, _42116_);
  nor (_42309_, _42308_, _42261_);
  and (_42310_, _42060_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  and (_42311_, _42065_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  nor (_42312_, _42311_, _42310_);
  and (_42313_, _42058_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  and (_42314_, _42054_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  nor (_42315_, _42314_, _42313_);
  and (_42316_, _42315_, _42312_);
  and (_42317_, _42047_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  and (_42318_, _42051_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  nor (_42319_, _42318_, _42317_);
  and (_42320_, _42063_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  and (_42321_, _42044_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  nor (_42322_, _42321_, _42320_);
  and (_42323_, _42322_, _42319_);
  and (_42324_, _42323_, _42316_);
  nor (_42325_, _42324_, _42041_);
  and (_42326_, _42041_, _39896_);
  nor (_42327_, _42326_, _42325_);
  not (_42328_, _42327_);
  and (_42329_, _42328_, _42142_);
  not (_42330_, _42329_);
  not (_42331_, _38253_);
  and (_42332_, _42331_, _38135_);
  not (_42333_, _42332_);
  not (_42334_, _42022_);
  and (_42335_, _42189_, _42334_);
  and (_42336_, _42079_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [3]);
  and (_42337_, _37078_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_42338_, _37133_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_42339_, _42338_, _42337_);
  and (_42340_, _37232_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_42341_, _37177_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_42342_, _42341_, _42340_);
  and (_42343_, _37210_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_42344_, _37045_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor (_42345_, _42344_, _42343_);
  and (_42346_, _42345_, _42342_);
  and (_42347_, _42346_, _42339_);
  nor (_42348_, _42347_, _42093_);
  nor (_42349_, _42348_, _42336_);
  not (_42350_, _42349_);
  and (_42351_, _42350_, _42078_);
  nor (_42352_, _42351_, _42335_);
  and (_42353_, _42352_, _42333_);
  and (_42354_, _42353_, _42330_);
  not (_42355_, _42354_);
  and (_42356_, _42355_, _42117_);
  and (_42357_, _42044_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  and (_42358_, _42047_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  nor (_42359_, _42358_, _42357_);
  and (_42360_, _42051_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  and (_42361_, _42058_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  nor (_42362_, _42361_, _42360_);
  and (_42363_, _42362_, _42359_);
  and (_42364_, _42054_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  and (_42365_, _42060_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  nor (_42366_, _42365_, _42364_);
  and (_42367_, _42063_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  and (_42368_, _42065_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  nor (_42369_, _42368_, _42367_);
  and (_42370_, _42369_, _42366_);
  and (_42371_, _42370_, _42363_);
  nor (_42372_, _42371_, _42041_);
  and (_42373_, _42041_, _38204_);
  nor (_42374_, _42373_, _42372_);
  not (_42375_, _42374_);
  and (_42376_, _42375_, _42142_);
  not (_42377_, _42376_);
  and (_42378_, _42079_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [0]);
  and (_42379_, _37078_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_42380_, _37133_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_42381_, _42380_, _42379_);
  and (_42382_, _37210_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_42383_, _37177_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_42384_, _42383_, _42382_);
  and (_42385_, _37045_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  and (_42386_, _37232_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nor (_42387_, _42386_, _42385_);
  and (_42388_, _42387_, _42384_);
  and (_42389_, _42388_, _42381_);
  nor (_42390_, _42389_, _42093_);
  nor (_42391_, _42390_, _42378_);
  not (_42392_, _42391_);
  and (_42393_, _42392_, _42078_);
  not (_42394_, _42393_);
  not (_42395_, _38235_);
  and (_42396_, _42395_, _38135_);
  and (_42397_, _42189_, _37657_);
  nor (_42398_, _42397_, _42396_);
  and (_42399_, _42398_, _42394_);
  and (_42400_, _42399_, _42377_);
  nor (_42401_, _42400_, _42116_);
  nor (_42402_, _42401_, _42356_);
  or (_42403_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  not (_42404_, _42402_);
  or (_42405_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  and (_42406_, _42405_, _42403_);
  or (_42407_, _42406_, _42309_);
  not (_42408_, _38271_);
  and (_42409_, _42408_, _38135_);
  not (_42410_, _42409_);
  and (_42411_, _42060_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  and (_42412_, _42051_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  nor (_42413_, _42412_, _42411_);
  and (_42414_, _42044_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  and (_42415_, _42054_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  nor (_42416_, _42415_, _42414_);
  and (_42417_, _42416_, _42413_);
  and (_42418_, _42058_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  and (_42419_, _42047_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  nor (_42420_, _42419_, _42418_);
  and (_42421_, _42063_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  and (_42422_, _42065_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  nor (_42423_, _42422_, _42421_);
  and (_42424_, _42423_, _42420_);
  and (_42425_, _42424_, _42417_);
  nor (_42426_, _42425_, _42041_);
  and (_42427_, _42041_, _39933_);
  nor (_42428_, _42427_, _42426_);
  not (_42429_, _42428_);
  and (_42430_, _42429_, _42142_);
  not (_42431_, _42430_);
  nor (_42432_, _42020_, _37999_);
  and (_42433_, _42079_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [6]);
  and (_42434_, _37078_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_42435_, _37133_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor (_42436_, _42435_, _42434_);
  and (_42437_, _37210_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_42438_, _37045_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor (_42439_, _42438_, _42437_);
  and (_42440_, _37232_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_42441_, _37177_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_42442_, _42441_, _42440_);
  and (_42443_, _42442_, _42439_);
  and (_42444_, _42443_, _42436_);
  nor (_42445_, _42444_, _42093_);
  nor (_42446_, _42445_, _42433_);
  not (_42447_, _42446_);
  and (_42448_, _42447_, _42077_);
  nor (_42449_, _42448_, _42432_);
  and (_42450_, _42449_, _42431_);
  and (_42451_, _42450_, _42410_);
  and (_42452_, _42451_, _42117_);
  nor (_42453_, _42355_, _42117_);
  nor (_42454_, _42453_, _42452_);
  not (_42455_, _42309_);
  or (_42456_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  or (_42457_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  and (_42458_, _42457_, _42456_);
  or (_42459_, _42458_, _42455_);
  and (_42460_, _42459_, _42454_);
  and (_42461_, _42460_, _42407_);
  and (_42462_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  and (_42463_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  or (_42464_, _42463_, _42455_);
  or (_42465_, _42464_, _42462_);
  not (_42466_, _42454_);
  and (_42467_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  and (_42468_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  or (_42469_, _42468_, _42309_);
  or (_42470_, _42469_, _42467_);
  and (_42471_, _42470_, _42466_);
  and (_42472_, _42471_, _42465_);
  or (_42473_, _42472_, _42461_);
  and (_42474_, _42473_, _42215_);
  nor (_42475_, _28244_, _27103_);
  nor (_42476_, _42475_, _31190_);
  and (_42477_, _28244_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_42478_, _42477_, _40289_);
  nor (_42479_, _27674_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_42480_, _42479_, _42478_);
  nand (_42481_, _42480_, _42309_);
  or (_42482_, _42480_, _42309_);
  and (_42483_, _42482_, _42481_);
  not (_42484_, _42483_);
  and (_42485_, _42477_, _31790_);
  nor (_42486_, _27795_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_42487_, _42486_, _42485_);
  not (_42488_, _42487_);
  and (_42489_, _42488_, _42402_);
  nor (_42490_, _42488_, _42402_);
  nor (_42491_, _42490_, _42489_);
  and (_42492_, _42491_, _42484_);
  and (_42493_, _42477_, _38138_);
  nor (_42494_, _42477_, _27948_);
  nor (_42495_, _42494_, _42493_);
  nor (_42496_, _42495_, _42454_);
  and (_42497_, _42495_, _42454_);
  nor (_42498_, _42497_, _42496_);
  and (_42499_, _42477_, _38613_);
  nor (_42500_, _28069_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_42501_, _42500_, _42499_);
  not (_42502_, _42501_);
  nor (_42503_, _42502_, _42214_);
  and (_42504_, _42502_, _42214_);
  nor (_42505_, _42504_, _42503_);
  and (_42506_, _42505_, _42498_);
  and (_42507_, _42506_, _42492_);
  and (_42508_, _42507_, _42476_);
  or (_42509_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  or (_42510_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  and (_42511_, _42510_, _42509_);
  or (_42512_, _42511_, _42309_);
  or (_42513_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  or (_42514_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  and (_42515_, _42514_, _42513_);
  or (_42516_, _42515_, _42455_);
  and (_42517_, _42516_, _42454_);
  and (_42518_, _42517_, _42512_);
  and (_42519_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  and (_42520_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  or (_42521_, _42520_, _42455_);
  or (_42522_, _42521_, _42519_);
  and (_42523_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  and (_42524_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  or (_42525_, _42524_, _42309_);
  or (_42526_, _42525_, _42523_);
  and (_42527_, _42526_, _42466_);
  and (_42528_, _42527_, _42522_);
  or (_42529_, _42528_, _42518_);
  and (_42530_, _42529_, _42214_);
  or (_42531_, _42530_, _42508_);
  or (_42532_, _42531_, _42474_);
  nor (_42533_, _42259_, _42117_);
  nor (_42534_, _42477_, _27542_);
  not (_42535_, _42534_);
  and (_42536_, _42535_, _42533_);
  nor (_42537_, _42535_, _42533_);
  nor (_42538_, _42537_, _42536_);
  nor (_42539_, _42165_, _42117_);
  nor (_42540_, _42477_, _38613_);
  not (_42541_, _42540_);
  nor (_42542_, _42541_, _42539_);
  and (_42543_, _42541_, _42539_);
  nor (_42544_, _42543_, _42542_);
  and (_42545_, _42544_, _42538_);
  nor (_42546_, _42100_, _31779_);
  and (_42547_, _42100_, _31779_);
  nor (_42548_, _42547_, _42546_);
  nor (_42549_, _42451_, _42117_);
  nor (_42550_, _42477_, _28376_);
  not (_42551_, _42550_);
  and (_42552_, _42551_, _42549_);
  nor (_42553_, _42551_, _42549_);
  nor (_42554_, _42553_, _42552_);
  and (_42555_, _42554_, _42548_);
  and (_42557_, _42555_, _42545_);
  and (_42558_, _42557_, _42508_);
  not (_42560_, _42558_);
  or (_42562_, _42560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  not (_42563_, _42508_);
  nor (_42565_, _42558_, _42563_);
  nor (_42567_, _42565_, rst);
  and (_42569_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  nand (_42571_, _42569_, _28935_);
  nor (_42572_, _42571_, _31757_);
  nand (_42573_, _28935_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_42574_, _20601_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_42575_, _42574_, _42573_);
  nor (_42576_, _38225_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  or (_42577_, _42576_, _42575_);
  or (_42578_, _42577_, _42572_);
  and (_39844_, _42578_, _42618_);
  or (_42579_, _39844_, _42567_);
  and (_42580_, _42579_, _42562_);
  and (_02564_, _42580_, _42532_);
  not (_42581_, _42476_);
  nor (_42582_, _42487_, _42581_);
  nor (_42583_, _42581_, _42480_);
  and (_42584_, _42583_, _42582_);
  nor (_42585_, _42495_, _42581_);
  nor (_42586_, _42581_, _42501_);
  and (_42587_, _42586_, _42585_);
  and (_42588_, _42587_, _42584_);
  and (_42589_, _42578_, _42476_);
  and (_42590_, _42589_, _42588_);
  not (_42591_, _42588_);
  and (_42592_, _42591_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  or (_02574_, _42592_, _42590_);
  nor (_42593_, _42586_, _42585_);
  nor (_42594_, _42583_, _42582_);
  and (_42595_, _42594_, _42476_);
  and (_42596_, _42595_, _42593_);
  not (_42597_, _42596_);
  and (_42598_, _42597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  and (_42599_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , _29012_);
  and (_42600_, _42599_, _28957_);
  not (_42601_, _42600_);
  nor (_42602_, _42601_, _31757_);
  not (_42603_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand (_42604_, _38203_, _42603_);
  or (_42606_, _19441_, _42603_);
  and (_42608_, _42606_, _42601_);
  and (_42610_, _42608_, _42604_);
  or (_42612_, _42610_, _42602_);
  and (_42614_, _42612_, _42596_);
  or (_02798_, _42614_, _42598_);
  and (_42617_, _42597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  nand (_42619_, _42599_, _28912_);
  nor (_42620_, _42619_, _31757_);
  nor (_42622_, _38191_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_42624_, _42599_, _28847_);
  and (_42625_, _42599_, _28935_);
  or (_42626_, _42625_, _42569_);
  or (_42627_, _42626_, _42624_);
  and (_42628_, _42627_, _20427_);
  or (_42629_, _42628_, _42622_);
  or (_42630_, _42629_, _42620_);
  and (_42631_, _42630_, _42596_);
  or (_02803_, _42631_, _42617_);
  and (_42632_, _42597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  nand (_42633_, _42599_, _28858_);
  nor (_42634_, _42633_, _31757_);
  nor (_42635_, _38184_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_42636_, _42599_, _28891_);
  or (_42637_, _42636_, _42626_);
  and (_42638_, _42637_, _19080_);
  or (_42639_, _42638_, _42635_);
  or (_42640_, _42639_, _42634_);
  and (_42641_, _42640_, _42596_);
  or (_02809_, _42641_, _42632_);
  and (_42642_, _42625_, _32410_);
  nor (_42643_, _38177_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  or (_42644_, _42624_, _42569_);
  or (_42645_, _42644_, _42636_);
  and (_42646_, _42645_, _20112_);
  or (_42647_, _42646_, _42643_);
  or (_42648_, _42647_, _42642_);
  and (_42649_, _42648_, _42596_);
  and (_42650_, _42597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  or (_02814_, _42650_, _42649_);
  nand (_42651_, _42569_, _28957_);
  nor (_42652_, _42651_, _31757_);
  nor (_42653_, _38169_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand (_42654_, _28957_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_42655_, _19277_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_42656_, _42655_, _42654_);
  or (_42657_, _42656_, _42653_);
  or (_42658_, _42657_, _42652_);
  and (_42659_, _42658_, _42596_);
  and (_42660_, _42597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  or (_02819_, _42660_, _42659_);
  nand (_42661_, _42569_, _28912_);
  nor (_42662_, _42661_, _31757_);
  nor (_42663_, _38162_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand (_42664_, _28912_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_42665_, _20264_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_42666_, _42665_, _42664_);
  or (_42667_, _42666_, _42663_);
  or (_42668_, _42667_, _42662_);
  and (_42669_, _42668_, _42596_);
  and (_42670_, _42597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  or (_02824_, _42670_, _42669_);
  and (_42671_, _42597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  nand (_42672_, _42569_, _28858_);
  nor (_42673_, _42672_, _31757_);
  nor (_42674_, _38155_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand (_42675_, _28858_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_42676_, _19615_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_42677_, _42676_, _42675_);
  or (_42678_, _42677_, _42674_);
  or (_42679_, _42678_, _42673_);
  and (_42680_, _42679_, _42596_);
  or (_02829_, _42680_, _42671_);
  and (_42681_, _42597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  and (_42682_, _42596_, _42578_);
  or (_02831_, _42682_, _42681_);
  and (_42683_, _42612_, _42476_);
  and (_42684_, _42582_, _42480_);
  and (_42685_, _42684_, _42593_);
  and (_42686_, _42685_, _42683_);
  not (_42687_, _42685_);
  and (_42688_, _42687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  or (_02839_, _42688_, _42686_);
  and (_42689_, _42630_, _42476_);
  and (_42690_, _42685_, _42689_);
  and (_42691_, _42687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  or (_02842_, _42691_, _42690_);
  and (_42692_, _42640_, _42476_);
  and (_42693_, _42685_, _42692_);
  and (_42694_, _42687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  or (_02846_, _42694_, _42693_);
  and (_42695_, _42648_, _42476_);
  and (_42696_, _42685_, _42695_);
  and (_42697_, _42687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  or (_02850_, _42697_, _42696_);
  and (_42698_, _42658_, _42476_);
  and (_42699_, _42685_, _42698_);
  and (_42700_, _42687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  or (_02853_, _42700_, _42699_);
  and (_42701_, _42668_, _42476_);
  and (_42702_, _42685_, _42701_);
  and (_42703_, _42687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  or (_02856_, _42703_, _42702_);
  and (_42704_, _42679_, _42476_);
  and (_42705_, _42685_, _42704_);
  and (_42706_, _42687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  or (_02860_, _42706_, _42705_);
  and (_42707_, _42685_, _42589_);
  and (_42708_, _42687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  or (_02862_, _42708_, _42707_);
  and (_42709_, _42583_, _42487_);
  and (_42710_, _42709_, _42593_);
  and (_42711_, _42710_, _42683_);
  not (_42712_, _42710_);
  and (_42713_, _42712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  or (_02868_, _42713_, _42711_);
  and (_42714_, _42710_, _42689_);
  and (_42715_, _42712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  or (_02873_, _42715_, _42714_);
  and (_42716_, _42710_, _42692_);
  and (_42717_, _42712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  or (_02876_, _42717_, _42716_);
  and (_42718_, _42710_, _42695_);
  and (_42719_, _42712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or (_02879_, _42719_, _42718_);
  and (_42720_, _42710_, _42698_);
  and (_42721_, _42712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  or (_02884_, _42721_, _42720_);
  and (_42722_, _42710_, _42701_);
  and (_42723_, _42712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  or (_02887_, _42723_, _42722_);
  and (_42724_, _42710_, _42704_);
  and (_42725_, _42712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  or (_02890_, _42725_, _42724_);
  and (_42726_, _42710_, _42589_);
  and (_42727_, _42712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  or (_02893_, _42727_, _42726_);
  and (_42728_, _42593_, _42584_);
  and (_42729_, _42728_, _42683_);
  not (_42730_, _42728_);
  and (_42731_, _42730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  or (_02898_, _42731_, _42729_);
  and (_42732_, _42728_, _42689_);
  and (_42733_, _42730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  or (_02902_, _42733_, _42732_);
  and (_42734_, _42728_, _42692_);
  and (_42735_, _42730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  or (_02905_, _42735_, _42734_);
  and (_42736_, _42728_, _42695_);
  and (_42737_, _42730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  or (_02908_, _42737_, _42736_);
  and (_42738_, _42728_, _42698_);
  and (_42739_, _42730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  or (_02911_, _42739_, _42738_);
  and (_42740_, _42728_, _42701_);
  and (_42741_, _42730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  or (_02915_, _42741_, _42740_);
  and (_42742_, _42728_, _42704_);
  and (_42743_, _42730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  or (_02918_, _42743_, _42742_);
  and (_42744_, _42728_, _42589_);
  and (_42745_, _42730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  or (_02921_, _42745_, _42744_);
  and (_42746_, _42586_, _42495_);
  and (_42747_, _42746_, _42594_);
  and (_42748_, _42747_, _42683_);
  not (_42749_, _42747_);
  and (_42750_, _42749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  or (_02929_, _42750_, _42748_);
  and (_42751_, _42747_, _42689_);
  and (_42752_, _42749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  or (_02933_, _42752_, _42751_);
  and (_42753_, _42747_, _42692_);
  and (_42754_, _42749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  or (_02937_, _42754_, _42753_);
  and (_42755_, _42747_, _42695_);
  and (_42756_, _42749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  or (_02941_, _42756_, _42755_);
  and (_42757_, _42747_, _42698_);
  and (_42758_, _42749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  or (_02945_, _42758_, _42757_);
  and (_42759_, _42747_, _42701_);
  and (_42760_, _42749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  or (_02948_, _42760_, _42759_);
  and (_42761_, _42747_, _42704_);
  and (_42762_, _42749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  or (_02952_, _42762_, _42761_);
  and (_42763_, _42747_, _42589_);
  and (_42764_, _42749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  or (_02956_, _42764_, _42763_);
  and (_42765_, _42746_, _42684_);
  and (_42766_, _42765_, _42683_);
  not (_42767_, _42765_);
  and (_42768_, _42767_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  or (_02960_, _42768_, _42766_);
  and (_42769_, _42765_, _42689_);
  and (_42770_, _42767_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  or (_02964_, _42770_, _42769_);
  and (_42771_, _42765_, _42692_);
  and (_42772_, _42767_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  or (_02969_, _42772_, _42771_);
  and (_42773_, _42765_, _42695_);
  and (_42774_, _42767_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  or (_02973_, _42774_, _42773_);
  and (_42775_, _42765_, _42698_);
  and (_42776_, _42767_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  or (_02977_, _42776_, _42775_);
  and (_42777_, _42765_, _42701_);
  and (_42778_, _42767_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  or (_02982_, _42778_, _42777_);
  and (_42779_, _42765_, _42704_);
  and (_42780_, _42767_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  or (_02986_, _42780_, _42779_);
  and (_42781_, _42765_, _42589_);
  and (_42782_, _42767_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  or (_02988_, _42782_, _42781_);
  and (_42783_, _42746_, _42709_);
  and (_42784_, _42783_, _42683_);
  not (_42785_, _42783_);
  and (_42786_, _42785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  or (_02993_, _42786_, _42784_);
  and (_42787_, _42783_, _42689_);
  and (_42788_, _42785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  or (_02998_, _42788_, _42787_);
  and (_42789_, _42783_, _42692_);
  and (_42790_, _42785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  or (_03002_, _42790_, _42789_);
  and (_42791_, _42783_, _42695_);
  and (_42792_, _42785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or (_03005_, _42792_, _42791_);
  and (_42793_, _42783_, _42698_);
  and (_42794_, _42785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  or (_03010_, _42794_, _42793_);
  and (_42795_, _42783_, _42701_);
  and (_42796_, _42785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  or (_03014_, _42796_, _42795_);
  and (_42797_, _42783_, _42704_);
  and (_42798_, _42785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  or (_03017_, _42798_, _42797_);
  and (_42799_, _42783_, _42589_);
  and (_42800_, _42785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  or (_03020_, _42800_, _42799_);
  and (_42801_, _42746_, _42584_);
  and (_42802_, _42801_, _42683_);
  not (_42803_, _42801_);
  and (_42804_, _42803_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  or (_03026_, _42804_, _42802_);
  and (_42805_, _42801_, _42689_);
  and (_42806_, _42803_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  or (_03030_, _42806_, _42805_);
  and (_42807_, _42801_, _42692_);
  and (_42808_, _42803_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  or (_03033_, _42808_, _42807_);
  and (_42809_, _42801_, _42695_);
  and (_42810_, _42803_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  or (_03037_, _42810_, _42809_);
  and (_42811_, _42801_, _42698_);
  and (_42812_, _42803_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  or (_03040_, _42812_, _42811_);
  and (_42813_, _42801_, _42701_);
  and (_42814_, _42803_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  or (_03043_, _42814_, _42813_);
  and (_42815_, _42801_, _42704_);
  and (_42816_, _42803_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  or (_03046_, _42816_, _42815_);
  and (_42817_, _42801_, _42589_);
  and (_42818_, _42803_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  or (_03049_, _42818_, _42817_);
  and (_42819_, _42585_, _42501_);
  and (_42820_, _42819_, _42594_);
  and (_42821_, _42820_, _42683_);
  not (_42822_, _42820_);
  and (_42823_, _42822_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  or (_03055_, _42823_, _42821_);
  and (_42824_, _42820_, _42689_);
  and (_42825_, _42822_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  or (_03058_, _42825_, _42824_);
  and (_42826_, _42820_, _42692_);
  and (_42827_, _42822_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  or (_03062_, _42827_, _42826_);
  and (_42828_, _42820_, _42695_);
  and (_42829_, _42822_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  or (_03065_, _42829_, _42828_);
  and (_42830_, _42820_, _42698_);
  and (_42831_, _42822_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  or (_03069_, _42831_, _42830_);
  and (_42832_, _42820_, _42701_);
  and (_42833_, _42822_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  or (_03072_, _42833_, _42832_);
  and (_42834_, _42820_, _42704_);
  and (_42835_, _42822_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  or (_03076_, _42835_, _42834_);
  and (_42836_, _42820_, _42589_);
  and (_42837_, _42822_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  or (_03079_, _42837_, _42836_);
  and (_42838_, _42819_, _42684_);
  and (_42839_, _42838_, _42683_);
  not (_42840_, _42838_);
  and (_42841_, _42840_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  or (_03083_, _42841_, _42839_);
  and (_42842_, _42838_, _42689_);
  and (_42843_, _42840_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  or (_03087_, _42843_, _42842_);
  and (_42844_, _42838_, _42692_);
  and (_42845_, _42840_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  or (_03090_, _42845_, _42844_);
  and (_42846_, _42838_, _42695_);
  and (_42847_, _42840_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  or (_03094_, _42847_, _42846_);
  and (_42848_, _42838_, _42698_);
  and (_42849_, _42840_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  or (_03097_, _42849_, _42848_);
  and (_42850_, _42838_, _42701_);
  and (_42851_, _42840_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  or (_03101_, _42851_, _42850_);
  and (_42852_, _42838_, _42704_);
  and (_42853_, _42840_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  or (_03104_, _42853_, _42852_);
  and (_42854_, _42838_, _42589_);
  and (_42855_, _42840_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  or (_03107_, _42855_, _42854_);
  and (_42856_, _42819_, _42709_);
  and (_42857_, _42856_, _42683_);
  not (_42858_, _42856_);
  and (_42859_, _42858_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  or (_03112_, _42859_, _42857_);
  and (_42860_, _42856_, _42689_);
  and (_42861_, _42858_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  or (_03115_, _42861_, _42860_);
  and (_42862_, _42856_, _42692_);
  and (_42863_, _42858_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  or (_03119_, _42863_, _42862_);
  and (_42864_, _42856_, _42695_);
  and (_42865_, _42858_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  or (_03122_, _42865_, _42864_);
  and (_42866_, _42856_, _42698_);
  and (_42867_, _42858_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  or (_03126_, _42867_, _42866_);
  and (_42868_, _42856_, _42701_);
  and (_42869_, _42858_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  or (_03130_, _42869_, _42868_);
  and (_42870_, _42856_, _42704_);
  and (_42871_, _42858_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  or (_03133_, _42871_, _42870_);
  and (_42872_, _42856_, _42589_);
  and (_42873_, _42858_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  or (_03136_, _42873_, _42872_);
  and (_42874_, _42819_, _42584_);
  and (_42875_, _42874_, _42683_);
  not (_42876_, _42874_);
  and (_42877_, _42876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  or (_03140_, _42877_, _42875_);
  and (_42878_, _42874_, _42689_);
  and (_42879_, _42876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  or (_03143_, _42879_, _42878_);
  and (_42880_, _42874_, _42692_);
  and (_42881_, _42876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  or (_03146_, _42881_, _42880_);
  and (_42882_, _42874_, _42695_);
  and (_42883_, _42876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  or (_03149_, _42883_, _42882_);
  and (_42884_, _42874_, _42698_);
  and (_42885_, _42876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  or (_03153_, _42885_, _42884_);
  and (_42886_, _42874_, _42701_);
  and (_42887_, _42876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  or (_03156_, _42887_, _42886_);
  and (_42888_, _42874_, _42704_);
  and (_42889_, _42876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  or (_03159_, _42889_, _42888_);
  and (_42890_, _42874_, _42589_);
  and (_42891_, _42876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  or (_03162_, _42891_, _42890_);
  and (_42892_, _42594_, _42587_);
  and (_42893_, _42892_, _42683_);
  not (_42894_, _42892_);
  and (_42895_, _42894_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  or (_03166_, _42895_, _42893_);
  and (_42896_, _42892_, _42689_);
  and (_42897_, _42894_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  or (_03170_, _42897_, _42896_);
  and (_42898_, _42892_, _42692_);
  and (_42899_, _42894_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  or (_03173_, _42899_, _42898_);
  and (_42900_, _42892_, _42695_);
  and (_42901_, _42894_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  or (_03176_, _42901_, _42900_);
  and (_42902_, _42892_, _42698_);
  and (_42903_, _42894_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  or (_03179_, _42903_, _42902_);
  and (_42904_, _42892_, _42701_);
  and (_42905_, _42894_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  or (_03183_, _42905_, _42904_);
  and (_42906_, _42892_, _42704_);
  and (_42907_, _42894_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  or (_03186_, _42907_, _42906_);
  and (_42908_, _42892_, _42589_);
  and (_42909_, _42894_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  or (_03188_, _42909_, _42908_);
  and (_42910_, _42684_, _42587_);
  and (_42911_, _42910_, _42683_);
  not (_42912_, _42910_);
  and (_42913_, _42912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  or (_03193_, _42913_, _42911_);
  and (_42914_, _42910_, _42689_);
  and (_42915_, _42912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  or (_03196_, _42915_, _42914_);
  and (_42916_, _42910_, _42692_);
  and (_42917_, _42912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  or (_03200_, _42917_, _42916_);
  and (_42918_, _42910_, _42695_);
  and (_42919_, _42912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  or (_03204_, _42919_, _42918_);
  and (_42920_, _42910_, _42698_);
  and (_42921_, _42912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  or (_03207_, _42921_, _42920_);
  and (_42922_, _42910_, _42701_);
  and (_42923_, _42912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  or (_03211_, _42923_, _42922_);
  and (_42924_, _42910_, _42704_);
  and (_42925_, _42912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  or (_03214_, _42925_, _42924_);
  and (_42926_, _42910_, _42589_);
  and (_42927_, _42912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  or (_03217_, _42927_, _42926_);
  and (_42928_, _42709_, _42587_);
  and (_42929_, _42928_, _42683_);
  not (_42930_, _42928_);
  and (_42931_, _42930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  or (_03221_, _42931_, _42929_);
  and (_42932_, _42928_, _42689_);
  and (_42933_, _42930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  or (_03225_, _42933_, _42932_);
  and (_42934_, _42928_, _42692_);
  and (_42935_, _42930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  or (_03228_, _42935_, _42934_);
  and (_42936_, _42928_, _42695_);
  and (_42937_, _42930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  or (_03232_, _42937_, _42936_);
  and (_42938_, _42928_, _42698_);
  and (_42939_, _42930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  or (_03235_, _42939_, _42938_);
  and (_42940_, _42928_, _42701_);
  and (_42941_, _42930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  or (_03238_, _42941_, _42940_);
  and (_42942_, _42928_, _42704_);
  and (_42943_, _42930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  or (_03242_, _42943_, _42942_);
  and (_42944_, _42928_, _42589_);
  and (_42945_, _42930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  or (_03244_, _42945_, _42944_);
  and (_42946_, _42683_, _42588_);
  and (_42947_, _42591_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  or (_03248_, _42947_, _42946_);
  and (_42948_, _42689_, _42588_);
  and (_42949_, _42591_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  or (_03251_, _42949_, _42948_);
  and (_42950_, _42692_, _42588_);
  and (_42951_, _42591_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  or (_03255_, _42951_, _42950_);
  and (_42952_, _42695_, _42588_);
  and (_42953_, _42591_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  or (_03258_, _42953_, _42952_);
  and (_42954_, _42698_, _42588_);
  and (_42955_, _42591_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  or (_03261_, _42955_, _42954_);
  and (_42956_, _42701_, _42588_);
  and (_42957_, _42591_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  or (_03264_, _42957_, _42956_);
  and (_42958_, _42704_, _42588_);
  and (_42959_, _42591_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  or (_03268_, _42959_, _42958_);
  and (_42960_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  and (_42961_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  or (_42962_, _42961_, _42309_);
  or (_42963_, _42962_, _42960_);
  and (_42964_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  and (_42965_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  or (_42966_, _42965_, _42455_);
  or (_42967_, _42966_, _42964_);
  and (_42968_, _42967_, _42963_);
  or (_42969_, _42968_, _42215_);
  and (_42970_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  and (_42971_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  or (_42972_, _42971_, _42309_);
  or (_42973_, _42972_, _42970_);
  and (_42974_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  and (_42975_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  or (_42976_, _42975_, _42455_);
  or (_42977_, _42976_, _42974_);
  and (_42978_, _42977_, _42973_);
  or (_42979_, _42978_, _42214_);
  and (_42980_, _42979_, _42466_);
  and (_42981_, _42980_, _42969_);
  or (_42982_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  or (_42983_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  and (_42984_, _42983_, _42982_);
  or (_42985_, _42984_, _42455_);
  or (_42986_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  or (_42987_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  and (_42988_, _42987_, _42986_);
  or (_42989_, _42988_, _42309_);
  and (_42990_, _42989_, _42985_);
  or (_42991_, _42990_, _42215_);
  or (_42992_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  or (_42993_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  and (_42994_, _42993_, _42992_);
  or (_42995_, _42994_, _42455_);
  or (_42996_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  or (_42997_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  and (_42998_, _42997_, _42996_);
  or (_42999_, _42998_, _42309_);
  and (_43000_, _42999_, _42995_);
  or (_43001_, _43000_, _42214_);
  and (_43002_, _43001_, _42454_);
  and (_43003_, _43002_, _42991_);
  or (_43004_, _43003_, _42981_);
  and (_43005_, _43004_, _42560_);
  and (_43006_, _42558_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  or (_43007_, _43006_, _42565_);
  or (_43008_, _43007_, _43005_);
  and (_39864_, _42612_, _42618_);
  or (_43009_, _39864_, _42567_);
  and (_05053_, _43009_, _43008_);
  and (_43010_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  and (_43011_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  or (_43012_, _43011_, _42309_);
  or (_43013_, _43012_, _43010_);
  and (_43014_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  and (_43015_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  or (_43016_, _43015_, _42455_);
  or (_43017_, _43016_, _43014_);
  and (_43018_, _43017_, _43013_);
  or (_43019_, _43018_, _42215_);
  and (_43020_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  and (_43021_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  or (_43022_, _43021_, _42309_);
  or (_43023_, _43022_, _43020_);
  and (_43024_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  and (_43025_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  or (_43026_, _43025_, _42455_);
  or (_43027_, _43026_, _43024_);
  and (_43028_, _43027_, _43023_);
  or (_43029_, _43028_, _42214_);
  and (_43030_, _43029_, _42466_);
  and (_43031_, _43030_, _43019_);
  or (_43032_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  or (_43033_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  and (_43034_, _43033_, _43032_);
  or (_43035_, _43034_, _42455_);
  or (_43036_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  or (_43037_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  and (_43038_, _43037_, _43036_);
  or (_43039_, _43038_, _42309_);
  and (_43040_, _43039_, _43035_);
  or (_43041_, _43040_, _42215_);
  or (_43042_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  or (_43043_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  and (_43044_, _43043_, _43042_);
  or (_43045_, _43044_, _42455_);
  or (_43046_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  or (_43047_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  and (_43048_, _43047_, _43046_);
  or (_43049_, _43048_, _42309_);
  and (_43050_, _43049_, _43045_);
  or (_43051_, _43050_, _42214_);
  and (_43052_, _43051_, _42454_);
  and (_43053_, _43052_, _43041_);
  or (_43054_, _43053_, _43031_);
  or (_43055_, _43054_, _42558_);
  or (_43056_, _42560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  and (_43057_, _43056_, _42567_);
  and (_43058_, _43057_, _43055_);
  and (_39865_, _42630_, _42618_);
  and (_43059_, _39865_, _42565_);
  or (_05055_, _43059_, _43058_);
  and (_43060_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  and (_43061_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  or (_43062_, _43061_, _42309_);
  or (_43063_, _43062_, _43060_);
  and (_43064_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  and (_43065_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  or (_43066_, _43065_, _42455_);
  or (_43067_, _43066_, _43064_);
  and (_43068_, _43067_, _43063_);
  or (_43069_, _43068_, _42215_);
  and (_43070_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  and (_43071_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  or (_43072_, _43071_, _42309_);
  or (_43073_, _43072_, _43070_);
  and (_43074_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  and (_43075_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  or (_43076_, _43075_, _42455_);
  or (_43077_, _43076_, _43074_);
  and (_43078_, _43077_, _43073_);
  or (_43079_, _43078_, _42214_);
  and (_43080_, _43079_, _42466_);
  and (_43081_, _43080_, _43069_);
  or (_43082_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  or (_43083_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  and (_43084_, _43083_, _43082_);
  or (_43085_, _43084_, _42455_);
  or (_43086_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  or (_43087_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  and (_43088_, _43087_, _43086_);
  or (_43089_, _43088_, _42309_);
  and (_43090_, _43089_, _43085_);
  or (_43091_, _43090_, _42215_);
  or (_43092_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  or (_43093_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  and (_43094_, _43093_, _43092_);
  or (_43095_, _43094_, _42455_);
  or (_43096_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  or (_43097_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  and (_43098_, _43097_, _43096_);
  or (_43099_, _43098_, _42309_);
  and (_43100_, _43099_, _43095_);
  or (_43101_, _43100_, _42214_);
  and (_43102_, _43101_, _42454_);
  and (_43103_, _43102_, _43091_);
  or (_43104_, _43103_, _43081_);
  or (_43105_, _43104_, _42558_);
  or (_43106_, _42560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  and (_43107_, _43106_, _42567_);
  and (_43108_, _43107_, _43105_);
  and (_39866_, _42640_, _42618_);
  and (_43109_, _39866_, _42565_);
  or (_05057_, _43109_, _43108_);
  and (_43110_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  and (_43111_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  or (_43112_, _43111_, _42455_);
  or (_43113_, _43112_, _43110_);
  and (_43114_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  and (_43115_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or (_43116_, _43115_, _42309_);
  or (_43117_, _43116_, _43114_);
  and (_43118_, _43117_, _43113_);
  or (_43119_, _43118_, _42215_);
  and (_43120_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  and (_43121_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or (_43122_, _43121_, _42309_);
  or (_43123_, _43122_, _43120_);
  and (_43124_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  and (_43125_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  or (_43126_, _43125_, _42455_);
  or (_43127_, _43126_, _43124_);
  and (_43128_, _43127_, _43123_);
  or (_43129_, _43128_, _42214_);
  and (_43130_, _43129_, _42466_);
  and (_43131_, _43130_, _43119_);
  and (_43132_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  and (_43133_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  or (_43134_, _43133_, _42309_);
  or (_43135_, _43134_, _43132_);
  and (_43136_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  and (_43137_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  or (_43138_, _43137_, _42455_);
  or (_43139_, _43138_, _43136_);
  and (_43140_, _43139_, _43135_);
  or (_43141_, _43140_, _42215_);
  and (_43142_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  and (_43143_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  or (_43144_, _43143_, _42309_);
  or (_43145_, _43144_, _43142_);
  and (_43146_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  and (_43147_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  or (_43148_, _43147_, _42455_);
  or (_43149_, _43148_, _43146_);
  and (_43150_, _43149_, _43145_);
  or (_43151_, _43150_, _42214_);
  and (_43152_, _43151_, _42454_);
  and (_43158_, _43152_, _43141_);
  or (_43162_, _43158_, _43131_);
  and (_43169_, _43162_, _42563_);
  and (_43177_, _42648_, _42565_);
  and (_43181_, _42558_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  or (_43186_, _43181_, _43177_);
  or (_43194_, _43186_, _43169_);
  and (_05059_, _43194_, _42618_);
  and (_43203_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  and (_43210_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  or (_43218_, _43210_, _42455_);
  or (_43222_, _43218_, _43203_);
  and (_43227_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  and (_43235_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  or (_43241_, _43235_, _42309_);
  or (_43244_, _43241_, _43227_);
  and (_43248_, _43244_, _43222_);
  or (_43259_, _43248_, _42215_);
  and (_43263_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  and (_43270_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  or (_43278_, _43270_, _42309_);
  or (_43282_, _43278_, _43263_);
  and (_43287_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  and (_43295_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  or (_43301_, _43295_, _42455_);
  or (_43305_, _43301_, _43287_);
  and (_43312_, _43305_, _43282_);
  or (_43320_, _43312_, _42214_);
  and (_43324_, _43320_, _42466_);
  and (_43329_, _43324_, _43259_);
  and (_43337_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  and (_43343_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  or (_43346_, _43343_, _42309_);
  or (_43347_, _43346_, _43337_);
  and (_43348_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  and (_43349_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  or (_43350_, _43349_, _42455_);
  or (_43351_, _43350_, _43348_);
  and (_43352_, _43351_, _43347_);
  or (_43353_, _43352_, _42215_);
  and (_43354_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  and (_43355_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  or (_43356_, _43355_, _42309_);
  or (_43357_, _43356_, _43354_);
  and (_43358_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  and (_43359_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  or (_43360_, _43359_, _42455_);
  or (_43361_, _43360_, _43358_);
  and (_43362_, _43361_, _43357_);
  or (_43363_, _43362_, _42214_);
  and (_43364_, _43363_, _42454_);
  and (_43365_, _43364_, _43353_);
  or (_43366_, _43365_, _43329_);
  and (_43367_, _43366_, _42563_);
  and (_43368_, _42658_, _42565_);
  and (_43369_, _42558_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  or (_43370_, _43369_, _43368_);
  or (_43371_, _43370_, _43367_);
  and (_05061_, _43371_, _42618_);
  and (_43372_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  and (_43373_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  or (_43374_, _43373_, _42309_);
  or (_43375_, _43374_, _43372_);
  and (_43376_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  and (_43377_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  or (_43378_, _43377_, _42455_);
  or (_43379_, _43378_, _43376_);
  and (_43380_, _43379_, _43375_);
  or (_43381_, _43380_, _42215_);
  and (_43382_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  and (_43383_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  or (_43384_, _43383_, _42309_);
  or (_43385_, _43384_, _43382_);
  and (_43386_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  and (_43387_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  or (_43388_, _43387_, _42455_);
  or (_43389_, _43388_, _43386_);
  and (_43390_, _43389_, _43385_);
  or (_43391_, _43390_, _42214_);
  and (_43392_, _43391_, _42466_);
  and (_43393_, _43392_, _43381_);
  or (_43394_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  or (_43395_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  and (_43396_, _43395_, _43394_);
  or (_43397_, _43396_, _42455_);
  or (_43398_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  or (_43399_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  and (_43400_, _43399_, _43398_);
  or (_43401_, _43400_, _42309_);
  and (_43402_, _43401_, _43397_);
  or (_43403_, _43402_, _42215_);
  or (_43404_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  or (_43405_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  and (_43406_, _43405_, _43404_);
  or (_43407_, _43406_, _42455_);
  or (_43408_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  or (_43409_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  and (_43410_, _43409_, _43408_);
  or (_43411_, _43410_, _42309_);
  and (_43412_, _43411_, _43407_);
  or (_43413_, _43412_, _42214_);
  and (_43414_, _43413_, _42454_);
  and (_43415_, _43414_, _43403_);
  or (_43416_, _43415_, _43393_);
  or (_43417_, _43416_, _42558_);
  or (_43418_, _42560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  and (_43419_, _43418_, _42567_);
  and (_43420_, _43419_, _43417_);
  and (_39869_, _42668_, _42618_);
  and (_43421_, _39869_, _42565_);
  or (_05063_, _43421_, _43420_);
  and (_43422_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  and (_43423_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  or (_43424_, _43423_, _42309_);
  or (_43425_, _43424_, _43422_);
  and (_43426_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  and (_43427_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  or (_43428_, _43427_, _42455_);
  or (_43429_, _43428_, _43426_);
  and (_43430_, _43429_, _43425_);
  or (_43431_, _43430_, _42215_);
  and (_43432_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  and (_43433_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  or (_43434_, _43433_, _42309_);
  or (_43435_, _43434_, _43432_);
  and (_43436_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  and (_43437_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  or (_43438_, _43437_, _42455_);
  or (_43439_, _43438_, _43436_);
  and (_43440_, _43439_, _43435_);
  or (_43441_, _43440_, _42214_);
  and (_43442_, _43441_, _42466_);
  and (_43443_, _43442_, _43431_);
  or (_43444_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  or (_43445_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  and (_43446_, _43445_, _43444_);
  or (_43447_, _43446_, _42455_);
  or (_43448_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  or (_43449_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  and (_43450_, _43449_, _43448_);
  or (_43451_, _43450_, _42309_);
  and (_43452_, _43451_, _43447_);
  or (_43453_, _43452_, _42215_);
  or (_43454_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  or (_43455_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  and (_43456_, _43455_, _43454_);
  or (_43457_, _43456_, _42455_);
  or (_43458_, _42402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  or (_43459_, _42404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  and (_43460_, _43459_, _43458_);
  or (_43461_, _43460_, _42309_);
  and (_43462_, _43461_, _43457_);
  or (_43463_, _43462_, _42214_);
  and (_43464_, _43463_, _42454_);
  and (_43465_, _43464_, _43453_);
  or (_43466_, _43465_, _43443_);
  or (_43467_, _43466_, _42558_);
  or (_43468_, _42560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  and (_43469_, _43468_, _42567_);
  and (_43470_, _43469_, _43467_);
  and (_39870_, _42679_, _42618_);
  and (_43471_, _39870_, _42565_);
  or (_05065_, _43471_, _43470_);
  or (_43472_, \oc8051_gm_cxrom_1.cell0.valid , word_in[7]);
  not (_43473_, \oc8051_gm_cxrom_1.cell0.valid );
  or (_43474_, _43473_, \oc8051_gm_cxrom_1.cell0.data [7]);
  nand (_43475_, _43474_, _43472_);
  nand (_43476_, _43475_, _42618_);
  or (_43477_, \oc8051_gm_cxrom_1.cell0.data [7], _42618_);
  and (_05073_, _43477_, _43476_);
  or (_43478_, word_in[0], \oc8051_gm_cxrom_1.cell0.valid );
  or (_43479_, \oc8051_gm_cxrom_1.cell0.data [0], _43473_);
  nand (_43480_, _43479_, _43478_);
  nand (_43481_, _43480_, _42618_);
  or (_43482_, \oc8051_gm_cxrom_1.cell0.data [0], _42618_);
  and (_05080_, _43482_, _43481_);
  or (_43483_, word_in[1], \oc8051_gm_cxrom_1.cell0.valid );
  or (_43484_, \oc8051_gm_cxrom_1.cell0.data [1], _43473_);
  nand (_43485_, _43484_, _43483_);
  nand (_43486_, _43485_, _42618_);
  or (_43487_, \oc8051_gm_cxrom_1.cell0.data [1], _42618_);
  and (_05083_, _43487_, _43486_);
  or (_43488_, word_in[2], \oc8051_gm_cxrom_1.cell0.valid );
  or (_43489_, \oc8051_gm_cxrom_1.cell0.data [2], _43473_);
  nand (_43490_, _43489_, _43488_);
  nand (_43491_, _43490_, _42618_);
  or (_43492_, \oc8051_gm_cxrom_1.cell0.data [2], _42618_);
  and (_05087_, _43492_, _43491_);
  or (_43493_, word_in[3], \oc8051_gm_cxrom_1.cell0.valid );
  or (_43494_, \oc8051_gm_cxrom_1.cell0.data [3], _43473_);
  nand (_43495_, _43494_, _43493_);
  nand (_43496_, _43495_, _42618_);
  or (_43497_, \oc8051_gm_cxrom_1.cell0.data [3], _42618_);
  and (_05091_, _43497_, _43496_);
  or (_43498_, word_in[4], \oc8051_gm_cxrom_1.cell0.valid );
  or (_43499_, \oc8051_gm_cxrom_1.cell0.data [4], _43473_);
  nand (_43500_, _43499_, _43498_);
  nand (_43501_, _43500_, _42618_);
  or (_43502_, \oc8051_gm_cxrom_1.cell0.data [4], _42618_);
  and (_05095_, _43502_, _43501_);
  or (_43503_, word_in[5], \oc8051_gm_cxrom_1.cell0.valid );
  or (_43504_, \oc8051_gm_cxrom_1.cell0.data [5], _43473_);
  nand (_43505_, _43504_, _43503_);
  nand (_43506_, _43505_, _42618_);
  or (_43507_, \oc8051_gm_cxrom_1.cell0.data [5], _42618_);
  and (_05099_, _43507_, _43506_);
  or (_43508_, word_in[6], \oc8051_gm_cxrom_1.cell0.valid );
  or (_43509_, \oc8051_gm_cxrom_1.cell0.data [6], _43473_);
  nand (_43510_, _43509_, _43508_);
  nand (_43511_, _43510_, _42618_);
  or (_43512_, \oc8051_gm_cxrom_1.cell0.data [6], _42618_);
  and (_05103_, _43512_, _43511_);
  or (_43513_, \oc8051_gm_cxrom_1.cell1.valid , word_in[15]);
  not (_43514_, \oc8051_gm_cxrom_1.cell1.valid );
  or (_43515_, _43514_, \oc8051_gm_cxrom_1.cell1.data [7]);
  nand (_43516_, _43515_, _43513_);
  nand (_43517_, _43516_, _42618_);
  or (_43518_, \oc8051_gm_cxrom_1.cell1.data [7], _42618_);
  and (_05124_, _43518_, _43517_);
  or (_43519_, word_in[8], \oc8051_gm_cxrom_1.cell1.valid );
  or (_43520_, \oc8051_gm_cxrom_1.cell1.data [0], _43514_);
  nand (_43521_, _43520_, _43519_);
  nand (_43522_, _43521_, _42618_);
  or (_43523_, \oc8051_gm_cxrom_1.cell1.data [0], _42618_);
  and (_05131_, _43523_, _43522_);
  or (_43524_, word_in[9], \oc8051_gm_cxrom_1.cell1.valid );
  or (_43525_, \oc8051_gm_cxrom_1.cell1.data [1], _43514_);
  nand (_43526_, _43525_, _43524_);
  nand (_43527_, _43526_, _42618_);
  or (_43528_, \oc8051_gm_cxrom_1.cell1.data [1], _42618_);
  and (_05135_, _43528_, _43527_);
  or (_43529_, word_in[10], \oc8051_gm_cxrom_1.cell1.valid );
  or (_43530_, \oc8051_gm_cxrom_1.cell1.data [2], _43514_);
  nand (_43531_, _43530_, _43529_);
  nand (_43532_, _43531_, _42618_);
  or (_43533_, \oc8051_gm_cxrom_1.cell1.data [2], _42618_);
  and (_05139_, _43533_, _43532_);
  or (_00001_, word_in[11], \oc8051_gm_cxrom_1.cell1.valid );
  or (_00002_, \oc8051_gm_cxrom_1.cell1.data [3], _43514_);
  nand (_00003_, _00002_, _00001_);
  nand (_00004_, _00003_, _42618_);
  or (_00005_, \oc8051_gm_cxrom_1.cell1.data [3], _42618_);
  and (_05143_, _00005_, _00004_);
  or (_00006_, word_in[12], \oc8051_gm_cxrom_1.cell1.valid );
  or (_00007_, \oc8051_gm_cxrom_1.cell1.data [4], _43514_);
  nand (_00008_, _00007_, _00006_);
  nand (_00009_, _00008_, _42618_);
  or (_00010_, \oc8051_gm_cxrom_1.cell1.data [4], _42618_);
  and (_05147_, _00010_, _00009_);
  or (_00011_, word_in[13], \oc8051_gm_cxrom_1.cell1.valid );
  or (_00012_, \oc8051_gm_cxrom_1.cell1.data [5], _43514_);
  nand (_00013_, _00012_, _00011_);
  nand (_00014_, _00013_, _42618_);
  or (_00015_, \oc8051_gm_cxrom_1.cell1.data [5], _42618_);
  and (_05151_, _00015_, _00014_);
  or (_00016_, word_in[14], \oc8051_gm_cxrom_1.cell1.valid );
  or (_00017_, \oc8051_gm_cxrom_1.cell1.data [6], _43514_);
  nand (_00018_, _00017_, _00016_);
  nand (_00019_, _00018_, _42618_);
  or (_00020_, \oc8051_gm_cxrom_1.cell1.data [6], _42618_);
  and (_05155_, _00020_, _00019_);
  or (_00021_, \oc8051_gm_cxrom_1.cell2.valid , word_in[23]);
  not (_00022_, \oc8051_gm_cxrom_1.cell2.valid );
  or (_00023_, _00022_, \oc8051_gm_cxrom_1.cell2.data [7]);
  nand (_00024_, _00023_, _00021_);
  nand (_00025_, _00024_, _42618_);
  or (_00026_, \oc8051_gm_cxrom_1.cell2.data [7], _42618_);
  and (_05176_, _00026_, _00025_);
  or (_00027_, word_in[16], \oc8051_gm_cxrom_1.cell2.valid );
  or (_00028_, \oc8051_gm_cxrom_1.cell2.data [0], _00022_);
  nand (_00029_, _00028_, _00027_);
  nand (_00030_, _00029_, _42618_);
  or (_00031_, \oc8051_gm_cxrom_1.cell2.data [0], _42618_);
  and (_05183_, _00031_, _00030_);
  or (_00032_, word_in[17], \oc8051_gm_cxrom_1.cell2.valid );
  or (_00033_, \oc8051_gm_cxrom_1.cell2.data [1], _00022_);
  nand (_00034_, _00033_, _00032_);
  nand (_00035_, _00034_, _42618_);
  or (_00036_, \oc8051_gm_cxrom_1.cell2.data [1], _42618_);
  and (_05187_, _00036_, _00035_);
  or (_00037_, word_in[18], \oc8051_gm_cxrom_1.cell2.valid );
  or (_00038_, \oc8051_gm_cxrom_1.cell2.data [2], _00022_);
  nand (_00039_, _00038_, _00037_);
  nand (_00040_, _00039_, _42618_);
  or (_00041_, \oc8051_gm_cxrom_1.cell2.data [2], _42618_);
  and (_05191_, _00041_, _00040_);
  or (_00042_, word_in[19], \oc8051_gm_cxrom_1.cell2.valid );
  or (_00043_, \oc8051_gm_cxrom_1.cell2.data [3], _00022_);
  nand (_00044_, _00043_, _00042_);
  nand (_00045_, _00044_, _42618_);
  or (_00046_, \oc8051_gm_cxrom_1.cell2.data [3], _42618_);
  and (_05194_, _00046_, _00045_);
  or (_00047_, word_in[20], \oc8051_gm_cxrom_1.cell2.valid );
  or (_00048_, \oc8051_gm_cxrom_1.cell2.data [4], _00022_);
  nand (_00049_, _00048_, _00047_);
  nand (_00050_, _00049_, _42618_);
  or (_00051_, \oc8051_gm_cxrom_1.cell2.data [4], _42618_);
  and (_05198_, _00051_, _00050_);
  or (_00052_, word_in[21], \oc8051_gm_cxrom_1.cell2.valid );
  or (_00053_, \oc8051_gm_cxrom_1.cell2.data [5], _00022_);
  nand (_00054_, _00053_, _00052_);
  nand (_00055_, _00054_, _42618_);
  or (_00056_, \oc8051_gm_cxrom_1.cell2.data [5], _42618_);
  and (_05202_, _00056_, _00055_);
  or (_00057_, word_in[22], \oc8051_gm_cxrom_1.cell2.valid );
  or (_00058_, \oc8051_gm_cxrom_1.cell2.data [6], _00022_);
  nand (_00059_, _00058_, _00057_);
  nand (_00060_, _00059_, _42618_);
  or (_00061_, \oc8051_gm_cxrom_1.cell2.data [6], _42618_);
  and (_05206_, _00061_, _00060_);
  or (_00062_, \oc8051_gm_cxrom_1.cell3.valid , word_in[31]);
  not (_00063_, \oc8051_gm_cxrom_1.cell3.valid );
  or (_00064_, _00063_, \oc8051_gm_cxrom_1.cell3.data [7]);
  nand (_00065_, _00064_, _00062_);
  nand (_00066_, _00065_, _42618_);
  or (_00067_, \oc8051_gm_cxrom_1.cell3.data [7], _42618_);
  and (_05227_, _00067_, _00066_);
  or (_00068_, word_in[24], \oc8051_gm_cxrom_1.cell3.valid );
  or (_00069_, \oc8051_gm_cxrom_1.cell3.data [0], _00063_);
  nand (_00070_, _00069_, _00068_);
  nand (_00071_, _00070_, _42618_);
  or (_00072_, \oc8051_gm_cxrom_1.cell3.data [0], _42618_);
  and (_05234_, _00072_, _00071_);
  or (_00073_, word_in[25], \oc8051_gm_cxrom_1.cell3.valid );
  or (_00074_, \oc8051_gm_cxrom_1.cell3.data [1], _00063_);
  nand (_00075_, _00074_, _00073_);
  nand (_00076_, _00075_, _42618_);
  or (_00077_, \oc8051_gm_cxrom_1.cell3.data [1], _42618_);
  and (_05238_, _00077_, _00076_);
  or (_00078_, word_in[26], \oc8051_gm_cxrom_1.cell3.valid );
  or (_00079_, \oc8051_gm_cxrom_1.cell3.data [2], _00063_);
  nand (_00080_, _00079_, _00078_);
  nand (_00081_, _00080_, _42618_);
  or (_00082_, \oc8051_gm_cxrom_1.cell3.data [2], _42618_);
  and (_05242_, _00082_, _00081_);
  or (_00083_, word_in[27], \oc8051_gm_cxrom_1.cell3.valid );
  or (_00084_, \oc8051_gm_cxrom_1.cell3.data [3], _00063_);
  nand (_00085_, _00084_, _00083_);
  nand (_00086_, _00085_, _42618_);
  or (_00087_, \oc8051_gm_cxrom_1.cell3.data [3], _42618_);
  and (_05246_, _00087_, _00086_);
  or (_00088_, word_in[28], \oc8051_gm_cxrom_1.cell3.valid );
  or (_00089_, \oc8051_gm_cxrom_1.cell3.data [4], _00063_);
  nand (_00090_, _00089_, _00088_);
  nand (_00091_, _00090_, _42618_);
  or (_00092_, \oc8051_gm_cxrom_1.cell3.data [4], _42618_);
  and (_05250_, _00092_, _00091_);
  or (_00093_, word_in[29], \oc8051_gm_cxrom_1.cell3.valid );
  or (_00094_, \oc8051_gm_cxrom_1.cell3.data [5], _00063_);
  nand (_00095_, _00094_, _00093_);
  nand (_00096_, _00095_, _42618_);
  or (_00097_, \oc8051_gm_cxrom_1.cell3.data [5], _42618_);
  and (_05254_, _00097_, _00096_);
  or (_00098_, word_in[30], \oc8051_gm_cxrom_1.cell3.valid );
  or (_00099_, \oc8051_gm_cxrom_1.cell3.data [6], _00063_);
  nand (_00100_, _00099_, _00098_);
  nand (_00101_, _00100_, _42618_);
  or (_00102_, \oc8051_gm_cxrom_1.cell3.data [6], _42618_);
  and (_05258_, _00102_, _00101_);
  or (_00103_, \oc8051_gm_cxrom_1.cell4.valid , word_in[39]);
  not (_00104_, \oc8051_gm_cxrom_1.cell4.valid );
  or (_00105_, _00104_, \oc8051_gm_cxrom_1.cell4.data [7]);
  nand (_00106_, _00105_, _00103_);
  nand (_00107_, _00106_, _42618_);
  or (_00108_, \oc8051_gm_cxrom_1.cell4.data [7], _42618_);
  and (_05279_, _00108_, _00107_);
  or (_00109_, word_in[32], \oc8051_gm_cxrom_1.cell4.valid );
  or (_00110_, \oc8051_gm_cxrom_1.cell4.data [0], _00104_);
  nand (_00111_, _00110_, _00109_);
  nand (_00112_, _00111_, _42618_);
  or (_00113_, \oc8051_gm_cxrom_1.cell4.data [0], _42618_);
  and (_05286_, _00113_, _00112_);
  or (_00114_, word_in[33], \oc8051_gm_cxrom_1.cell4.valid );
  or (_00115_, \oc8051_gm_cxrom_1.cell4.data [1], _00104_);
  nand (_00116_, _00115_, _00114_);
  nand (_00117_, _00116_, _42618_);
  or (_00118_, \oc8051_gm_cxrom_1.cell4.data [1], _42618_);
  and (_05290_, _00118_, _00117_);
  or (_00119_, word_in[34], \oc8051_gm_cxrom_1.cell4.valid );
  or (_00120_, \oc8051_gm_cxrom_1.cell4.data [2], _00104_);
  nand (_00121_, _00120_, _00119_);
  nand (_00122_, _00121_, _42618_);
  or (_00123_, \oc8051_gm_cxrom_1.cell4.data [2], _42618_);
  and (_05294_, _00123_, _00122_);
  or (_00124_, word_in[35], \oc8051_gm_cxrom_1.cell4.valid );
  or (_00125_, \oc8051_gm_cxrom_1.cell4.data [3], _00104_);
  nand (_00126_, _00125_, _00124_);
  nand (_00127_, _00126_, _42618_);
  or (_00128_, \oc8051_gm_cxrom_1.cell4.data [3], _42618_);
  and (_05298_, _00128_, _00127_);
  or (_00129_, word_in[36], \oc8051_gm_cxrom_1.cell4.valid );
  or (_00131_, \oc8051_gm_cxrom_1.cell4.data [4], _00104_);
  nand (_00133_, _00131_, _00129_);
  nand (_00135_, _00133_, _42618_);
  or (_00137_, \oc8051_gm_cxrom_1.cell4.data [4], _42618_);
  and (_05301_, _00137_, _00135_);
  or (_00140_, word_in[37], \oc8051_gm_cxrom_1.cell4.valid );
  or (_00142_, \oc8051_gm_cxrom_1.cell4.data [5], _00104_);
  nand (_00144_, _00142_, _00140_);
  nand (_00146_, _00144_, _42618_);
  or (_00148_, \oc8051_gm_cxrom_1.cell4.data [5], _42618_);
  and (_05305_, _00148_, _00146_);
  or (_00151_, word_in[38], \oc8051_gm_cxrom_1.cell4.valid );
  or (_00153_, \oc8051_gm_cxrom_1.cell4.data [6], _00104_);
  nand (_00155_, _00153_, _00151_);
  nand (_00157_, _00155_, _42618_);
  or (_00159_, \oc8051_gm_cxrom_1.cell4.data [6], _42618_);
  and (_05309_, _00159_, _00157_);
  or (_00162_, \oc8051_gm_cxrom_1.cell5.valid , word_in[47]);
  not (_00164_, \oc8051_gm_cxrom_1.cell5.valid );
  or (_00166_, _00164_, \oc8051_gm_cxrom_1.cell5.data [7]);
  nand (_00168_, _00166_, _00162_);
  nand (_00170_, _00168_, _42618_);
  or (_00172_, \oc8051_gm_cxrom_1.cell5.data [7], _42618_);
  and (_05331_, _00172_, _00170_);
  or (_00175_, word_in[40], \oc8051_gm_cxrom_1.cell5.valid );
  or (_00177_, \oc8051_gm_cxrom_1.cell5.data [0], _00164_);
  nand (_00179_, _00177_, _00175_);
  nand (_00181_, _00179_, _42618_);
  or (_00183_, \oc8051_gm_cxrom_1.cell5.data [0], _42618_);
  and (_05337_, _00183_, _00181_);
  or (_00186_, word_in[41], \oc8051_gm_cxrom_1.cell5.valid );
  or (_00187_, \oc8051_gm_cxrom_1.cell5.data [1], _00164_);
  nand (_00188_, _00187_, _00186_);
  nand (_00189_, _00188_, _42618_);
  or (_00190_, \oc8051_gm_cxrom_1.cell5.data [1], _42618_);
  and (_05341_, _00190_, _00189_);
  or (_00191_, word_in[42], \oc8051_gm_cxrom_1.cell5.valid );
  or (_00192_, \oc8051_gm_cxrom_1.cell5.data [2], _00164_);
  nand (_00193_, _00192_, _00191_);
  nand (_00194_, _00193_, _42618_);
  or (_00195_, \oc8051_gm_cxrom_1.cell5.data [2], _42618_);
  and (_05345_, _00195_, _00194_);
  or (_00196_, word_in[43], \oc8051_gm_cxrom_1.cell5.valid );
  or (_00197_, \oc8051_gm_cxrom_1.cell5.data [3], _00164_);
  nand (_00198_, _00197_, _00196_);
  nand (_00199_, _00198_, _42618_);
  or (_00200_, \oc8051_gm_cxrom_1.cell5.data [3], _42618_);
  and (_05349_, _00200_, _00199_);
  or (_00201_, word_in[44], \oc8051_gm_cxrom_1.cell5.valid );
  or (_00202_, \oc8051_gm_cxrom_1.cell5.data [4], _00164_);
  nand (_00203_, _00202_, _00201_);
  nand (_00204_, _00203_, _42618_);
  or (_00205_, \oc8051_gm_cxrom_1.cell5.data [4], _42618_);
  and (_05353_, _00205_, _00204_);
  or (_00206_, word_in[45], \oc8051_gm_cxrom_1.cell5.valid );
  or (_00207_, \oc8051_gm_cxrom_1.cell5.data [5], _00164_);
  nand (_00208_, _00207_, _00206_);
  nand (_00209_, _00208_, _42618_);
  or (_00210_, \oc8051_gm_cxrom_1.cell5.data [5], _42618_);
  and (_05357_, _00210_, _00209_);
  or (_00211_, word_in[46], \oc8051_gm_cxrom_1.cell5.valid );
  or (_00212_, \oc8051_gm_cxrom_1.cell5.data [6], _00164_);
  nand (_00213_, _00212_, _00211_);
  nand (_00214_, _00213_, _42618_);
  or (_00215_, \oc8051_gm_cxrom_1.cell5.data [6], _42618_);
  and (_05361_, _00215_, _00214_);
  or (_00216_, \oc8051_gm_cxrom_1.cell6.valid , word_in[55]);
  not (_00217_, \oc8051_gm_cxrom_1.cell6.valid );
  or (_00218_, _00217_, \oc8051_gm_cxrom_1.cell6.data [7]);
  nand (_00219_, _00218_, _00216_);
  nand (_00220_, _00219_, _42618_);
  or (_00221_, \oc8051_gm_cxrom_1.cell6.data [7], _42618_);
  and (_05382_, _00221_, _00220_);
  or (_00222_, word_in[48], \oc8051_gm_cxrom_1.cell6.valid );
  or (_00223_, \oc8051_gm_cxrom_1.cell6.data [0], _00217_);
  nand (_00224_, _00223_, _00222_);
  nand (_00225_, _00224_, _42618_);
  or (_00226_, \oc8051_gm_cxrom_1.cell6.data [0], _42618_);
  and (_05389_, _00226_, _00225_);
  or (_00227_, word_in[49], \oc8051_gm_cxrom_1.cell6.valid );
  or (_00228_, \oc8051_gm_cxrom_1.cell6.data [1], _00217_);
  nand (_00229_, _00228_, _00227_);
  nand (_00230_, _00229_, _42618_);
  or (_00231_, \oc8051_gm_cxrom_1.cell6.data [1], _42618_);
  and (_05393_, _00231_, _00230_);
  or (_00232_, word_in[50], \oc8051_gm_cxrom_1.cell6.valid );
  or (_00233_, \oc8051_gm_cxrom_1.cell6.data [2], _00217_);
  nand (_00234_, _00233_, _00232_);
  nand (_00235_, _00234_, _42618_);
  or (_00236_, \oc8051_gm_cxrom_1.cell6.data [2], _42618_);
  and (_05397_, _00236_, _00235_);
  or (_00237_, word_in[51], \oc8051_gm_cxrom_1.cell6.valid );
  or (_00238_, \oc8051_gm_cxrom_1.cell6.data [3], _00217_);
  nand (_00239_, _00238_, _00237_);
  nand (_00240_, _00239_, _42618_);
  or (_00241_, \oc8051_gm_cxrom_1.cell6.data [3], _42618_);
  and (_05401_, _00241_, _00240_);
  or (_00242_, word_in[52], \oc8051_gm_cxrom_1.cell6.valid );
  or (_00243_, \oc8051_gm_cxrom_1.cell6.data [4], _00217_);
  nand (_00244_, _00243_, _00242_);
  nand (_00245_, _00244_, _42618_);
  or (_00246_, \oc8051_gm_cxrom_1.cell6.data [4], _42618_);
  and (_05405_, _00246_, _00245_);
  or (_00247_, word_in[53], \oc8051_gm_cxrom_1.cell6.valid );
  or (_00248_, \oc8051_gm_cxrom_1.cell6.data [5], _00217_);
  nand (_00249_, _00248_, _00247_);
  nand (_00250_, _00249_, _42618_);
  or (_00251_, \oc8051_gm_cxrom_1.cell6.data [5], _42618_);
  and (_05409_, _00251_, _00250_);
  or (_00252_, word_in[54], \oc8051_gm_cxrom_1.cell6.valid );
  or (_00253_, \oc8051_gm_cxrom_1.cell6.data [6], _00217_);
  nand (_00254_, _00253_, _00252_);
  nand (_00255_, _00254_, _42618_);
  or (_00256_, \oc8051_gm_cxrom_1.cell6.data [6], _42618_);
  and (_05412_, _00256_, _00255_);
  or (_00257_, \oc8051_gm_cxrom_1.cell7.valid , word_in[63]);
  not (_00258_, \oc8051_gm_cxrom_1.cell7.valid );
  or (_00259_, _00258_, \oc8051_gm_cxrom_1.cell7.data [7]);
  nand (_00260_, _00259_, _00257_);
  nand (_00261_, _00260_, _42618_);
  or (_00262_, \oc8051_gm_cxrom_1.cell7.data [7], _42618_);
  and (_05434_, _00262_, _00261_);
  or (_00263_, word_in[56], \oc8051_gm_cxrom_1.cell7.valid );
  or (_00264_, \oc8051_gm_cxrom_1.cell7.data [0], _00258_);
  nand (_00265_, _00264_, _00263_);
  nand (_00266_, _00265_, _42618_);
  or (_00267_, \oc8051_gm_cxrom_1.cell7.data [0], _42618_);
  and (_05441_, _00267_, _00266_);
  or (_00268_, word_in[57], \oc8051_gm_cxrom_1.cell7.valid );
  or (_00269_, \oc8051_gm_cxrom_1.cell7.data [1], _00258_);
  nand (_00270_, _00269_, _00268_);
  nand (_00271_, _00270_, _42618_);
  or (_00272_, \oc8051_gm_cxrom_1.cell7.data [1], _42618_);
  and (_05445_, _00272_, _00271_);
  or (_00273_, word_in[58], \oc8051_gm_cxrom_1.cell7.valid );
  or (_00274_, \oc8051_gm_cxrom_1.cell7.data [2], _00258_);
  nand (_00275_, _00274_, _00273_);
  nand (_00276_, _00275_, _42618_);
  or (_00277_, \oc8051_gm_cxrom_1.cell7.data [2], _42618_);
  and (_05448_, _00277_, _00276_);
  or (_00278_, word_in[59], \oc8051_gm_cxrom_1.cell7.valid );
  or (_00279_, \oc8051_gm_cxrom_1.cell7.data [3], _00258_);
  nand (_00280_, _00279_, _00278_);
  nand (_00281_, _00280_, _42618_);
  or (_00282_, \oc8051_gm_cxrom_1.cell7.data [3], _42618_);
  and (_05452_, _00282_, _00281_);
  or (_00283_, word_in[60], \oc8051_gm_cxrom_1.cell7.valid );
  or (_00284_, \oc8051_gm_cxrom_1.cell7.data [4], _00258_);
  nand (_00285_, _00284_, _00283_);
  nand (_00286_, _00285_, _42618_);
  or (_00287_, \oc8051_gm_cxrom_1.cell7.data [4], _42618_);
  and (_05456_, _00287_, _00286_);
  or (_00288_, word_in[61], \oc8051_gm_cxrom_1.cell7.valid );
  or (_00289_, \oc8051_gm_cxrom_1.cell7.data [5], _00258_);
  nand (_00290_, _00289_, _00288_);
  nand (_00291_, _00290_, _42618_);
  or (_00292_, \oc8051_gm_cxrom_1.cell7.data [5], _42618_);
  and (_05460_, _00292_, _00291_);
  or (_00293_, word_in[62], \oc8051_gm_cxrom_1.cell7.valid );
  or (_00294_, \oc8051_gm_cxrom_1.cell7.data [6], _00258_);
  nand (_00295_, _00294_, _00293_);
  nand (_00296_, _00295_, _42618_);
  or (_00297_, \oc8051_gm_cxrom_1.cell7.data [6], _42618_);
  and (_05464_, _00297_, _00296_);
  or (_00298_, \oc8051_gm_cxrom_1.cell8.valid , word_in[71]);
  not (_00299_, \oc8051_gm_cxrom_1.cell8.valid );
  or (_00300_, _00299_, \oc8051_gm_cxrom_1.cell8.data [7]);
  nand (_00301_, _00300_, _00298_);
  nand (_00302_, _00301_, _42618_);
  or (_00303_, \oc8051_gm_cxrom_1.cell8.data [7], _42618_);
  and (_05485_, _00303_, _00302_);
  or (_00304_, word_in[64], \oc8051_gm_cxrom_1.cell8.valid );
  or (_00305_, \oc8051_gm_cxrom_1.cell8.data [0], _00299_);
  nand (_00306_, _00305_, _00304_);
  nand (_00307_, _00306_, _42618_);
  or (_00308_, \oc8051_gm_cxrom_1.cell8.data [0], _42618_);
  and (_05492_, _00308_, _00307_);
  or (_00309_, word_in[65], \oc8051_gm_cxrom_1.cell8.valid );
  or (_00310_, \oc8051_gm_cxrom_1.cell8.data [1], _00299_);
  nand (_00311_, _00310_, _00309_);
  nand (_00312_, _00311_, _42618_);
  or (_00313_, \oc8051_gm_cxrom_1.cell8.data [1], _42618_);
  and (_05496_, _00313_, _00312_);
  or (_00314_, word_in[66], \oc8051_gm_cxrom_1.cell8.valid );
  or (_00315_, \oc8051_gm_cxrom_1.cell8.data [2], _00299_);
  nand (_00316_, _00315_, _00314_);
  nand (_00317_, _00316_, _42618_);
  or (_00318_, \oc8051_gm_cxrom_1.cell8.data [2], _42618_);
  and (_05500_, _00318_, _00317_);
  or (_00319_, word_in[67], \oc8051_gm_cxrom_1.cell8.valid );
  or (_00320_, \oc8051_gm_cxrom_1.cell8.data [3], _00299_);
  nand (_00321_, _00320_, _00319_);
  nand (_00322_, _00321_, _42618_);
  or (_00323_, \oc8051_gm_cxrom_1.cell8.data [3], _42618_);
  and (_05504_, _00323_, _00322_);
  or (_00324_, word_in[68], \oc8051_gm_cxrom_1.cell8.valid );
  or (_00325_, \oc8051_gm_cxrom_1.cell8.data [4], _00299_);
  nand (_00326_, _00325_, _00324_);
  nand (_00327_, _00326_, _42618_);
  or (_00328_, \oc8051_gm_cxrom_1.cell8.data [4], _42618_);
  and (_05508_, _00328_, _00327_);
  or (_00329_, word_in[69], \oc8051_gm_cxrom_1.cell8.valid );
  or (_00330_, \oc8051_gm_cxrom_1.cell8.data [5], _00299_);
  nand (_00331_, _00330_, _00329_);
  nand (_00332_, _00331_, _42618_);
  or (_00333_, \oc8051_gm_cxrom_1.cell8.data [5], _42618_);
  and (_05512_, _00333_, _00332_);
  or (_00334_, word_in[70], \oc8051_gm_cxrom_1.cell8.valid );
  or (_00335_, \oc8051_gm_cxrom_1.cell8.data [6], _00299_);
  nand (_00336_, _00335_, _00334_);
  nand (_00337_, _00336_, _42618_);
  or (_00338_, \oc8051_gm_cxrom_1.cell8.data [6], _42618_);
  and (_05516_, _00338_, _00337_);
  or (_00339_, \oc8051_gm_cxrom_1.cell9.valid , word_in[79]);
  not (_00340_, \oc8051_gm_cxrom_1.cell9.valid );
  or (_00341_, _00340_, \oc8051_gm_cxrom_1.cell9.data [7]);
  nand (_00342_, _00341_, _00339_);
  nand (_00343_, _00342_, _42618_);
  or (_00344_, \oc8051_gm_cxrom_1.cell9.data [7], _42618_);
  and (_05537_, _00344_, _00343_);
  or (_00345_, word_in[72], \oc8051_gm_cxrom_1.cell9.valid );
  or (_00346_, \oc8051_gm_cxrom_1.cell9.data [0], _00340_);
  nand (_00347_, _00346_, _00345_);
  nand (_00348_, _00347_, _42618_);
  or (_00349_, \oc8051_gm_cxrom_1.cell9.data [0], _42618_);
  and (_05544_, _00349_, _00348_);
  or (_00350_, word_in[73], \oc8051_gm_cxrom_1.cell9.valid );
  or (_00351_, \oc8051_gm_cxrom_1.cell9.data [1], _00340_);
  nand (_00352_, _00351_, _00350_);
  nand (_00353_, _00352_, _42618_);
  or (_00354_, \oc8051_gm_cxrom_1.cell9.data [1], _42618_);
  and (_05548_, _00354_, _00353_);
  or (_00355_, word_in[74], \oc8051_gm_cxrom_1.cell9.valid );
  or (_00356_, \oc8051_gm_cxrom_1.cell9.data [2], _00340_);
  nand (_00357_, _00356_, _00355_);
  nand (_00358_, _00357_, _42618_);
  or (_00359_, \oc8051_gm_cxrom_1.cell9.data [2], _42618_);
  and (_05552_, _00359_, _00358_);
  or (_00360_, word_in[75], \oc8051_gm_cxrom_1.cell9.valid );
  or (_00361_, \oc8051_gm_cxrom_1.cell9.data [3], _00340_);
  nand (_00362_, _00361_, _00360_);
  nand (_00363_, _00362_, _42618_);
  or (_00364_, \oc8051_gm_cxrom_1.cell9.data [3], _42618_);
  and (_05555_, _00364_, _00363_);
  or (_00365_, word_in[76], \oc8051_gm_cxrom_1.cell9.valid );
  or (_00366_, \oc8051_gm_cxrom_1.cell9.data [4], _00340_);
  nand (_00367_, _00366_, _00365_);
  nand (_00368_, _00367_, _42618_);
  or (_00369_, \oc8051_gm_cxrom_1.cell9.data [4], _42618_);
  and (_05559_, _00369_, _00368_);
  or (_00370_, word_in[77], \oc8051_gm_cxrom_1.cell9.valid );
  or (_00371_, \oc8051_gm_cxrom_1.cell9.data [5], _00340_);
  nand (_00372_, _00371_, _00370_);
  nand (_00373_, _00372_, _42618_);
  or (_00374_, \oc8051_gm_cxrom_1.cell9.data [5], _42618_);
  and (_05563_, _00374_, _00373_);
  or (_00375_, word_in[78], \oc8051_gm_cxrom_1.cell9.valid );
  or (_00376_, \oc8051_gm_cxrom_1.cell9.data [6], _00340_);
  nand (_00377_, _00376_, _00375_);
  nand (_00378_, _00377_, _42618_);
  or (_00379_, \oc8051_gm_cxrom_1.cell9.data [6], _42618_);
  and (_05567_, _00379_, _00378_);
  or (_00380_, \oc8051_gm_cxrom_1.cell10.valid , word_in[87]);
  not (_00381_, \oc8051_gm_cxrom_1.cell10.valid );
  or (_00382_, _00381_, \oc8051_gm_cxrom_1.cell10.data [7]);
  nand (_00383_, _00382_, _00380_);
  nand (_00384_, _00383_, _42618_);
  or (_00385_, \oc8051_gm_cxrom_1.cell10.data [7], _42618_);
  and (_05589_, _00385_, _00384_);
  or (_00386_, word_in[80], \oc8051_gm_cxrom_1.cell10.valid );
  or (_00387_, \oc8051_gm_cxrom_1.cell10.data [0], _00381_);
  nand (_00388_, _00387_, _00386_);
  nand (_00389_, _00388_, _42618_);
  or (_00390_, \oc8051_gm_cxrom_1.cell10.data [0], _42618_);
  and (_05595_, _00390_, _00389_);
  or (_00391_, word_in[81], \oc8051_gm_cxrom_1.cell10.valid );
  or (_00392_, \oc8051_gm_cxrom_1.cell10.data [1], _00381_);
  nand (_00393_, _00392_, _00391_);
  nand (_00394_, _00393_, _42618_);
  or (_00395_, \oc8051_gm_cxrom_1.cell10.data [1], _42618_);
  and (_05599_, _00395_, _00394_);
  or (_00396_, word_in[82], \oc8051_gm_cxrom_1.cell10.valid );
  or (_00397_, \oc8051_gm_cxrom_1.cell10.data [2], _00381_);
  nand (_00398_, _00397_, _00396_);
  nand (_00399_, _00398_, _42618_);
  or (_00400_, \oc8051_gm_cxrom_1.cell10.data [2], _42618_);
  and (_05603_, _00400_, _00399_);
  or (_00401_, word_in[83], \oc8051_gm_cxrom_1.cell10.valid );
  or (_00402_, \oc8051_gm_cxrom_1.cell10.data [3], _00381_);
  nand (_00403_, _00402_, _00401_);
  nand (_00404_, _00403_, _42618_);
  or (_00405_, \oc8051_gm_cxrom_1.cell10.data [3], _42618_);
  and (_05607_, _00405_, _00404_);
  or (_00406_, word_in[84], \oc8051_gm_cxrom_1.cell10.valid );
  or (_00407_, \oc8051_gm_cxrom_1.cell10.data [4], _00381_);
  nand (_00408_, _00407_, _00406_);
  nand (_00409_, _00408_, _42618_);
  or (_00410_, \oc8051_gm_cxrom_1.cell10.data [4], _42618_);
  and (_05611_, _00410_, _00409_);
  or (_00411_, word_in[85], \oc8051_gm_cxrom_1.cell10.valid );
  or (_00412_, \oc8051_gm_cxrom_1.cell10.data [5], _00381_);
  nand (_00413_, _00412_, _00411_);
  nand (_00414_, _00413_, _42618_);
  or (_00415_, \oc8051_gm_cxrom_1.cell10.data [5], _42618_);
  and (_05615_, _00415_, _00414_);
  or (_00416_, word_in[86], \oc8051_gm_cxrom_1.cell10.valid );
  or (_00417_, \oc8051_gm_cxrom_1.cell10.data [6], _00381_);
  nand (_00418_, _00417_, _00416_);
  nand (_00419_, _00418_, _42618_);
  or (_00420_, \oc8051_gm_cxrom_1.cell10.data [6], _42618_);
  and (_05619_, _00420_, _00419_);
  or (_00421_, \oc8051_gm_cxrom_1.cell11.valid , word_in[95]);
  not (_00422_, \oc8051_gm_cxrom_1.cell11.valid );
  or (_00423_, _00422_, \oc8051_gm_cxrom_1.cell11.data [7]);
  nand (_00424_, _00423_, _00421_);
  nand (_00425_, _00424_, _42618_);
  or (_00426_, \oc8051_gm_cxrom_1.cell11.data [7], _42618_);
  and (_05641_, _00426_, _00425_);
  or (_00427_, word_in[88], \oc8051_gm_cxrom_1.cell11.valid );
  or (_00428_, \oc8051_gm_cxrom_1.cell11.data [0], _00422_);
  nand (_00429_, _00428_, _00427_);
  nand (_00430_, _00429_, _42618_);
  or (_00431_, \oc8051_gm_cxrom_1.cell11.data [0], _42618_);
  and (_05648_, _00431_, _00430_);
  or (_00432_, word_in[89], \oc8051_gm_cxrom_1.cell11.valid );
  or (_00433_, \oc8051_gm_cxrom_1.cell11.data [1], _00422_);
  nand (_00434_, _00433_, _00432_);
  nand (_00435_, _00434_, _42618_);
  or (_00436_, \oc8051_gm_cxrom_1.cell11.data [1], _42618_);
  and (_05652_, _00436_, _00435_);
  or (_00437_, word_in[90], \oc8051_gm_cxrom_1.cell11.valid );
  or (_00438_, \oc8051_gm_cxrom_1.cell11.data [2], _00422_);
  nand (_00439_, _00438_, _00437_);
  nand (_00440_, _00439_, _42618_);
  or (_00441_, \oc8051_gm_cxrom_1.cell11.data [2], _42618_);
  and (_05656_, _00441_, _00440_);
  or (_00442_, word_in[91], \oc8051_gm_cxrom_1.cell11.valid );
  or (_00443_, \oc8051_gm_cxrom_1.cell11.data [3], _00422_);
  nand (_00444_, _00443_, _00442_);
  nand (_00445_, _00444_, _42618_);
  or (_00446_, \oc8051_gm_cxrom_1.cell11.data [3], _42618_);
  and (_05660_, _00446_, _00445_);
  or (_00447_, word_in[92], \oc8051_gm_cxrom_1.cell11.valid );
  or (_00448_, \oc8051_gm_cxrom_1.cell11.data [4], _00422_);
  nand (_00449_, _00448_, _00447_);
  nand (_00450_, _00449_, _42618_);
  or (_00451_, \oc8051_gm_cxrom_1.cell11.data [4], _42618_);
  and (_05664_, _00451_, _00450_);
  or (_00452_, word_in[93], \oc8051_gm_cxrom_1.cell11.valid );
  or (_00453_, \oc8051_gm_cxrom_1.cell11.data [5], _00422_);
  nand (_00454_, _00453_, _00452_);
  nand (_00455_, _00454_, _42618_);
  or (_00456_, \oc8051_gm_cxrom_1.cell11.data [5], _42618_);
  and (_05668_, _00456_, _00455_);
  or (_00457_, word_in[94], \oc8051_gm_cxrom_1.cell11.valid );
  or (_00458_, \oc8051_gm_cxrom_1.cell11.data [6], _00422_);
  nand (_00459_, _00458_, _00457_);
  nand (_00460_, _00459_, _42618_);
  or (_00461_, \oc8051_gm_cxrom_1.cell11.data [6], _42618_);
  and (_05672_, _00461_, _00460_);
  or (_00462_, \oc8051_gm_cxrom_1.cell12.valid , word_in[103]);
  not (_00463_, \oc8051_gm_cxrom_1.cell12.valid );
  or (_00464_, _00463_, \oc8051_gm_cxrom_1.cell12.data [7]);
  nand (_00465_, _00464_, _00462_);
  nand (_00466_, _00465_, _42618_);
  or (_00467_, \oc8051_gm_cxrom_1.cell12.data [7], _42618_);
  and (_05694_, _00467_, _00466_);
  or (_00468_, word_in[96], \oc8051_gm_cxrom_1.cell12.valid );
  or (_00469_, \oc8051_gm_cxrom_1.cell12.data [0], _00463_);
  nand (_00470_, _00469_, _00468_);
  nand (_00471_, _00470_, _42618_);
  or (_00472_, \oc8051_gm_cxrom_1.cell12.data [0], _42618_);
  and (_05701_, _00472_, _00471_);
  or (_00473_, word_in[97], \oc8051_gm_cxrom_1.cell12.valid );
  or (_00474_, \oc8051_gm_cxrom_1.cell12.data [1], _00463_);
  nand (_00475_, _00474_, _00473_);
  nand (_00476_, _00475_, _42618_);
  or (_00477_, \oc8051_gm_cxrom_1.cell12.data [1], _42618_);
  and (_05705_, _00477_, _00476_);
  or (_00478_, word_in[98], \oc8051_gm_cxrom_1.cell12.valid );
  or (_00479_, \oc8051_gm_cxrom_1.cell12.data [2], _00463_);
  nand (_00480_, _00479_, _00478_);
  nand (_00481_, _00480_, _42618_);
  or (_00482_, \oc8051_gm_cxrom_1.cell12.data [2], _42618_);
  and (_05709_, _00482_, _00481_);
  or (_00483_, word_in[99], \oc8051_gm_cxrom_1.cell12.valid );
  or (_00484_, \oc8051_gm_cxrom_1.cell12.data [3], _00463_);
  nand (_00485_, _00484_, _00483_);
  nand (_00486_, _00485_, _42618_);
  or (_00487_, \oc8051_gm_cxrom_1.cell12.data [3], _42618_);
  and (_05713_, _00487_, _00486_);
  or (_00488_, word_in[100], \oc8051_gm_cxrom_1.cell12.valid );
  or (_00489_, \oc8051_gm_cxrom_1.cell12.data [4], _00463_);
  nand (_00490_, _00489_, _00488_);
  nand (_00491_, _00490_, _42618_);
  or (_00492_, \oc8051_gm_cxrom_1.cell12.data [4], _42618_);
  and (_05717_, _00492_, _00491_);
  or (_00493_, word_in[101], \oc8051_gm_cxrom_1.cell12.valid );
  or (_00494_, \oc8051_gm_cxrom_1.cell12.data [5], _00463_);
  nand (_00495_, _00494_, _00493_);
  nand (_00496_, _00495_, _42618_);
  or (_00497_, \oc8051_gm_cxrom_1.cell12.data [5], _42618_);
  and (_05721_, _00497_, _00496_);
  or (_00498_, word_in[102], \oc8051_gm_cxrom_1.cell12.valid );
  or (_00499_, \oc8051_gm_cxrom_1.cell12.data [6], _00463_);
  nand (_00500_, _00499_, _00498_);
  nand (_00501_, _00500_, _42618_);
  or (_00502_, \oc8051_gm_cxrom_1.cell12.data [6], _42618_);
  and (_05725_, _00502_, _00501_);
  or (_00503_, \oc8051_gm_cxrom_1.cell13.valid , word_in[111]);
  not (_00504_, \oc8051_gm_cxrom_1.cell13.valid );
  or (_00505_, _00504_, \oc8051_gm_cxrom_1.cell13.data [7]);
  nand (_00506_, _00505_, _00503_);
  nand (_00507_, _00506_, _42618_);
  or (_00508_, \oc8051_gm_cxrom_1.cell13.data [7], _42618_);
  and (_05747_, _00508_, _00507_);
  or (_00509_, word_in[104], \oc8051_gm_cxrom_1.cell13.valid );
  or (_00510_, \oc8051_gm_cxrom_1.cell13.data [0], _00504_);
  nand (_00511_, _00510_, _00509_);
  nand (_00512_, _00511_, _42618_);
  or (_00513_, \oc8051_gm_cxrom_1.cell13.data [0], _42618_);
  and (_05754_, _00513_, _00512_);
  or (_00514_, word_in[105], \oc8051_gm_cxrom_1.cell13.valid );
  or (_00515_, \oc8051_gm_cxrom_1.cell13.data [1], _00504_);
  nand (_00516_, _00515_, _00514_);
  nand (_00517_, _00516_, _42618_);
  or (_00518_, \oc8051_gm_cxrom_1.cell13.data [1], _42618_);
  and (_05758_, _00518_, _00517_);
  or (_00519_, word_in[106], \oc8051_gm_cxrom_1.cell13.valid );
  or (_00520_, \oc8051_gm_cxrom_1.cell13.data [2], _00504_);
  nand (_00521_, _00520_, _00519_);
  nand (_00522_, _00521_, _42618_);
  or (_00523_, \oc8051_gm_cxrom_1.cell13.data [2], _42618_);
  and (_05762_, _00523_, _00522_);
  or (_00524_, word_in[107], \oc8051_gm_cxrom_1.cell13.valid );
  or (_00525_, \oc8051_gm_cxrom_1.cell13.data [3], _00504_);
  nand (_00526_, _00525_, _00524_);
  nand (_00527_, _00526_, _42618_);
  or (_00528_, \oc8051_gm_cxrom_1.cell13.data [3], _42618_);
  and (_05766_, _00528_, _00527_);
  or (_00529_, word_in[108], \oc8051_gm_cxrom_1.cell13.valid );
  or (_00530_, \oc8051_gm_cxrom_1.cell13.data [4], _00504_);
  nand (_00531_, _00530_, _00529_);
  nand (_00532_, _00531_, _42618_);
  or (_00533_, \oc8051_gm_cxrom_1.cell13.data [4], _42618_);
  and (_05770_, _00533_, _00532_);
  or (_00534_, word_in[109], \oc8051_gm_cxrom_1.cell13.valid );
  or (_00535_, \oc8051_gm_cxrom_1.cell13.data [5], _00504_);
  nand (_00536_, _00535_, _00534_);
  nand (_00537_, _00536_, _42618_);
  or (_00538_, \oc8051_gm_cxrom_1.cell13.data [5], _42618_);
  and (_05774_, _00538_, _00537_);
  or (_00539_, word_in[110], \oc8051_gm_cxrom_1.cell13.valid );
  or (_00540_, \oc8051_gm_cxrom_1.cell13.data [6], _00504_);
  nand (_00541_, _00540_, _00539_);
  nand (_00542_, _00541_, _42618_);
  or (_00544_, \oc8051_gm_cxrom_1.cell13.data [6], _42618_);
  and (_05778_, _00544_, _00542_);
  or (_00546_, \oc8051_gm_cxrom_1.cell14.valid , word_in[119]);
  not (_00547_, \oc8051_gm_cxrom_1.cell14.valid );
  or (_00549_, _00547_, \oc8051_gm_cxrom_1.cell14.data [7]);
  nand (_00550_, _00549_, _00546_);
  nand (_00552_, _00550_, _42618_);
  or (_00553_, \oc8051_gm_cxrom_1.cell14.data [7], _42618_);
  and (_05800_, _00553_, _00552_);
  or (_00555_, word_in[112], \oc8051_gm_cxrom_1.cell14.valid );
  or (_00557_, \oc8051_gm_cxrom_1.cell14.data [0], _00547_);
  nand (_00558_, _00557_, _00555_);
  nand (_00560_, _00558_, _42618_);
  or (_00561_, \oc8051_gm_cxrom_1.cell14.data [0], _42618_);
  and (_05807_, _00561_, _00560_);
  or (_00563_, word_in[113], \oc8051_gm_cxrom_1.cell14.valid );
  or (_00565_, \oc8051_gm_cxrom_1.cell14.data [1], _00547_);
  nand (_00566_, _00565_, _00563_);
  nand (_00568_, _00566_, _42618_);
  or (_00569_, \oc8051_gm_cxrom_1.cell14.data [1], _42618_);
  and (_05811_, _00569_, _00568_);
  or (_00571_, word_in[114], \oc8051_gm_cxrom_1.cell14.valid );
  or (_00573_, \oc8051_gm_cxrom_1.cell14.data [2], _00547_);
  nand (_00574_, _00573_, _00571_);
  nand (_00576_, _00574_, _42618_);
  or (_00577_, \oc8051_gm_cxrom_1.cell14.data [2], _42618_);
  and (_05815_, _00577_, _00576_);
  or (_00579_, word_in[115], \oc8051_gm_cxrom_1.cell14.valid );
  or (_00581_, \oc8051_gm_cxrom_1.cell14.data [3], _00547_);
  nand (_00582_, _00581_, _00579_);
  nand (_00584_, _00582_, _42618_);
  or (_00585_, \oc8051_gm_cxrom_1.cell14.data [3], _42618_);
  and (_05819_, _00585_, _00584_);
  or (_00587_, word_in[116], \oc8051_gm_cxrom_1.cell14.valid );
  or (_00589_, \oc8051_gm_cxrom_1.cell14.data [4], _00547_);
  nand (_00590_, _00589_, _00587_);
  nand (_00592_, _00590_, _42618_);
  or (_00593_, \oc8051_gm_cxrom_1.cell14.data [4], _42618_);
  and (_05823_, _00593_, _00592_);
  or (_00594_, word_in[117], \oc8051_gm_cxrom_1.cell14.valid );
  or (_00595_, \oc8051_gm_cxrom_1.cell14.data [5], _00547_);
  nand (_00596_, _00595_, _00594_);
  nand (_00597_, _00596_, _42618_);
  or (_00598_, \oc8051_gm_cxrom_1.cell14.data [5], _42618_);
  and (_05827_, _00598_, _00597_);
  or (_00599_, word_in[118], \oc8051_gm_cxrom_1.cell14.valid );
  or (_00600_, \oc8051_gm_cxrom_1.cell14.data [6], _00547_);
  nand (_00601_, _00600_, _00599_);
  nand (_00602_, _00601_, _42618_);
  or (_00603_, \oc8051_gm_cxrom_1.cell14.data [6], _42618_);
  and (_05831_, _00603_, _00602_);
  or (_00604_, \oc8051_gm_cxrom_1.cell15.valid , word_in[127]);
  not (_00605_, \oc8051_gm_cxrom_1.cell15.valid );
  or (_00606_, _00605_, \oc8051_gm_cxrom_1.cell15.data [7]);
  nand (_00607_, _00606_, _00604_);
  nand (_00608_, _00607_, _42618_);
  or (_00609_, \oc8051_gm_cxrom_1.cell15.data [7], _42618_);
  and (_05853_, _00609_, _00608_);
  or (_00610_, word_in[120], \oc8051_gm_cxrom_1.cell15.valid );
  or (_00611_, \oc8051_gm_cxrom_1.cell15.data [0], _00605_);
  nand (_00612_, _00611_, _00610_);
  nand (_00613_, _00612_, _42618_);
  or (_00614_, \oc8051_gm_cxrom_1.cell15.data [0], _42618_);
  and (_05860_, _00614_, _00613_);
  or (_00615_, word_in[121], \oc8051_gm_cxrom_1.cell15.valid );
  or (_00616_, \oc8051_gm_cxrom_1.cell15.data [1], _00605_);
  nand (_00617_, _00616_, _00615_);
  nand (_00618_, _00617_, _42618_);
  or (_00619_, \oc8051_gm_cxrom_1.cell15.data [1], _42618_);
  and (_05864_, _00619_, _00618_);
  or (_00620_, word_in[122], \oc8051_gm_cxrom_1.cell15.valid );
  or (_00621_, \oc8051_gm_cxrom_1.cell15.data [2], _00605_);
  nand (_00622_, _00621_, _00620_);
  nand (_00623_, _00622_, _42618_);
  or (_00624_, \oc8051_gm_cxrom_1.cell15.data [2], _42618_);
  and (_05868_, _00624_, _00623_);
  or (_00625_, word_in[123], \oc8051_gm_cxrom_1.cell15.valid );
  or (_00626_, \oc8051_gm_cxrom_1.cell15.data [3], _00605_);
  nand (_00627_, _00626_, _00625_);
  nand (_00628_, _00627_, _42618_);
  or (_00629_, \oc8051_gm_cxrom_1.cell15.data [3], _42618_);
  and (_05872_, _00629_, _00628_);
  or (_00630_, word_in[124], \oc8051_gm_cxrom_1.cell15.valid );
  or (_00631_, \oc8051_gm_cxrom_1.cell15.data [4], _00605_);
  nand (_00632_, _00631_, _00630_);
  nand (_00633_, _00632_, _42618_);
  or (_00634_, \oc8051_gm_cxrom_1.cell15.data [4], _42618_);
  and (_05876_, _00634_, _00633_);
  or (_00635_, word_in[125], \oc8051_gm_cxrom_1.cell15.valid );
  or (_00636_, \oc8051_gm_cxrom_1.cell15.data [5], _00605_);
  nand (_00637_, _00636_, _00635_);
  nand (_00638_, _00637_, _42618_);
  or (_00639_, \oc8051_gm_cxrom_1.cell15.data [5], _42618_);
  and (_05880_, _00639_, _00638_);
  or (_00640_, word_in[126], \oc8051_gm_cxrom_1.cell15.valid );
  or (_00641_, \oc8051_gm_cxrom_1.cell15.data [6], _00605_);
  nand (_00642_, _00641_, _00640_);
  nand (_00643_, _00642_, _42618_);
  or (_00644_, \oc8051_gm_cxrom_1.cell15.data [6], _42618_);
  and (_05884_, _00644_, _00643_);
  nor (_09659_, _37997_, rst);
  and (_00645_, _38048_, _37987_);
  and (_00646_, _00645_, _37890_);
  not (_00647_, _00646_);
  and (_00648_, _37970_, _37866_);
  and (_00649_, _38049_, _38005_);
  nor (_00650_, _00649_, _00648_);
  and (_00651_, _00650_, _00647_);
  and (_00652_, _38048_, _37889_);
  or (_00653_, _37987_, _38005_);
  nand (_00654_, _00653_, _00652_);
  and (_00655_, _00654_, _00651_);
  and (_00656_, _36958_, _42618_);
  not (_00657_, _00656_);
  or (_00658_, _00657_, _00648_);
  or (_09662_, _00658_, _00655_);
  not (_00659_, _37858_);
  and (_00660_, _00659_, _37602_);
  and (_00661_, _37832_, _37330_);
  and (_00662_, _00661_, _00660_);
  not (_00663_, _37954_);
  and (_00664_, _00663_, _37931_);
  and (_00665_, _00664_, _37884_);
  and (_00666_, _00665_, _00662_);
  nor (_00667_, _37858_, _37832_);
  and (_00668_, _00667_, _37330_);
  and (_00669_, _00668_, _37602_);
  not (_00670_, _37884_);
  nor (_00671_, _00663_, _37931_);
  and (_00672_, _00671_, _00670_);
  and (_00673_, _00672_, _00669_);
  and (_00674_, _37908_, _37884_);
  nor (_00675_, _37954_, _37931_);
  and (_00676_, _00675_, _00674_);
  not (_00677_, _37602_);
  and (_00678_, _00668_, _00677_);
  and (_00679_, _00678_, _00676_);
  or (_00680_, _00679_, _00673_);
  or (_00681_, _00680_, _00666_);
  nor (_00682_, _37908_, _00670_);
  and (_00683_, _00671_, _00682_);
  and (_00684_, _00683_, _00668_);
  and (_00685_, _37858_, _37832_);
  and (_00686_, _37330_, _37602_);
  and (_00687_, _00686_, _00685_);
  not (_00688_, _00674_);
  and (_00689_, _37954_, _37931_);
  and (_00690_, _00689_, _00688_);
  and (_00691_, _00690_, _00687_);
  or (_00692_, _00691_, _00684_);
  and (_00693_, _00671_, _37908_);
  and (_00694_, _00685_, _37330_);
  and (_00695_, _00694_, _00677_);
  and (_00696_, _00695_, _00693_);
  not (_00697_, _37330_);
  and (_00698_, _00676_, _00697_);
  or (_00699_, _00698_, _00696_);
  or (_00700_, _00699_, _00692_);
  and (_00701_, _00682_, _00664_);
  and (_00702_, _00695_, _00701_);
  and (_00703_, _37908_, _00670_);
  and (_00704_, _00703_, _00671_);
  and (_00705_, _00704_, _00662_);
  or (_00706_, _00705_, _00702_);
  nor (_00707_, _00659_, _37832_);
  nor (_00708_, _00707_, _00697_);
  not (_00709_, _00708_);
  and (_00710_, _00709_, _00683_);
  not (_00711_, _37908_);
  and (_00712_, _00675_, _00711_);
  and (_00713_, _00712_, _00662_);
  or (_00714_, _00713_, _00710_);
  or (_00715_, _00714_, _00706_);
  or (_00716_, _00715_, _00700_);
  or (_00717_, _00716_, _00681_);
  nor (_00718_, _37908_, _37884_);
  and (_00719_, _00718_, _00664_);
  nor (_00720_, _00719_, _00677_);
  and (_00721_, _00661_, _00659_);
  not (_00722_, _00721_);
  nor (_00723_, _00722_, _00720_);
  not (_00724_, _00723_);
  and (_00725_, _00703_, _00664_);
  and (_00726_, _00725_, _00662_);
  and (_00727_, _00689_, _00682_);
  and (_00728_, _00727_, _00662_);
  nor (_00729_, _00728_, _00726_);
  and (_00730_, _00729_, _00724_);
  and (_00731_, _00712_, _00694_);
  not (_00732_, _00662_);
  and (_00733_, _00689_, _00674_);
  and (_00734_, _00689_, _00718_);
  nor (_00735_, _00734_, _00733_);
  nor (_00736_, _00735_, _00732_);
  and (_00737_, _00733_, _00687_);
  or (_00738_, _00737_, _00736_);
  nor (_00739_, _00738_, _00731_);
  nand (_00740_, _00739_, _00730_);
  or (_00741_, _00740_, _00717_);
  and (_00742_, _00741_, _36969_);
  not (_00743_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_00744_, _36947_, _18772_);
  and (_00745_, _00744_, _37988_);
  nor (_00746_, _00745_, _00743_);
  or (_00747_, _00746_, rst);
  or (_09665_, _00747_, _00742_);
  nand (_00748_, _37931_, _36893_);
  or (_00749_, _36893_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and (_00750_, _00749_, _42618_);
  and (_09668_, _00750_, _00748_);
  and (_00751_, \oc8051_top_1.oc8051_sfr1.wait_data , _42618_);
  and (_00752_, _00751_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  or (_00753_, _38034_, _38007_);
  and (_00754_, _37866_, _38003_);
  or (_00755_, _00754_, _00753_);
  and (_00756_, _37978_, _38049_);
  and (_00757_, _00648_, _37890_);
  or (_00758_, _00757_, _00756_);
  and (_00759_, _37985_, _37987_);
  and (_00760_, _37975_, _37987_);
  or (_00761_, _00760_, _00759_);
  or (_00762_, _00761_, _00758_);
  nor (_00763_, _00762_, _00755_);
  nand (_00764_, _00763_, _38045_);
  and (_00765_, _00764_, _00656_);
  or (_09671_, _00765_, _00752_);
  and (_00766_, _37971_, _37987_);
  or (_00767_, _00766_, _37963_);
  and (_00768_, _37395_, _37890_);
  and (_00769_, _00768_, _38002_);
  or (_00770_, _00769_, _38112_);
  and (_00771_, _37977_, _38013_);
  and (_00772_, _00771_, _38003_);
  or (_00773_, _00772_, _00770_);
  or (_00774_, _00773_, _00767_);
  and (_00775_, _00774_, _36958_);
  and (_00776_, _38092_, _00743_);
  not (_00777_, _37981_);
  and (_00778_, _00777_, _00776_);
  and (_00779_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_00780_, _00779_, _00778_);
  or (_00781_, _00780_, _00775_);
  and (_09674_, _00781_, _42618_);
  and (_00782_, _00751_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and (_00783_, _37978_, _38046_);
  or (_00784_, _38046_, _38020_);
  and (_00785_, _00784_, _38015_);
  or (_00786_, _00785_, _00783_);
  and (_00787_, _00771_, _38024_);
  or (_00788_, _00787_, _00786_);
  not (_00789_, _38105_);
  and (_00790_, _00784_, _37395_);
  and (_00791_, _37395_, _37889_);
  and (_00792_, _00791_, _38023_);
  or (_00793_, _00792_, _00790_);
  or (_00794_, _00793_, _00789_);
  not (_00795_, _38084_);
  and (_00796_, _37978_, _00795_);
  and (_00797_, _38008_, _37395_);
  or (_00798_, _00797_, _00767_);
  or (_00799_, _00798_, _00796_);
  or (_00800_, _00799_, _00794_);
  or (_00801_, _00800_, _00788_);
  and (_00802_, _00801_, _00656_);
  or (_09677_, _00802_, _00782_);
  and (_00803_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_00804_, _38081_, _36958_);
  or (_00805_, _00804_, _00803_);
  or (_00806_, _00805_, _00778_);
  and (_09680_, _00806_, _42618_);
  and (_00807_, _38024_, _38006_);
  and (_00808_, _38014_, _37986_);
  and (_00809_, _00808_, _37889_);
  or (_00810_, _00809_, _00807_);
  or (_00811_, _00810_, _00757_);
  and (_00812_, _00810_, _37990_);
  or (_00813_, _00812_, _36903_);
  and (_00814_, _00813_, _00811_);
  not (_00815_, _00651_);
  and (_00816_, _00815_, _00776_);
  or (_00817_, _00816_, \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_00818_, _00817_, _00814_);
  or (_00819_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2], _18772_);
  and (_00820_, _00819_, _42618_);
  and (_09683_, _00820_, _00818_);
  and (_00821_, _00751_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  or (_00822_, _00769_, _38066_);
  and (_00823_, _00791_, _38002_);
  or (_00824_, _00792_, _00823_);
  or (_00825_, _37963_, _38021_);
  or (_00826_, _00825_, _00824_);
  or (_00827_, _00826_, _00822_);
  and (_00828_, _38052_, _38003_);
  and (_00829_, _38102_, _38023_);
  or (_00830_, _00787_, _00829_);
  or (_00831_, _00830_, _00828_);
  or (_00832_, _38034_, _38033_);
  or (_00833_, _00832_, _38010_);
  or (_00834_, _00833_, _00831_);
  or (_00835_, _00834_, _00827_);
  and (_00836_, _00835_, _00656_);
  or (_09686_, _00836_, _00821_);
  and (_00837_, _00751_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and (_00838_, _00771_, _38064_);
  and (_00839_, _37866_, _38022_);
  or (_00840_, _00839_, _00772_);
  or (_00841_, _00840_, _00838_);
  or (_00842_, _00841_, _00793_);
  not (_00843_, _38029_);
  and (_00844_, _37978_, _38017_);
  or (_00845_, _00844_, _00843_);
  and (_00846_, _38053_, _38001_);
  or (_00847_, _00846_, _38118_);
  and (_00848_, _38052_, _38020_);
  or (_00849_, _00848_, _00847_);
  or (_00850_, _00849_, _00845_);
  or (_00851_, _00850_, _00842_);
  and (_00852_, _00768_, _38001_);
  and (_00853_, _00768_, _37966_);
  or (_00854_, _00853_, _00852_);
  nor (_00855_, _38104_, _38069_);
  nand (_00856_, _00855_, _38019_);
  or (_00857_, _00856_, _00854_);
  or (_00858_, _00857_, _00788_);
  or (_00859_, _00858_, _00851_);
  and (_00860_, _00859_, _00656_);
  or (_09689_, _00860_, _00837_);
  and (_00861_, _37971_, _37395_);
  or (_00862_, _00861_, _38110_);
  and (_00863_, _37971_, _38052_);
  and (_00864_, _38037_, _37395_);
  and (_00865_, _00771_, _38037_);
  or (_00866_, _00865_, _00864_);
  or (_00867_, _00866_, _00863_);
  or (_00868_, _00867_, _00862_);
  and (_00869_, _00771_, _37971_);
  or (_00870_, _00869_, _00868_);
  and (_00871_, _00870_, _36958_);
  and (_00872_, \oc8051_top_1.oc8051_sfr1.wait_data , \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or (_00873_, _00872_, _37994_);
  or (_00874_, _00873_, _00871_);
  and (_09692_, _00874_, _42618_);
  nand (_00875_, _38082_, _38070_);
  or (_00876_, _00875_, _00785_);
  or (_00877_, _38066_, _38035_);
  and (_00878_, _37965_, _37889_);
  and (_00879_, _00878_, _38015_);
  nor (_00880_, _00879_, _38028_);
  nor (_00881_, _00807_, _38025_);
  and (_00882_, _00881_, _00880_);
  nand (_00883_, _00882_, _38011_);
  or (_00884_, _00883_, _00877_);
  or (_00885_, _00884_, _00876_);
  and (_00886_, _00791_, _37965_);
  or (_00887_, _00886_, _38077_);
  and (_00888_, _00768_, _37970_);
  or (_00889_, _00888_, _00809_);
  or (_00890_, _00889_, _00770_);
  or (_00891_, _00890_, _00887_);
  and (_00892_, _00878_, _38052_);
  or (_00893_, _00892_, _38104_);
  or (_00894_, _00893_, _38054_);
  or (_00895_, _38106_, _38074_);
  or (_00896_, _00895_, _00894_);
  or (_00897_, _00896_, _00891_);
  or (_00898_, _00897_, _00793_);
  or (_00899_, _00898_, _00885_);
  and (_00900_, _00899_, _36958_);
  and (_00901_, \oc8051_top_1.oc8051_decoder1.wr , \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_00902_, _00812_, _00778_);
  and (_00903_, _37990_, _38043_);
  or (_00904_, _00903_, _00902_);
  or (_00905_, _00904_, _00901_);
  or (_00906_, _00905_, _00900_);
  and (_09695_, _00906_, _42618_);
  nor (_09754_, _38131_, rst);
  nor (_09756_, _38097_, rst);
  or (_09759_, _00657_, _00651_);
  nor (_00907_, _00648_, _00645_);
  or (_09762_, _00907_, _00657_);
  and (_00908_, _00689_, _00711_);
  and (_00909_, _00908_, _00687_);
  or (_00910_, _00909_, _00673_);
  or (_00911_, _00696_, \oc8051_top_1.oc8051_decoder1.state [1]);
  or (_00912_, _00911_, _00910_);
  and (_00913_, _00912_, _00745_);
  nor (_00914_, _00744_, _37988_);
  or (_00915_, _00914_, rst);
  or (_09765_, _00915_, _00913_);
  nand (_00916_, _37602_, _36893_);
  or (_00917_, _36893_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and (_00918_, _00917_, _42618_);
  and (_09768_, _00918_, _00916_);
  or (_00919_, _37858_, _37993_);
  or (_00920_, _36893_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and (_00921_, _00920_, _42618_);
  and (_09771_, _00921_, _00919_);
  nand (_00922_, _37832_, _36893_);
  or (_00923_, _36893_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and (_00924_, _00923_, _42618_);
  and (_09774_, _00924_, _00922_);
  nand (_00926_, _37330_, _36893_);
  or (_00927_, _36893_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and (_00928_, _00927_, _42618_);
  and (_09777_, _00928_, _00926_);
  or (_00929_, _37884_, _37993_);
  or (_00930_, _36893_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and (_00931_, _00930_, _42618_);
  and (_09780_, _00931_, _00929_);
  nand (_00932_, _37908_, _36893_);
  or (_00933_, _36893_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and (_00934_, _00933_, _42618_);
  and (_09783_, _00934_, _00932_);
  nand (_00935_, _37954_, _36893_);
  or (_00936_, _36893_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and (_00937_, _00936_, _42618_);
  and (_09786_, _00937_, _00935_);
  or (_00938_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], _18772_);
  and (_00939_, _00938_, _42618_);
  and (_00940_, _00939_, _00817_);
  not (_00941_, _38061_);
  and (_00942_, _00771_, _00941_);
  and (_00943_, _00771_, _38017_);
  or (_00944_, _00943_, _00766_);
  or (_00945_, _00771_, _37395_);
  or (_00946_, _38064_, _38049_);
  and (_00947_, _00946_, _00945_);
  or (_00948_, _00947_, _00944_);
  or (_00949_, _00948_, _00942_);
  or (_00950_, _38123_, _00863_);
  and (_00952_, _38060_, _38052_);
  or (_00953_, _00952_, _38118_);
  or (_00954_, _00953_, _00950_);
  and (_00955_, _00768_, _38016_);
  or (_00956_, _00955_, _00839_);
  or (_00957_, _00956_, _37963_);
  or (_00958_, _00957_, _00862_);
  or (_00959_, _00958_, _00954_);
  nor (_00960_, _38061_, _37406_);
  or (_00961_, _00960_, _00869_);
  or (_00962_, _38023_, _38020_);
  or (_00963_, _00962_, _00878_);
  and (_00964_, _00963_, _37978_);
  or (_00965_, _00964_, _00961_);
  or (_00966_, _00965_, _00959_);
  or (_00967_, _00966_, _00949_);
  and (_00968_, _00967_, _00656_);
  or (_09789_, _00968_, _00940_);
  and (_00969_, _00751_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  or (_00970_, _38064_, _38017_);
  and (_00972_, _00970_, _38006_);
  and (_00973_, _00791_, _37961_);
  nor (_00974_, _00973_, _38103_);
  nand (_00975_, _37978_, _00941_);
  nand (_00976_, _00975_, _00974_);
  or (_00977_, _00976_, _00972_);
  or (_00978_, _00796_, _00758_);
  or (_00979_, _00944_, _00854_);
  or (_00980_, _00979_, _00978_);
  not (_00981_, _38067_);
  and (_00982_, _37978_, _38064_);
  or (_00983_, _00982_, _00981_);
  or (_00984_, _00983_, _00849_);
  or (_00985_, _00984_, _00980_);
  or (_00986_, _00985_, _00977_);
  and (_00987_, _00986_, _00656_);
  or (_34182_, _00987_, _00969_);
  or (_00988_, _00895_, _00889_);
  or (_00989_, _00988_, _00885_);
  and (_00990_, _00989_, _36958_);
  and (_00991_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_00992_, _00991_, _00904_);
  or (_00993_, _00992_, _00990_);
  and (_34184_, _00993_, _42618_);
  and (_00994_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_00995_, _00994_, _00902_);
  and (_00996_, _00995_, _42618_);
  and (_00997_, _38068_, _37890_);
  or (_00998_, _00997_, _38112_);
  or (_00999_, _00998_, _00810_);
  or (_01000_, _00999_, _00894_);
  and (_01001_, _01000_, _00656_);
  or (_34187_, _01001_, _00996_);
  or (_01002_, _00648_, _37980_);
  and (_01003_, _00771_, _38060_);
  and (_01004_, _00865_, _37889_);
  or (_01005_, _01004_, _01003_);
  or (_01006_, _01005_, _01002_);
  or (_01007_, _00861_, _38111_);
  and (_01008_, _00652_, _38015_);
  and (_01009_, _37978_, _37967_);
  and (_01010_, _38060_, _38006_);
  or (_01011_, _01010_, _01009_);
  or (_01012_, _01011_, _01008_);
  or (_01013_, _01012_, _01007_);
  or (_01014_, _01013_, _01006_);
  and (_01015_, _00771_, _38008_);
  or (_01016_, _01015_, _00756_);
  and (_01017_, _00652_, _37978_);
  or (_01018_, _01017_, _37979_);
  or (_01019_, _01018_, _01016_);
  and (_01020_, _00962_, _37978_);
  or (_01021_, _01020_, _01019_);
  and (_01022_, _37978_, _38003_);
  or (_01023_, _00839_, _01022_);
  or (_01024_, _01023_, _00961_);
  or (_01025_, _00844_, _00863_);
  and (_01026_, _00865_, _37890_);
  or (_01027_, _01026_, _00982_);
  or (_01028_, _01027_, _01025_);
  or (_01029_, _00892_, _00886_);
  or (_01030_, _01029_, _37968_);
  or (_01031_, _01030_, _00810_);
  or (_01032_, _01031_, _01028_);
  or (_01033_, _01032_, _01024_);
  or (_01034_, _01033_, _01021_);
  or (_01035_, _01034_, _01014_);
  and (_01036_, _01035_, _36958_);
  and (_01037_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_01038_, _00816_, _37995_);
  or (_01039_, _01038_, _01037_);
  or (_01040_, _01039_, _01036_);
  and (_34189_, _01040_, _42618_);
  and (_01041_, _00791_, _38048_);
  or (_01042_, _01041_, _00879_);
  nor (_01043_, _01042_, _00863_);
  nand (_01044_, _01043_, _37973_);
  and (_01045_, _00970_, _37866_);
  or (_01046_, _01045_, _38062_);
  or (_01047_, _01046_, _01044_);
  or (_01048_, _37980_, _38074_);
  and (_01049_, _00652_, _38052_);
  or (_01050_, _01049_, _00766_);
  or (_01051_, _01050_, _01048_);
  or (_01052_, _01051_, _01007_);
  or (_01053_, _01052_, _01047_);
  or (_01054_, _01024_, _01021_);
  or (_01055_, _01054_, _01053_);
  and (_01056_, _01055_, _36958_);
  and (_01057_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_01058_, _01057_, _01038_);
  or (_01059_, _01058_, _01056_);
  and (_34191_, _01059_, _42618_);
  and (_01060_, _00751_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  or (_01061_, _00828_, _00829_);
  or (_01062_, _01061_, _01004_);
  nor (_01063_, _00863_, _38080_);
  nand (_01064_, _01063_, _42104_);
  or (_01065_, _01064_, _01062_);
  not (_01066_, _42102_);
  or (_01067_, _00869_, _01066_);
  or (_01068_, _01067_, _00877_);
  or (_01069_, _01068_, _01065_);
  or (_01070_, _00861_, _00769_);
  or (_01071_, _38051_, _37395_);
  or (_01072_, _01071_, _37866_);
  and (_01073_, _01072_, _38038_);
  and (_01074_, _38009_, _37657_);
  or (_01075_, _01074_, _01073_);
  or (_01076_, _01075_, _01070_);
  or (_01077_, _38024_, _38020_);
  and (_01078_, _01077_, _37866_);
  and (_01079_, _37978_, _38020_);
  or (_01080_, _01079_, _00787_);
  or (_01081_, _01080_, _01078_);
  or (_01082_, _01081_, _00826_);
  or (_01083_, _01082_, _01076_);
  or (_01084_, _01083_, _01069_);
  and (_01085_, _01084_, _00656_);
  or (_34193_, _01085_, _01060_);
  and (_01086_, _00751_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_01087_, _37866_, _38024_);
  or (_01088_, _01026_, _00848_);
  or (_01089_, _01088_, _01087_);
  or (_01090_, _01089_, _00845_);
  or (_01091_, _01090_, _01006_);
  and (_01092_, _38038_, _37866_);
  or (_01093_, _01092_, _01079_);
  not (_01094_, _38075_);
  or (_01095_, _00960_, _01094_);
  or (_01096_, _01095_, _01093_);
  or (_01097_, _37968_, _38018_);
  or (_01098_, _00846_, _00772_);
  or (_01099_, _01098_, _01097_);
  or (_01100_, _00852_, _36914_);
  or (_01101_, _01100_, _37963_);
  or (_01102_, _01101_, _38111_);
  or (_01103_, _01102_, _01099_);
  or (_01104_, _01103_, _01096_);
  or (_01105_, _01104_, _01091_);
  or (_01106_, _37980_, _36903_);
  nor (_01107_, \oc8051_top_1.oc8051_sfr1.wait_data , rst);
  and (_01108_, _01107_, _01106_);
  and (_01109_, _01108_, _01105_);
  or (_34195_, _01109_, _01086_);
  and (_01110_, _00751_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  not (_01111_, _01003_);
  and (_01112_, _01111_, _38075_);
  and (_01113_, _38060_, _37395_);
  or (_01114_, _01113_, _00869_);
  or (_01115_, _01114_, _00952_);
  nor (_01116_, _01115_, _00786_);
  nand (_01117_, _01116_, _01112_);
  or (_01118_, _01017_, _38009_);
  or (_01119_, _01070_, _01016_);
  or (_01120_, _01119_, _01118_);
  or (_01121_, _00772_, _42103_);
  or (_01122_, _00797_, _00787_);
  or (_01123_, _01122_, _01121_);
  and (_01124_, _38037_, _37866_);
  or (_01125_, _01124_, _37980_);
  or (_01126_, _01125_, _38115_);
  or (_01127_, _01126_, _01123_);
  or (_01128_, _01127_, _01120_);
  or (_01129_, _01128_, _00794_);
  or (_01130_, _01129_, _01117_);
  and (_01131_, _01130_, _01108_);
  or (_34197_, _01131_, _01110_);
  or (_01132_, _01080_, _00822_);
  or (_01133_, _01132_, _01118_);
  and (_01134_, _01071_, _38060_);
  or (_01135_, _01003_, _38074_);
  or (_01136_, _01135_, _01134_);
  and (_01137_, _37866_, _38023_);
  or (_01138_, _38112_, _38104_);
  nor (_01139_, _01138_, _01137_);
  nand (_01140_, _01139_, _42102_);
  or (_01141_, _01140_, _01136_);
  or (_01142_, _00793_, _00786_);
  or (_01143_, _01142_, _01141_);
  or (_01144_, _01143_, _01133_);
  and (_01145_, _01144_, _36958_);
  and (_01146_, \oc8051_top_1.oc8051_decoder1.alu_op [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_01147_, _37979_, _18772_);
  or (_01148_, _01147_, _01146_);
  or (_01149_, _01148_, _01145_);
  and (_34199_, _01149_, _42618_);
  and (_01150_, _00751_, \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  or (_01151_, _01078_, _42105_);
  or (_01152_, _01093_, _01074_);
  or (_01153_, _01152_, _01151_);
  or (_01154_, _00754_, _38033_);
  not (_01155_, _37986_);
  and (_01156_, _38008_, _01155_);
  or (_01157_, _01156_, _01154_);
  or (_01158_, _01157_, _00868_);
  or (_01159_, _01158_, _01067_);
  or (_01160_, _01159_, _01153_);
  and (_01161_, _01160_, _00656_);
  or (_34201_, _01161_, _01150_);
  nor (_38643_, _37931_, rst);
  nor (_38644_, _42095_, rst);
  and (_01162_, _42079_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [7]);
  and (_01163_, _37012_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  and (_01164_, _37210_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and (_01165_, _37177_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor (_01166_, _01165_, _01164_);
  and (_01167_, _37078_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_01168_, _37045_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_01169_, _01168_, _01167_);
  and (_01170_, _37232_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_01171_, _37133_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor (_01172_, _01171_, _01170_);
  and (_01173_, _01172_, _01169_);
  and (_01174_, _01173_, _01166_);
  nor (_01175_, _01174_, _37012_);
  nor (_01176_, _01175_, _01163_);
  nor (_01177_, _01176_, _42079_);
  nor (_01178_, _01177_, _01162_);
  nor (_38646_, _01178_, rst);
  nor (_38656_, _37602_, rst);
  and (_38658_, _37858_, _42618_);
  nor (_38659_, _37832_, rst);
  nor (_38660_, _37330_, rst);
  and (_38661_, _37884_, _42618_);
  nor (_38662_, _37908_, rst);
  nor (_38663_, _37954_, rst);
  nor (_38664_, _42391_, rst);
  nor (_38665_, _42298_, rst);
  nor (_38667_, _42207_, rst);
  nor (_38668_, _42349_, rst);
  nor (_38669_, _42253_, rst);
  nor (_38670_, _42131_, rst);
  nor (_38671_, _42446_, rst);
  and (_01179_, _42079_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [0]);
  and (_01180_, _37012_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  and (_01181_, _37232_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_01182_, _37045_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_01183_, _01182_, _01181_);
  and (_01184_, _37210_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and (_01185_, _37133_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor (_01186_, _01185_, _01184_);
  and (_01187_, _37177_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  and (_01188_, _37078_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nor (_01189_, _01188_, _01187_);
  and (_01190_, _01189_, _01186_);
  and (_01191_, _01190_, _01183_);
  nor (_01192_, _01191_, _37012_);
  nor (_01193_, _01192_, _01180_);
  nor (_01194_, _01193_, _42079_);
  nor (_01195_, _01194_, _01179_);
  nor (_38673_, _01195_, rst);
  and (_01196_, _42079_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [1]);
  and (_01197_, _37012_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  and (_01198_, _37078_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_01199_, _37177_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_01200_, _01199_, _01198_);
  and (_01201_, _37232_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_01202_, _37133_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nor (_01203_, _01202_, _01201_);
  and (_01204_, _01203_, _01200_);
  and (_01205_, _37210_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and (_01207_, _37045_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_01209_, _01207_, _01205_);
  and (_01211_, _01209_, _01204_);
  nor (_01213_, _01211_, _37012_);
  nor (_01215_, _01213_, _01197_);
  nor (_01217_, _01215_, _42079_);
  nor (_01219_, _01217_, _01196_);
  nor (_38674_, _01219_, rst);
  and (_01222_, _42079_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [2]);
  and (_01224_, _37012_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  and (_01226_, _37078_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_01228_, _37177_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_01230_, _01228_, _01226_);
  and (_01232_, _37232_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_01234_, _37133_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor (_01236_, _01234_, _01232_);
  and (_01238_, _01236_, _01230_);
  and (_01240_, _37210_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and (_01242_, _37045_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_01244_, _01242_, _01240_);
  and (_01246_, _01244_, _01238_);
  nor (_01248_, _01246_, _37012_);
  nor (_01250_, _01248_, _01224_);
  nor (_01252_, _01250_, _42079_);
  nor (_01254_, _01252_, _01222_);
  nor (_38675_, _01254_, rst);
  and (_01257_, _42079_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [3]);
  and (_01259_, _37012_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  and (_01261_, _37210_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and (_01263_, _37177_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_01265_, _01263_, _01261_);
  and (_01267_, _37078_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_01269_, _37045_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_01271_, _01269_, _01267_);
  and (_01273_, _37232_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_01275_, _37133_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor (_01277_, _01275_, _01273_);
  and (_01279_, _01277_, _01271_);
  and (_01281_, _01279_, _01265_);
  nor (_01283_, _01281_, _37012_);
  nor (_01285_, _01283_, _01259_);
  nor (_01287_, _01285_, _42079_);
  nor (_01289_, _01287_, _01257_);
  nor (_38676_, _01289_, rst);
  and (_01292_, _42079_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [4]);
  and (_01294_, _37012_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  and (_01296_, _37078_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_01298_, _37177_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_01300_, _01298_, _01296_);
  and (_01301_, _37232_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_01302_, _37133_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor (_01303_, _01302_, _01301_);
  and (_01304_, _01303_, _01300_);
  and (_01305_, _37210_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and (_01306_, _37045_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_01307_, _01306_, _01305_);
  and (_01308_, _01307_, _01304_);
  nor (_01309_, _01308_, _37012_);
  nor (_01310_, _01309_, _01294_);
  nor (_01311_, _01310_, _42079_);
  nor (_01312_, _01311_, _01292_);
  nor (_38677_, _01312_, rst);
  and (_01313_, _42079_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [5]);
  and (_01314_, _37012_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  and (_01315_, _37078_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_01316_, _37177_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_01317_, _01316_, _01315_);
  and (_01318_, _37232_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_01319_, _37133_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor (_01320_, _01319_, _01318_);
  and (_01321_, _01320_, _01317_);
  and (_01322_, _37210_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and (_01323_, _37045_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_01324_, _01323_, _01322_);
  and (_01325_, _01324_, _01321_);
  nor (_01326_, _01325_, _37012_);
  nor (_01327_, _01326_, _01314_);
  nor (_01328_, _01327_, _42079_);
  nor (_01329_, _01328_, _01313_);
  nor (_38679_, _01329_, rst);
  and (_01330_, _42079_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [6]);
  and (_01331_, _37012_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  and (_01332_, _37232_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_01333_, _37045_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_01334_, _01333_, _01332_);
  and (_01335_, _37210_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and (_01336_, _37133_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor (_01337_, _01336_, _01335_);
  and (_01338_, _37177_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  and (_01339_, _37078_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nor (_01340_, _01339_, _01338_);
  and (_01341_, _01340_, _01337_);
  and (_01342_, _01341_, _01334_);
  nor (_01343_, _01342_, _37012_);
  nor (_01344_, _01343_, _01331_);
  nor (_01345_, _01344_, _42079_);
  nor (_01346_, _01345_, _01330_);
  nor (_38680_, _01346_, rst);
  and (_01347_, _36969_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  or (_01348_, _01347_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nand (_01349_, _01347_, _38317_);
  and (_01350_, _01349_, _42618_);
  and (_38705_, _01350_, _01348_);
  not (_01351_, _01347_);
  or (_01352_, _01351_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  and (_01353_, _36969_, _42618_);
  and (_01354_, _01353_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  and (_01355_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _42618_);
  or (_01356_, _01355_, _01354_);
  and (_38706_, _01356_, _01352_);
  nor (_38741_, _42100_, rst);
  nor (_38744_, _42072_, rst);
  nor (_01357_, _42354_, _27948_);
  and (_01358_, _42354_, _27948_);
  nor (_01359_, _01358_, _01357_);
  not (_01360_, _01359_);
  nor (_01361_, _42451_, _28376_);
  and (_01362_, _42451_, _28376_);
  nor (_01363_, _01362_, _01361_);
  not (_01364_, _01363_);
  and (_01365_, _01364_, _42548_);
  nor (_01366_, _42259_, _27542_);
  and (_01367_, _42259_, _27542_);
  nor (_01368_, _01367_, _01366_);
  nor (_01369_, _42164_, _27345_);
  and (_01370_, _42164_, _27345_);
  nor (_01371_, _01370_, _01369_);
  nor (_01372_, _01371_, _01368_);
  and (_01373_, _01372_, _01365_);
  and (_01374_, _01373_, _01360_);
  nor (_01375_, _42307_, _33107_);
  and (_01376_, _42307_, _33107_);
  or (_01377_, _01376_, _01375_);
  nor (_01378_, _01377_, _38947_);
  nor (_01379_, _42400_, _27795_);
  and (_01380_, _42400_, _27795_);
  nor (_01381_, _01380_, _01379_);
  nor (_01382_, _42212_, _28069_);
  and (_01383_, _42212_, _28069_);
  nor (_01384_, _01383_, _01382_);
  nor (_01385_, _01384_, _01381_);
  and (_01386_, _01385_, _01378_);
  and (_01387_, _01386_, _01374_);
  nor (_01388_, _28244_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_01389_, _01388_, _01387_);
  not (_01390_, _01389_);
  nor (_01391_, _38045_, _38092_);
  nor (_01392_, _31855_, _39551_);
  and (_01393_, _01392_, _01374_);
  and (_01394_, _01393_, _01391_);
  and (_01395_, _38023_, _38006_);
  nor (_01396_, _01395_, _00808_);
  nor (_01397_, _01396_, _36914_);
  and (_01398_, _33379_, _29987_);
  nand (_01399_, _01398_, _34064_);
  nor (_01400_, _01399_, _34760_);
  and (_01401_, _01400_, _35577_);
  nand (_01402_, _01401_, _36295_);
  nor (_01403_, _01402_, _31996_);
  nor (_01404_, _01391_, _37992_);
  and (_01405_, _01404_, _01403_);
  and (_01406_, _01405_, _30173_);
  not (_01407_, _01406_);
  and (_01408_, _01391_, _29143_);
  not (_01409_, _01408_);
  not (_01410_, _37992_);
  nor (_01411_, _01391_, _38016_);
  nor (_01412_, _01411_, _01410_);
  and (_01413_, _01412_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_01414_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_01415_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_01416_, _01415_, _01414_);
  nor (_01417_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor (_01418_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_01419_, _01418_, _01417_);
  and (_01420_, _01419_, _01416_);
  and (_01421_, _01420_, _38129_);
  nor (_01422_, _01421_, _01413_);
  and (_01423_, _01422_, _01409_);
  and (_01424_, _01423_, _01407_);
  and (_01425_, _00759_, _37890_);
  not (_01426_, _01425_);
  and (_01427_, _01426_, _38044_);
  nor (_01428_, _01427_, _01424_);
  not (_01429_, _01428_);
  not (_01430_, _37987_);
  or (_01431_, _38038_, _37967_);
  nor (_01432_, _01431_, _38060_);
  nor (_01433_, _01432_, _01430_);
  not (_01434_, _01433_);
  nor (_01435_, _01015_, _38021_);
  not (_01436_, _01435_);
  nor (_01437_, _01436_, _00823_);
  and (_01438_, _01437_, _00974_);
  and (_01439_, _01438_, _01434_);
  not (_01440_, _01439_);
  and (_01441_, _01440_, _01424_);
  or (_01442_, _37968_, _38076_);
  or (_01443_, _01442_, _00760_);
  nor (_01444_, _01443_, _01441_);
  and (_01445_, _01444_, _01429_);
  nor (_01446_, _37990_, _38094_);
  nor (_01447_, _01446_, _01445_);
  nor (_01448_, _01447_, _01397_);
  not (_01449_, _38889_);
  and (_01450_, _01449_, _38129_);
  nor (_01451_, _38624_, _38616_);
  and (_01452_, _01451_, _38638_);
  not (_01453_, _01452_);
  and (_01454_, _01453_, _01412_);
  nor (_01455_, _01454_, _01450_);
  not (_01456_, _01455_);
  nor (_01457_, _01456_, _01448_);
  not (_01458_, _01457_);
  nor (_01459_, _01458_, _01394_);
  and (_01460_, _01459_, _01390_);
  nor (_01461_, _38094_, rst);
  and (_38748_, _01461_, _01460_);
  and (_38749_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _42618_);
  and (_38750_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [7], _42618_);
  and (_01462_, _38094_, _31147_);
  not (_01463_, _38368_);
  and (_01464_, _37968_, _37990_);
  and (_01465_, _01464_, _01463_);
  nand (_01466_, _00974_, _38045_);
  or (_01467_, _01466_, _01436_);
  and (_01468_, _01467_, _37990_);
  and (_01469_, _01395_, _36903_);
  not (_01470_, _01469_);
  and (_01471_, _38037_, _36903_);
  and (_01472_, _01471_, _37987_);
  nor (_01473_, _01472_, _38094_);
  and (_01474_, _01473_, _01470_);
  not (_01475_, _01474_);
  nor (_01476_, _01475_, _01468_);
  nor (_01477_, _01464_, _01397_);
  nor (_01478_, _00761_, _37968_);
  nand (_01479_, _01478_, _01437_);
  or (_01480_, _01479_, _01466_);
  and (_01481_, _01480_, _37990_);
  nor (_01482_, _01481_, _01472_);
  and (_01483_, _01482_, _01477_);
  and (_01484_, _01483_, _01476_);
  and (_01485_, _01484_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_01486_, _01469_, _42096_);
  or (_01487_, _01486_, _01485_);
  or (_01488_, _01487_, _01465_);
  or (_01489_, _01488_, _01462_);
  and (_01490_, _01476_, _42095_);
  not (_01491_, _01178_);
  nor (_01492_, _01476_, _01491_);
  nor (_01493_, _01492_, _01490_);
  and (_01494_, _01493_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor (_01495_, _01493_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_01496_, _01476_, _42446_);
  not (_01497_, _01346_);
  nor (_01498_, _01476_, _01497_);
  nor (_01499_, _01498_, _01496_);
  nand (_01500_, _01499_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  or (_01501_, _01499_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_01502_, _01501_, _01500_);
  and (_01503_, _01476_, _42131_);
  not (_01504_, _01329_);
  nor (_01505_, _01476_, _01504_);
  nor (_01506_, _01505_, _01503_);
  and (_01507_, _01506_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nor (_01508_, _01506_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_01509_, _01476_, _42253_);
  not (_01510_, _01312_);
  nor (_01511_, _01476_, _01510_);
  nor (_01512_, _01511_, _01509_);
  nand (_01513_, _01512_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_01514_, _01476_, _42349_);
  not (_01515_, _01289_);
  nor (_01516_, _01476_, _01515_);
  nor (_01517_, _01516_, _01514_);
  and (_01518_, _01517_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nor (_01519_, _01517_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_01520_, _01476_, _42207_);
  not (_01521_, _01254_);
  nor (_01522_, _01476_, _01521_);
  nor (_01523_, _01522_, _01520_);
  and (_01524_, _01523_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_01525_, _01476_, _42298_);
  not (_01526_, _01219_);
  nor (_01527_, _01476_, _01526_);
  nor (_01528_, _01527_, _01525_);
  and (_01529_, _01528_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_01530_, _01476_, _42391_);
  not (_01531_, _01195_);
  nor (_01532_, _01476_, _01531_);
  nor (_01533_, _01532_, _01530_);
  and (_01534_, _01533_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor (_01535_, _01528_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nor (_01536_, _01535_, _01529_);
  and (_01537_, _01536_, _01534_);
  nor (_01538_, _01537_, _01529_);
  not (_01539_, _01538_);
  nor (_01540_, _01523_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nor (_01541_, _01540_, _01524_);
  and (_01542_, _01541_, _01539_);
  nor (_01543_, _01542_, _01524_);
  nor (_01544_, _01543_, _01519_);
  or (_01545_, _01544_, _01518_);
  or (_01546_, _01512_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_01547_, _01546_, _01513_);
  nand (_01548_, _01547_, _01545_);
  and (_01549_, _01548_, _01513_);
  nor (_01550_, _01549_, _01508_);
  or (_01551_, _01550_, _01507_);
  nand (_01552_, _01551_, _01502_);
  and (_01553_, _01552_, _01500_);
  nor (_01554_, _01553_, _01495_);
  or (_01555_, _01554_, _01494_);
  and (_01556_, \oc8051_top_1.oc8051_memory_interface1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_01557_, _01556_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_01558_, _01557_, _01555_);
  and (_01559_, _01558_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_01560_, \oc8051_top_1.oc8051_memory_interface1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_01561_, _01560_, _01559_);
  nor (_01562_, _01561_, _01493_);
  not (_01563_, _01493_);
  nor (_01564_, _01555_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_01565_, _01564_, _38291_);
  and (_01566_, _01565_, _38296_);
  and (_01567_, _01566_, _38281_);
  nor (_01568_, \oc8051_top_1.oc8051_memory_interface1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_01569_, _01568_, _01567_);
  nor (_01570_, _01569_, _01563_);
  nor (_01571_, _01570_, _01562_);
  or (_01572_, _01493_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand (_01573_, _01493_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_01574_, _01573_, _01572_);
  and (_01575_, _01574_, _01571_);
  or (_01576_, _01575_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nand (_01577_, _01575_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  not (_01578_, _01477_);
  and (_01579_, _01578_, _01476_);
  and (_01580_, _37987_, _36903_);
  and (_01581_, _01580_, _38037_);
  nor (_01582_, _01481_, _01581_);
  nor (_01583_, _01582_, _01579_);
  and (_01584_, _01583_, _01577_);
  and (_01585_, _01584_, _01576_);
  or (_01586_, _01585_, _01489_);
  and (_01587_, _01482_, _01579_);
  and (_01588_, \oc8051_top_1.oc8051_memory_interface1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_01589_, _01588_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_01590_, \oc8051_top_1.oc8051_memory_interface1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_01591_, \oc8051_top_1.oc8051_memory_interface1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_01592_, _01591_, _01590_);
  and (_01593_, _01592_, _01589_);
  and (_01594_, _01593_, _01557_);
  and (_01595_, _01594_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_01596_, _01595_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_01597_, _01596_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nand (_01598_, _01597_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand (_01599_, _01598_, _38317_);
  or (_01600_, _01598_, _38317_);
  and (_01601_, _01600_, _01599_);
  nand (_01602_, _01601_, _01587_);
  nand (_01603_, _01602_, _01460_);
  or (_01604_, _01603_, _01586_);
  and (_01605_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12], \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor (_01606_, _37067_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_01607_, _01606_, _42079_);
  nor (_01608_, _01607_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  and (_01609_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and (_01610_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5], \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and (_01611_, _01610_, _01609_);
  not (_01612_, _01611_);
  nor (_01613_, _01612_, _01608_);
  and (_01614_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7], \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_01615_, _01614_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_01616_, _01615_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and (_01617_, _01616_, _01613_);
  and (_01618_, _01617_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_01619_, _01618_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and (_01620_, _01619_, _01605_);
  and (_01621_, _01620_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or (_01622_, _01621_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nand (_01623_, _01621_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_01624_, _01623_, _01622_);
  or (_01625_, _01624_, _01460_);
  and (_01627_, _01625_, _42618_);
  and (_38751_, _01627_, _01604_);
  and (_01629_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _42618_);
  and (_01630_, _01629_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  not (_01632_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_01633_, _36958_, _01632_);
  not (_01635_, _01633_);
  not (_01636_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  and (_01638_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_01639_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_01641_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_01642_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  nor (_01644_, _01642_, _01639_);
  and (_01645_, _01644_, _01641_);
  nor (_01647_, _01645_, _01639_);
  nor (_01648_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_01650_, _01648_, _01638_);
  not (_01651_, _01650_);
  nor (_01653_, _01651_, _01647_);
  nor (_01654_, _01653_, _01638_);
  not (_01656_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  not (_01657_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  not (_01658_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  not (_01659_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  not (_01660_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  not (_01661_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  not (_01662_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  not (_01663_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  not (_01664_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_01665_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4], \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_01666_, _01665_, _01664_);
  and (_01667_, _01666_, _01663_);
  and (_01668_, _01667_, _01662_);
  and (_01669_, _01668_, _01661_);
  and (_01670_, _01669_, _01660_);
  and (_01671_, _01670_, _01659_);
  and (_01672_, _01671_, _01658_);
  and (_01673_, _01672_, _01657_);
  and (_01674_, _01673_, _01656_);
  and (_01675_, _01674_, _01654_);
  and (_01676_, _01675_, _01636_);
  nor (_01677_, _01676_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_01678_, _01676_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nor (_01679_, _01678_, _01677_);
  not (_01680_, _01679_);
  nor (_01681_, _01675_, _01636_);
  nor (_01682_, _01681_, _01676_);
  not (_01683_, _01682_);
  and (_01684_, _01673_, _01654_);
  nor (_01685_, _01684_, _01656_);
  or (_01686_, _01685_, _01675_);
  and (_01687_, _01672_, _01654_);
  nor (_01688_, _01687_, _01657_);
  nor (_01689_, _01688_, _01684_);
  not (_01690_, _01689_);
  and (_01691_, _01670_, _01654_);
  and (_01692_, _01691_, _01659_);
  nor (_01693_, _01692_, _01658_);
  nor (_01694_, _01693_, _01687_);
  not (_01695_, _01694_);
  nor (_01696_, _01691_, _01659_);
  nor (_01697_, _01696_, _01692_);
  not (_01698_, _01697_);
  and (_01699_, _01669_, _01654_);
  nor (_01700_, _01699_, _01660_);
  nor (_01701_, _01700_, _01691_);
  not (_01702_, _01701_);
  and (_01703_, _01667_, _01654_);
  nor (_01704_, _01703_, _01662_);
  and (_01705_, _01668_, _01654_);
  nor (_01706_, _01705_, _01704_);
  not (_01707_, _01706_);
  and (_01708_, _01666_, _01654_);
  nor (_01709_, _01708_, _01663_);
  nor (_01710_, _01709_, _01703_);
  not (_01711_, _01710_);
  and (_01712_, _01665_, _01654_);
  nor (_01713_, _01712_, _01664_);
  nor (_01714_, _01713_, _01708_);
  not (_01715_, _01714_);
  not (_01716_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_01717_, _01654_, _01716_);
  nor (_01718_, _01654_, _01716_);
  nor (_01719_, _01718_, _01717_);
  not (_01720_, _01719_);
  not (_01721_, _00730_);
  not (_01722_, _00687_);
  and (_01723_, _00675_, _00703_);
  not (_01724_, _01723_);
  nor (_01725_, _00683_, _00676_);
  and (_01726_, _01725_, _01724_);
  and (_01727_, _00718_, _00671_);
  and (_01728_, _00671_, _00674_);
  or (_01729_, _01728_, _01727_);
  nor (_01730_, _00704_, _00701_);
  not (_01731_, _01730_);
  nor (_01732_, _01731_, _01729_);
  and (_01733_, _01732_, _01726_);
  nor (_01734_, _01733_, _01722_);
  nor (_01735_, _01734_, _01721_);
  and (_01736_, _00683_, _00669_);
  not (_01737_, _01736_);
  nor (_01738_, _00736_, _00679_);
  and (_01739_, _01738_, _01737_);
  not (_01740_, _01739_);
  or (_01741_, _01728_, _00719_);
  nor (_01742_, _01730_, _37602_);
  or (_01743_, _01742_, _01741_);
  and (_01744_, _01743_, _00668_);
  nor (_01745_, _01744_, _01740_);
  and (_01746_, _01745_, _01735_);
  nor (_01747_, _00710_, _00698_);
  and (_01748_, _00675_, _00718_);
  and (_01749_, _01748_, _00678_);
  nor (_01750_, _01749_, _00666_);
  and (_01751_, _01750_, _01747_);
  and (_01752_, _00683_, _00678_);
  and (_01753_, _00674_, _00664_);
  and (_01754_, _00695_, _01753_);
  nor (_01755_, _01754_, _01752_);
  and (_01756_, _00689_, _37908_);
  and (_01757_, _01756_, _00687_);
  nor (_01758_, _01757_, _00705_);
  and (_01759_, _01758_, _01755_);
  and (_01760_, _01759_, _01751_);
  not (_01761_, _00678_);
  and (_01762_, _00675_, _00682_);
  not (_01763_, _01762_);
  nor (_01764_, _01723_, _00725_);
  and (_01765_, _01764_, _01763_);
  nor (_01766_, _01765_, _01761_);
  not (_01767_, _01766_);
  and (_01768_, _00719_, _00694_);
  and (_01769_, _00725_, _00695_);
  nor (_01770_, _01769_, _01768_);
  and (_01771_, _00704_, _00697_);
  and (_01772_, _00689_, _00678_);
  nor (_01773_, _01772_, _01771_);
  and (_01774_, _01773_, _01770_);
  and (_01775_, _01774_, _01767_);
  and (_01776_, _01775_, _01760_);
  nor (_01777_, _00672_, _00701_);
  and (_01778_, _00707_, _37330_);
  not (_01779_, _01778_);
  nor (_01780_, _01779_, _01777_);
  not (_01781_, _01780_);
  not (_01782_, _01753_);
  nor (_01783_, _00687_, _00668_);
  nor (_01784_, _01783_, _01782_);
  and (_01785_, _00671_, _00662_);
  and (_01786_, _01785_, _37884_);
  nor (_01787_, _01786_, _01784_);
  and (_01788_, _01787_, _01781_);
  not (_01789_, _00725_);
  nor (_01790_, _00687_, _00669_);
  nor (_01791_, _01790_, _01789_);
  not (_01792_, _00669_);
  nor (_01793_, _00908_, _00701_);
  nor (_01794_, _01793_, _01792_);
  nor (_01795_, _01794_, _01791_);
  nor (_01796_, _01727_, _00701_);
  nor (_01797_, _01796_, _37330_);
  and (_01798_, _00675_, _37908_);
  nor (_01799_, _01798_, _01727_);
  nor (_01800_, _01799_, _00732_);
  nor (_01801_, _01800_, _01797_);
  and (_01802_, _01801_, _01795_);
  and (_01803_, _01802_, _01788_);
  and (_01804_, _01803_, _01776_);
  and (_01805_, _01804_, _01746_);
  nor (_01806_, _01644_, _01641_);
  nor (_01807_, _01806_, _01645_);
  not (_01808_, _01807_);
  nor (_01809_, _01808_, _01805_);
  and (_01810_, _01755_, _01739_);
  nor (_01811_, _01730_, _01761_);
  not (_01812_, _01811_);
  nor (_01813_, _01757_, _00710_);
  and (_01814_, _01813_, _01812_);
  nor (_01815_, _01769_, _00728_);
  and (_01816_, _01728_, _00662_);
  and (_01817_, _00719_, _00695_);
  nor (_01818_, _01817_, _01816_);
  and (_01819_, _01818_, _01815_);
  and (_01820_, _01819_, _01814_);
  and (_01821_, _01820_, _01810_);
  not (_01822_, _01821_);
  nor (_01823_, _01822_, _01805_);
  not (_01824_, _01823_);
  nor (_01825_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_01826_, _01825_, _01641_);
  and (_01827_, _01826_, _01824_);
  and (_01828_, _01808_, _01805_);
  nor (_01829_, _01828_, _01809_);
  and (_01830_, _01829_, _01827_);
  nor (_01831_, _01830_, _01809_);
  not (_01832_, _01831_);
  and (_01833_, _01651_, _01647_);
  nor (_01834_, _01833_, _01653_);
  and (_01835_, _01834_, _01832_);
  and (_01836_, _01835_, _01720_);
  not (_01837_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_01838_, _01717_, _01837_);
  or (_01839_, _01838_, _01712_);
  and (_01840_, _01839_, _01836_);
  and (_01841_, _01840_, _01715_);
  and (_01842_, _01841_, _01711_);
  and (_01843_, _01842_, _01707_);
  nor (_01844_, _01705_, _01661_);
  or (_01845_, _01844_, _01699_);
  and (_01846_, _01845_, _01843_);
  and (_01847_, _01846_, _01702_);
  and (_01848_, _01847_, _01698_);
  and (_01849_, _01848_, _01695_);
  and (_01850_, _01849_, _01690_);
  and (_01851_, _01850_, _01686_);
  nand (_01852_, _01851_, _01683_);
  nand (_01853_, _01852_, _01680_);
  or (_01854_, _01852_, _01680_);
  and (_01855_, _01854_, _01853_);
  or (_01856_, _01855_, _01635_);
  or (_01857_, _01633_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor (_01858_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , rst);
  and (_01859_, _01858_, _01857_);
  and (_01860_, _01859_, _01856_);
  or (_38753_, _01860_, _01630_);
  nor (_01861_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , rst);
  and (_38754_, _01861_, \oc8051_top_1.oc8051_memory_interface1.int_ack_buff );
  and (_38755_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , _42618_);
  nor (_01862_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  nor (_01863_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_01864_, _01863_, _01862_);
  nor (_01865_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  nor (_01866_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and (_01867_, _01866_, _01865_);
  and (_01868_, _01867_, _01864_);
  nor (_01869_, _01868_, rst);
  and (_01870_, \oc8051_top_1.oc8051_rom1.ea_int , _36925_);
  nand (_01871_, _01870_, _36958_);
  and (_01872_, _01871_, _38755_);
  or (_38756_, _01872_, _01869_);
  and (_01873_, _01868_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  or (_01874_, _01873_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  and (_38758_, _01874_, _42618_);
  nor (_01875_, _01608_, _42079_);
  nor (_01876_, _01805_, _37155_);
  nor (_01877_, _01823_, _37111_);
  and (_01878_, _01805_, _37155_);
  nor (_01879_, _01878_, _01876_);
  and (_01880_, _01879_, _01877_);
  nor (_01881_, _01880_, _01876_);
  nor (_01882_, _01881_, _42079_);
  and (_01883_, _01882_, _37023_);
  nor (_01884_, _01882_, _37023_);
  nor (_01885_, _01884_, _01883_);
  nor (_01886_, _01885_, _01875_);
  and (_01887_, _37166_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nand (_01888_, _01887_, _01875_);
  nor (_01889_, _01888_, _01821_);
  or (_01890_, _01889_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_01891_, _01890_, _01886_);
  and (_38759_, _01891_, _42618_);
  or (_01892_, _37559_, _37927_);
  nor (_01893_, _01892_, _37286_);
  not (_01894_, _37852_);
  and (_01895_, _01894_, _37950_);
  and (_01896_, _01895_, _37820_);
  not (_01897_, _01353_);
  nor (_01898_, _01897_, _37878_);
  and (_01899_, _01898_, _37904_);
  and (_01900_, _01899_, _01896_);
  and (_38762_, _01900_, _01893_);
  nor (_01901_, \oc8051_top_1.oc8051_memory_interface1.istb_t , rst);
  and (_01902_, _01901_, \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  and (_01903_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [7]);
  and (_38765_, \oc8051_top_1.oc8051_memory_interface1.istb_t , _42618_);
  and (_01904_, _38765_, _01903_);
  or (_38763_, _01904_, _01902_);
  not (_01905_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and (_01906_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_01907_, _01906_, _01905_);
  and (_01908_, _01906_, _01905_);
  nor (_01909_, _01908_, _01907_);
  not (_01910_, _01909_);
  and (_01911_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and (_01912_, _01911_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_01913_, _01911_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_01914_, _01913_, _01912_);
  or (_01915_, _01914_, _01906_);
  and (_01916_, _01915_, _01910_);
  nor (_01917_, _01907_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and (_01918_, _01907_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  or (_01919_, _01918_, _01917_);
  or (_01920_, _01912_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  and (_38767_, _01920_, _42618_);
  and (_01921_, _38767_, _01919_);
  and (_38766_, _01921_, _01916_);
  not (_01922_, \oc8051_top_1.oc8051_rom1.ea_int );
  nor (_01923_, _01608_, _01922_);
  and (_01924_, _01923_, \oc8051_top_1.oc8051_rom1.data_o [31]);
  not (_01925_, _01923_);
  and (_01926_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  or (_01927_, _01926_, _01924_);
  and (_38768_, _01927_, _42618_);
  and (_01928_, _01923_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and (_01929_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  or (_01930_, _01929_, _01928_);
  and (_38769_, _01930_, _42618_);
  and (_01931_, \oc8051_top_1.oc8051_decoder1.mem_act [2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  not (_01932_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_01933_, \oc8051_top_1.oc8051_decoder1.mem_act [0], _01932_);
  and (_01934_, _01933_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_01935_, _01934_, _01931_);
  and (_38770_, _01935_, _42618_);
  and (_01936_, \oc8051_top_1.oc8051_memory_interface1.dwe_o , \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_01937_, _01936_, _01933_);
  and (_38771_, _01937_, _42618_);
  or (_01938_, _01932_, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  and (_38773_, _01938_, _42618_);
  not (_01939_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  and (_01940_, _01939_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_01941_, _01940_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_01942_, _01932_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  and (_01943_, _01942_, _42618_);
  and (_38774_, _01943_, _01941_);
  or (_01944_, _01932_, \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and (_38775_, _01944_, _42618_);
  nor (_01945_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  and (_01946_, _01945_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_01947_, _01946_, _42618_);
  and (_01948_, _38765_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or (_38776_, _01948_, _01947_);
  and (_01949_, _01922_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or (_01950_, _01949_, _01946_);
  and (_38777_, _01950_, _42618_);
  nand (_01951_, _01946_, _38368_);
  or (_01952_, _01946_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [15]);
  and (_01953_, _01952_, _42618_);
  and (_38778_, _01953_, _01951_);
  nand (_01954_, _37999_, _42618_);
  nor (_38779_, _01954_, _38133_);
  or (_01955_, _01347_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  not (_01956_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nand (_01957_, _01347_, _01956_);
  and (_01958_, _01957_, _42618_);
  and (_38816_, _01958_, _01955_);
  or (_01959_, _01347_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  not (_01960_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nand (_01961_, _01347_, _01960_);
  and (_01962_, _01961_, _42618_);
  and (_38817_, _01962_, _01959_);
  or (_01963_, _01347_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  not (_01964_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nand (_01965_, _01347_, _01964_);
  and (_01966_, _01965_, _42618_);
  and (_38818_, _01966_, _01963_);
  or (_01967_, _01347_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  not (_01968_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nand (_01969_, _01347_, _01968_);
  and (_01970_, _01969_, _42618_);
  and (_38819_, _01970_, _01967_);
  or (_01971_, _01347_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  or (_01972_, _01351_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_01973_, _01972_, _42618_);
  and (_38820_, _01973_, _01971_);
  or (_01974_, _01347_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  not (_01975_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nand (_01976_, _01347_, _01975_);
  and (_01977_, _01976_, _42618_);
  and (_38822_, _01977_, _01974_);
  or (_01978_, _01347_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  not (_01979_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nand (_01980_, _01347_, _01979_);
  and (_01981_, _01980_, _42618_);
  and (_38823_, _01981_, _01978_);
  or (_01982_, _01347_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  not (_01983_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nand (_01984_, _01347_, _01983_);
  and (_01985_, _01984_, _42618_);
  and (_38824_, _01985_, _01982_);
  or (_01986_, _01347_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nand (_01987_, _01347_, _38285_);
  and (_01988_, _01987_, _42618_);
  and (_38825_, _01988_, _01986_);
  or (_01989_, _01347_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nand (_01990_, _01347_, _38291_);
  and (_01991_, _01990_, _42618_);
  and (_38826_, _01991_, _01989_);
  or (_01992_, _01347_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nand (_01993_, _01347_, _38296_);
  and (_01994_, _01993_, _42618_);
  and (_38827_, _01994_, _01992_);
  or (_01995_, _01347_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nand (_01996_, _01347_, _38281_);
  and (_01997_, _01996_, _42618_);
  and (_38828_, _01997_, _01995_);
  or (_01998_, _01347_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nand (_01999_, _01347_, _38302_);
  and (_02000_, _01999_, _42618_);
  and (_38829_, _02000_, _01998_);
  or (_02001_, _01347_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nand (_02002_, _01347_, _38307_);
  and (_02003_, _02002_, _42618_);
  and (_38830_, _02003_, _02001_);
  or (_02004_, _01347_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nand (_02005_, _01347_, _38312_);
  and (_02006_, _02005_, _42618_);
  and (_38831_, _02006_, _02004_);
  and (_02007_, _01347_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_02008_, _01351_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  or (_02009_, _02008_, _02007_);
  and (_38836_, _02009_, _42618_);
  and (_02010_, _01347_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_02011_, _01351_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  or (_02012_, _02011_, _02010_);
  and (_38837_, _02012_, _42618_);
  and (_02013_, _01347_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_02014_, _01351_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  or (_02015_, _02014_, _02013_);
  and (_38838_, _02015_, _42618_);
  and (_02016_, _01347_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_02017_, _01351_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or (_02018_, _02017_, _02016_);
  and (_38839_, _02018_, _42618_);
  and (_02019_, _01347_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  and (_02020_, _01351_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  or (_02021_, _02020_, _02019_);
  and (_38840_, _02021_, _42618_);
  and (_02022_, _01347_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  and (_02023_, _01351_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  or (_02024_, _02023_, _02022_);
  and (_38841_, _02024_, _42618_);
  and (_02025_, _01347_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  and (_02026_, _01351_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  or (_02027_, _02026_, _02025_);
  and (_38842_, _02027_, _42618_);
  and (_02028_, _01347_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  and (_02029_, _01351_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  or (_02030_, _02029_, _02028_);
  and (_38843_, _02030_, _42618_);
  and (_02031_, _01347_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  and (_02032_, _01351_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  or (_02033_, _02032_, _02031_);
  and (_38844_, _02033_, _42618_);
  and (_02034_, _01347_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and (_02035_, _01351_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  or (_02036_, _02035_, _02034_);
  and (_38845_, _02036_, _42618_);
  and (_02037_, _01347_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  and (_02038_, _01351_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  or (_02039_, _02038_, _02037_);
  and (_38847_, _02039_, _42618_);
  and (_02040_, _01347_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and (_02041_, _01351_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  or (_02042_, _02041_, _02040_);
  and (_38848_, _02042_, _42618_);
  and (_02043_, _01347_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  and (_02044_, _01351_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  or (_02045_, _02044_, _02043_);
  and (_38849_, _02045_, _42618_);
  and (_02046_, _01347_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and (_02047_, _01351_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  or (_02048_, _02047_, _02046_);
  and (_38850_, _02048_, _42618_);
  and (_02049_, _01347_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  and (_02050_, _01351_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  or (_02051_, _02050_, _02049_);
  and (_38851_, _02051_, _42618_);
  and (_39027_, _37657_, _42618_);
  and (_39028_, _37863_, _42618_);
  and (_39029_, _37837_, _42618_);
  nor (_39030_, _42022_, rst);
  and (_02052_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_02053_, _01923_, \oc8051_top_1.oc8051_rom1.data_o [0]);
  or (_02054_, _02053_, _02052_);
  and (_39031_, _02054_, _42618_);
  and (_02055_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_02056_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [1]);
  and (_02057_, _02056_, _01923_);
  or (_02058_, _02057_, _02055_);
  and (_39032_, _02058_, _42618_);
  and (_02059_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_02060_, _01923_, \oc8051_top_1.oc8051_rom1.data_o [2]);
  or (_02061_, _02060_, _02059_);
  and (_39033_, _02061_, _42618_);
  and (_02062_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_02063_, _01923_, \oc8051_top_1.oc8051_rom1.data_o [3]);
  or (_02064_, _02063_, _02062_);
  and (_39034_, _02064_, _42618_);
  and (_02065_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_02066_, _01923_, \oc8051_top_1.oc8051_rom1.data_o [4]);
  or (_02067_, _02066_, _02065_);
  and (_39036_, _02067_, _42618_);
  and (_02068_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_02069_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [5]);
  and (_02070_, _02069_, _01923_);
  or (_02071_, _02070_, _02068_);
  and (_39037_, _02071_, _42618_);
  and (_02072_, _01923_, \oc8051_top_1.oc8051_rom1.data_o [6]);
  and (_02073_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  or (_02074_, _02073_, _02072_);
  and (_39038_, _02074_, _42618_);
  and (_02075_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_02076_, _01923_, \oc8051_top_1.oc8051_rom1.data_o [7]);
  or (_02077_, _02076_, _02075_);
  and (_39039_, _02077_, _42618_);
  and (_02078_, _01923_, \oc8051_top_1.oc8051_rom1.data_o [8]);
  and (_02079_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  or (_02080_, _02079_, _02078_);
  and (_39040_, _02080_, _42618_);
  and (_02081_, _01923_, \oc8051_top_1.oc8051_rom1.data_o [9]);
  and (_02082_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  or (_02083_, _02082_, _02081_);
  and (_39041_, _02083_, _42618_);
  and (_02084_, _01923_, \oc8051_top_1.oc8051_rom1.data_o [10]);
  and (_02085_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  or (_02086_, _02085_, _02084_);
  and (_39042_, _02086_, _42618_);
  and (_02087_, _01923_, \oc8051_top_1.oc8051_rom1.data_o [11]);
  and (_02088_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  or (_02089_, _02088_, _02087_);
  and (_39043_, _02089_, _42618_);
  and (_02090_, _01923_, \oc8051_top_1.oc8051_rom1.data_o [12]);
  and (_02091_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  or (_02092_, _02091_, _02090_);
  and (_39044_, _02092_, _42618_);
  and (_02093_, _01923_, \oc8051_top_1.oc8051_rom1.data_o [13]);
  and (_02094_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  or (_02095_, _02094_, _02093_);
  and (_39045_, _02095_, _42618_);
  and (_02096_, _01923_, \oc8051_top_1.oc8051_rom1.data_o [14]);
  and (_02097_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  or (_02098_, _02097_, _02096_);
  and (_39047_, _02098_, _42618_);
  and (_02099_, _01923_, \oc8051_top_1.oc8051_rom1.data_o [15]);
  and (_02100_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  or (_02101_, _02100_, _02099_);
  and (_39048_, _02101_, _42618_);
  and (_02102_, _01923_, \oc8051_top_1.oc8051_rom1.data_o [16]);
  and (_02103_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  or (_02104_, _02103_, _02102_);
  and (_39049_, _02104_, _42618_);
  and (_02105_, _01923_, \oc8051_top_1.oc8051_rom1.data_o [17]);
  and (_02106_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  or (_02107_, _02106_, _02105_);
  and (_39050_, _02107_, _42618_);
  and (_02108_, _01923_, \oc8051_top_1.oc8051_rom1.data_o [18]);
  and (_02109_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  or (_02110_, _02109_, _02108_);
  and (_39051_, _02110_, _42618_);
  and (_02112_, _01923_, \oc8051_top_1.oc8051_rom1.data_o [19]);
  and (_02114_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  or (_02116_, _02114_, _02112_);
  and (_39052_, _02116_, _42618_);
  and (_02119_, _01923_, \oc8051_top_1.oc8051_rom1.data_o [20]);
  and (_02121_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  or (_02123_, _02121_, _02119_);
  and (_39053_, _02123_, _42618_);
  and (_02126_, _01923_, \oc8051_top_1.oc8051_rom1.data_o [21]);
  and (_02128_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  or (_02130_, _02128_, _02126_);
  and (_39054_, _02130_, _42618_);
  and (_02133_, _01923_, \oc8051_top_1.oc8051_rom1.data_o [22]);
  and (_02135_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  or (_02137_, _02135_, _02133_);
  and (_39055_, _02137_, _42618_);
  and (_02140_, _01923_, \oc8051_top_1.oc8051_rom1.data_o [23]);
  and (_02142_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  or (_02144_, _02142_, _02140_);
  and (_39056_, _02144_, _42618_);
  and (_02147_, _01923_, \oc8051_top_1.oc8051_rom1.data_o [24]);
  and (_02149_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  or (_02151_, _02149_, _02147_);
  and (_39058_, _02151_, _42618_);
  and (_02154_, _01923_, \oc8051_top_1.oc8051_rom1.data_o [25]);
  and (_02156_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  or (_02158_, _02156_, _02154_);
  and (_39059_, _02158_, _42618_);
  and (_02161_, _01923_, \oc8051_top_1.oc8051_rom1.data_o [26]);
  and (_02163_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  or (_02165_, _02163_, _02161_);
  and (_39060_, _02165_, _42618_);
  and (_02168_, _01923_, \oc8051_top_1.oc8051_rom1.data_o [27]);
  and (_02170_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  or (_02172_, _02170_, _02168_);
  and (_39061_, _02172_, _42618_);
  and (_02173_, _01923_, \oc8051_top_1.oc8051_rom1.data_o [28]);
  and (_02174_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  or (_02175_, _02174_, _02173_);
  and (_39062_, _02175_, _42618_);
  and (_02176_, _01923_, \oc8051_top_1.oc8051_rom1.data_o [29]);
  and (_02177_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  or (_02178_, _02177_, _02176_);
  and (_39063_, _02178_, _42618_);
  and (_02179_, _01923_, \oc8051_top_1.oc8051_rom1.data_o [30]);
  and (_02180_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  or (_02181_, _02180_, _02179_);
  and (_39064_, _02181_, _42618_);
  nor (_39065_, _42374_, rst);
  nor (_39067_, _42280_, rst);
  nor (_39068_, _42184_, rst);
  nor (_39069_, _42327_, rst);
  nor (_39070_, _42233_, rst);
  nor (_39071_, _42160_, rst);
  nor (_39073_, _42428_, rst);
  and (_39089_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], _42618_);
  and (_39090_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _42618_);
  and (_39091_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], _42618_);
  and (_39092_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], _42618_);
  and (_39093_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _42618_);
  and (_39095_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], _42618_);
  and (_39096_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], _42618_);
  or (_02182_, _01484_, _01464_);
  and (_02183_, _02182_, _32334_);
  and (_02184_, _01587_, _42392_);
  and (_02185_, _01469_, _01531_);
  and (_02186_, _38094_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  or (_02187_, _02186_, _02185_);
  or (_02188_, _02187_, _02184_);
  nor (_02189_, _01533_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor (_02190_, _02189_, _01534_);
  and (_02191_, _02190_, _01583_);
  nor (_02192_, _02191_, _02188_);
  nand (_02193_, _02192_, _01460_);
  or (_02194_, _02193_, _02183_);
  or (_02195_, _01460_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and (_02196_, _02195_, _42618_);
  and (_39097_, _02196_, _02194_);
  and (_02197_, _02182_, _33031_);
  and (_02198_, _01587_, _42299_);
  and (_02199_, _01469_, _01526_);
  and (_02200_, _38094_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or (_02201_, _02200_, _02199_);
  or (_02202_, _02201_, _02198_);
  or (_02203_, _02202_, _02197_);
  nor (_02204_, _01536_, _01534_);
  nor (_02205_, _02204_, _01537_);
  nand (_02206_, _02205_, _01583_);
  nand (_02207_, _02206_, _01460_);
  or (_02208_, _02207_, _02203_);
  or (_02209_, _01460_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  and (_02210_, _02209_, _42618_);
  and (_39098_, _02210_, _02208_);
  and (_02211_, _02182_, _33728_);
  and (_02212_, _01587_, _42208_);
  and (_02213_, _01469_, _01521_);
  or (_02214_, _02213_, _02212_);
  or (_02215_, _01541_, _01539_);
  not (_02216_, _01542_);
  and (_02217_, _01583_, _02216_);
  and (_02218_, _02217_, _02215_);
  or (_02219_, _02218_, _02214_);
  or (_02220_, _02219_, _02211_);
  nand (_02221_, _38094_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nand (_02222_, _02221_, _01460_);
  or (_02223_, _02222_, _02220_);
  not (_02224_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_02225_, _01608_, _02224_);
  and (_02226_, _01608_, _02224_);
  nor (_02227_, _02226_, _02225_);
  or (_02228_, _02227_, _01460_);
  and (_02229_, _02228_, _42618_);
  and (_39099_, _02229_, _02223_);
  and (_02230_, _02182_, _34489_);
  and (_02231_, _01587_, _42350_);
  and (_02232_, _01469_, _01515_);
  or (_02233_, _02232_, _02231_);
  or (_02234_, _01519_, _01518_);
  or (_02235_, _02234_, _01543_);
  nand (_02236_, _02234_, _01543_);
  and (_02237_, _02236_, _01583_);
  and (_02238_, _02237_, _02235_);
  or (_02239_, _02238_, _02233_);
  or (_02240_, _02239_, _02230_);
  nand (_02241_, _38094_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nand (_02242_, _02241_, _01460_);
  or (_02243_, _02242_, _02240_);
  and (_02244_, _02225_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_02245_, _02225_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_02246_, _02245_, _02244_);
  or (_02247_, _02246_, _01460_);
  and (_02248_, _02247_, _42618_);
  and (_39100_, _02248_, _02243_);
  and (_02249_, _02182_, _35251_);
  and (_02250_, _01469_, _01510_);
  and (_02251_, _01587_, _42254_);
  or (_02252_, _02251_, _02250_);
  or (_02253_, _01547_, _01545_);
  and (_02254_, _01583_, _01548_);
  and (_02255_, _02254_, _02253_);
  or (_02256_, _02255_, _02252_);
  or (_02257_, _02256_, _02249_);
  nand (_02258_, _38094_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nand (_02259_, _02258_, _01460_);
  or (_02260_, _02259_, _02257_);
  and (_02261_, _02244_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_02262_, _02244_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_02263_, _02262_, _02261_);
  or (_02264_, _02263_, _01460_);
  and (_02265_, _02264_, _42618_);
  and (_39101_, _02265_, _02260_);
  and (_02266_, _02182_, _36057_);
  and (_02267_, _01587_, _42132_);
  and (_02268_, _01469_, _01504_);
  and (_02269_, _38094_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  or (_02270_, _02269_, _02268_);
  or (_02271_, _02270_, _02267_);
  or (_02272_, _02271_, _02266_);
  or (_02273_, _01508_, _01507_);
  or (_02274_, _02273_, _01549_);
  nand (_02275_, _02273_, _01549_);
  and (_02276_, _02275_, _02274_);
  nand (_02277_, _02276_, _01583_);
  nand (_02278_, _02277_, _01460_);
  or (_02279_, _02278_, _02272_);
  nor (_02280_, _02261_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_02281_, _02280_, _01613_);
  or (_02282_, _02281_, _01460_);
  and (_02283_, _02282_, _42618_);
  and (_39102_, _02283_, _02279_);
  nor (_02284_, _01613_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_02285_, _01613_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor (_02286_, _02285_, _02284_);
  or (_02287_, _02286_, _01460_);
  and (_02288_, _02287_, _42618_);
  not (_02289_, _01460_);
  and (_02290_, _38094_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_02291_, _02182_, _36698_);
  and (_02292_, _01469_, _01497_);
  and (_02293_, _01587_, _42447_);
  or (_02294_, _02293_, _02292_);
  or (_02295_, _01551_, _01502_);
  and (_02296_, _01583_, _01552_);
  and (_02297_, _02296_, _02295_);
  or (_02298_, _02297_, _02294_);
  or (_02299_, _02298_, _02291_);
  or (_02300_, _02299_, _02290_);
  or (_02301_, _02300_, _02289_);
  and (_39103_, _02301_, _02288_);
  or (_02302_, _01494_, _01495_);
  or (_02303_, _02302_, _01553_);
  nand (_02304_, _02302_, _01553_);
  and (_02305_, _02304_, _02303_);
  and (_02306_, _02305_, _01583_);
  and (_02307_, _02182_, _31147_);
  and (_02308_, _38094_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and (_02309_, _01469_, _01491_);
  and (_02310_, _01587_, _42096_);
  or (_02311_, _02310_, _02309_);
  or (_02312_, _02311_, _02308_);
  or (_02313_, _02312_, _02307_);
  or (_02314_, _02313_, _02306_);
  or (_02315_, _02314_, _02289_);
  nor (_02316_, _02285_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and (_02317_, _02285_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor (_02318_, _02317_, _02316_);
  or (_02319_, _02318_, _01460_);
  and (_02320_, _02319_, _42618_);
  and (_39104_, _02320_, _02315_);
  and (_02321_, _38094_, _32334_);
  and (_02322_, _01555_, _38285_);
  nor (_02323_, _01555_, _38285_);
  nor (_02324_, _02323_, _02322_);
  nor (_02325_, _02324_, _01493_);
  and (_02326_, _02324_, _01493_);
  or (_02327_, _02326_, _02325_);
  and (_02328_, _02327_, _01583_);
  not (_02329_, _38405_);
  and (_02330_, _01464_, _02329_);
  and (_02331_, _01587_, _00711_);
  and (_02332_, _01469_, _42392_);
  or (_02333_, _02332_, _02331_);
  and (_02334_, _01484_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  or (_02335_, _02334_, _02333_);
  or (_02336_, _02335_, _02330_);
  or (_02337_, _02336_, _02328_);
  or (_02338_, _02337_, _02321_);
  or (_02339_, _02338_, _02289_);
  or (_02340_, _02317_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nand (_02341_, _01615_, _01613_);
  and (_02342_, _02341_, _02340_);
  or (_02343_, _02342_, _01460_);
  and (_02344_, _02343_, _42618_);
  and (_39106_, _02344_, _02339_);
  and (_02345_, _38094_, _33031_);
  not (_02346_, _38436_);
  and (_02347_, _01464_, _02346_);
  and (_02348_, _01587_, _00663_);
  and (_02349_, _01469_, _42299_);
  or (_02350_, _02349_, _02348_);
  and (_02351_, _01484_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  or (_02352_, _02351_, _02350_);
  or (_02353_, _02352_, _02347_);
  and (_02355_, _01555_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_02356_, _02355_, _01563_);
  and (_02357_, _01564_, _01493_);
  nor (_02358_, _02357_, _02356_);
  nand (_02359_, _02358_, _38291_);
  or (_02360_, _02358_, _38291_);
  and (_02361_, _02360_, _02359_);
  and (_02362_, _02361_, _01583_);
  or (_02363_, _02362_, _02353_);
  or (_02364_, _02363_, _02289_);
  or (_02365_, _02364_, _02345_);
  nand (_02366_, _02341_, _01660_);
  or (_02367_, _02341_, _01660_);
  and (_02368_, _02367_, _02366_);
  or (_02369_, _02368_, _01460_);
  and (_02370_, _02369_, _42618_);
  and (_39107_, _02370_, _02365_);
  and (_02371_, _38094_, _33728_);
  not (_02372_, _38466_);
  and (_02373_, _01464_, _02372_);
  and (_02374_, _01469_, _42208_);
  not (_02375_, _37931_);
  and (_02376_, _01587_, _02375_);
  and (_02377_, _01484_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  or (_02378_, _02377_, _02376_);
  or (_02379_, _02378_, _02374_);
  or (_02380_, _02379_, _02373_);
  and (_02381_, _01565_, _01493_);
  and (_02382_, _02356_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor (_02383_, _02382_, _02381_);
  nand (_02384_, _02383_, _38296_);
  or (_02385_, _02383_, _38296_);
  and (_02386_, _02385_, _02384_);
  and (_02387_, _02386_, _01583_);
  or (_02388_, _02387_, _02380_);
  or (_02389_, _02388_, _02371_);
  or (_02390_, _02389_, _02289_);
  nor (_02391_, _01617_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor (_02392_, _02391_, _01618_);
  or (_02393_, _02392_, _01460_);
  and (_02394_, _02393_, _42618_);
  and (_39108_, _02394_, _02390_);
  and (_02395_, _01558_, _01563_);
  and (_02396_, _01566_, _01493_);
  nor (_02397_, _02396_, _02395_);
  nand (_02398_, _02397_, _38281_);
  or (_02399_, _02397_, _38281_);
  and (_02400_, _02399_, _02398_);
  and (_02401_, _02400_, _01583_);
  and (_02402_, _38094_, _34489_);
  not (_02403_, _38497_);
  and (_02404_, _01464_, _02403_);
  and (_02405_, _01484_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor (_02406_, _01594_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_02407_, _02406_, _01595_);
  and (_02408_, _02407_, _01587_);
  and (_02409_, _01469_, _42350_);
  or (_02410_, _02409_, _02408_);
  or (_02411_, _02410_, _02405_);
  or (_02412_, _02411_, _02404_);
  or (_02413_, _02412_, _02402_);
  or (_02414_, _02413_, _02401_);
  or (_02415_, _02414_, _02289_);
  nor (_02416_, _01618_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor (_02417_, _02416_, _01619_);
  or (_02418_, _02417_, _01460_);
  and (_02419_, _02418_, _42618_);
  and (_39109_, _02419_, _02415_);
  nor (_02420_, _01595_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_02421_, _02420_, _01596_);
  and (_02422_, _02421_, _01587_);
  and (_02423_, _01559_, _01563_);
  and (_02424_, _01567_, _01493_);
  nor (_02425_, _02424_, _02423_);
  or (_02426_, _02425_, _38302_);
  nand (_02427_, _02425_, _38302_);
  and (_02428_, _02427_, _01583_);
  and (_02429_, _02428_, _02426_);
  and (_02430_, _38094_, _35251_);
  not (_02431_, _38528_);
  and (_02432_, _01464_, _02431_);
  and (_02433_, _01484_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and (_02434_, _01469_, _42254_);
  or (_02435_, _02434_, _02433_);
  or (_02436_, _02435_, _02432_);
  or (_02437_, _02436_, _02430_);
  or (_02438_, _02437_, _02429_);
  or (_02439_, _02438_, _02422_);
  or (_02440_, _02439_, _02289_);
  nor (_02441_, _01619_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and (_02442_, _01619_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor (_02443_, _02442_, _02441_);
  or (_02444_, _02443_, _01460_);
  and (_02445_, _02444_, _42618_);
  and (_39110_, _02445_, _02440_);
  nor (_02446_, _01596_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_02447_, _02446_, _01597_);
  and (_02448_, _02447_, _01587_);
  and (_02449_, _38094_, _36057_);
  not (_02450_, _38561_);
  and (_02451_, _01464_, _02450_);
  and (_02452_, _01484_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and (_02453_, _01469_, _42132_);
  or (_02454_, _02453_, _02452_);
  or (_02455_, _02454_, _02451_);
  or (_02456_, _02455_, _02449_);
  or (_02457_, _02456_, _02448_);
  and (_02458_, _02423_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_02459_, _02424_, _38302_);
  nor (_02460_, _02459_, _02458_);
  or (_02461_, _02460_, _38307_);
  nand (_02462_, _02460_, _38307_);
  and (_02463_, _02462_, _01583_);
  and (_02464_, _02463_, _02461_);
  or (_02465_, _02464_, _02289_);
  or (_02466_, _02465_, _02457_);
  or (_02467_, _02442_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nand (_02468_, _02442_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and (_02469_, _02468_, _02467_);
  or (_02470_, _02469_, _01460_);
  and (_02471_, _02470_, _42618_);
  and (_39111_, _02471_, _02466_);
  or (_02472_, _01597_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_02473_, _02472_, _01598_);
  and (_02474_, _02473_, _01587_);
  and (_02475_, _38094_, _36698_);
  and (_02476_, _01464_, _38589_);
  and (_02477_, _01469_, _42447_);
  and (_02478_, _01484_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or (_02479_, _02478_, _02477_);
  or (_02480_, _02479_, _02476_);
  or (_02481_, _02480_, _02475_);
  or (_02482_, _01571_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand (_02483_, _01571_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_02484_, _02483_, _01583_);
  and (_02485_, _02484_, _02482_);
  or (_02486_, _02485_, _02481_);
  or (_02487_, _02486_, _02474_);
  or (_02488_, _02487_, _02289_);
  nor (_02489_, _01620_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor (_02490_, _02489_, _01621_);
  or (_02491_, _02490_, _01460_);
  and (_02492_, _02491_, _42618_);
  and (_39112_, _02492_, _02488_);
  and (_02493_, _01629_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nor (_02494_, _01826_, _01824_);
  nor (_02495_, _02494_, _01827_);
  or (_02496_, _02495_, _01635_);
  or (_02497_, _01633_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_02498_, _02497_, _01858_);
  and (_02499_, _02498_, _02496_);
  or (_39113_, _02499_, _02493_);
  nor (_02500_, _01829_, _01827_);
  nor (_02501_, _02500_, _01830_);
  or (_02502_, _02501_, _01635_);
  or (_02503_, _01633_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_02504_, _02503_, _01858_);
  and (_02505_, _02504_, _02502_);
  and (_02506_, _01629_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or (_39114_, _02506_, _02505_);
  and (_02507_, _01629_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_02508_, _01834_, _01832_);
  nor (_02509_, _02508_, _01835_);
  or (_02510_, _02509_, _01635_);
  or (_02511_, _01633_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_02512_, _02511_, _01858_);
  and (_02513_, _02512_, _02510_);
  or (_39115_, _02513_, _02507_);
  and (_02514_, _01629_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_02515_, _01835_, _01720_);
  nor (_02516_, _02515_, _01836_);
  or (_02517_, _02516_, _01635_);
  or (_02518_, _01633_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_02519_, _02518_, _01858_);
  and (_02520_, _02519_, _02517_);
  or (_39117_, _02520_, _02514_);
  and (_02521_, _01629_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_02522_, _01839_, _01836_);
  nor (_02523_, _02522_, _01840_);
  or (_02524_, _02523_, _01635_);
  or (_02525_, _01633_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_02526_, _02525_, _01858_);
  and (_02527_, _02526_, _02524_);
  or (_39118_, _02527_, _02521_);
  and (_02528_, _01629_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_02529_, _01840_, _01715_);
  nor (_02530_, _02529_, _01841_);
  or (_02531_, _02530_, _01635_);
  or (_02532_, _01633_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_02533_, _02532_, _01858_);
  and (_02534_, _02533_, _02531_);
  or (_39119_, _02534_, _02528_);
  nor (_02535_, _01841_, _01711_);
  nor (_02536_, _02535_, _01842_);
  or (_02537_, _02536_, _01635_);
  or (_02538_, _01633_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_02539_, _02538_, _01858_);
  and (_02540_, _02539_, _02537_);
  and (_02541_, _01629_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or (_39120_, _02541_, _02540_);
  nor (_02543_, _01842_, _01707_);
  nor (_02544_, _02543_, _01843_);
  or (_02545_, _02544_, _01635_);
  or (_02546_, _01633_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_02547_, _02546_, _01858_);
  and (_02548_, _02547_, _02545_);
  and (_02549_, _01629_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  or (_39121_, _02549_, _02548_);
  and (_02550_, _01629_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor (_02551_, _01845_, _01843_);
  nor (_02552_, _02551_, _01846_);
  or (_02553_, _02552_, _01635_);
  or (_02554_, _01633_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_02555_, _02554_, _01858_);
  and (_02556_, _02555_, _02553_);
  or (_39122_, _02556_, _02550_);
  nor (_02557_, _01846_, _01702_);
  nor (_02558_, _02557_, _01847_);
  or (_02559_, _02558_, _01635_);
  or (_02560_, _01633_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_02561_, _02560_, _01858_);
  and (_02562_, _02561_, _02559_);
  and (_02563_, _01629_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  or (_39123_, _02563_, _02562_);
  nor (_02565_, _01847_, _01698_);
  nor (_02566_, _02565_, _01848_);
  or (_02567_, _02566_, _01635_);
  or (_02568_, _01633_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_02569_, _02568_, _01858_);
  and (_02570_, _02569_, _02567_);
  and (_02571_, _01629_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  or (_39124_, _02571_, _02570_);
  nor (_02572_, _01848_, _01695_);
  nor (_02573_, _02572_, _01849_);
  or (_02575_, _02573_, _01635_);
  or (_02576_, _01633_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_02577_, _02576_, _01858_);
  and (_02578_, _02577_, _02575_);
  and (_02579_, _01629_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  or (_39125_, _02579_, _02578_);
  or (_02580_, _01849_, _01690_);
  nor (_02581_, _01850_, _01635_);
  and (_02582_, _02581_, _02580_);
  nor (_02583_, _01633_, _38302_);
  or (_02584_, _02583_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_02585_, _02584_, _02582_);
  or (_02586_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12], _36925_);
  and (_02587_, _02586_, _42618_);
  and (_39126_, _02587_, _02585_);
  nor (_02588_, _01850_, _01686_);
  nor (_02589_, _02588_, _01851_);
  or (_02590_, _02589_, _01635_);
  or (_02591_, _01633_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_02592_, _02591_, _01858_);
  and (_02593_, _02592_, _02590_);
  and (_02594_, _01629_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or (_39128_, _02594_, _02593_);
  or (_02595_, _01851_, _01683_);
  and (_02596_, _02595_, _01852_);
  or (_02597_, _02596_, _01635_);
  or (_02598_, _01633_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_02599_, _02598_, _01858_);
  and (_02600_, _02599_, _02597_);
  and (_02601_, _01629_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or (_39129_, _02601_, _02600_);
  and (_02602_, _01868_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  or (_02603_, _02602_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  and (_39130_, _02603_, _42618_);
  and (_02604_, _01868_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  or (_02605_, _02604_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and (_39131_, _02605_, _42618_);
  and (_02606_, _01868_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  or (_02607_, _02606_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  and (_39132_, _02607_, _42618_);
  and (_02608_, _01868_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  or (_02609_, _02608_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_39133_, _02609_, _42618_);
  and (_02610_, _01868_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  or (_02611_, _02610_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and (_39134_, _02611_, _42618_);
  and (_02612_, _01868_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  or (_02613_, _02612_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  and (_39135_, _02613_, _42618_);
  and (_02614_, _01868_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  or (_02615_, _02614_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  and (_39136_, _02615_, _42618_);
  nor (_02616_, _01823_, _42079_);
  nand (_02617_, _02616_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  or (_02618_, _02616_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_02619_, _02618_, _01858_);
  and (_39137_, _02619_, _02617_);
  nor (_02620_, _01879_, _01877_);
  nor (_02621_, _02620_, _01880_);
  or (_02622_, _02621_, _42079_);
  or (_02623_, _36958_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_02624_, _02623_, _01858_);
  and (_39139_, _02624_, _02622_);
  and (_02625_, _01901_, \oc8051_top_1.oc8051_memory_interface1.cdata [0]);
  and (_02626_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [0]);
  and (_02627_, _02626_, _38765_);
  or (_39155_, _02627_, _02625_);
  and (_02628_, _01901_, \oc8051_top_1.oc8051_memory_interface1.cdata [1]);
  and (_02629_, _02056_, _38765_);
  or (_39156_, _02629_, _02628_);
  and (_02630_, _01901_, \oc8051_top_1.oc8051_memory_interface1.cdata [2]);
  and (_02631_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [2]);
  and (_02632_, _02631_, _38765_);
  or (_39157_, _02632_, _02630_);
  and (_02633_, _01901_, \oc8051_top_1.oc8051_memory_interface1.cdata [3]);
  and (_02634_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [3]);
  and (_02635_, _02634_, _38765_);
  or (_39158_, _02635_, _02633_);
  and (_02636_, _01901_, \oc8051_top_1.oc8051_memory_interface1.cdata [4]);
  and (_02637_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [4]);
  and (_02638_, _02637_, _38765_);
  or (_39159_, _02638_, _02636_);
  and (_02639_, _01901_, \oc8051_top_1.oc8051_memory_interface1.cdata [5]);
  and (_02640_, _02069_, _38765_);
  or (_39161_, _02640_, _02639_);
  and (_02641_, _01901_, \oc8051_top_1.oc8051_memory_interface1.cdata [6]);
  and (_02642_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [6]);
  and (_02643_, _02642_, _38765_);
  or (_39162_, _02643_, _02641_);
  and (_39163_, _01909_, _42618_);
  nor (_39164_, _01919_, rst);
  and (_39165_, _01915_, _42618_);
  and (_02644_, _01923_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_02645_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  or (_02646_, _02645_, _02644_);
  and (_39166_, _02646_, _42618_);
  and (_02647_, _01923_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_02648_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  or (_02649_, _02648_, _02647_);
  and (_39167_, _02649_, _42618_);
  and (_02650_, _01923_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_02651_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  or (_02652_, _02651_, _02650_);
  and (_39168_, _02652_, _42618_);
  and (_02653_, _01923_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_02654_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  or (_02655_, _02654_, _02653_);
  and (_39169_, _02655_, _42618_);
  and (_02656_, _01923_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_02657_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  or (_02658_, _02657_, _02656_);
  and (_39170_, _02658_, _42618_);
  and (_02659_, _01923_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_02660_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  or (_02661_, _02660_, _02659_);
  and (_39171_, _02661_, _42618_);
  and (_02662_, _01923_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_02663_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  or (_02664_, _02663_, _02662_);
  and (_39172_, _02664_, _42618_);
  and (_02665_, _01923_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_02666_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  or (_02667_, _02666_, _02665_);
  and (_39173_, _02667_, _42618_);
  and (_02668_, _01923_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_02669_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  or (_02670_, _02669_, _02668_);
  and (_39174_, _02670_, _42618_);
  and (_02671_, _01923_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_02672_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  or (_02673_, _02672_, _02671_);
  and (_39175_, _02673_, _42618_);
  and (_02674_, _01923_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_02675_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  or (_02676_, _02675_, _02674_);
  and (_39176_, _02676_, _42618_);
  and (_02677_, _01923_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_02678_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  or (_02679_, _02678_, _02677_);
  and (_39177_, _02679_, _42618_);
  and (_02680_, _01923_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_02681_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  or (_02682_, _02681_, _02680_);
  and (_39178_, _02682_, _42618_);
  and (_02683_, _01923_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_02684_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  or (_02685_, _02684_, _02683_);
  and (_39179_, _02685_, _42618_);
  and (_02686_, _01923_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_02687_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  or (_02688_, _02687_, _02686_);
  and (_39180_, _02688_, _42618_);
  and (_02689_, _01923_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_02690_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  or (_02691_, _02690_, _02689_);
  and (_39182_, _02691_, _42618_);
  and (_02692_, _01923_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_02693_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  or (_02694_, _02693_, _02692_);
  and (_39183_, _02694_, _42618_);
  and (_02695_, _01923_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_02696_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  or (_02697_, _02696_, _02695_);
  and (_39184_, _02697_, _42618_);
  and (_02698_, _01923_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_02699_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  or (_02701_, _02699_, _02698_);
  and (_39185_, _02701_, _42618_);
  and (_02702_, _01923_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_02703_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  or (_02704_, _02703_, _02702_);
  and (_39186_, _02704_, _42618_);
  and (_02705_, _01923_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_02706_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  or (_02707_, _02706_, _02705_);
  and (_39187_, _02707_, _42618_);
  and (_02708_, _01923_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_02709_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  or (_02710_, _02709_, _02708_);
  and (_39188_, _02710_, _42618_);
  and (_02711_, _01923_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_02712_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  or (_02713_, _02712_, _02711_);
  and (_39189_, _02713_, _42618_);
  and (_02714_, _01923_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_02715_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  or (_02716_, _02715_, _02714_);
  and (_39190_, _02716_, _42618_);
  and (_02717_, _01923_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and (_02718_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  or (_02719_, _02718_, _02717_);
  and (_39191_, _02719_, _42618_);
  and (_02720_, _01923_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and (_02721_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  or (_02722_, _02721_, _02720_);
  and (_39193_, _02722_, _42618_);
  and (_02723_, _01923_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and (_02724_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  or (_02725_, _02724_, _02723_);
  and (_39194_, _02725_, _42618_);
  and (_02726_, _01923_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and (_02727_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  or (_02728_, _02727_, _02726_);
  and (_39195_, _02728_, _42618_);
  and (_02729_, _01923_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and (_02730_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  or (_02731_, _02730_, _02729_);
  and (_39196_, _02731_, _42618_);
  and (_02732_, _01923_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and (_02733_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  or (_02734_, _02733_, _02732_);
  and (_39197_, _02734_, _42618_);
  and (_02735_, _01923_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and (_02736_, _01925_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  or (_02737_, _02736_, _02735_);
  and (_39198_, _02737_, _42618_);
  and (_02738_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [0], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_02739_, _01933_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_02740_, _02739_, _02738_);
  and (_39199_, _02740_, _42618_);
  and (_02741_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [1], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_02742_, _01933_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_02743_, _02742_, _02741_);
  and (_39200_, _02743_, _42618_);
  and (_02744_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_02745_, _01933_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_02746_, _02745_, _02744_);
  and (_39201_, _02746_, _42618_);
  and (_02747_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [3], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_02748_, _01933_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_02749_, _02748_, _02747_);
  and (_39202_, _02749_, _42618_);
  and (_02750_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [4], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_02751_, _01933_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or (_02752_, _02751_, _02750_);
  and (_39204_, _02752_, _42618_);
  and (_02753_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [5], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_02754_, _01933_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or (_02755_, _02754_, _02753_);
  and (_39205_, _02755_, _42618_);
  and (_02756_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [6], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_02757_, _01933_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_02758_, _02757_, _02756_);
  and (_39206_, _02758_, _42618_);
  and (_02759_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_02760_, _42374_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_02761_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_02762_, _02761_, _01932_);
  and (_02763_, _02762_, _02760_);
  or (_02764_, _02763_, _02759_);
  and (_39207_, _02764_, _42618_);
  and (_02765_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_02766_, _42280_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_02767_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_02768_, _02767_, _01932_);
  and (_02769_, _02768_, _02766_);
  or (_02770_, _02769_, _02765_);
  and (_39208_, _02770_, _42618_);
  and (_02771_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_02772_, _42184_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_02773_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_02774_, _02773_, _01932_);
  and (_02775_, _02774_, _02772_);
  or (_02776_, _02775_, _02771_);
  and (_39209_, _02776_, _42618_);
  and (_02777_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_02778_, _42327_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_02779_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_02780_, _02779_, _01932_);
  and (_02781_, _02780_, _02778_);
  or (_02782_, _02781_, _02777_);
  and (_39210_, _02782_, _42618_);
  and (_02783_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_02784_, _42233_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_02785_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_02786_, _02785_, _01932_);
  and (_02787_, _02786_, _02784_);
  or (_02788_, _02787_, _02783_);
  and (_39211_, _02788_, _42618_);
  and (_02789_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_02790_, _42160_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_02791_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_02792_, _02791_, _01932_);
  and (_02793_, _02792_, _02790_);
  or (_02794_, _02793_, _02789_);
  and (_39212_, _02794_, _42618_);
  and (_02795_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_02796_, _42428_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_02797_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_02799_, _02797_, _01932_);
  and (_02800_, _02799_, _02796_);
  or (_02801_, _02800_, _02795_);
  and (_39213_, _02801_, _42618_);
  and (_02802_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_02804_, _42072_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_02805_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_02806_, _02805_, _01932_);
  and (_02807_, _02806_, _02804_);
  or (_02808_, _02807_, _02802_);
  and (_39215_, _02808_, _42618_);
  and (_02810_, _01939_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or (_02811_, _02810_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_02812_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8], _01932_);
  and (_02813_, _02812_, _42618_);
  and (_39216_, _02813_, _02811_);
  and (_02815_, _01939_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_02816_, _02815_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_02817_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9], _01932_);
  and (_02818_, _02817_, _42618_);
  and (_39217_, _02818_, _02816_);
  and (_02820_, _01939_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_02821_, _02820_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_02822_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10], _01932_);
  and (_02823_, _02822_, _42618_);
  and (_39218_, _02823_, _02821_);
  and (_02825_, _01939_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_02826_, _02825_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_02827_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11], _01932_);
  and (_02828_, _02827_, _42618_);
  and (_39219_, _02828_, _02826_);
  and (_02830_, _01939_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or (_02832_, _02830_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_02833_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12], _01932_);
  and (_02834_, _02833_, _42618_);
  and (_39220_, _02834_, _02832_);
  and (_02835_, _01939_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or (_02837_, _02835_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_02838_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13], _01932_);
  and (_02840_, _02838_, _42618_);
  and (_39221_, _02840_, _02837_);
  and (_02841_, _01939_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_02843_, _02841_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_02844_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14], _01932_);
  and (_02845_, _02844_, _42618_);
  and (_39222_, _02845_, _02843_);
  nand (_02847_, _01946_, _32323_);
  or (_02849_, _01946_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  and (_02851_, _02849_, _42618_);
  and (_39223_, _02851_, _02847_);
  nand (_02852_, _01946_, _33020_);
  or (_02854_, _01946_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1]);
  and (_02855_, _02854_, _42618_);
  and (_39224_, _02855_, _02852_);
  nand (_02857_, _01946_, _33717_);
  or (_02858_, _01946_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2]);
  and (_02859_, _02858_, _42618_);
  and (_39226_, _02859_, _02857_);
  nand (_02861_, _01946_, _34478_);
  or (_02863_, _01946_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3]);
  and (_02864_, _02863_, _42618_);
  and (_39227_, _02864_, _02861_);
  nand (_02865_, _01946_, _35240_);
  or (_02866_, _01946_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [4]);
  and (_02867_, _02866_, _42618_);
  and (_39228_, _02867_, _02865_);
  nand (_02869_, _01946_, _36046_);
  or (_02871_, _01946_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [5]);
  and (_02872_, _02871_, _42618_);
  and (_39229_, _02872_, _02869_);
  not (_02874_, _01946_);
  or (_02875_, _02874_, _36698_);
  or (_02877_, _01946_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [6]);
  and (_02878_, _02877_, _42618_);
  and (_39230_, _02878_, _02875_);
  nand (_02880_, _01946_, _31136_);
  or (_02881_, _01946_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [7]);
  and (_02883_, _02881_, _42618_);
  and (_39231_, _02883_, _02880_);
  nand (_02885_, _01946_, _38405_);
  or (_02886_, _01946_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [8]);
  and (_02888_, _02886_, _42618_);
  and (_39232_, _02888_, _02885_);
  nand (_02889_, _01946_, _38436_);
  or (_02891_, _01946_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [9]);
  and (_02892_, _02891_, _42618_);
  and (_39233_, _02892_, _02889_);
  nand (_02895_, _01946_, _38466_);
  or (_02896_, _01946_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [10]);
  and (_02897_, _02896_, _42618_);
  and (_39234_, _02897_, _02895_);
  nand (_02899_, _01946_, _38497_);
  or (_02900_, _01946_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [11]);
  and (_02901_, _02900_, _42618_);
  and (_39235_, _02901_, _02899_);
  nand (_02903_, _01946_, _38528_);
  or (_02904_, _01946_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [12]);
  and (_02906_, _02904_, _42618_);
  and (_39237_, _02906_, _02903_);
  nand (_02907_, _01946_, _38561_);
  or (_02909_, _01946_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [13]);
  and (_02910_, _02909_, _42618_);
  and (_39238_, _02910_, _02907_);
  or (_02912_, _02874_, _38589_);
  or (_02913_, _01946_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [14]);
  and (_02914_, _02913_, _42618_);
  and (_39239_, _02914_, _02912_);
  nor (_39457_, _42115_, rst);
  and (_02917_, _42030_, _38137_);
  and (_02919_, _02917_, _28091_);
  and (_02920_, _02919_, _42032_);
  nand (_02922_, _02920_, _38225_);
  or (_02923_, _02920_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  and (_02924_, _02923_, _42618_);
  and (_39458_, _02924_, _02922_);
  and (_02925_, _02917_, _39011_);
  not (_02926_, _02925_);
  nor (_02928_, _02926_, _38225_);
  not (_02930_, _42032_);
  and (_02931_, _02926_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  or (_02932_, _02931_, _02930_);
  or (_02934_, _02932_, _02928_);
  or (_02935_, _42032_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  and (_02936_, _02935_, _42618_);
  and (_39459_, _02936_, _02934_);
  and (_02938_, _38813_, _31790_);
  and (_02939_, _02917_, _02938_);
  and (_02942_, _02939_, _42032_);
  nand (_02943_, _02942_, _38225_);
  or (_02944_, _02942_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  and (_02946_, _02944_, _42618_);
  and (_39460_, _02946_, _02943_);
  and (_02947_, _02917_, _41127_);
  and (_02949_, _02947_, _42032_);
  not (_02950_, _02949_);
  nor (_02951_, _02950_, _38225_);
  and (_02953_, _02950_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  or (_02955_, _02953_, _02951_);
  and (_39462_, _02955_, _42618_);
  and (_02957_, _42030_, _38629_);
  and (_02958_, _02957_, _28091_);
  and (_02959_, _02958_, _42032_);
  not (_02961_, _02959_);
  nor (_02962_, _02961_, _38225_);
  nor (_02963_, _02925_, _02919_);
  not (_02965_, _02939_);
  and (_02966_, _02965_, _02963_);
  not (_02968_, _02947_);
  and (_02970_, _02968_, _02966_);
  not (_02971_, _02958_);
  and (_02972_, _02971_, _02970_);
  or (_02974_, _02972_, _02930_);
  or (_02975_, _02974_, _02919_);
  and (_02976_, _02975_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  or (_02978_, _02947_, _02939_);
  or (_02979_, _02978_, _02925_);
  and (_02980_, _42032_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  and (_02983_, _02980_, _02979_);
  or (_02984_, _02983_, _02976_);
  or (_02985_, _02984_, _02962_);
  and (_39463_, _02985_, _42618_);
  and (_02987_, _02957_, _39011_);
  nor (_02989_, _02987_, _02958_);
  and (_02990_, _02989_, _02968_);
  and (_02991_, _02990_, _02966_);
  or (_02992_, _02958_, _02978_);
  and (_02994_, _02992_, _42032_);
  nand (_02996_, _02963_, _42032_);
  or (_02997_, _02996_, _02994_);
  or (_02999_, _02997_, _02991_);
  and (_03000_, _02999_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  and (_03001_, _02987_, _42032_);
  and (_03003_, _03001_, _41608_);
  or (_03004_, _03003_, _03000_);
  and (_39464_, _03004_, _42618_);
  and (_03006_, _02957_, _02938_);
  and (_03007_, _03006_, _42032_);
  not (_03009_, _03007_);
  and (_03011_, _03009_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  nor (_03012_, _03009_, _38225_);
  or (_03013_, _03012_, _03011_);
  and (_39465_, _03013_, _42618_);
  and (_03015_, _02957_, _41127_);
  and (_03016_, _03015_, _42032_);
  not (_03018_, _03016_);
  nor (_03019_, _03018_, _38225_);
  not (_03021_, _03006_);
  and (_03023_, _03021_, _02989_);
  nor (_03024_, _03015_, _03006_);
  and (_03025_, _03024_, _02991_);
  nand (_03027_, _02970_, _42032_);
  nor (_03028_, _03027_, _03025_);
  nand (_03029_, _03028_, _03023_);
  and (_03031_, _03029_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  or (_03032_, _03031_, _03019_);
  and (_39466_, _03032_, _42618_);
  nand (_03034_, _02920_, _38203_);
  or (_03035_, _02920_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  and (_03036_, _03035_, _42618_);
  and (_39555_, _03036_, _03034_);
  nand (_03038_, _02920_, _38191_);
  or (_03039_, _02920_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  and (_03041_, _03039_, _42618_);
  and (_39556_, _03041_, _03038_);
  nand (_03042_, _02920_, _38184_);
  or (_03044_, _02920_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  and (_03045_, _03044_, _42618_);
  and (_39557_, _03045_, _03042_);
  nand (_03047_, _02920_, _38177_);
  or (_03048_, _02920_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  and (_03050_, _03048_, _42618_);
  and (_39558_, _03050_, _03047_);
  nand (_03051_, _02920_, _38169_);
  or (_03052_, _02920_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  and (_03053_, _03052_, _42618_);
  and (_39559_, _03053_, _03051_);
  nand (_03054_, _02920_, _38162_);
  or (_03056_, _02920_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  and (_03057_, _03056_, _42618_);
  and (_39560_, _03057_, _03054_);
  nand (_03059_, _02920_, _38155_);
  or (_03060_, _02920_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  and (_03061_, _03060_, _42618_);
  and (_39561_, _03061_, _03059_);
  and (_03063_, _02926_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  nor (_03064_, _02926_, _38203_);
  or (_03066_, _03064_, _02930_);
  or (_03067_, _03066_, _03063_);
  or (_03068_, _42032_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  and (_03070_, _03068_, _42618_);
  and (_39562_, _03070_, _03067_);
  nor (_03071_, _02926_, _38191_);
  and (_03073_, _02926_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  or (_03074_, _03073_, _02930_);
  or (_03075_, _03074_, _03071_);
  or (_03077_, _42032_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  and (_03078_, _03077_, _42618_);
  and (_39563_, _03078_, _03075_);
  nor (_03080_, _02926_, _38184_);
  and (_03081_, _02926_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  or (_03082_, _03081_, _02930_);
  or (_03084_, _03082_, _03080_);
  or (_03085_, _42032_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  and (_03086_, _03085_, _42618_);
  and (_39564_, _03086_, _03084_);
  nor (_03088_, _02926_, _38177_);
  and (_03089_, _02926_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  or (_03091_, _03089_, _02930_);
  or (_03092_, _03091_, _03088_);
  or (_03093_, _42032_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  and (_03095_, _03093_, _42618_);
  and (_39566_, _03095_, _03092_);
  nor (_03096_, _02926_, _38169_);
  and (_03098_, _02926_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  or (_03099_, _03098_, _02930_);
  or (_03100_, _03099_, _03096_);
  or (_03102_, _42032_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  and (_03103_, _03102_, _42618_);
  and (_39567_, _03103_, _03100_);
  nor (_03105_, _02926_, _38162_);
  and (_03106_, _02926_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  or (_03108_, _03106_, _02930_);
  or (_03109_, _03108_, _03105_);
  or (_03110_, _42032_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  and (_03111_, _03110_, _42618_);
  and (_39568_, _03111_, _03109_);
  nor (_03113_, _02926_, _38155_);
  and (_03114_, _02926_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  or (_03116_, _03114_, _02930_);
  or (_03117_, _03116_, _03113_);
  or (_03118_, _42032_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  and (_03120_, _03118_, _42618_);
  and (_39569_, _03120_, _03117_);
  nand (_03121_, _02942_, _38203_);
  or (_03123_, _02942_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  and (_03124_, _03123_, _03121_);
  and (_39570_, _03124_, _42618_);
  not (_03127_, _02942_);
  nor (_03128_, _03127_, _38191_);
  and (_03129_, _03127_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  or (_03131_, _03129_, _03128_);
  and (_39571_, _03131_, _42618_);
  nor (_03132_, _03127_, _38184_);
  and (_03134_, _03127_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  or (_03135_, _03134_, _03132_);
  and (_39572_, _03135_, _42618_);
  nor (_03137_, _03127_, _38177_);
  and (_03138_, _03127_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  or (_03139_, _03138_, _03137_);
  and (_39573_, _03139_, _42618_);
  nand (_03141_, _02942_, _38169_);
  or (_03142_, _02942_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  and (_03144_, _03142_, _42618_);
  and (_39574_, _03144_, _03141_);
  nor (_03145_, _03127_, _38162_);
  and (_03147_, _03127_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  or (_03148_, _03147_, _03145_);
  and (_39575_, _03148_, _42618_);
  nor (_03150_, _03127_, _38155_);
  and (_03151_, _03127_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  or (_03152_, _03151_, _03150_);
  and (_39577_, _03152_, _42618_);
  and (_03154_, _02949_, _38204_);
  and (_03155_, _02950_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  or (_03157_, _03155_, _03154_);
  and (_39578_, _03157_, _42618_);
  nor (_03158_, _02950_, _38191_);
  and (_03160_, _02950_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  or (_03161_, _03160_, _03158_);
  and (_39579_, _03161_, _42618_);
  and (_03163_, _02950_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  nor (_03164_, _02950_, _38184_);
  or (_03165_, _03164_, _03163_);
  and (_39580_, _03165_, _42618_);
  nor (_03167_, _02950_, _38177_);
  and (_03168_, _02950_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  or (_03169_, _03168_, _03167_);
  and (_39581_, _03169_, _42618_);
  nor (_03171_, _02950_, _38169_);
  and (_03172_, _02950_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  or (_03174_, _03172_, _03171_);
  and (_39582_, _03174_, _42618_);
  nor (_03175_, _02950_, _38162_);
  and (_03177_, _02950_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  or (_03178_, _03177_, _03175_);
  and (_39583_, _03178_, _42618_);
  nor (_03180_, _02950_, _38155_);
  and (_03181_, _02950_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  or (_03182_, _03181_, _03180_);
  and (_39584_, _03182_, _42618_);
  and (_03184_, _02959_, _38204_);
  and (_03185_, _02961_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  or (_03187_, _03185_, _03184_);
  and (_39585_, _03187_, _42618_);
  and (_03189_, _02971_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  nor (_03190_, _02971_, _38191_);
  or (_03191_, _03190_, _03189_);
  or (_03192_, _03191_, _02930_);
  or (_03194_, _42032_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  and (_03195_, _03194_, _42618_);
  and (_39586_, _03195_, _03192_);
  nor (_03197_, _02971_, _38184_);
  and (_03198_, _02971_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  or (_03199_, _03198_, _02930_);
  or (_03201_, _03199_, _03197_);
  or (_03202_, _42032_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  and (_03203_, _03202_, _42618_);
  and (_39588_, _03203_, _03201_);
  and (_03205_, _02975_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  and (_03206_, _42032_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  and (_03208_, _03206_, _02979_);
  nor (_03209_, _02961_, _38177_);
  or (_03210_, _03209_, _03208_);
  or (_03212_, _03210_, _03205_);
  and (_39589_, _03212_, _42618_);
  and (_03213_, _02975_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  and (_03215_, _42032_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  and (_03216_, _03215_, _02979_);
  nor (_03218_, _02961_, _38169_);
  or (_03219_, _03218_, _03216_);
  or (_03220_, _03219_, _03213_);
  and (_39590_, _03220_, _42618_);
  nor (_03222_, _02961_, _38162_);
  and (_03223_, _02961_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  or (_03224_, _03223_, _03222_);
  and (_39591_, _03224_, _42618_);
  nor (_03226_, _02961_, _38155_);
  and (_03227_, _02975_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  and (_03229_, _42032_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  and (_03230_, _03229_, _02979_);
  or (_03231_, _03230_, _03227_);
  or (_03233_, _03231_, _03226_);
  and (_39592_, _03233_, _42618_);
  and (_03234_, _02999_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  and (_03236_, _03001_, _38204_);
  or (_03237_, _03236_, _03234_);
  and (_39593_, _03237_, _42618_);
  and (_03239_, _02999_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  and (_03240_, _03001_, _42278_);
  or (_03241_, _03240_, _03239_);
  and (_39594_, _03241_, _42618_);
  and (_03243_, _02999_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  and (_03245_, _03001_, _39884_);
  or (_03246_, _03245_, _03243_);
  and (_39595_, _03246_, _42618_);
  and (_03247_, _02999_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  and (_03249_, _03001_, _39896_);
  or (_03250_, _03249_, _03247_);
  and (_39596_, _03250_, _42618_);
  and (_03252_, _02999_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  and (_03253_, _03001_, _39907_);
  or (_03254_, _03253_, _03252_);
  and (_39597_, _03254_, _42618_);
  and (_03256_, _02999_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  and (_03257_, _03001_, _39920_);
  or (_03259_, _03257_, _03256_);
  and (_39599_, _03259_, _42618_);
  and (_03260_, _02999_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  and (_03262_, _03001_, _39933_);
  or (_03263_, _03262_, _03260_);
  and (_39600_, _03263_, _42618_);
  and (_03265_, _03009_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  and (_03266_, _03007_, _38204_);
  or (_03267_, _03266_, _03265_);
  and (_39601_, _03267_, _42618_);
  and (_03269_, _03023_, _02970_);
  nor (_03270_, _03269_, _02930_);
  nand (_03271_, _03270_, _02966_);
  and (_03272_, _03271_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  nor (_03273_, _03009_, _38191_);
  nand (_03274_, _42032_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  nor (_03275_, _03274_, _02990_);
  or (_03276_, _03275_, _03273_);
  or (_03277_, _03276_, _03272_);
  and (_39602_, _03277_, _42618_);
  nor (_03278_, _03009_, _38184_);
  and (_03279_, _03009_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  or (_03280_, _03279_, _03278_);
  and (_39603_, _03280_, _42618_);
  nor (_03281_, _03009_, _38177_);
  and (_03282_, _03009_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  or (_03283_, _03282_, _03281_);
  and (_39604_, _03283_, _42618_);
  nor (_03284_, _03009_, _38169_);
  and (_03285_, _03009_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  or (_03286_, _03285_, _03284_);
  and (_39605_, _03286_, _42618_);
  nor (_03287_, _03009_, _38162_);
  and (_03288_, _03009_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  or (_03289_, _03288_, _03287_);
  and (_39606_, _03289_, _42618_);
  nor (_03290_, _03009_, _38155_);
  and (_03291_, _03009_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  or (_03292_, _03291_, _03290_);
  and (_39607_, _03292_, _42618_);
  and (_03293_, _03024_, _02989_);
  or (_03294_, _03293_, _02930_);
  and (_03295_, _03294_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  and (_03296_, _03016_, _38204_);
  nand (_03297_, _42032_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  nor (_03298_, _03297_, _03023_);
  or (_03299_, _03298_, _03296_);
  or (_03300_, _03299_, _03295_);
  and (_39608_, _03300_, _42618_);
  and (_03301_, _03029_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  nor (_03302_, _03018_, _38191_);
  or (_03303_, _03302_, _03301_);
  and (_39610_, _03303_, _42618_);
  and (_03304_, _03294_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  nor (_03305_, _03018_, _38184_);
  nand (_03306_, _42032_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  nor (_03307_, _03306_, _03023_);
  or (_03308_, _03307_, _03305_);
  or (_03309_, _03308_, _03304_);
  and (_39611_, _03309_, _42618_);
  and (_03310_, _03294_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  nor (_03311_, _03018_, _38177_);
  nand (_03312_, _42032_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  nor (_03313_, _03312_, _03023_);
  or (_03314_, _03313_, _03311_);
  or (_03315_, _03314_, _03310_);
  and (_39612_, _03315_, _42618_);
  nor (_03316_, _03018_, _38169_);
  and (_03317_, _03018_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  or (_03318_, _03317_, _03316_);
  and (_39613_, _03318_, _42618_);
  and (_03319_, _03018_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  nor (_03320_, _03018_, _38162_);
  or (_03321_, _03320_, _03319_);
  and (_39614_, _03321_, _42618_);
  and (_03322_, _03294_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  nor (_03323_, _03018_, _38155_);
  nand (_03324_, _42032_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  nor (_03325_, _03324_, _03023_);
  or (_03326_, _03325_, _03323_);
  or (_03327_, _03326_, _03322_);
  and (_39615_, _03327_, _42618_);
  not (_03329_, \oc8051_top_1.oc8051_sfr1.prescaler [2]);
  and (_03330_, \oc8051_top_1.oc8051_sfr1.prescaler [0], \oc8051_top_1.oc8051_sfr1.prescaler [1]);
  and (_03331_, _03330_, _03329_);
  and (_03332_, \oc8051_top_1.oc8051_sfr1.prescaler [3], _42618_);
  and (_39679_, _03332_, _03331_);
  nor (_03333_, _03331_, rst);
  nand (_03334_, _03330_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  or (_03335_, _03330_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  and (_03336_, _03335_, _03334_);
  and (_39681_, _03336_, _03333_);
  nor (_03337_, _42451_, _42164_);
  not (_03338_, _42100_);
  and (_03339_, _42259_, _03338_);
  and (_03340_, _03339_, _42354_);
  and (_03341_, _03340_, _03337_);
  and (_03342_, _03341_, _38785_);
  nor (_03343_, _03342_, _01393_);
  nor (_03344_, _42212_, _38162_);
  and (_03345_, _42212_, _42278_);
  or (_03346_, _03345_, _03344_);
  not (_03347_, _42400_);
  and (_03348_, _03347_, _42307_);
  and (_03349_, _03348_, _03346_);
  or (_03350_, _42212_, _39933_);
  nor (_03351_, _03347_, _42307_);
  nand (_03352_, _42212_, _38184_);
  and (_03353_, _03352_, _03351_);
  and (_03354_, _03353_, _03350_);
  nor (_03355_, _42212_, _38225_);
  and (_03356_, _42212_, _39896_);
  or (_03357_, _03356_, _03355_);
  nor (_03358_, _42400_, _42307_);
  and (_03359_, _03358_, _03357_);
  nand (_03360_, _42212_, _38203_);
  and (_03361_, _42400_, _42307_);
  or (_03362_, _42212_, _39907_);
  and (_03363_, _03362_, _03361_);
  and (_03364_, _03363_, _03360_);
  or (_03365_, _03364_, _03359_);
  or (_03366_, _03365_, _03354_);
  nor (_03367_, _03366_, _03349_);
  nor (_03368_, _03367_, _03343_);
  nor (_03369_, _42451_, _42165_);
  nor (_03370_, _42259_, _42100_);
  and (_03371_, _03370_, _42354_);
  and (_03372_, _03371_, _03369_);
  nor (_03373_, _38899_, _38887_);
  and (_03374_, _38899_, _38887_);
  nor (_03375_, _03374_, _03373_);
  and (_03376_, _38872_, _38857_);
  nor (_03377_, _38872_, _38857_);
  or (_03378_, _03377_, _03376_);
  nor (_03379_, _03378_, _03375_);
  and (_03380_, _03378_, _03375_);
  nor (_03381_, _03380_, _03379_);
  nor (_03382_, _38923_, _38911_);
  and (_03383_, _38923_, _38911_);
  nor (_03384_, _03383_, _03382_);
  not (_03385_, _38809_);
  nor (_03386_, _38933_, _03385_);
  and (_03387_, _38933_, _03385_);
  nor (_03388_, _03387_, _03386_);
  nor (_03389_, _03388_, _03384_);
  and (_03390_, _03388_, _03384_);
  or (_03391_, _03390_, _03389_);
  nor (_03392_, _03391_, _03381_);
  and (_03393_, _03391_, _03381_);
  nor (_03394_, _03393_, _03392_);
  nand (_03395_, _03394_, _42212_);
  or (_03396_, _42212_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_03397_, _03396_, _03361_);
  and (_03398_, _03397_, _03395_);
  not (_03399_, _42212_);
  and (_03400_, _03348_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_03401_, _03358_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or (_03402_, _03401_, _03400_);
  and (_03403_, _03402_, _03399_);
  nor (_03404_, _42212_, _34086_);
  and (_03405_, _42212_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_03406_, _03405_, _03404_);
  and (_03407_, _03406_, _03351_);
  and (_03408_, _03348_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_03409_, _03358_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  or (_03410_, _03409_, _03408_);
  and (_03411_, _03410_, _42212_);
  or (_03412_, _03411_, _03407_);
  or (_03413_, _03412_, _03403_);
  or (_03414_, _03413_, _03398_);
  and (_03415_, _03414_, _03372_);
  and (_03416_, _01387_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_03417_, _03358_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_03418_, _03348_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or (_03419_, _03418_, _03417_);
  and (_03420_, _03419_, _03399_);
  or (_03421_, _42212_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nand (_03422_, _42212_, _38815_);
  and (_03423_, _03422_, _03361_);
  and (_03424_, _03423_, _03421_);
  and (_03425_, _03399_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_03426_, _42212_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_03427_, _03426_, _03425_);
  and (_03428_, _03427_, _03351_);
  or (_03429_, _03428_, _03424_);
  and (_03430_, _03358_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_03431_, _03348_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_03432_, _03431_, _03430_);
  and (_03433_, _03432_, _42212_);
  or (_03434_, _03433_, _03429_);
  or (_03435_, _03434_, _03420_);
  and (_03436_, _03435_, _03341_);
  or (_03437_, _03436_, _03416_);
  and (_03438_, _03369_, _03339_);
  and (_03439_, _03438_, _42355_);
  and (_03440_, _03361_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and (_03441_, _03351_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or (_03442_, _03441_, _03440_);
  and (_03443_, _03442_, _03399_);
  and (_03444_, _42212_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and (_03445_, _03399_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  or (_03446_, _03445_, _03444_);
  and (_03447_, _03446_, _03358_);
  and (_03448_, _42212_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  nor (_03449_, _42212_, _41014_);
  or (_03450_, _03449_, _03448_);
  and (_03451_, _03450_, _03348_);
  or (_03452_, _03451_, _03447_);
  and (_03453_, _03361_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and (_03454_, _03351_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or (_03455_, _03454_, _03453_);
  and (_03456_, _03455_, _42212_);
  or (_03457_, _03456_, _03452_);
  or (_03458_, _03457_, _03443_);
  and (_03459_, _03458_, _03439_);
  and (_03460_, _42451_, _42164_);
  and (_03461_, _03460_, _03340_);
  nor (_03462_, _00790_, _38035_);
  and (_03463_, _03462_, _00855_);
  nor (_03464_, _00853_, _38109_);
  and (_03465_, _38053_, _37985_);
  not (_03466_, _03465_);
  and (_03467_, _03466_, _03464_);
  and (_03468_, _38016_, _37395_);
  nor (_03469_, _03468_, _38065_);
  nor (_03470_, _00792_, _38047_);
  and (_03471_, _03470_, _03469_);
  and (_03472_, _03471_, _03467_);
  and (_03473_, _03472_, _01112_);
  and (_03474_, _03473_, _03463_);
  and (_03475_, _03474_, _38032_);
  nor (_03476_, _03475_, _36914_);
  nor (_03477_, _03476_, p0_in[0]);
  and (_03478_, _03476_, _39007_);
  nor (_03479_, _03478_, _03477_);
  or (_03480_, _03479_, _03399_);
  nor (_03481_, _03476_, p0_in[4]);
  and (_03482_, _03476_, _39258_);
  nor (_03483_, _03482_, _03481_);
  or (_03484_, _03483_, _42212_);
  and (_03485_, _03484_, _03361_);
  and (_03486_, _03485_, _03480_);
  or (_03487_, _03476_, p0_in[3]);
  not (_03488_, _03476_);
  or (_03489_, _03488_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_03490_, _03489_, _03487_);
  or (_03491_, _03490_, _03399_);
  or (_03492_, _03476_, p0_in[7]);
  or (_03493_, _03488_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_03494_, _03493_, _03492_);
  or (_03495_, _03494_, _42212_);
  and (_03496_, _03495_, _03358_);
  and (_03497_, _03496_, _03491_);
  or (_03498_, _03497_, _03486_);
  or (_03499_, _03476_, p0_in[5]);
  or (_03500_, _03488_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_03501_, _03500_, _03499_);
  and (_03502_, _03501_, _03399_);
  or (_03503_, _03476_, p0_in[1]);
  or (_03504_, _03488_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_03505_, _03504_, _03503_);
  and (_03506_, _03505_, _42212_);
  or (_03507_, _03506_, _03502_);
  and (_03508_, _03507_, _03348_);
  or (_03509_, _03476_, p0_in[2]);
  nand (_03510_, _03476_, _39024_);
  and (_03511_, _03510_, _03509_);
  or (_03512_, _03511_, _03399_);
  or (_03513_, _03476_, p0_in[6]);
  or (_03514_, _03488_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_03515_, _03514_, _03513_);
  or (_03516_, _03515_, _42212_);
  and (_03517_, _03516_, _03351_);
  and (_03518_, _03517_, _03512_);
  or (_03519_, _03518_, _03508_);
  or (_03520_, _03519_, _03498_);
  and (_03521_, _03520_, _03461_);
  or (_03522_, _03521_, _03459_);
  or (_03523_, _03522_, _03437_);
  and (_03524_, _42451_, _42165_);
  and (_03525_, _03370_, _42355_);
  or (_03526_, _42212_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  nand (_03528_, _42212_, _40470_);
  and (_03529_, _03528_, _03358_);
  and (_03530_, _03529_, _03526_);
  and (_03531_, _03399_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and (_03532_, _42212_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_03533_, _03532_, _03531_);
  and (_03534_, _03533_, _03351_);
  or (_03535_, _03534_, _03530_);
  and (_03536_, _42212_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  nor (_03537_, _42212_, _40465_);
  or (_03538_, _03537_, _03536_);
  and (_03539_, _03538_, _03361_);
  and (_03540_, _42212_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  nor (_03541_, _42212_, _40467_);
  or (_03542_, _03541_, _03540_);
  and (_03543_, _03542_, _03348_);
  or (_03544_, _03543_, _03539_);
  or (_03545_, _03544_, _03535_);
  and (_03546_, _03545_, _03525_);
  or (_03547_, _03476_, p2_in[3]);
  or (_03548_, _03488_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_03549_, _03548_, _03547_);
  or (_03550_, _03549_, _03399_);
  or (_03551_, _03476_, p2_in[7]);
  or (_03552_, _03488_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_03553_, _03552_, _03551_);
  or (_03554_, _03553_, _42212_);
  and (_03555_, _03554_, _03358_);
  and (_03556_, _03555_, _03550_);
  or (_03557_, _03476_, p2_in[6]);
  or (_03558_, _03488_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_03559_, _03558_, _03557_);
  and (_03560_, _03559_, _03399_);
  or (_03561_, _03476_, p2_in[2]);
  or (_03562_, _03488_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_03563_, _03562_, _03561_);
  and (_03564_, _03563_, _42212_);
  or (_03565_, _03564_, _03560_);
  and (_03566_, _03565_, _03351_);
  or (_03567_, _03566_, _03556_);
  nor (_03568_, _03476_, p2_in[0]);
  and (_03569_, _03476_, _39376_);
  nor (_03570_, _03569_, _03568_);
  or (_03571_, _03570_, _03399_);
  nor (_03572_, _03476_, p2_in[4]);
  and (_03573_, _03476_, _39425_);
  nor (_03574_, _03573_, _03572_);
  or (_03575_, _03574_, _42212_);
  and (_03576_, _03575_, _03361_);
  and (_03577_, _03576_, _03571_);
  or (_03578_, _03476_, p2_in[5]);
  or (_03579_, _03488_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_03580_, _03579_, _03578_);
  and (_03581_, _03580_, _03399_);
  or (_03582_, _03476_, p2_in[1]);
  or (_03583_, _03488_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_03584_, _03583_, _03582_);
  and (_03585_, _03584_, _42212_);
  or (_03586_, _03585_, _03581_);
  and (_03587_, _03586_, _03348_);
  or (_03588_, _03587_, _03577_);
  or (_03589_, _03588_, _03567_);
  and (_03590_, _03589_, _03340_);
  or (_03591_, _03590_, _03546_);
  and (_03592_, _03591_, _03524_);
  and (_03593_, _03525_, _03460_);
  and (_03594_, _42212_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  nor (_03595_, _42212_, _41017_);
  or (_03596_, _03595_, _03594_);
  and (_03597_, _03596_, _03358_);
  and (_03598_, _42212_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  nor (_03599_, _42212_, _41443_);
  or (_03600_, _03599_, _03598_);
  and (_03601_, _03600_, _03348_);
  or (_03602_, _03601_, _03597_);
  and (_03603_, _42212_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  nor (_03604_, _42212_, _41042_);
  or (_03605_, _03604_, _03603_);
  and (_03606_, _03605_, _03361_);
  and (_03607_, _03399_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  and (_03608_, _42212_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  or (_03609_, _03608_, _03607_);
  and (_03610_, _03609_, _03351_);
  or (_03611_, _03610_, _03606_);
  or (_03612_, _03611_, _03602_);
  and (_03613_, _03612_, _03593_);
  nor (_03614_, _03439_, _03371_);
  not (_03615_, _03369_);
  nand (_03616_, _03615_, _03340_);
  and (_03617_, _42451_, _03338_);
  nand (_03618_, _03617_, _42355_);
  and (_03619_, _03618_, \oc8051_top_1.oc8051_sfr1.bit_out );
  and (_03620_, _03619_, _03616_);
  and (_03621_, _03620_, _03614_);
  and (_03622_, _03524_, _03371_);
  or (_03623_, _03476_, p3_in[3]);
  or (_03624_, _03488_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_03625_, _03624_, _03623_);
  or (_03626_, _03625_, _03399_);
  or (_03627_, _03476_, p3_in[7]);
  or (_03628_, _03488_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and (_03629_, _03628_, _03627_);
  or (_03630_, _03629_, _42212_);
  and (_03631_, _03630_, _03358_);
  and (_03632_, _03631_, _03626_);
  or (_03633_, _03476_, p3_in[5]);
  or (_03634_, _03488_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_03635_, _03634_, _03633_);
  and (_03636_, _03635_, _03399_);
  or (_03637_, _03476_, p3_in[1]);
  or (_03638_, _03488_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_03639_, _03638_, _03637_);
  and (_03640_, _03639_, _42212_);
  or (_03641_, _03640_, _03636_);
  and (_03642_, _03641_, _03348_);
  or (_03643_, _03642_, _03632_);
  nor (_03644_, _03476_, p3_in[0]);
  and (_03645_, _03476_, _39471_);
  nor (_03646_, _03645_, _03644_);
  or (_03647_, _03646_, _03399_);
  nor (_03648_, _03476_, p3_in[4]);
  and (_03649_, _03476_, _39520_);
  nor (_03650_, _03649_, _03648_);
  or (_03651_, _03650_, _42212_);
  and (_03652_, _03651_, _03361_);
  and (_03653_, _03652_, _03647_);
  or (_03654_, _03476_, p3_in[6]);
  or (_03655_, _03488_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and (_03656_, _03655_, _03654_);
  and (_03657_, _03656_, _03399_);
  or (_03658_, _03476_, p3_in[2]);
  or (_03659_, _03488_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_03660_, _03659_, _03658_);
  and (_03661_, _03660_, _42212_);
  or (_03662_, _03661_, _03657_);
  and (_03663_, _03662_, _03351_);
  or (_03664_, _03663_, _03653_);
  or (_03665_, _03664_, _03643_);
  and (_03666_, _03665_, _03622_);
  or (_03667_, _03666_, _03621_);
  or (_03668_, _03667_, _03613_);
  or (_03669_, _03668_, _03592_);
  or (_03670_, _03669_, _03523_);
  and (_03671_, _03339_, _42355_);
  and (_03672_, _42212_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  nor (_03673_, _42212_, _39713_);
  or (_03674_, _03673_, _03672_);
  and (_03675_, _03674_, _03361_);
  or (_03676_, _42212_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or (_03677_, _03399_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and (_03678_, _03677_, _03358_);
  and (_03679_, _03678_, _03676_);
  or (_03680_, _03679_, _03675_);
  and (_03681_, _42212_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  and (_03682_, _03399_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or (_03683_, _03682_, _03681_);
  and (_03684_, _03683_, _03348_);
  nand (_03685_, _42212_, _40896_);
  or (_03686_, _42212_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and (_03687_, _03686_, _03351_);
  and (_03688_, _03687_, _03685_);
  or (_03689_, _03688_, _03684_);
  or (_03690_, _03689_, _03680_);
  and (_03691_, _03690_, _03460_);
  and (_03692_, _42212_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  nor (_03693_, _42212_, _40446_);
  or (_03694_, _03693_, _03692_);
  and (_03695_, _03694_, _03361_);
  or (_03696_, _42212_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  or (_03697_, _03399_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_03698_, _03697_, _03358_);
  and (_03699_, _03698_, _03696_);
  or (_03700_, _03699_, _03695_);
  and (_03701_, _42212_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  nor (_03702_, _42212_, _40450_);
  or (_03703_, _03702_, _03701_);
  and (_03704_, _03703_, _03348_);
  or (_03705_, _03399_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_03706_, _42212_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_03707_, _03706_, _03351_);
  and (_03708_, _03707_, _03705_);
  or (_03709_, _03708_, _03704_);
  or (_03710_, _03709_, _03700_);
  and (_03711_, _03710_, _03524_);
  or (_03712_, _03711_, _03691_);
  and (_03713_, _03712_, _03671_);
  and (_03714_, _42212_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nor (_03715_, _42212_, _35273_);
  or (_03716_, _03715_, _03714_);
  and (_03717_, _03716_, _03361_);
  and (_03718_, _42212_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  nor (_03719_, _42212_, _36078_);
  or (_03720_, _03719_, _03718_);
  and (_03721_, _03720_, _03348_);
  or (_03722_, _03721_, _03717_);
  and (_03723_, _42212_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nor (_03724_, _42212_, _31233_);
  or (_03725_, _03724_, _03723_);
  and (_03726_, _03725_, _03358_);
  nor (_03727_, _42212_, _36719_);
  and (_03729_, _42212_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or (_03730_, _03729_, _03727_);
  and (_03731_, _03730_, _03351_);
  or (_03732_, _03731_, _03726_);
  or (_03733_, _03732_, _03722_);
  and (_03734_, _03733_, _03337_);
  or (_03735_, _03476_, p1_in[5]);
  or (_03736_, _03488_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_03737_, _03736_, _03735_);
  and (_03738_, _03737_, _03399_);
  or (_03739_, _03476_, p1_in[1]);
  or (_03740_, _03488_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_03741_, _03740_, _03739_);
  and (_03742_, _03741_, _42212_);
  or (_03743_, _03742_, _03738_);
  and (_03744_, _03743_, _03348_);
  or (_03745_, _03476_, p1_in[2]);
  or (_03746_, _03488_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_03747_, _03746_, _03745_);
  or (_03748_, _03747_, _03399_);
  or (_03749_, _03476_, p1_in[6]);
  or (_03750_, _03488_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_03751_, _03750_, _03749_);
  or (_03752_, _03751_, _42212_);
  and (_03753_, _03752_, _03351_);
  and (_03754_, _03753_, _03748_);
  or (_03755_, _03476_, p1_in[3]);
  or (_03756_, _03488_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_03757_, _03756_, _03755_);
  or (_03758_, _03757_, _03399_);
  or (_03759_, _03476_, p1_in[7]);
  or (_03760_, _03488_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_03761_, _03760_, _03759_);
  or (_03762_, _03761_, _42212_);
  and (_03763_, _03762_, _03358_);
  and (_03764_, _03763_, _03758_);
  nor (_03765_, _03476_, p1_in[0]);
  and (_03766_, _03476_, _39294_);
  nor (_03767_, _03766_, _03765_);
  or (_03768_, _03767_, _03399_);
  nor (_03769_, _03476_, p1_in[4]);
  and (_03770_, _03476_, _39343_);
  nor (_03771_, _03770_, _03769_);
  or (_03772_, _03771_, _42212_);
  and (_03773_, _03772_, _03361_);
  and (_03774_, _03773_, _03768_);
  or (_03775_, _03774_, _03764_);
  or (_03776_, _03775_, _03754_);
  or (_03777_, _03776_, _03744_);
  and (_03778_, _03777_, _03460_);
  or (_03779_, _03778_, _03734_);
  and (_03780_, _03779_, _03371_);
  or (_03781_, _03780_, _03713_);
  or (_03782_, _03781_, _03670_);
  or (_03783_, _03782_, _03415_);
  nand (_03784_, _03416_, _31757_);
  and (_03785_, _03784_, _03343_);
  and (_03786_, _03785_, _03783_);
  or (_03787_, _03786_, _03368_);
  and (_39682_, _03787_, _42618_);
  and (_03788_, _42354_, _42212_);
  and (_03789_, _03788_, _03361_);
  and (_03790_, _03339_, _03337_);
  and (_03791_, _03790_, _03789_);
  and (_03792_, _03791_, _38785_);
  and (_03793_, _03358_, _03399_);
  not (_03794_, _03793_);
  and (_03795_, _03794_, _38795_);
  and (_03796_, _03795_, _01374_);
  nor (_03797_, _03796_, _03792_);
  and (_03798_, _03797_, _01390_);
  and (_03799_, _03460_, _03339_);
  and (_03800_, _03788_, _03358_);
  and (_03801_, _03800_, _03799_);
  and (_03802_, _03801_, _38276_);
  not (_03803_, _03802_);
  and (_03804_, _03791_, _38782_);
  nor (_03805_, _42451_, _42100_);
  and (_03806_, _42260_, _42164_);
  and (_03807_, _03806_, _03805_);
  and (_03808_, _03807_, _03789_);
  and (_03809_, _03808_, _38624_);
  nor (_03810_, _03809_, _03804_);
  and (_03811_, _03810_, _03803_);
  nor (_03812_, _03811_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_03813_, _03812_);
  and (_03814_, _03813_, _03798_);
  and (_03815_, _03788_, _03351_);
  and (_03816_, _03815_, _03799_);
  and (_03817_, _03816_, _38276_);
  or (_03818_, _03817_, rst);
  nor (_39683_, _03818_, _03814_);
  nand (_03819_, _03817_, _31136_);
  and (_03820_, _42355_, _42212_);
  and (_03821_, _03820_, _03358_);
  and (_03822_, _03821_, _03438_);
  and (_03823_, _03822_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  and (_03824_, _03820_, _03361_);
  and (_03825_, _03824_, _03799_);
  and (_03826_, _03825_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or (_03827_, _03826_, _03823_);
  and (_03828_, _03524_, _03339_);
  and (_03829_, _03828_, _03824_);
  and (_03830_, _03829_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_03831_, _03793_, _42354_);
  nor (_03832_, _42259_, _42164_);
  and (_03833_, _03832_, _03617_);
  and (_03834_, _03833_, _03831_);
  and (_03835_, _03834_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  or (_03836_, _03835_, _03830_);
  or (_03837_, _03836_, _03827_);
  nor (_03838_, _42354_, _42212_);
  and (_03839_, _03838_, _03361_);
  and (_03840_, _03839_, _03438_);
  and (_03841_, _03840_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and (_03842_, _03824_, _03438_);
  and (_03843_, _03842_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  or (_03844_, _03843_, _03841_);
  and (_03845_, _03838_, _03348_);
  and (_03846_, _03845_, _03438_);
  and (_03847_, _03846_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  and (_03848_, _03820_, _03351_);
  and (_03849_, _03848_, _03438_);
  and (_03850_, _03849_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  or (_03851_, _03850_, _03847_);
  or (_03852_, _03851_, _03844_);
  or (_03853_, _03852_, _03837_);
  and (_03854_, _03460_, _03370_);
  and (_03855_, _03820_, _03348_);
  and (_03856_, _03855_, _03854_);
  and (_03857_, _03856_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  and (_03858_, _03854_, _03824_);
  and (_03859_, _03858_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  or (_03860_, _03859_, _03857_);
  and (_03861_, _03839_, _03799_);
  and (_03862_, _03861_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and (_03863_, _03831_, _03799_);
  and (_03864_, _03863_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or (_03865_, _03864_, _03862_);
  or (_03866_, _03865_, _03860_);
  and (_03867_, _03821_, _03799_);
  and (_03868_, _03867_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and (_03869_, _03855_, _03799_);
  and (_03870_, _03869_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  or (_03871_, _03870_, _03868_);
  and (_03872_, _03845_, _03799_);
  and (_03873_, _03872_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and (_03874_, _03848_, _03799_);
  and (_03875_, _03874_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  or (_03876_, _03875_, _03873_);
  or (_03877_, _03876_, _03871_);
  or (_03878_, _03877_, _03866_);
  or (_03879_, _03878_, _03853_);
  and (_03880_, _03801_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  and (_03881_, _03816_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  or (_03882_, _03881_, _03880_);
  and (_03883_, _03832_, _03805_);
  and (_03884_, _03883_, _03789_);
  and (_03885_, _03884_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_03886_, _03788_, _03348_);
  and (_03887_, _03886_, _03799_);
  and (_03888_, _03887_, _38227_);
  or (_03889_, _03888_, _03885_);
  or (_03890_, _03889_, _03882_);
  and (_03891_, _03828_, _03789_);
  and (_03892_, _03891_, _03553_);
  and (_03893_, _03833_, _03789_);
  and (_03894_, _03893_, _03629_);
  or (_03895_, _03894_, _03892_);
  and (_03896_, _03799_, _03789_);
  and (_03897_, _03896_, _03494_);
  and (_03898_, _03854_, _03789_);
  and (_03899_, _03898_, _03761_);
  or (_03900_, _03899_, _03897_);
  or (_03901_, _03900_, _03895_);
  or (_03902_, _03901_, _03890_);
  and (_03903_, _03791_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_03904_, _03808_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or (_03905_, _03904_, _03903_);
  or (_03906_, _03905_, _03902_);
  or (_03907_, _03906_, _03879_);
  and (_03908_, _03907_, _03814_);
  not (_03909_, _03814_);
  nor (_03910_, _03842_, _03840_);
  nor (_03911_, _03849_, _03846_);
  and (_03912_, _03911_, _03910_);
  nor (_03913_, _03825_, _03822_);
  nor (_03914_, _03834_, _03829_);
  and (_03915_, _03914_, _03913_);
  and (_03916_, _03915_, _03912_);
  nor (_03917_, _03869_, _03867_);
  nor (_03918_, _03874_, _03872_);
  and (_03919_, _03918_, _03917_);
  nor (_03920_, _03863_, _03861_);
  nor (_03921_, _03858_, _03856_);
  and (_03922_, _03921_, _03920_);
  and (_03923_, _03922_, _03919_);
  and (_03924_, _03923_, _03916_);
  nor (_03925_, _03816_, _03801_);
  nor (_03926_, _03887_, _03884_);
  and (_03928_, _03926_, _03925_);
  nor (_03929_, _03893_, _03891_);
  nor (_03930_, _03898_, _03896_);
  and (_03931_, _03930_, _03929_);
  and (_03932_, _03931_, _03928_);
  nor (_03933_, _03808_, _03791_);
  and (_03934_, _03933_, _03932_);
  and (_03935_, _03934_, _03924_);
  or (_03936_, _03935_, _03909_);
  and (_03937_, _03936_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  or (_03938_, _03937_, _03908_);
  or (_03939_, _03938_, _03817_);
  and (_03940_, _03939_, _42618_);
  and (_39684_, _03940_, _03819_);
  nor (_39764_, \oc8051_top_1.oc8051_sfr1.prescaler [0], rst);
  or (_03941_, \oc8051_top_1.oc8051_sfr1.prescaler [0], \oc8051_top_1.oc8051_sfr1.prescaler [1]);
  nor (_03942_, _03330_, rst);
  and (_39765_, _03942_, _03941_);
  nor (_03943_, _03330_, _03329_);
  or (_03944_, _03943_, _03331_);
  and (_03945_, _03334_, _42618_);
  and (_39766_, _03945_, _03944_);
  nand (_03946_, _03840_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  nand (_03947_, _03842_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and (_03948_, _03947_, _03946_);
  nand (_03949_, _03846_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nand (_03950_, _03849_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  and (_03951_, _03950_, _03949_);
  and (_03952_, _03951_, _03948_);
  nand (_03953_, _03825_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  nand (_03954_, _03822_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  and (_03955_, _03954_, _03953_);
  nand (_03956_, _03829_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  nand (_03957_, _03834_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_03958_, _03957_, _03956_);
  and (_03959_, _03958_, _03955_);
  and (_03960_, _03959_, _03952_);
  nand (_03961_, _03867_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nand (_03962_, _03869_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_03963_, _03962_, _03961_);
  nand (_03964_, _03872_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  nand (_03965_, _03874_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and (_03966_, _03965_, _03964_);
  and (_03967_, _03966_, _03963_);
  nand (_03968_, _03861_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand (_03969_, _03863_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  and (_03970_, _03969_, _03968_);
  nand (_03971_, _03856_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  nand (_03972_, _03858_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  and (_03973_, _03972_, _03971_);
  and (_03974_, _03973_, _03970_);
  and (_03975_, _03974_, _03967_);
  and (_03976_, _03975_, _03960_);
  nand (_03977_, _03816_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  nand (_03978_, _03801_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and (_03979_, _03978_, _03977_);
  nand (_03980_, _03884_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nand (_03981_, _03887_, _42395_);
  and (_03982_, _03981_, _03980_);
  and (_03983_, _03982_, _03979_);
  nand (_03984_, _03891_, _03570_);
  nand (_03985_, _03893_, _03646_);
  and (_03986_, _03985_, _03984_);
  nand (_03987_, _03898_, _03767_);
  nand (_03988_, _03896_, _03479_);
  and (_03989_, _03988_, _03987_);
  and (_03990_, _03989_, _03986_);
  and (_03991_, _03990_, _03983_);
  not (_03992_, _03808_);
  or (_03993_, _03992_, _03394_);
  nand (_03994_, _03791_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and (_03995_, _03994_, _03993_);
  and (_03996_, _03995_, _03991_);
  and (_03997_, _03996_, _03976_);
  nor (_03998_, _03997_, _03909_);
  not (_03999_, _03817_);
  nand (_04000_, _03936_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  nand (_04001_, _04000_, _03999_);
  or (_04002_, _04001_, _03998_);
  nand (_04003_, _03817_, _32323_);
  and (_04004_, _04003_, _42618_);
  and (_39768_, _04004_, _04002_);
  nand (_04005_, _03817_, _33020_);
  or (_04006_, _03798_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  and (_04007_, _03840_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and (_04008_, _03842_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or (_04009_, _04008_, _04007_);
  and (_04010_, _03849_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and (_04011_, _03846_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  or (_04012_, _04011_, _04010_);
  or (_04013_, _04012_, _04009_);
  and (_04014_, _03825_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  and (_04015_, _03822_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  or (_04016_, _04015_, _04014_);
  and (_04017_, _03829_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_04018_, _03834_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  or (_04019_, _04018_, _04017_);
  or (_04020_, _04019_, _04016_);
  or (_04021_, _04020_, _04013_);
  and (_04022_, _03867_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  and (_04024_, _03869_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  or (_04025_, _04024_, _04022_);
  and (_04026_, _03872_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and (_04027_, _03874_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  or (_04028_, _04027_, _04026_);
  or (_04029_, _04028_, _04025_);
  and (_04030_, _03856_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  and (_04031_, _03858_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  or (_04032_, _04031_, _04030_);
  and (_04033_, _03861_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and (_04034_, _03863_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  or (_04035_, _04034_, _04033_);
  or (_04036_, _04035_, _04032_);
  or (_04037_, _04036_, _04029_);
  or (_04038_, _04037_, _04021_);
  and (_04039_, _03801_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  and (_04040_, _03816_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  or (_04041_, _04040_, _04039_);
  and (_04042_, _03884_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_04043_, _03887_, _42302_);
  or (_04044_, _04043_, _04042_);
  or (_04045_, _04044_, _04041_);
  and (_04046_, _03891_, _03584_);
  and (_04047_, _03893_, _03639_);
  or (_04048_, _04047_, _04046_);
  and (_04049_, _03896_, _03505_);
  and (_04050_, _03898_, _03741_);
  or (_04051_, _04050_, _04049_);
  or (_04052_, _04051_, _04048_);
  or (_04053_, _04052_, _04045_);
  and (_04054_, _03791_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_04055_, _03808_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  or (_04056_, _04055_, _04054_);
  or (_04057_, _04056_, _04053_);
  or (_04058_, _04057_, _04038_);
  and (_04059_, _04058_, _03813_);
  and (_04060_, _03936_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  or (_04061_, _04060_, _04059_);
  and (_04062_, _04061_, _04006_);
  or (_04063_, _04062_, _03817_);
  and (_04064_, _04063_, _42618_);
  and (_39769_, _04064_, _04005_);
  nand (_04065_, _03817_, _33717_);
  or (_04066_, _03798_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  and (_04067_, _03858_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  and (_04068_, _03856_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  or (_04069_, _04068_, _04067_);
  and (_04070_, _03861_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_04071_, _03863_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  or (_04072_, _04071_, _04070_);
  or (_04073_, _04072_, _04069_);
  and (_04074_, _03867_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  and (_04075_, _03869_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  or (_04076_, _04075_, _04074_);
  and (_04077_, _03872_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_04078_, _03874_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  or (_04079_, _04078_, _04077_);
  or (_04080_, _04079_, _04076_);
  or (_04081_, _04080_, _04073_);
  and (_04082_, _03842_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and (_04083_, _03840_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or (_04084_, _04083_, _04082_);
  and (_04085_, _03846_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and (_04086_, _03849_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  or (_04087_, _04086_, _04085_);
  or (_04088_, _04087_, _04084_);
  and (_04089_, _03825_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and (_04090_, _03822_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  or (_04091_, _04090_, _04089_);
  and (_04092_, _03829_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and (_04093_, _03834_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_04094_, _04093_, _04092_);
  or (_04095_, _04094_, _04091_);
  or (_04096_, _04095_, _04088_);
  or (_04097_, _04096_, _04081_);
  and (_04098_, _03801_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  and (_04099_, _03816_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  or (_04100_, _04099_, _04098_);
  and (_04101_, _03884_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_04102_, _03887_, _42192_);
  or (_04103_, _04102_, _04101_);
  or (_04104_, _04103_, _04100_);
  and (_04105_, _03891_, _03563_);
  and (_04106_, _03893_, _03660_);
  or (_04107_, _04106_, _04105_);
  and (_04108_, _03898_, _03747_);
  and (_04109_, _03896_, _03511_);
  or (_04110_, _04109_, _04108_);
  or (_04111_, _04110_, _04107_);
  or (_04112_, _04111_, _04104_);
  and (_04113_, _03808_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  and (_04114_, _03791_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_04115_, _04114_, _04113_);
  or (_04116_, _04115_, _04112_);
  or (_04117_, _04116_, _04097_);
  and (_04118_, _04117_, _03813_);
  and (_04119_, _03936_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  or (_04120_, _04119_, _04118_);
  and (_04121_, _04120_, _04066_);
  or (_04122_, _04121_, _03817_);
  and (_04124_, _04122_, _42618_);
  and (_39770_, _04124_, _04065_);
  nand (_04125_, _03817_, _34478_);
  and (_04126_, _03840_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and (_04127_, _03842_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  or (_04128_, _04127_, _04126_);
  and (_04129_, _03846_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and (_04130_, _03849_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  or (_04131_, _04130_, _04129_);
  or (_04132_, _04131_, _04128_);
  and (_04133_, _03825_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and (_04134_, _03822_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  or (_04135_, _04134_, _04133_);
  and (_04136_, _03829_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_04137_, _03834_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  or (_04138_, _04137_, _04136_);
  or (_04139_, _04138_, _04135_);
  or (_04140_, _04139_, _04132_);
  and (_04141_, _03867_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  and (_04142_, _03869_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  or (_04143_, _04142_, _04141_);
  and (_04144_, _03872_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and (_04145_, _03874_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  or (_04146_, _04145_, _04144_);
  or (_04147_, _04146_, _04143_);
  and (_04148_, _03856_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  and (_04149_, _03858_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  or (_04150_, _04149_, _04148_);
  and (_04151_, _03861_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_04152_, _03863_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  or (_04153_, _04152_, _04151_);
  or (_04154_, _04153_, _04150_);
  or (_04155_, _04154_, _04147_);
  or (_04156_, _04155_, _04140_);
  and (_04157_, _03816_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_04158_, _03801_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_04159_, _04158_, _04157_);
  and (_04160_, _03884_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_04161_, _03887_, _42331_);
  or (_04162_, _04161_, _04160_);
  or (_04163_, _04162_, _04159_);
  and (_04164_, _03891_, _03549_);
  and (_04165_, _03893_, _03625_);
  or (_04166_, _04165_, _04164_);
  and (_04167_, _03896_, _03490_);
  and (_04168_, _03898_, _03757_);
  or (_04169_, _04168_, _04167_);
  or (_04170_, _04169_, _04166_);
  or (_04171_, _04170_, _04163_);
  and (_04172_, _03791_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_04173_, _03808_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  or (_04174_, _04173_, _04172_);
  or (_04175_, _04174_, _04171_);
  or (_04176_, _04175_, _04156_);
  and (_04177_, _04176_, _03814_);
  and (_04178_, _03936_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  or (_04179_, _04178_, _04177_);
  or (_04180_, _04179_, _03817_);
  and (_04181_, _04180_, _42618_);
  and (_39771_, _04181_, _04125_);
  nand (_04182_, _03817_, _35240_);
  nand (_04183_, _03842_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  nand (_04184_, _03840_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and (_04185_, _04184_, _04183_);
  nand (_04186_, _03846_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  nand (_04187_, _03849_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and (_04188_, _04187_, _04186_);
  and (_04189_, _04188_, _04185_);
  nand (_04190_, _03822_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  nand (_04191_, _03825_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and (_04192_, _04191_, _04190_);
  nand (_04193_, _03829_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  nand (_04194_, _03834_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_04195_, _04194_, _04193_);
  and (_04196_, _04195_, _04192_);
  and (_04197_, _04196_, _04189_);
  nand (_04198_, _03869_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  nand (_04199_, _03867_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and (_04200_, _04199_, _04198_);
  nand (_04201_, _03872_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nand (_04202_, _03874_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and (_04203_, _04202_, _04201_);
  and (_04204_, _04203_, _04200_);
  nand (_04205_, _03858_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  nand (_04206_, _03856_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  and (_04207_, _04206_, _04205_);
  nand (_04208_, _03861_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nand (_04209_, _03863_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  and (_04210_, _04209_, _04208_);
  and (_04211_, _04210_, _04207_);
  and (_04212_, _04211_, _04204_);
  and (_04213_, _04212_, _04197_);
  nand (_04214_, _03801_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  nand (_04215_, _03816_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_04216_, _04215_, _04214_);
  nand (_04217_, _03884_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nand (_04218_, _03887_, _42237_);
  and (_04219_, _04218_, _04217_);
  and (_04220_, _04219_, _04216_);
  nand (_04221_, _03891_, _03574_);
  nand (_04223_, _03893_, _03650_);
  and (_04224_, _04223_, _04221_);
  nand (_04225_, _03896_, _03483_);
  nand (_04226_, _03898_, _03771_);
  and (_04227_, _04226_, _04225_);
  and (_04228_, _04227_, _04224_);
  and (_04229_, _04228_, _04220_);
  nand (_04230_, _03791_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nand (_04231_, _03808_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_04232_, _04231_, _04230_);
  and (_04233_, _04232_, _04229_);
  nand (_04234_, _04233_, _04213_);
  and (_04235_, _04234_, _03814_);
  and (_04236_, _03936_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  or (_04237_, _04236_, _03817_);
  or (_04238_, _04237_, _04235_);
  and (_04239_, _04238_, _42618_);
  and (_39772_, _04239_, _04182_);
  nand (_04240_, _03817_, _36046_);
  and (_04241_, _03856_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  and (_04242_, _03858_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  or (_04243_, _04242_, _04241_);
  and (_04244_, _03861_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_04245_, _03863_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  or (_04246_, _04245_, _04244_);
  or (_04247_, _04246_, _04243_);
  and (_04248_, _03867_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and (_04249_, _03869_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  or (_04250_, _04249_, _04248_);
  and (_04251_, _03872_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and (_04252_, _03874_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  or (_04253_, _04252_, _04251_);
  or (_04254_, _04253_, _04250_);
  or (_04255_, _04254_, _04247_);
  and (_04256_, _03825_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and (_04257_, _03822_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  or (_04258_, _04257_, _04256_);
  and (_04259_, _03829_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and (_04260_, _03834_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  or (_04261_, _04260_, _04259_);
  or (_04262_, _04261_, _04258_);
  and (_04263_, _03842_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and (_04264_, _03840_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or (_04265_, _04264_, _04263_);
  and (_04266_, _03846_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  and (_04267_, _03849_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  or (_04268_, _04267_, _04266_);
  or (_04269_, _04268_, _04265_);
  or (_04270_, _04269_, _04262_);
  or (_04271_, _04270_, _04255_);
  and (_04272_, _03801_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  and (_04273_, _03816_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  or (_04274_, _04273_, _04272_);
  and (_04275_, _03884_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_04276_, _03887_, _42137_);
  or (_04277_, _04276_, _04275_);
  or (_04278_, _04277_, _04274_);
  and (_04279_, _03891_, _03580_);
  and (_04280_, _03893_, _03635_);
  or (_04281_, _04280_, _04279_);
  and (_04282_, _03898_, _03737_);
  and (_04283_, _03896_, _03501_);
  or (_04284_, _04283_, _04282_);
  or (_04285_, _04284_, _04281_);
  or (_04286_, _04285_, _04278_);
  and (_04287_, _03791_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_04288_, _03808_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  or (_04289_, _04288_, _04287_);
  or (_04290_, _04289_, _04286_);
  or (_04291_, _04290_, _04271_);
  and (_04292_, _04291_, _03814_);
  and (_04293_, _03936_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  or (_04294_, _04293_, _04292_);
  or (_04295_, _04294_, _03817_);
  and (_04296_, _04295_, _42618_);
  and (_39773_, _04296_, _04240_);
  and (_04297_, _03936_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  and (_04298_, _03856_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  and (_04299_, _03858_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  or (_04300_, _04299_, _04298_);
  and (_04301_, _03863_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  and (_04302_, _03861_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or (_04303_, _04302_, _04301_);
  or (_04304_, _04303_, _04300_);
  and (_04305_, _03867_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and (_04306_, _03869_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  or (_04307_, _04306_, _04305_);
  and (_04308_, _03872_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and (_04309_, _03874_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  or (_04310_, _04309_, _04308_);
  or (_04311_, _04310_, _04307_);
  or (_04312_, _04311_, _04304_);
  and (_04313_, _03840_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and (_04314_, _03842_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or (_04315_, _04314_, _04313_);
  and (_04316_, _03849_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and (_04317_, _03846_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or (_04318_, _04317_, _04316_);
  or (_04319_, _04318_, _04315_);
  and (_04320_, _03825_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and (_04322_, _03822_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  or (_04323_, _04322_, _04320_);
  and (_04324_, _03829_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_04325_, _03834_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  or (_04326_, _04325_, _04324_);
  or (_04327_, _04326_, _04323_);
  or (_04328_, _04327_, _04319_);
  or (_04329_, _04328_, _04312_);
  and (_04330_, _03801_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  and (_04331_, _03816_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  or (_04332_, _04331_, _04330_);
  and (_04333_, _03884_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_04334_, _03887_, _42408_);
  or (_04335_, _04334_, _04333_);
  or (_04336_, _04335_, _04332_);
  and (_04337_, _03891_, _03559_);
  and (_04338_, _03893_, _03656_);
  or (_04339_, _04338_, _04337_);
  and (_04340_, _03896_, _03515_);
  and (_04341_, _03898_, _03751_);
  or (_04342_, _04341_, _04340_);
  or (_04343_, _04342_, _04339_);
  or (_04344_, _04343_, _04336_);
  and (_04345_, _03808_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_04346_, _03791_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_04347_, _04346_, _04345_);
  or (_04348_, _04347_, _04344_);
  or (_04349_, _04348_, _04329_);
  and (_04350_, _04349_, _03814_);
  or (_04351_, _04350_, _04297_);
  and (_04352_, _04351_, _03999_);
  and (_04353_, _03817_, _36698_);
  or (_04354_, _04353_, _04352_);
  and (_39774_, _04354_, _42618_);
  and (_39843_, _42558_, _42618_);
  nor (_39846_, _42212_, rst);
  and (_39867_, _42648_, _42618_);
  and (_39868_, _42658_, _42618_);
  nor (_39871_, _42400_, rst);
  nor (_39872_, _42307_, rst);
  not (_04355_, _00342_);
  nor (_04356_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  not (_04357_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_04358_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _04357_);
  nor (_04359_, _04358_, _04356_);
  nor (_04360_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_04361_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _04357_);
  nor (_04362_, _04361_, _04360_);
  nor (_04363_, _04362_, _04359_);
  and (_04364_, _04362_, _04359_);
  nor (_04365_, _02227_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_04366_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _04357_);
  nor (_04367_, _04366_, _04365_);
  and (_04368_, _04367_, _04364_);
  nor (_04369_, _04367_, _04364_);
  nor (_04370_, _04369_, _04368_);
  nor (_04371_, _02246_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_04372_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _04357_);
  nor (_04373_, _04372_, _04371_);
  not (_04374_, _04373_);
  and (_04375_, _04374_, _04368_);
  nor (_04376_, _04374_, _04368_);
  nor (_04377_, _04376_, _04375_);
  nor (_04378_, _04377_, _04370_);
  and (_04379_, _04378_, _04363_);
  and (_04380_, _04379_, _04355_);
  not (_04381_, _43516_);
  not (_04382_, _04370_);
  and (_04383_, _04377_, _04382_);
  and (_04384_, _04383_, _04363_);
  and (_04385_, _04384_, _04381_);
  or (_04386_, _04385_, _04380_);
  not (_04387_, _00424_);
  not (_04388_, _04359_);
  and (_04389_, _04362_, _04388_);
  and (_04390_, _04378_, _04389_);
  and (_04391_, _04390_, _04387_);
  not (_04392_, _00065_);
  and (_04393_, _04383_, _04389_);
  and (_04394_, _04393_, _04392_);
  or (_04395_, _04394_, _04391_);
  or (_04396_, _04395_, _04386_);
  not (_04397_, _00168_);
  and (_04398_, _04374_, _04370_);
  and (_04399_, _04398_, _04363_);
  and (_04400_, _04399_, _04397_);
  not (_04401_, _00550_);
  nor (_04402_, _04362_, _04388_);
  and (_04403_, _04373_, _04370_);
  and (_04404_, _04403_, _04402_);
  and (_04405_, _04404_, _04401_);
  not (_04406_, _00106_);
  and (_04407_, _04398_, _04364_);
  and (_04408_, _04407_, _04406_);
  or (_04409_, _04408_, _04405_);
  or (_04410_, _04409_, _04400_);
  not (_04411_, _00465_);
  and (_04412_, _04376_, _04364_);
  and (_04413_, _04412_, _04411_);
  not (_04415_, _00260_);
  and (_04416_, _04367_, _04389_);
  and (_04417_, _04416_, _04374_);
  and (_04418_, _04417_, _04415_);
  not (_04419_, _43475_);
  and (_04420_, _04373_, _04368_);
  and (_04421_, _04420_, _04419_);
  or (_04422_, _04421_, _04418_);
  not (_04423_, _00607_);
  and (_04424_, _04416_, _04373_);
  and (_04425_, _04424_, _04423_);
  not (_04426_, _00301_);
  and (_04427_, _04375_, _04426_);
  or (_04428_, _04427_, _04425_);
  or (_04429_, _04428_, _04422_);
  or (_04430_, _04429_, _04413_);
  not (_04431_, _00506_);
  and (_04432_, _04403_, _04363_);
  and (_04433_, _04432_, _04431_);
  not (_04434_, _00219_);
  and (_04435_, _04398_, _04402_);
  and (_04436_, _04435_, _04434_);
  or (_04437_, _04436_, _04433_);
  or (_04438_, _04437_, _04430_);
  not (_04439_, _00383_);
  and (_04440_, _04378_, _04402_);
  and (_04441_, _04440_, _04439_);
  not (_04442_, _00024_);
  and (_04443_, _04383_, _04402_);
  and (_04444_, _04443_, _04442_);
  or (_04445_, _04444_, _04441_);
  or (_04446_, _04445_, _04438_);
  or (_04447_, _04446_, _04410_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [15], _04447_, _04396_);
  and (_04448_, _04393_, _04406_);
  and (_04449_, _04384_, _04442_);
  or (_04450_, _04449_, _04448_);
  and (_04451_, _04440_, _04387_);
  and (_04452_, _04443_, _04392_);
  or (_04453_, _04452_, _04451_);
  or (_04454_, _04453_, _04450_);
  and (_04455_, _04404_, _04423_);
  and (_04456_, _04432_, _04401_);
  and (_04457_, _04435_, _04415_);
  or (_04458_, _04457_, _04456_);
  or (_04459_, _04458_, _04455_);
  and (_04460_, _04407_, _04397_);
  and (_04461_, _04399_, _04434_);
  or (_04462_, _04461_, _04460_);
  and (_04463_, _04412_, _04431_);
  and (_04464_, _04375_, _04355_);
  and (_04465_, _04424_, _04419_);
  or (_04466_, _04465_, _04464_);
  and (_04467_, _04417_, _04426_);
  and (_04468_, _04420_, _04381_);
  or (_04469_, _04468_, _04467_);
  or (_04470_, _04469_, _04466_);
  or (_04471_, _04470_, _04463_);
  or (_04472_, _04471_, _04462_);
  and (_04473_, _04390_, _04411_);
  and (_04474_, _04379_, _04439_);
  or (_04475_, _04474_, _04473_);
  or (_04476_, _04475_, _04472_);
  or (_04477_, _04476_, _04459_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [23], _04477_, _04454_);
  and (_04478_, _04379_, _04387_);
  and (_04479_, _04384_, _04392_);
  or (_04480_, _04479_, _04478_);
  and (_04481_, _04393_, _04397_);
  and (_04482_, _04443_, _04406_);
  or (_04483_, _04482_, _04481_);
  or (_04484_, _04483_, _04480_);
  and (_04485_, _04435_, _04426_);
  and (_04486_, _04407_, _04434_);
  and (_04487_, _04404_, _04419_);
  or (_04488_, _04487_, _04486_);
  or (_04489_, _04488_, _04485_);
  and (_04490_, _04412_, _04401_);
  and (_04491_, _04417_, _04355_);
  and (_04492_, _04420_, _04442_);
  or (_04493_, _04492_, _04491_);
  and (_04494_, _04375_, _04439_);
  and (_04495_, _04424_, _04381_);
  or (_04496_, _04495_, _04494_);
  or (_04497_, _04496_, _04493_);
  or (_04498_, _04497_, _04490_);
  and (_04499_, _04432_, _04423_);
  and (_04500_, _04399_, _04415_);
  or (_04501_, _04500_, _04499_);
  or (_04502_, _04501_, _04498_);
  and (_04503_, _04440_, _04411_);
  and (_04504_, _04390_, _04431_);
  or (_04505_, _04504_, _04503_);
  or (_04506_, _04505_, _04502_);
  or (_04507_, _04506_, _04489_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [31], _04507_, _04484_);
  and (_04508_, _04440_, _04355_);
  and (_04509_, _04384_, _04419_);
  or (_04510_, _04509_, _04508_);
  and (_04511_, _04379_, _04426_);
  and (_04513_, _04443_, _04381_);
  or (_04514_, _04513_, _04511_);
  or (_04515_, _04514_, _04510_);
  and (_04516_, _04407_, _04392_);
  and (_04517_, _04399_, _04406_);
  or (_04518_, _04517_, _04516_);
  and (_04519_, _04435_, _04397_);
  or (_04520_, _04519_, _04518_);
  and (_04521_, _04412_, _04387_);
  and (_04522_, _04424_, _04401_);
  and (_04523_, _04375_, _04415_);
  or (_04524_, _04523_, _04522_);
  and (_04525_, _04420_, _04423_);
  and (_04526_, _04417_, _04434_);
  or (_04527_, _04526_, _04525_);
  or (_04528_, _04527_, _04524_);
  or (_04529_, _04528_, _04521_);
  and (_04530_, _04404_, _04431_);
  and (_04531_, _04432_, _04411_);
  or (_04532_, _04531_, _04530_);
  or (_04533_, _04532_, _04529_);
  and (_04534_, _04390_, _04439_);
  and (_04535_, _04393_, _04442_);
  or (_04536_, _04535_, _04534_);
  or (_04537_, _04536_, _04533_);
  or (_04538_, _04537_, _04520_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [7], _04538_, _04515_);
  not (_04539_, _00029_);
  and (_04540_, _04393_, _04539_);
  not (_04541_, _00388_);
  and (_04542_, _04390_, _04541_);
  or (_04543_, _04542_, _04540_);
  not (_04544_, _43480_);
  and (_04545_, _04384_, _04544_);
  not (_04546_, _00306_);
  and (_04547_, _04379_, _04546_);
  or (_04548_, _04547_, _04545_);
  or (_04549_, _04548_, _04543_);
  not (_04550_, _00470_);
  and (_04551_, _04432_, _04550_);
  not (_04552_, _00179_);
  and (_04553_, _04435_, _04552_);
  not (_04554_, _00511_);
  and (_04555_, _04404_, _04554_);
  or (_04556_, _04555_, _04553_);
  or (_04557_, _04556_, _04551_);
  not (_04558_, _00070_);
  and (_04559_, _04407_, _04558_);
  not (_04560_, _00111_);
  and (_04561_, _04399_, _04560_);
  or (_04562_, _04561_, _04559_);
  not (_04563_, _00429_);
  and (_04564_, _04412_, _04563_);
  not (_04565_, _00612_);
  and (_04566_, _04420_, _04565_);
  not (_04567_, _00265_);
  and (_04568_, _04375_, _04567_);
  or (_04569_, _04568_, _04566_);
  not (_04570_, _00224_);
  and (_04571_, _04417_, _04570_);
  not (_04572_, _00558_);
  and (_04573_, _04424_, _04572_);
  or (_04574_, _04573_, _04571_);
  or (_04575_, _04574_, _04569_);
  or (_04576_, _04575_, _04564_);
  or (_04577_, _04576_, _04562_);
  not (_04578_, _43521_);
  and (_04579_, _04443_, _04578_);
  not (_04580_, _00347_);
  and (_04581_, _04440_, _04580_);
  or (_04582_, _04581_, _04579_);
  or (_04583_, _04582_, _04577_);
  or (_04584_, _04583_, _04557_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [0], _04584_, _04549_);
  not (_04585_, _00352_);
  and (_04586_, _04440_, _04585_);
  not (_04587_, _00311_);
  and (_04588_, _04379_, _04587_);
  or (_04589_, _04588_, _04586_);
  not (_04590_, _43485_);
  and (_04591_, _04384_, _04590_);
  not (_04592_, _00393_);
  and (_04593_, _04390_, _04592_);
  or (_04594_, _04593_, _04591_);
  or (_04595_, _04594_, _04589_);
  not (_04596_, _00516_);
  and (_04597_, _04404_, _04596_);
  not (_04598_, _00075_);
  and (_04599_, _04407_, _04598_);
  not (_04600_, _00475_);
  and (_04601_, _04432_, _04600_);
  or (_04602_, _04601_, _04599_);
  or (_04603_, _04602_, _04597_);
  not (_04604_, _43526_);
  and (_04605_, _04443_, _04604_);
  not (_04606_, _00034_);
  and (_04607_, _04393_, _04606_);
  or (_04608_, _04607_, _04605_);
  not (_04609_, _00434_);
  and (_04610_, _04412_, _04609_);
  not (_04612_, _00617_);
  and (_04613_, _04420_, _04612_);
  not (_04614_, _00270_);
  and (_04615_, _04375_, _04614_);
  or (_04616_, _04615_, _04613_);
  not (_04617_, _00229_);
  and (_04618_, _04417_, _04617_);
  not (_04619_, _00566_);
  and (_04620_, _04424_, _04619_);
  or (_04621_, _04620_, _04618_);
  or (_04622_, _04621_, _04616_);
  or (_04623_, _04622_, _04610_);
  not (_04624_, _00188_);
  and (_04625_, _04435_, _04624_);
  not (_04626_, _00116_);
  and (_04627_, _04399_, _04626_);
  or (_04628_, _04627_, _04625_);
  or (_04629_, _04628_, _04623_);
  or (_04630_, _04629_, _04608_);
  or (_04631_, _04630_, _04603_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [1], _04631_, _04595_);
  not (_04632_, _00316_);
  and (_04633_, _04379_, _04632_);
  not (_04634_, _43531_);
  and (_04635_, _04443_, _04634_);
  or (_04636_, _04635_, _04633_);
  not (_04637_, _00357_);
  and (_04638_, _04440_, _04637_);
  not (_04639_, _43490_);
  and (_04640_, _04384_, _04639_);
  or (_04641_, _04640_, _04638_);
  or (_04642_, _04641_, _04636_);
  not (_04643_, _00121_);
  and (_04644_, _04399_, _04643_);
  not (_04645_, _00521_);
  and (_04646_, _04404_, _04645_);
  not (_04647_, _00080_);
  and (_04648_, _04407_, _04647_);
  or (_04649_, _04648_, _04646_);
  or (_04650_, _04649_, _04644_);
  not (_04651_, _00439_);
  and (_04652_, _04412_, _04651_);
  not (_04653_, _00574_);
  and (_04654_, _04424_, _04653_);
  not (_04655_, _00275_);
  and (_04656_, _04375_, _04655_);
  or (_04657_, _04656_, _04654_);
  not (_04658_, _00622_);
  and (_04659_, _04420_, _04658_);
  not (_04660_, _00234_);
  and (_04661_, _04417_, _04660_);
  or (_04662_, _04661_, _04659_);
  or (_04663_, _04662_, _04657_);
  or (_04664_, _04663_, _04652_);
  not (_04665_, _00480_);
  and (_04666_, _04432_, _04665_);
  not (_04667_, _00193_);
  and (_04668_, _04435_, _04667_);
  or (_04669_, _04668_, _04666_);
  or (_04670_, _04669_, _04664_);
  not (_04671_, _00398_);
  and (_04672_, _04390_, _04671_);
  not (_04673_, _00039_);
  and (_04674_, _04393_, _04673_);
  or (_04675_, _04674_, _04672_);
  or (_04676_, _04675_, _04670_);
  or (_04677_, _04676_, _04650_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [2], _04677_, _04642_);
  not (_04678_, _00403_);
  and (_04679_, _04390_, _04678_);
  not (_04680_, _00003_);
  and (_04681_, _04443_, _04680_);
  or (_04682_, _04681_, _04679_);
  not (_04683_, _00321_);
  and (_04684_, _04379_, _04683_);
  not (_04685_, _43495_);
  and (_04686_, _04384_, _04685_);
  or (_04687_, _04686_, _04684_);
  or (_04688_, _04687_, _04682_);
  not (_04689_, _00526_);
  and (_04690_, _04404_, _04689_);
  not (_04691_, _00485_);
  and (_04692_, _04432_, _04691_);
  not (_04693_, _00085_);
  and (_04694_, _04407_, _04693_);
  or (_04695_, _04694_, _04692_);
  or (_04696_, _04695_, _04690_);
  not (_04697_, _00444_);
  and (_04698_, _04412_, _04697_);
  not (_04699_, _00627_);
  and (_04700_, _04420_, _04699_);
  not (_04701_, _00239_);
  and (_04702_, _04417_, _04701_);
  or (_04703_, _04702_, _04700_);
  not (_04704_, _00582_);
  and (_04705_, _04424_, _04704_);
  not (_04706_, _00280_);
  and (_04707_, _04375_, _04706_);
  or (_04708_, _04707_, _04705_);
  or (_04709_, _04708_, _04703_);
  or (_04710_, _04709_, _04698_);
  not (_04711_, _00198_);
  and (_04712_, _04435_, _04711_);
  not (_04713_, _00126_);
  and (_04714_, _04399_, _04713_);
  or (_04715_, _04714_, _04712_);
  or (_04716_, _04715_, _04710_);
  not (_04717_, _00362_);
  and (_04718_, _04440_, _04717_);
  not (_04719_, _00044_);
  and (_04720_, _04393_, _04719_);
  or (_04721_, _04720_, _04718_);
  or (_04722_, _04721_, _04716_);
  or (_04723_, _04722_, _04696_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [3], _04723_, _04688_);
  not (_04724_, _00326_);
  and (_04725_, _04379_, _04724_);
  not (_04726_, _00008_);
  and (_04727_, _04443_, _04726_);
  or (_04728_, _04727_, _04725_);
  not (_04729_, _00367_);
  and (_04730_, _04440_, _04729_);
  not (_04731_, _43500_);
  and (_04732_, _04384_, _04731_);
  or (_04733_, _04732_, _04730_);
  or (_04734_, _04733_, _04728_);
  not (_04735_, _00133_);
  and (_04736_, _04399_, _04735_);
  not (_04737_, _00531_);
  and (_04738_, _04404_, _04737_);
  not (_04739_, _00090_);
  and (_04740_, _04407_, _04739_);
  or (_04741_, _04740_, _04738_);
  or (_04742_, _04741_, _04736_);
  not (_04743_, _00449_);
  and (_04744_, _04412_, _04743_);
  not (_04745_, _00590_);
  and (_04746_, _04424_, _04745_);
  not (_04747_, _00285_);
  and (_04748_, _04375_, _04747_);
  or (_04749_, _04748_, _04746_);
  not (_04750_, _00632_);
  and (_04751_, _04420_, _04750_);
  not (_04752_, _00244_);
  and (_04753_, _04417_, _04752_);
  or (_04754_, _04753_, _04751_);
  or (_04755_, _04754_, _04749_);
  or (_04756_, _04755_, _04744_);
  not (_04757_, _00490_);
  and (_04758_, _04432_, _04757_);
  not (_04759_, _00203_);
  and (_04760_, _04435_, _04759_);
  or (_04761_, _04760_, _04758_);
  or (_04762_, _04761_, _04756_);
  not (_04763_, _00408_);
  and (_04764_, _04390_, _04763_);
  not (_04765_, _00049_);
  and (_04766_, _04393_, _04765_);
  or (_04767_, _04766_, _04764_);
  or (_04768_, _04767_, _04762_);
  or (_04769_, _04768_, _04742_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [4], _04769_, _04734_);
  not (_04770_, _00331_);
  and (_04771_, _04379_, _04770_);
  not (_04772_, _00013_);
  and (_04773_, _04443_, _04772_);
  or (_04774_, _04773_, _04771_);
  not (_04775_, _00372_);
  and (_04776_, _04440_, _04775_);
  not (_04777_, _43505_);
  and (_04778_, _04384_, _04777_);
  or (_04779_, _04778_, _04776_);
  or (_04780_, _04779_, _04774_);
  not (_04781_, _00095_);
  and (_04782_, _04407_, _04781_);
  not (_04783_, _00536_);
  and (_04784_, _04404_, _04783_);
  not (_04785_, _00495_);
  and (_04786_, _04432_, _04785_);
  or (_04787_, _04786_, _04784_);
  or (_04788_, _04787_, _04782_);
  not (_04789_, _00454_);
  and (_04790_, _04412_, _04789_);
  not (_04791_, _00596_);
  and (_04792_, _04424_, _04791_);
  not (_04793_, _00290_);
  and (_04794_, _04375_, _04793_);
  or (_04795_, _04794_, _04792_);
  not (_04796_, _00637_);
  and (_04797_, _04420_, _04796_);
  not (_04798_, _00249_);
  and (_04799_, _04417_, _04798_);
  or (_04800_, _04799_, _04797_);
  or (_04801_, _04800_, _04795_);
  or (_04802_, _04801_, _04790_);
  not (_04803_, _00208_);
  and (_04804_, _04435_, _04803_);
  not (_04805_, _00144_);
  and (_04806_, _04399_, _04805_);
  or (_04807_, _04806_, _04804_);
  or (_04808_, _04807_, _04802_);
  not (_04809_, _00413_);
  and (_04810_, _04390_, _04809_);
  not (_04811_, _00054_);
  and (_04812_, _04393_, _04811_);
  or (_04813_, _04812_, _04810_);
  or (_04814_, _04813_, _04808_);
  or (_04815_, _04814_, _04788_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [5], _04815_, _04780_);
  not (_04816_, _00336_);
  and (_04817_, _04379_, _04816_);
  not (_04818_, _00018_);
  and (_04819_, _04443_, _04818_);
  or (_04820_, _04819_, _04817_);
  not (_04821_, _00377_);
  and (_04822_, _04440_, _04821_);
  not (_04823_, _43510_);
  and (_04824_, _04384_, _04823_);
  or (_04825_, _04824_, _04822_);
  or (_04826_, _04825_, _04820_);
  not (_04827_, _00155_);
  and (_04828_, _04399_, _04827_);
  not (_04829_, _00541_);
  and (_04830_, _04404_, _04829_);
  not (_04831_, _00100_);
  and (_04832_, _04407_, _04831_);
  or (_04833_, _04832_, _04830_);
  or (_04834_, _04833_, _04828_);
  not (_04835_, _00459_);
  and (_04836_, _04412_, _04835_);
  not (_04837_, _00601_);
  and (_04838_, _04424_, _04837_);
  not (_04839_, _00295_);
  and (_04840_, _04375_, _04839_);
  or (_04841_, _04840_, _04838_);
  not (_04842_, _00642_);
  and (_04843_, _04420_, _04842_);
  not (_04844_, _00254_);
  and (_04845_, _04417_, _04844_);
  or (_04846_, _04845_, _04843_);
  or (_04847_, _04846_, _04841_);
  or (_04848_, _04847_, _04836_);
  not (_04849_, _00500_);
  and (_04850_, _04432_, _04849_);
  not (_04851_, _00213_);
  and (_04852_, _04435_, _04851_);
  or (_04853_, _04852_, _04850_);
  or (_04854_, _04853_, _04848_);
  not (_04855_, _00418_);
  and (_04856_, _04390_, _04855_);
  not (_04857_, _00059_);
  and (_04858_, _04393_, _04857_);
  or (_04859_, _04858_, _04856_);
  or (_04860_, _04859_, _04854_);
  or (_04861_, _04860_, _04834_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [6], _04861_, _04826_);
  and (_04862_, _04393_, _04552_);
  and (_04863_, _04384_, _04558_);
  or (_04864_, _04863_, _04862_);
  and (_04865_, _04390_, _04554_);
  and (_04866_, _04379_, _04563_);
  or (_04867_, _04866_, _04865_);
  or (_04868_, _04867_, _04864_);
  and (_04869_, _04404_, _04544_);
  and (_04870_, _04432_, _04565_);
  and (_04871_, _04435_, _04546_);
  or (_04872_, _04871_, _04870_);
  or (_04873_, _04872_, _04869_);
  and (_04874_, _04399_, _04567_);
  and (_04875_, _04407_, _04570_);
  or (_04876_, _04875_, _04874_);
  and (_04877_, _04412_, _04572_);
  and (_04878_, _04417_, _04580_);
  and (_04879_, _04420_, _04539_);
  or (_04880_, _04879_, _04878_);
  and (_04881_, _04375_, _04541_);
  and (_04882_, _04424_, _04578_);
  or (_04883_, _04882_, _04881_);
  or (_04884_, _04883_, _04880_);
  or (_04885_, _04884_, _04877_);
  or (_04886_, _04885_, _04876_);
  and (_04887_, _04440_, _04550_);
  and (_04888_, _04443_, _04560_);
  or (_04889_, _04888_, _04887_);
  or (_04890_, _04889_, _04886_);
  or (_04891_, _04890_, _04873_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [24], _04891_, _04868_);
  and (_04892_, _04384_, _04598_);
  and (_04893_, _04443_, _04626_);
  or (_04894_, _04893_, _04892_);
  and (_04895_, _04390_, _04596_);
  and (_04896_, _04393_, _04624_);
  or (_04897_, _04896_, _04895_);
  or (_04898_, _04897_, _04894_);
  and (_04899_, _04404_, _04590_);
  and (_04900_, _04432_, _04612_);
  and (_04901_, _04435_, _04587_);
  or (_04902_, _04901_, _04900_);
  or (_04903_, _04902_, _04899_);
  and (_04904_, _04440_, _04600_);
  and (_04905_, _04379_, _04609_);
  or (_04906_, _04905_, _04904_);
  and (_04907_, _04399_, _04614_);
  and (_04908_, _04407_, _04617_);
  or (_04909_, _04908_, _04907_);
  and (_04910_, _04412_, _04619_);
  and (_04911_, _04417_, _04585_);
  and (_04912_, _04375_, _04592_);
  or (_04913_, _04912_, _04911_);
  and (_04914_, _04424_, _04604_);
  and (_04915_, _04420_, _04606_);
  or (_04916_, _04915_, _04914_);
  or (_04917_, _04916_, _04913_);
  or (_04918_, _04917_, _04910_);
  or (_04919_, _04918_, _04909_);
  or (_04920_, _04919_, _04906_);
  or (_04921_, _04920_, _04903_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [25], _04921_, _04898_);
  and (_04922_, _04443_, _04643_);
  and (_04923_, _04384_, _04647_);
  or (_04924_, _04923_, _04922_);
  and (_04925_, _04390_, _04645_);
  and (_04926_, _04379_, _04651_);
  or (_04927_, _04926_, _04925_);
  or (_04928_, _04927_, _04924_);
  and (_04929_, _04435_, _04632_);
  and (_04930_, _04399_, _04655_);
  and (_04931_, _04404_, _04639_);
  or (_04932_, _04931_, _04930_);
  or (_04933_, _04932_, _04929_);
  and (_04934_, _04412_, _04653_);
  and (_04935_, _04375_, _04671_);
  and (_04936_, _04424_, _04634_);
  or (_04937_, _04936_, _04935_);
  and (_04938_, _04417_, _04637_);
  and (_04939_, _04420_, _04673_);
  or (_04940_, _04939_, _04938_);
  or (_04941_, _04940_, _04937_);
  or (_04942_, _04941_, _04934_);
  and (_04943_, _04432_, _04658_);
  and (_04944_, _04407_, _04660_);
  or (_04945_, _04944_, _04943_);
  or (_04946_, _04945_, _04942_);
  and (_04947_, _04440_, _04665_);
  and (_04948_, _04393_, _04667_);
  or (_04949_, _04948_, _04947_);
  or (_04950_, _04949_, _04946_);
  or (_04951_, _04950_, _04933_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [26], _04951_, _04928_);
  and (_04952_, _04440_, _04691_);
  and (_04953_, _04384_, _04693_);
  or (_04954_, _04953_, _04952_);
  and (_04955_, _04379_, _04697_);
  and (_04956_, _04443_, _04713_);
  or (_04957_, _04956_, _04955_);
  or (_04958_, _04957_, _04954_);
  and (_04959_, _04432_, _04699_);
  and (_04960_, _04435_, _04683_);
  and (_04961_, _04404_, _04685_);
  or (_04962_, _04961_, _04960_);
  or (_04963_, _04962_, _04959_);
  and (_04964_, _04399_, _04706_);
  and (_04965_, _04407_, _04701_);
  or (_04966_, _04965_, _04964_);
  and (_04967_, _04412_, _04704_);
  and (_04968_, _04417_, _04717_);
  and (_04969_, _04420_, _04719_);
  or (_04970_, _04969_, _04968_);
  and (_04971_, _04375_, _04678_);
  and (_04972_, _04424_, _04680_);
  or (_04973_, _04972_, _04971_);
  or (_04974_, _04973_, _04970_);
  or (_04975_, _04974_, _04967_);
  or (_04976_, _04975_, _04966_);
  and (_04977_, _04390_, _04689_);
  and (_04978_, _04393_, _04711_);
  or (_04979_, _04978_, _04977_);
  or (_04980_, _04979_, _04976_);
  or (_04981_, _04980_, _04963_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [27], _04981_, _04958_);
  and (_04982_, _04379_, _04743_);
  and (_04983_, _04384_, _04739_);
  or (_04984_, _04983_, _04982_);
  and (_04985_, _04393_, _04759_);
  and (_04986_, _04443_, _04735_);
  or (_04987_, _04986_, _04985_);
  or (_04988_, _04987_, _04984_);
  and (_04989_, _04435_, _04724_);
  and (_04990_, _04407_, _04752_);
  and (_04991_, _04404_, _04731_);
  or (_04992_, _04991_, _04990_);
  or (_04993_, _04992_, _04989_);
  and (_04994_, _04412_, _04745_);
  and (_04995_, _04417_, _04729_);
  and (_04996_, _04420_, _04765_);
  or (_04997_, _04996_, _04995_);
  and (_04998_, _04375_, _04763_);
  and (_04999_, _04424_, _04726_);
  or (_05000_, _04999_, _04998_);
  or (_05001_, _05000_, _04997_);
  or (_05002_, _05001_, _04994_);
  and (_05003_, _04432_, _04750_);
  and (_05004_, _04399_, _04747_);
  or (_05005_, _05004_, _05003_);
  or (_05006_, _05005_, _05002_);
  and (_05007_, _04440_, _04757_);
  and (_05008_, _04390_, _04737_);
  or (_05009_, _05008_, _05007_);
  or (_05010_, _05009_, _05006_);
  or (_05011_, _05010_, _04993_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [28], _05011_, _04988_);
  and (_05012_, _04443_, _04805_);
  and (_05013_, _04384_, _04781_);
  or (_05014_, _05013_, _05012_);
  and (_05015_, _04440_, _04785_);
  and (_05016_, _04393_, _04803_);
  or (_05017_, _05016_, _05015_);
  or (_05018_, _05017_, _05014_);
  and (_05019_, _04407_, _04798_);
  and (_05020_, _04435_, _04770_);
  and (_05021_, _04404_, _04777_);
  or (_05022_, _05021_, _05020_);
  or (_05023_, _05022_, _05019_);
  and (_05024_, _04412_, _04791_);
  and (_05025_, _04375_, _04809_);
  and (_05026_, _04424_, _04772_);
  or (_05027_, _05026_, _05025_);
  and (_05028_, _04417_, _04775_);
  and (_05029_, _04420_, _04811_);
  or (_05030_, _05029_, _05028_);
  or (_05031_, _05030_, _05027_);
  or (_05032_, _05031_, _05024_);
  and (_05033_, _04432_, _04796_);
  and (_05034_, _04399_, _04793_);
  or (_05035_, _05034_, _05033_);
  or (_05036_, _05035_, _05032_);
  and (_05037_, _04379_, _04789_);
  and (_05038_, _04390_, _04783_);
  or (_05039_, _05038_, _05037_);
  or (_05040_, _05039_, _05036_);
  or (_05041_, _05040_, _05023_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [29], _05041_, _05018_);
  and (_05042_, _04443_, _04827_);
  and (_05043_, _04384_, _04831_);
  or (_05044_, _05043_, _05042_);
  and (_05045_, _04390_, _04829_);
  and (_05046_, _04379_, _04835_);
  or (_05047_, _05046_, _05045_);
  or (_05048_, _05047_, _05044_);
  and (_05049_, _04407_, _04844_);
  and (_05050_, _04432_, _04842_);
  and (_05051_, _04404_, _04823_);
  or (_05052_, _05051_, _05050_);
  or (_05054_, _05052_, _05049_);
  and (_05056_, _04399_, _04839_);
  and (_05058_, _04435_, _04816_);
  or (_05060_, _05058_, _05056_);
  and (_05062_, _04412_, _04837_);
  and (_05064_, _04417_, _04821_);
  and (_05066_, _04420_, _04857_);
  or (_05067_, _05066_, _05064_);
  and (_05068_, _04375_, _04855_);
  and (_05069_, _04424_, _04818_);
  or (_05070_, _05069_, _05068_);
  or (_05071_, _05070_, _05067_);
  or (_05072_, _05071_, _05062_);
  or (_05074_, _05072_, _05060_);
  and (_05075_, _04440_, _04849_);
  and (_05077_, _04393_, _04851_);
  or (_05078_, _05077_, _05075_);
  or (_05079_, _05078_, _05074_);
  or (_05081_, _05079_, _05054_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [30], _05081_, _05048_);
  and (_05082_, _04390_, _04563_);
  and (_05084_, _04393_, _04558_);
  or (_05085_, _05084_, _05082_);
  and (_05086_, _04379_, _04580_);
  and (_05088_, _04384_, _04578_);
  or (_05089_, _05088_, _05086_);
  or (_05090_, _05089_, _05085_);
  and (_05092_, _04407_, _04560_);
  and (_05093_, _04404_, _04572_);
  and (_05094_, _04435_, _04570_);
  or (_05096_, _05094_, _05093_);
  or (_05097_, _05096_, _05092_);
  and (_05098_, _04412_, _04550_);
  and (_05100_, _04375_, _04546_);
  and (_05101_, _04417_, _04567_);
  or (_05102_, _05101_, _05100_);
  and (_05104_, _04424_, _04565_);
  and (_05105_, _04420_, _04544_);
  or (_05106_, _05105_, _05104_);
  or (_05107_, _05106_, _05102_);
  or (_05108_, _05107_, _05098_);
  and (_05109_, _04432_, _04554_);
  and (_05110_, _04399_, _04552_);
  or (_05111_, _05110_, _05109_);
  or (_05112_, _05111_, _05108_);
  and (_05113_, _04440_, _04541_);
  and (_05114_, _04443_, _04539_);
  or (_05115_, _05114_, _05113_);
  or (_05116_, _05115_, _05112_);
  or (_05117_, _05116_, _05097_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [8], _05117_, _05090_);
  and (_05118_, _04390_, _04609_);
  and (_05119_, _04393_, _04598_);
  or (_05120_, _05119_, _05118_);
  and (_05121_, _04379_, _04585_);
  and (_05122_, _04384_, _04604_);
  or (_05123_, _05122_, _05121_);
  or (_05125_, _05123_, _05120_);
  and (_05126_, _04435_, _04617_);
  and (_05128_, _04404_, _04619_);
  and (_05129_, _04407_, _04626_);
  or (_05130_, _05129_, _05128_);
  or (_05132_, _05130_, _05126_);
  and (_05133_, _04412_, _04600_);
  and (_05134_, _04375_, _04587_);
  and (_05136_, _04417_, _04614_);
  or (_05137_, _05136_, _05134_);
  and (_05138_, _04424_, _04612_);
  and (_05140_, _04420_, _04590_);
  or (_05141_, _05140_, _05138_);
  or (_05142_, _05141_, _05137_);
  or (_05144_, _05142_, _05133_);
  and (_05145_, _04432_, _04596_);
  and (_05146_, _04399_, _04624_);
  or (_05148_, _05146_, _05145_);
  or (_05149_, _05148_, _05144_);
  and (_05150_, _04440_, _04592_);
  and (_05152_, _04443_, _04606_);
  or (_05153_, _05152_, _05150_);
  or (_05154_, _05153_, _05149_);
  or (_05156_, _05154_, _05132_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [9], _05156_, _05125_);
  and (_05157_, _04379_, _04637_);
  and (_05158_, _04384_, _04634_);
  or (_05159_, _05158_, _05157_);
  and (_05160_, _04390_, _04651_);
  and (_05161_, _04393_, _04647_);
  or (_05162_, _05161_, _05160_);
  or (_05163_, _05162_, _05159_);
  and (_05164_, _04432_, _04645_);
  and (_05165_, _04399_, _04667_);
  and (_05166_, _04435_, _04660_);
  or (_05167_, _05166_, _05165_);
  or (_05168_, _05167_, _05164_);
  and (_05169_, _04412_, _04665_);
  and (_05170_, _04417_, _04655_);
  and (_05171_, _04420_, _04639_);
  or (_05172_, _05171_, _05170_);
  and (_05173_, _04424_, _04658_);
  and (_05174_, _04375_, _04632_);
  or (_05175_, _05174_, _05173_);
  or (_05177_, _05175_, _05172_);
  or (_05178_, _05177_, _05169_);
  and (_05180_, _04404_, _04653_);
  and (_05181_, _04407_, _04643_);
  or (_05182_, _05181_, _05180_);
  or (_05184_, _05182_, _05178_);
  and (_05185_, _04440_, _04671_);
  and (_05186_, _04443_, _04673_);
  or (_05188_, _05186_, _05185_);
  or (_05189_, _05188_, _05184_);
  or (_05190_, _05189_, _05168_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [10], _05190_, _05163_);
  and (_05192_, _04443_, _04719_);
  and (_05193_, _04384_, _04680_);
  or (_05195_, _05193_, _05192_);
  and (_05196_, _04390_, _04697_);
  and (_05197_, _04393_, _04693_);
  or (_05199_, _05197_, _05196_);
  or (_05200_, _05199_, _05195_);
  and (_05201_, _04407_, _04713_);
  and (_05203_, _04399_, _04711_);
  and (_05204_, _04435_, _04701_);
  or (_05205_, _05204_, _05203_);
  or (_05207_, _05205_, _05201_);
  and (_05208_, _04440_, _04678_);
  and (_05209_, _04379_, _04717_);
  or (_05210_, _05209_, _05208_);
  and (_05211_, _04404_, _04704_);
  and (_05212_, _04432_, _04689_);
  or (_05213_, _05212_, _05211_);
  and (_05214_, _04412_, _04691_);
  and (_05215_, _04424_, _04699_);
  and (_05216_, _04417_, _04706_);
  or (_05217_, _05216_, _05215_);
  and (_05218_, _04375_, _04683_);
  and (_05219_, _04420_, _04685_);
  or (_05220_, _05219_, _05218_);
  or (_05221_, _05220_, _05217_);
  or (_05222_, _05221_, _05214_);
  or (_05223_, _05222_, _05213_);
  or (_05224_, _05223_, _05210_);
  or (_05225_, _05224_, _05207_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [11], _05225_, _05200_);
  and (_05226_, _04379_, _04729_);
  and (_05228_, _04384_, _04726_);
  or (_05229_, _05228_, _05226_);
  and (_05231_, _04390_, _04743_);
  and (_05232_, _04443_, _04765_);
  or (_05233_, _05232_, _05231_);
  or (_05235_, _05233_, _05229_);
  and (_05236_, _04404_, _04745_);
  and (_05237_, _04432_, _04737_);
  and (_05239_, _04399_, _04759_);
  or (_05240_, _05239_, _05237_);
  or (_05241_, _05240_, _05236_);
  and (_05243_, _04412_, _04757_);
  and (_05244_, _04417_, _04747_);
  and (_05245_, _04420_, _04731_);
  or (_05247_, _05245_, _05244_);
  and (_05248_, _04424_, _04750_);
  and (_05249_, _04375_, _04724_);
  or (_05251_, _05249_, _05248_);
  or (_05252_, _05251_, _05247_);
  or (_05253_, _05252_, _05243_);
  and (_05255_, _04435_, _04752_);
  and (_05256_, _04407_, _04735_);
  or (_05257_, _05256_, _05255_);
  or (_05259_, _05257_, _05253_);
  and (_05260_, _04440_, _04763_);
  and (_05261_, _04393_, _04739_);
  or (_05262_, _05261_, _05260_);
  or (_05263_, _05262_, _05259_);
  or (_05264_, _05263_, _05241_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [12], _05264_, _05235_);
  and (_05265_, _04390_, _04789_);
  and (_05266_, _04440_, _04809_);
  or (_05267_, _05266_, _05265_);
  and (_05268_, _04393_, _04781_);
  and (_05269_, _04384_, _04772_);
  or (_05270_, _05269_, _05268_);
  or (_05271_, _05270_, _05267_);
  and (_05272_, _04407_, _04805_);
  and (_05273_, _04404_, _04791_);
  and (_05274_, _04435_, _04798_);
  or (_05275_, _05274_, _05273_);
  or (_05276_, _05275_, _05272_);
  and (_05277_, _04412_, _04785_);
  and (_05278_, _04424_, _04796_);
  and (_05280_, _04375_, _04770_);
  or (_05281_, _05280_, _05278_);
  and (_05283_, _04417_, _04793_);
  and (_05284_, _04420_, _04777_);
  or (_05285_, _05284_, _05283_);
  or (_05287_, _05285_, _05281_);
  or (_05288_, _05287_, _05277_);
  and (_05289_, _04432_, _04783_);
  and (_05291_, _04399_, _04803_);
  or (_05292_, _05291_, _05289_);
  or (_05293_, _05292_, _05288_);
  and (_05295_, _04379_, _04775_);
  and (_05296_, _04443_, _04811_);
  or (_05297_, _05296_, _05295_);
  or (_05299_, _05297_, _05293_);
  or (_05300_, _05299_, _05276_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [13], _05300_, _05271_);
  and (_05302_, _04379_, _04821_);
  and (_05303_, _04384_, _04818_);
  or (_05304_, _05303_, _05302_);
  and (_05306_, _04390_, _04835_);
  and (_05307_, _04393_, _04831_);
  or (_05308_, _05307_, _05306_);
  or (_05310_, _05308_, _05304_);
  and (_05311_, _04404_, _04837_);
  and (_05312_, _04432_, _04829_);
  and (_05313_, _04407_, _04827_);
  or (_05314_, _05313_, _05312_);
  or (_05315_, _05314_, _05311_);
  and (_05316_, _04435_, _04844_);
  and (_05317_, _04399_, _04851_);
  or (_05318_, _05317_, _05316_);
  and (_05319_, _04412_, _04849_);
  and (_05320_, _04375_, _04816_);
  and (_05321_, _04417_, _04839_);
  or (_05322_, _05321_, _05320_);
  and (_05323_, _04424_, _04842_);
  and (_05324_, _04420_, _04823_);
  or (_05325_, _05324_, _05323_);
  or (_05326_, _05325_, _05322_);
  or (_05327_, _05326_, _05319_);
  or (_05328_, _05327_, _05318_);
  and (_05329_, _04440_, _04855_);
  and (_05330_, _04443_, _04857_);
  or (_05332_, _05330_, _05329_);
  or (_05333_, _05332_, _05328_);
  or (_05335_, _05333_, _05315_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [14], _05335_, _05310_);
  and (_05336_, _04379_, _04541_);
  and (_05338_, _04384_, _04539_);
  or (_05339_, _05338_, _05336_);
  and (_05340_, _04390_, _04550_);
  and (_05342_, _04393_, _04560_);
  or (_05343_, _05342_, _05340_);
  or (_05344_, _05343_, _05339_);
  and (_05346_, _04432_, _04572_);
  and (_05347_, _04435_, _04567_);
  and (_05348_, _04399_, _04570_);
  or (_05350_, _05348_, _05347_);
  or (_05351_, _05350_, _05346_);
  and (_05352_, _04412_, _04554_);
  and (_05354_, _04417_, _04546_);
  and (_05355_, _04420_, _04578_);
  or (_05356_, _05355_, _05354_);
  and (_05358_, _04375_, _04580_);
  and (_05359_, _04424_, _04544_);
  or (_05360_, _05359_, _05358_);
  or (_05362_, _05360_, _05356_);
  or (_05363_, _05362_, _05352_);
  and (_05364_, _04404_, _04565_);
  and (_05365_, _04407_, _04552_);
  or (_05366_, _05365_, _05364_);
  or (_05367_, _05366_, _05363_);
  and (_05368_, _04440_, _04563_);
  and (_05369_, _04443_, _04558_);
  or (_05370_, _05369_, _05368_);
  or (_05371_, _05370_, _05367_);
  or (_05372_, _05371_, _05351_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [16], _05372_, _05344_);
  and (_05373_, _04440_, _04609_);
  and (_05374_, _04393_, _04626_);
  or (_05375_, _05374_, _05373_);
  and (_05376_, _04390_, _04600_);
  and (_05377_, _04384_, _04606_);
  or (_05378_, _05377_, _05376_);
  or (_05379_, _05378_, _05375_);
  and (_05380_, _04407_, _04624_);
  and (_05381_, _04432_, _04619_);
  and (_05383_, _04399_, _04617_);
  or (_05384_, _05383_, _05381_);
  or (_05386_, _05384_, _05380_);
  and (_05387_, _04412_, _04596_);
  and (_05388_, _04417_, _04587_);
  and (_05390_, _04420_, _04604_);
  or (_05391_, _05390_, _05388_);
  and (_05392_, _04375_, _04585_);
  and (_05394_, _04424_, _04590_);
  or (_05395_, _05394_, _05392_);
  or (_05396_, _05395_, _05391_);
  or (_05398_, _05396_, _05387_);
  and (_05399_, _04404_, _04612_);
  and (_05400_, _04435_, _04614_);
  or (_05402_, _05400_, _05399_);
  or (_05403_, _05402_, _05398_);
  and (_05404_, _04379_, _04592_);
  and (_05406_, _04443_, _04598_);
  or (_05407_, _05406_, _05404_);
  or (_05408_, _05407_, _05403_);
  or (_05410_, _05408_, _05386_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [17], _05410_, _05379_);
  and (_05411_, _04393_, _04643_);
  and (_05413_, _04384_, _04673_);
  or (_05414_, _05413_, _05411_);
  and (_05415_, _04390_, _04665_);
  and (_05416_, _04379_, _04671_);
  or (_05417_, _05416_, _05415_);
  or (_05418_, _05417_, _05414_);
  and (_05419_, _04399_, _04660_);
  and (_05420_, _04435_, _04655_);
  and (_05421_, _04407_, _04667_);
  or (_05422_, _05421_, _05420_);
  or (_05423_, _05422_, _05419_);
  and (_05424_, _04412_, _04645_);
  and (_05425_, _04417_, _04632_);
  and (_05426_, _04420_, _04634_);
  or (_05427_, _05426_, _05425_);
  and (_05428_, _04375_, _04637_);
  and (_05429_, _04424_, _04639_);
  or (_05430_, _05429_, _05428_);
  or (_05431_, _05430_, _05427_);
  or (_05432_, _05431_, _05424_);
  and (_05433_, _04404_, _04658_);
  and (_05435_, _04432_, _04653_);
  or (_05436_, _05435_, _05433_);
  or (_05438_, _05436_, _05432_);
  and (_05439_, _04440_, _04651_);
  and (_05440_, _04443_, _04647_);
  or (_05442_, _05440_, _05439_);
  or (_05443_, _05442_, _05438_);
  or (_05444_, _05443_, _05423_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [18], _05444_, _05418_);
  and (_05446_, _04379_, _04678_);
  and (_05447_, _04384_, _04719_);
  or (_05449_, _05447_, _05446_);
  and (_05450_, _04390_, _04691_);
  and (_05451_, _04393_, _04713_);
  or (_05453_, _05451_, _05450_);
  or (_05454_, _05453_, _05449_);
  and (_05455_, _04435_, _04706_);
  and (_05457_, _04404_, _04699_);
  and (_05458_, _04399_, _04701_);
  or (_05459_, _05458_, _05457_);
  or (_05461_, _05459_, _05455_);
  and (_05462_, _04412_, _04689_);
  and (_05463_, _04417_, _04683_);
  and (_05465_, _04420_, _04680_);
  or (_05466_, _05465_, _05463_);
  and (_05467_, _04375_, _04717_);
  and (_05468_, _04424_, _04685_);
  or (_05469_, _05468_, _05467_);
  or (_05470_, _05469_, _05466_);
  or (_05471_, _05470_, _05462_);
  and (_05472_, _04432_, _04704_);
  and (_05473_, _04407_, _04711_);
  or (_05474_, _05473_, _05472_);
  or (_05475_, _05474_, _05471_);
  and (_05476_, _04440_, _04697_);
  and (_05477_, _04443_, _04693_);
  or (_05478_, _05477_, _05476_);
  or (_05479_, _05478_, _05475_);
  or (_05480_, _05479_, _05461_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [19], _05480_, _05454_);
  and (_05481_, _04379_, _04763_);
  and (_05482_, _04384_, _04765_);
  or (_05483_, _05482_, _05481_);
  and (_05484_, _04390_, _04757_);
  and (_05486_, _04393_, _04735_);
  or (_05487_, _05486_, _05484_);
  or (_05489_, _05487_, _05483_);
  and (_05490_, _04435_, _04747_);
  and (_05491_, _04404_, _04750_);
  and (_05493_, _04399_, _04752_);
  or (_05494_, _05493_, _05491_);
  or (_05495_, _05494_, _05490_);
  and (_05497_, _04412_, _04737_);
  and (_05498_, _04417_, _04724_);
  and (_05499_, _04420_, _04726_);
  or (_05501_, _05499_, _05498_);
  and (_05502_, _04375_, _04729_);
  and (_05503_, _04424_, _04731_);
  or (_05505_, _05503_, _05502_);
  or (_05506_, _05505_, _05501_);
  or (_05507_, _05506_, _05497_);
  and (_05509_, _04432_, _04745_);
  and (_05510_, _04407_, _04759_);
  or (_05511_, _05510_, _05509_);
  or (_05513_, _05511_, _05507_);
  and (_05514_, _04440_, _04743_);
  and (_05515_, _04443_, _04739_);
  or (_05517_, _05515_, _05514_);
  or (_05518_, _05517_, _05513_);
  or (_05519_, _05518_, _05495_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [20], _05519_, _05489_);
  and (_05520_, _04390_, _04785_);
  and (_05521_, _04393_, _04805_);
  or (_05522_, _05521_, _05520_);
  and (_05523_, _04379_, _04809_);
  and (_05524_, _04384_, _04811_);
  or (_05525_, _05524_, _05523_);
  or (_05526_, _05525_, _05522_);
  and (_05527_, _04435_, _04793_);
  and (_05528_, _04404_, _04796_);
  and (_05529_, _04407_, _04803_);
  or (_05530_, _05529_, _05528_);
  or (_05531_, _05530_, _05527_);
  and (_05532_, _04412_, _04783_);
  and (_05533_, _04375_, _04775_);
  and (_05534_, _04417_, _04770_);
  or (_05535_, _05534_, _05533_);
  and (_05536_, _04424_, _04777_);
  and (_05538_, _04420_, _04772_);
  or (_05539_, _05538_, _05536_);
  or (_05541_, _05539_, _05535_);
  or (_05542_, _05541_, _05532_);
  and (_05543_, _04432_, _04791_);
  and (_05545_, _04399_, _04798_);
  or (_05546_, _05545_, _05543_);
  or (_05547_, _05546_, _05542_);
  and (_05549_, _04440_, _04789_);
  and (_05550_, _04443_, _04781_);
  or (_05551_, _05550_, _05549_);
  or (_05553_, _05551_, _05547_);
  or (_05554_, _05553_, _05531_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [21], _05554_, _05526_);
  and (_05556_, _04393_, _04827_);
  and (_05557_, _04384_, _04857_);
  or (_05558_, _05557_, _05556_);
  and (_05560_, _04390_, _04849_);
  and (_05561_, _04379_, _04855_);
  or (_05562_, _05561_, _05560_);
  or (_05564_, _05562_, _05558_);
  and (_05565_, _04435_, _04839_);
  and (_05566_, _04404_, _04842_);
  and (_05568_, _04399_, _04844_);
  or (_05569_, _05568_, _05566_);
  or (_05570_, _05569_, _05565_);
  and (_05571_, _04412_, _04829_);
  and (_05572_, _04375_, _04821_);
  and (_05573_, _04420_, _04818_);
  or (_05574_, _05573_, _05572_);
  and (_05575_, _04417_, _04816_);
  and (_05576_, _04424_, _04823_);
  or (_05577_, _05576_, _05575_);
  or (_05578_, _05577_, _05574_);
  or (_05579_, _05578_, _05571_);
  and (_05580_, _04432_, _04837_);
  and (_05581_, _04407_, _04851_);
  or (_05582_, _05581_, _05580_);
  or (_05583_, _05582_, _05579_);
  and (_05584_, _04440_, _04835_);
  and (_05585_, _04443_, _04831_);
  or (_05586_, _05585_, _05584_);
  or (_05587_, _05586_, _05583_);
  or (_05588_, _05587_, _05570_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [22], _05588_, _05564_);
  nand (_05590_, \oc8051_golden_model_1.PC [1], \oc8051_golden_model_1.PC [0]);
  not (_05592_, \oc8051_golden_model_1.PC [3]);
  or (_05593_, \oc8051_golden_model_1.PC [2], _05592_);
  or (_05594_, _05593_, _05590_);
  or (_05596_, _05594_, _00459_);
  not (_05597_, \oc8051_golden_model_1.PC [1]);
  or (_05598_, _05597_, \oc8051_golden_model_1.PC [0]);
  or (_05600_, _05598_, _05593_);
  or (_05601_, _05600_, _00418_);
  and (_05602_, _05601_, _05596_);
  not (_05604_, \oc8051_golden_model_1.PC [2]);
  or (_05605_, _05604_, \oc8051_golden_model_1.PC [3]);
  or (_05606_, _05605_, _05590_);
  or (_05608_, _05606_, _00295_);
  or (_05609_, _05605_, _05598_);
  or (_05610_, _05609_, _00254_);
  and (_05612_, _05610_, _05608_);
  and (_05613_, _05612_, _05602_);
  nand (_05614_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [3]);
  or (_05616_, _05614_, _05590_);
  or (_05617_, _05616_, _00642_);
  or (_05618_, _05614_, _05598_);
  or (_05620_, _05618_, _00601_);
  and (_05621_, _05620_, _05617_);
  or (_05622_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [3]);
  or (_05623_, _05622_, _05590_);
  or (_05624_, _05623_, _00100_);
  or (_05625_, _05622_, _05598_);
  or (_05626_, _05625_, _00059_);
  and (_05627_, _05626_, _05624_);
  and (_05628_, _05627_, _05621_);
  and (_05629_, _05628_, _05613_);
  not (_05630_, \oc8051_golden_model_1.PC [0]);
  or (_05631_, \oc8051_golden_model_1.PC [1], _05630_);
  or (_05632_, _05631_, _05614_);
  or (_05633_, _05632_, _00541_);
  or (_05634_, \oc8051_golden_model_1.PC [1], \oc8051_golden_model_1.PC [0]);
  or (_05635_, _05634_, _05614_);
  or (_05636_, _05635_, _00500_);
  and (_05637_, _05636_, _05633_);
  or (_05638_, _05622_, _05634_);
  or (_05639_, _05638_, _43510_);
  or (_05640_, _05622_, _05631_);
  or (_05642_, _05640_, _00018_);
  and (_05643_, _05642_, _05639_);
  and (_05645_, _05643_, _05637_);
  or (_05646_, _05631_, _05593_);
  or (_05647_, _05646_, _00377_);
  or (_05649_, _05634_, _05593_);
  or (_05650_, _05649_, _00336_);
  and (_05651_, _05650_, _05647_);
  or (_05653_, _05631_, _05605_);
  or (_05654_, _05653_, _00213_);
  or (_05655_, _05634_, _05605_);
  or (_05657_, _05655_, _00155_);
  and (_05658_, _05657_, _05654_);
  and (_05659_, _05658_, _05651_);
  and (_05661_, _05659_, _05645_);
  nand (_05662_, _05661_, _05629_);
  or (_05663_, _05594_, _00424_);
  or (_05665_, _05600_, _00383_);
  and (_05666_, _05665_, _05663_);
  or (_05667_, _05606_, _00260_);
  or (_05669_, _05609_, _00219_);
  and (_05670_, _05669_, _05667_);
  and (_05671_, _05670_, _05666_);
  or (_05673_, _05616_, _00607_);
  or (_05674_, _05618_, _00550_);
  and (_05675_, _05674_, _05673_);
  or (_05676_, _05623_, _00065_);
  or (_05677_, _05625_, _00024_);
  and (_05678_, _05677_, _05676_);
  and (_05679_, _05678_, _05675_);
  and (_05680_, _05679_, _05671_);
  or (_05681_, _05632_, _00506_);
  or (_05682_, _05635_, _00465_);
  and (_05683_, _05682_, _05681_);
  or (_05684_, _05638_, _43475_);
  or (_05685_, _05640_, _43516_);
  and (_05686_, _05685_, _05684_);
  and (_05687_, _05686_, _05683_);
  or (_05688_, _05646_, _00342_);
  or (_05689_, _05649_, _00301_);
  and (_05690_, _05689_, _05688_);
  or (_05691_, _05653_, _00168_);
  or (_05692_, _05655_, _00106_);
  and (_05693_, _05692_, _05691_);
  and (_05695_, _05693_, _05690_);
  and (_05696_, _05695_, _05687_);
  nand (_05698_, _05696_, _05680_);
  or (_05699_, _05698_, _05662_);
  or (_05700_, _05594_, _00449_);
  or (_05702_, _05600_, _00408_);
  and (_05703_, _05702_, _05700_);
  or (_05704_, _05606_, _00285_);
  or (_05706_, _05609_, _00244_);
  and (_05707_, _05706_, _05704_);
  and (_05708_, _05707_, _05703_);
  or (_05710_, _05616_, _00632_);
  or (_05711_, _05618_, _00590_);
  and (_05712_, _05711_, _05710_);
  or (_05714_, _05623_, _00090_);
  or (_05715_, _05625_, _00049_);
  and (_05716_, _05715_, _05714_);
  and (_05718_, _05716_, _05712_);
  and (_05719_, _05718_, _05708_);
  or (_05720_, _05632_, _00531_);
  or (_05722_, _05635_, _00490_);
  and (_05723_, _05722_, _05720_);
  or (_05724_, _05638_, _43500_);
  or (_05726_, _05640_, _00008_);
  and (_05727_, _05726_, _05724_);
  and (_05728_, _05727_, _05723_);
  or (_05729_, _05646_, _00367_);
  or (_05730_, _05649_, _00326_);
  and (_05731_, _05730_, _05729_);
  or (_05732_, _05653_, _00203_);
  or (_05733_, _05655_, _00133_);
  and (_05734_, _05733_, _05732_);
  and (_05735_, _05734_, _05731_);
  and (_05736_, _05735_, _05728_);
  and (_05737_, _05736_, _05719_);
  or (_05738_, _05594_, _00454_);
  or (_05739_, _05600_, _00413_);
  and (_05740_, _05739_, _05738_);
  or (_05741_, _05606_, _00290_);
  or (_05742_, _05609_, _00249_);
  and (_05743_, _05742_, _05741_);
  and (_05744_, _05743_, _05740_);
  or (_05745_, _05616_, _00637_);
  or (_05746_, _05618_, _00596_);
  and (_05748_, _05746_, _05745_);
  or (_05749_, _05623_, _00095_);
  or (_05751_, _05625_, _00054_);
  and (_05752_, _05751_, _05749_);
  and (_05753_, _05752_, _05748_);
  and (_05755_, _05753_, _05744_);
  or (_05756_, _05632_, _00536_);
  or (_05757_, _05635_, _00495_);
  and (_05759_, _05757_, _05756_);
  or (_05760_, _05638_, _43505_);
  or (_05761_, _05640_, _00013_);
  and (_05763_, _05761_, _05760_);
  and (_05764_, _05763_, _05759_);
  or (_05765_, _05646_, _00372_);
  or (_05767_, _05649_, _00331_);
  and (_05768_, _05767_, _05765_);
  or (_05769_, _05653_, _00208_);
  or (_05771_, _05655_, _00144_);
  and (_05772_, _05771_, _05769_);
  and (_05773_, _05772_, _05768_);
  and (_05775_, _05773_, _05764_);
  nand (_05776_, _05775_, _05755_);
  or (_05777_, _05776_, _05737_);
  nor (_05779_, _05777_, _05699_);
  or (_05780_, _05594_, _00429_);
  or (_05781_, _05600_, _00388_);
  and (_05782_, _05781_, _05780_);
  or (_05783_, _05606_, _00265_);
  or (_05784_, _05609_, _00224_);
  and (_05785_, _05784_, _05783_);
  and (_05786_, _05785_, _05782_);
  or (_05787_, _05616_, _00612_);
  or (_05788_, _05618_, _00558_);
  and (_05789_, _05788_, _05787_);
  or (_05790_, _05623_, _00070_);
  or (_05791_, _05625_, _00029_);
  and (_05792_, _05791_, _05790_);
  and (_05793_, _05792_, _05789_);
  and (_05794_, _05793_, _05786_);
  or (_05795_, _05632_, _00511_);
  or (_05796_, _05635_, _00470_);
  and (_05797_, _05796_, _05795_);
  or (_05798_, _05638_, _43480_);
  or (_05799_, _05640_, _43521_);
  and (_05801_, _05799_, _05798_);
  and (_05802_, _05801_, _05797_);
  or (_05804_, _05646_, _00347_);
  or (_05805_, _05649_, _00306_);
  and (_05806_, _05805_, _05804_);
  or (_05808_, _05653_, _00179_);
  or (_05809_, _05655_, _00111_);
  and (_05810_, _05809_, _05808_);
  and (_05812_, _05810_, _05806_);
  and (_05813_, _05812_, _05802_);
  and (_05814_, _05813_, _05794_);
  or (_05816_, _05594_, _00434_);
  or (_05817_, _05600_, _00393_);
  and (_05818_, _05817_, _05816_);
  or (_05820_, _05606_, _00270_);
  or (_05821_, _05609_, _00229_);
  and (_05822_, _05821_, _05820_);
  and (_05824_, _05822_, _05818_);
  or (_05825_, _05616_, _00617_);
  or (_05826_, _05618_, _00566_);
  and (_05828_, _05826_, _05825_);
  or (_05829_, _05623_, _00075_);
  or (_05830_, _05625_, _00034_);
  and (_05832_, _05830_, _05829_);
  and (_05833_, _05832_, _05828_);
  and (_05834_, _05833_, _05824_);
  or (_05835_, _05632_, _00516_);
  or (_05836_, _05635_, _00475_);
  and (_05837_, _05836_, _05835_);
  or (_05838_, _05638_, _43485_);
  or (_05839_, _05640_, _43526_);
  and (_05840_, _05839_, _05838_);
  and (_05841_, _05840_, _05837_);
  or (_05842_, _05646_, _00352_);
  or (_05843_, _05649_, _00311_);
  and (_05844_, _05843_, _05842_);
  or (_05845_, _05653_, _00188_);
  or (_05846_, _05655_, _00116_);
  and (_05847_, _05846_, _05845_);
  and (_05848_, _05847_, _05844_);
  and (_05849_, _05848_, _05841_);
  nand (_05850_, _05849_, _05834_);
  not (_05851_, _05850_);
  and (_05852_, _05851_, _05814_);
  or (_05854_, _05594_, _00439_);
  or (_05855_, _05600_, _00398_);
  and (_05857_, _05855_, _05854_);
  or (_05858_, _05606_, _00275_);
  or (_05859_, _05609_, _00234_);
  and (_05861_, _05859_, _05858_);
  and (_05862_, _05861_, _05857_);
  or (_05863_, _05616_, _00622_);
  or (_05865_, _05618_, _00574_);
  and (_05866_, _05865_, _05863_);
  or (_05867_, _05623_, _00080_);
  or (_05869_, _05625_, _00039_);
  and (_05870_, _05869_, _05867_);
  and (_05871_, _05870_, _05866_);
  and (_05873_, _05871_, _05862_);
  or (_05874_, _05632_, _00521_);
  or (_05875_, _05635_, _00480_);
  and (_05877_, _05875_, _05874_);
  or (_05878_, _05638_, _43490_);
  or (_05879_, _05640_, _43531_);
  and (_05881_, _05879_, _05878_);
  and (_05882_, _05881_, _05877_);
  or (_05883_, _05646_, _00357_);
  or (_05885_, _05649_, _00316_);
  and (_05886_, _05885_, _05883_);
  or (_05887_, _05653_, _00193_);
  or (_05888_, _05655_, _00121_);
  and (_05889_, _05888_, _05887_);
  and (_05890_, _05889_, _05886_);
  and (_05891_, _05890_, _05882_);
  nand (_05892_, _05891_, _05873_);
  or (_05893_, _05594_, _00444_);
  or (_05894_, _05600_, _00403_);
  and (_05895_, _05894_, _05893_);
  or (_05896_, _05606_, _00280_);
  or (_05897_, _05609_, _00239_);
  and (_05898_, _05897_, _05896_);
  and (_05899_, _05898_, _05895_);
  or (_05900_, _05616_, _00627_);
  or (_05901_, _05618_, _00582_);
  and (_05902_, _05901_, _05900_);
  or (_05903_, _05623_, _00085_);
  or (_05904_, _05625_, _00044_);
  and (_05905_, _05904_, _05903_);
  and (_05906_, _05905_, _05902_);
  and (_05907_, _05906_, _05899_);
  or (_05908_, _05632_, _00526_);
  or (_05909_, _05635_, _00485_);
  and (_05910_, _05909_, _05908_);
  or (_05911_, _05638_, _43495_);
  or (_05912_, _05640_, _00003_);
  and (_05913_, _05912_, _05911_);
  and (_05914_, _05913_, _05910_);
  or (_05915_, _05646_, _00362_);
  or (_05916_, _05649_, _00321_);
  and (_05917_, _05916_, _05915_);
  or (_05918_, _05653_, _00198_);
  or (_05919_, _05655_, _00126_);
  and (_05920_, _05919_, _05918_);
  and (_05921_, _05920_, _05917_);
  and (_05922_, _05921_, _05914_);
  nand (_05923_, _05922_, _05907_);
  or (_05924_, _05923_, _05892_);
  not (_05925_, _05924_);
  and (_05926_, _05925_, _05852_);
  and (_05927_, _05926_, _05779_);
  not (_05928_, _05927_);
  nor (_05929_, _05614_, _05597_);
  and (_05930_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [1]);
  nor (_05931_, _05930_, \oc8051_golden_model_1.PC [3]);
  nor (_05932_, _05931_, _05929_);
  or (_05933_, _05850_, _05814_);
  or (_05934_, _05933_, _05924_);
  not (_05935_, _05934_);
  nand (_05936_, _05736_, _05719_);
  or (_05937_, _05776_, _05936_);
  nor (_05938_, _05937_, _05699_);
  and (_05939_, _05938_, _05935_);
  and (_05940_, _05935_, _05779_);
  nor (_05941_, _05940_, _05939_);
  and (_05942_, _05696_, _05680_);
  or (_05943_, _05942_, _05662_);
  nor (_05944_, _05943_, _05937_);
  not (_05945_, _05944_);
  or (_05946_, _05945_, _05934_);
  and (_05947_, _05661_, _05629_);
  or (_05948_, _05698_, _05947_);
  and (_05949_, _05775_, _05755_);
  or (_05950_, _05949_, _05737_);
  or (_05951_, _05950_, _05948_);
  or (_05952_, _05951_, _05934_);
  or (_05953_, _05949_, _05936_);
  or (_05954_, _05948_, _05953_);
  or (_05955_, _05954_, _05934_);
  and (_05956_, _05955_, _05952_);
  and (_05957_, _05956_, _05946_);
  or (_05958_, _05950_, _05699_);
  or (_05959_, _05958_, _05934_);
  or (_05960_, _05948_, _05777_);
  or (_05961_, _05960_, _05934_);
  and (_05962_, _05961_, _05959_);
  or (_05963_, _05953_, _05699_);
  or (_05964_, _05963_, _05934_);
  or (_05965_, _05948_, _05937_);
  or (_05966_, _05965_, _05934_);
  and (_05967_, _05966_, _05964_);
  and (_05968_, _05967_, _05962_);
  and (_05969_, _05968_, _05957_);
  and (_05970_, _05969_, _05941_);
  or (_05971_, _05970_, _05932_);
  or (_05972_, _05851_, _05814_);
  or (_05973_, _05972_, _05924_);
  nor (_05974_, _05973_, _05945_);
  not (_05975_, _05974_);
  nor (_05976_, _05943_, _05777_);
  not (_05977_, _05976_);
  or (_05978_, _05977_, _05934_);
  not (_05979_, _05892_);
  or (_05980_, _05923_, _05979_);
  or (_05981_, _05980_, _05933_);
  or (_05982_, _05981_, _05945_);
  and (_05983_, _05982_, _05978_);
  or (_05984_, _05977_, _05973_);
  and (_05985_, \oc8051_golden_model_1.DPL [2], \oc8051_golden_model_1.ACC [2]);
  and (_05986_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.ACC [1]);
  and (_05987_, \oc8051_golden_model_1.DPL [0], \oc8051_golden_model_1.ACC [0]);
  nor (_05988_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.ACC [1]);
  nor (_05989_, _05988_, _05986_);
  and (_05990_, _05989_, _05987_);
  nor (_05991_, _05990_, _05986_);
  nor (_05992_, \oc8051_golden_model_1.DPL [2], \oc8051_golden_model_1.ACC [2]);
  nor (_05993_, _05992_, _05985_);
  not (_05994_, _05993_);
  nor (_05995_, _05994_, _05991_);
  nor (_05996_, _05995_, _05985_);
  and (_05997_, \oc8051_golden_model_1.DPL [3], \oc8051_golden_model_1.ACC [3]);
  nor (_05998_, \oc8051_golden_model_1.DPL [3], \oc8051_golden_model_1.ACC [3]);
  nor (_05999_, _05998_, _05997_);
  not (_06000_, _05999_);
  nor (_06001_, _06000_, _05996_);
  and (_06002_, _06000_, _05996_);
  nor (_06003_, _06002_, _06001_);
  not (_06004_, _06003_);
  or (_06005_, _06004_, _05984_);
  or (_06006_, _05943_, _05950_);
  or (_06007_, _06006_, _05934_);
  or (_06008_, _05942_, _05947_);
  or (_06009_, _06008_, _05777_);
  or (_06010_, _06009_, _05934_);
  and (_06011_, _06010_, _06007_);
  or (_06012_, _06008_, _05937_);
  or (_06013_, _06012_, _05934_);
  or (_06014_, _06008_, _05953_);
  or (_06015_, _06014_, _05934_);
  and (_06016_, _06015_, _06013_);
  or (_06017_, _06008_, _05950_);
  or (_06018_, _06017_, _05934_);
  or (_06019_, _05943_, _05953_);
  or (_06020_, _06019_, _05934_);
  and (_06021_, _06020_, _06018_);
  and (_06022_, _06021_, _06016_);
  and (_06023_, _06022_, _06011_);
  not (_06024_, _05606_);
  nor (_06025_, _05590_, _05604_);
  nor (_06026_, _06025_, _05592_);
  nor (_06027_, _06026_, _06024_);
  not (_06028_, _06027_);
  and (_06029_, _05984_, _06028_);
  nand (_06030_, _06029_, _06023_);
  nand (_06031_, _06030_, _06005_);
  nand (_06032_, _06031_, _05983_);
  not (_06033_, _05932_);
  and (_06034_, _06023_, _05983_);
  or (_06035_, _06034_, _06033_);
  nand (_06036_, _06035_, _06032_);
  nand (_06037_, _06036_, _05975_);
  not (_06038_, _05970_);
  and (_06039_, _05590_, _05604_);
  nor (_06040_, _06039_, _06025_);
  and (_06041_, _06040_, \oc8051_golden_model_1.ACC [2]);
  not (_06042_, \oc8051_golden_model_1.ACC [1]);
  and (_06043_, _05631_, _05598_);
  nor (_06044_, _06043_, _06042_);
  and (_06045_, \oc8051_golden_model_1.ACC [0], _05630_);
  and (_06046_, _06043_, _06042_);
  nor (_06047_, _06046_, _06044_);
  and (_06048_, _06047_, _06045_);
  nor (_06049_, _06048_, _06044_);
  nor (_06050_, _06040_, \oc8051_golden_model_1.ACC [2]);
  nor (_06051_, _06050_, _06041_);
  not (_06052_, _06051_);
  nor (_06053_, _06052_, _06049_);
  nor (_06054_, _06053_, _06041_);
  not (_06055_, \oc8051_golden_model_1.ACC [3]);
  nor (_06056_, _06027_, _06055_);
  and (_06057_, _06027_, _06055_);
  nor (_06058_, _06057_, _06056_);
  and (_06059_, _06058_, _06054_);
  nor (_06060_, _06058_, _06054_);
  nor (_06061_, _06060_, _06059_);
  nor (_06062_, _06061_, _05975_);
  nor (_06063_, _06062_, _06038_);
  nand (_06064_, _06063_, _06037_);
  nand (_06065_, _06064_, _05971_);
  and (_06066_, _06052_, _06049_);
  nor (_06067_, _06066_, _06053_);
  and (_06068_, _06067_, _05974_);
  and (_06069_, _05994_, _05991_);
  nor (_06070_, _06069_, _05995_);
  not (_06071_, _06070_);
  or (_06072_, _06071_, _05984_);
  and (_06073_, _06072_, _05983_);
  not (_06074_, _06040_);
  nand (_06075_, _06074_, _06023_);
  nand (_06076_, _06075_, _05984_);
  nand (_06077_, _06076_, _06073_);
  nor (_06078_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [1]);
  nor (_06079_, _06078_, _05930_);
  or (_06080_, _06079_, _06034_);
  and (_06081_, _06080_, _05975_);
  and (_06082_, _06081_, _06077_);
  or (_06083_, _06082_, _06068_);
  nand (_06084_, _06083_, _05970_);
  not (_06085_, _06079_);
  or (_06086_, _06085_, _05970_);
  and (_06087_, _06086_, _06084_);
  or (_06088_, _06087_, _06065_);
  nor (_06089_, \oc8051_golden_model_1.DPL [0], \oc8051_golden_model_1.ACC [0]);
  nor (_06090_, _06089_, _05987_);
  or (_06091_, _06090_, _05984_);
  and (_06092_, _05984_, \oc8051_golden_model_1.PC [0]);
  nand (_06093_, _06092_, _06023_);
  nand (_06094_, _06093_, _06091_);
  and (_06095_, _05983_, _05975_);
  and (_06096_, _06095_, _06094_);
  not (_06097_, \oc8051_golden_model_1.ACC [0]);
  and (_06098_, _06097_, \oc8051_golden_model_1.PC [0]);
  nor (_06099_, _06098_, _06045_);
  nor (_06100_, _06099_, _05975_);
  or (_06101_, _06100_, _06096_);
  nand (_06102_, _06101_, _05970_);
  nand (_06103_, _06034_, _05970_);
  nand (_06104_, _06103_, _05630_);
  nand (_06105_, _06104_, _06102_);
  or (_06106_, _06034_, \oc8051_golden_model_1.PC [1]);
  nor (_06107_, _05989_, _05987_);
  nor (_06108_, _06107_, _05990_);
  not (_06109_, _06108_);
  or (_06110_, _06109_, _05984_);
  not (_06111_, _06043_);
  and (_06112_, _06111_, _05984_);
  nand (_06113_, _06112_, _06023_);
  nand (_06114_, _06113_, _06110_);
  and (_06115_, _05983_, _05970_);
  nand (_06116_, _06115_, _06114_);
  nand (_06117_, _06116_, _06106_);
  nand (_06118_, _06117_, _05975_);
  nor (_06119_, _06047_, _06045_);
  nor (_06120_, _06119_, _06048_);
  and (_06121_, _06120_, _05974_);
  nor (_06122_, _05970_, \oc8051_golden_model_1.PC [1]);
  nor (_06123_, _06122_, _06121_);
  and (_06124_, _06123_, _06118_);
  or (_06125_, _06124_, _06105_);
  or (_06126_, _06125_, _06088_);
  or (_06127_, _06126_, _00607_);
  nand (_06128_, _06123_, _06118_);
  or (_06129_, _06128_, _06105_);
  and (_06130_, _06064_, _05971_);
  nand (_06131_, _06086_, _06084_);
  or (_06132_, _06131_, _06130_);
  or (_06133_, _06132_, _06129_);
  or (_06134_, _06133_, _43516_);
  and (_06135_, _06134_, _06127_);
  or (_06136_, _06131_, _06065_);
  or (_06137_, _06136_, _06125_);
  or (_06138_, _06137_, _00424_);
  or (_06139_, _06132_, _06125_);
  or (_06140_, _06139_, _00065_);
  and (_06141_, _06140_, _06138_);
  and (_06142_, _06141_, _06135_);
  or (_06143_, _06136_, _06129_);
  or (_06144_, _06143_, _00342_);
  and (_06145_, _06104_, _06102_);
  or (_06146_, _06124_, _06145_);
  or (_06147_, _06132_, _06146_);
  or (_06148_, _06147_, _00024_);
  and (_06149_, _06148_, _06144_);
  or (_06150_, _06087_, _06130_);
  or (_06151_, _06150_, _06125_);
  or (_06152_, _06151_, _00260_);
  or (_06153_, _06150_, _06129_);
  or (_06154_, _06153_, _00168_);
  and (_06155_, _06154_, _06152_);
  and (_06156_, _06155_, _06149_);
  and (_06157_, _06156_, _06142_);
  or (_06158_, _06128_, _06145_);
  or (_06159_, _06150_, _06158_);
  or (_06160_, _06159_, _00106_);
  or (_06161_, _06132_, _06158_);
  or (_06162_, _06161_, _43475_);
  and (_06163_, _06162_, _06160_);
  or (_06164_, _06146_, _06088_);
  or (_06165_, _06164_, _00550_);
  or (_06166_, _06136_, _06146_);
  or (_06167_, _06166_, _00383_);
  and (_06168_, _06167_, _06165_);
  and (_06169_, _06168_, _06163_);
  or (_06170_, _06129_, _06088_);
  or (_06171_, _06170_, _00506_);
  or (_06172_, _06158_, _06136_);
  or (_06173_, _06172_, _00301_);
  and (_06174_, _06173_, _06171_);
  or (_06175_, _06158_, _06088_);
  or (_06176_, _06175_, _00465_);
  or (_06177_, _06150_, _06146_);
  or (_06178_, _06177_, _00219_);
  and (_06179_, _06178_, _06176_);
  and (_06180_, _06179_, _06174_);
  and (_06181_, _06180_, _06169_);
  nand (_06182_, _06181_, _06157_);
  or (_06183_, _06151_, _00280_);
  or (_06184_, _06139_, _00085_);
  and (_06185_, _06184_, _06183_);
  or (_06186_, _06170_, _00526_);
  or (_06187_, _06175_, _00485_);
  and (_06188_, _06187_, _06186_);
  and (_06189_, _06188_, _06185_);
  or (_06190_, _06147_, _00044_);
  or (_06191_, _06133_, _00003_);
  and (_06192_, _06191_, _06190_);
  or (_06193_, _06153_, _00198_);
  or (_06194_, _06159_, _00126_);
  and (_06195_, _06194_, _06193_);
  and (_06196_, _06195_, _06192_);
  and (_06197_, _06196_, _06189_);
  or (_06198_, _06137_, _00444_);
  or (_06199_, _06166_, _00403_);
  and (_06200_, _06199_, _06198_);
  or (_06201_, _06126_, _00627_);
  or (_06202_, _06143_, _00362_);
  and (_06203_, _06202_, _06201_);
  and (_06204_, _06203_, _06200_);
  or (_06205_, _06177_, _00239_);
  or (_06206_, _06161_, _43495_);
  and (_06207_, _06206_, _06205_);
  or (_06208_, _06164_, _00582_);
  or (_06209_, _06172_, _00321_);
  and (_06210_, _06209_, _06208_);
  and (_06211_, _06210_, _06207_);
  and (_06212_, _06211_, _06204_);
  and (_06213_, _06212_, _06197_);
  or (_06214_, _06213_, _06182_);
  nor (_06215_, _06214_, _05928_);
  nor (_06216_, _05959_, \oc8051_golden_model_1.SP [0]);
  not (_06217_, _05952_);
  nor (_06218_, _05981_, _05951_);
  not (_06219_, _06218_);
  nor (_06220_, _06219_, _06182_);
  or (_06221_, _06177_, _00224_);
  or (_06222_, _06153_, _00179_);
  and (_06223_, _06222_, _06221_);
  or (_06224_, _06139_, _00070_);
  or (_06225_, _06147_, _00029_);
  and (_06226_, _06225_, _06224_);
  and (_06227_, _06226_, _06223_);
  or (_06228_, _06143_, _00347_);
  or (_06229_, _06172_, _00306_);
  and (_06230_, _06229_, _06228_);
  or (_06231_, _06170_, _00511_);
  or (_06232_, _06175_, _00470_);
  and (_06233_, _06232_, _06231_);
  and (_06234_, _06233_, _06230_);
  and (_06235_, _06234_, _06227_);
  or (_06236_, _06161_, _43480_);
  or (_06237_, _06133_, _43521_);
  and (_06238_, _06237_, _06236_);
  or (_06239_, _06151_, _00265_);
  or (_06240_, _06159_, _00111_);
  and (_06241_, _06240_, _06239_);
  and (_06242_, _06241_, _06238_);
  or (_06243_, _06126_, _00612_);
  or (_06244_, _06164_, _00558_);
  and (_06245_, _06244_, _06243_);
  or (_06246_, _06137_, _00429_);
  or (_06247_, _06166_, _00388_);
  and (_06248_, _06247_, _06246_);
  and (_06249_, _06248_, _06245_);
  and (_06250_, _06249_, _06242_);
  and (_06251_, _06250_, _06235_);
  not (_06252_, _06251_);
  and (_06253_, _06252_, _06220_);
  not (_06254_, _05978_);
  and (_06255_, _05850_, _05814_);
  and (_06256_, _06255_, _05925_);
  and (_06257_, _06256_, _05976_);
  not (_06258_, _06257_);
  nor (_06259_, _06258_, _06214_);
  not (_06260_, _06006_);
  and (_06261_, _06256_, _06260_);
  not (_06262_, _06261_);
  nor (_06263_, _06262_, _06214_);
  nor (_06264_, _06262_, _06182_);
  not (_06265_, _06264_);
  not (_06266_, _06012_);
  and (_06267_, _06266_, _05926_);
  and (_06268_, _06256_, _06266_);
  not (_06269_, _06268_);
  nor (_06270_, _06269_, _06214_);
  not (_06271_, _06009_);
  and (_06272_, _06256_, _06271_);
  not (_06273_, _06272_);
  or (_06274_, _06273_, _06214_);
  nor (_06275_, _06273_, _06182_);
  not (_06276_, _06018_);
  not (_06277_, _05938_);
  nor (_06278_, _05981_, _06277_);
  not (_06279_, _06278_);
  not (_06280_, _05963_);
  and (_06281_, _06256_, _06280_);
  not (_06282_, _06281_);
  nor (_06283_, _05981_, _05963_);
  and (_06284_, _06283_, _06213_);
  not (_06285_, _06283_);
  not (_06286_, _06182_);
  nor (_06287_, _06151_, _00295_);
  nor (_06288_, _06139_, _00100_);
  nor (_06289_, _06288_, _06287_);
  nor (_06290_, _06170_, _00541_);
  nor (_06291_, _06175_, _00500_);
  nor (_06292_, _06291_, _06290_);
  and (_06293_, _06292_, _06289_);
  nor (_06294_, _06177_, _00254_);
  nor (_06295_, _06153_, _00213_);
  nor (_06296_, _06295_, _06294_);
  nor (_06297_, _06147_, _00059_);
  nor (_06298_, _06133_, _00018_);
  nor (_06299_, _06298_, _06297_);
  and (_06300_, _06299_, _06296_);
  and (_06301_, _06300_, _06293_);
  nor (_06302_, _06137_, _00459_);
  nor (_06303_, _06166_, _00418_);
  nor (_06304_, _06303_, _06302_);
  nor (_06305_, _06126_, _00642_);
  nor (_06306_, _06172_, _00336_);
  nor (_06307_, _06306_, _06305_);
  and (_06308_, _06307_, _06304_);
  nor (_06309_, _06159_, _00155_);
  nor (_06310_, _06161_, _43510_);
  nor (_06311_, _06310_, _06309_);
  nor (_06312_, _06164_, _00601_);
  nor (_06313_, _06143_, _00377_);
  nor (_06314_, _06313_, _06312_);
  and (_06315_, _06314_, _06311_);
  and (_06316_, _06315_, _06308_);
  and (_06317_, _06316_, _06301_);
  and (_06318_, _06317_, _06286_);
  and (_06319_, _06213_, _06182_);
  nor (_06320_, _06319_, _06318_);
  not (_06321_, _05951_);
  and (_06322_, _06256_, _06321_);
  and (_06323_, _06256_, _05944_);
  nor (_06324_, _06323_, _06322_);
  nor (_06325_, _06324_, _06320_);
  not (_06326_, _05981_);
  and (_06327_, _05923_, _05892_);
  and (_06328_, _06327_, _06255_);
  nor (_06329_, _06328_, _06326_);
  nor (_06330_, _06329_, _06006_);
  not (_06331_, _05933_);
  and (_06332_, _06327_, _06331_);
  not (_06333_, _06332_);
  not (_06334_, _05972_);
  and (_06335_, _06327_, _06334_);
  and (_06336_, _05923_, _05979_);
  and (_06337_, _06336_, _05852_);
  nor (_06338_, _06337_, _06335_);
  and (_06339_, _06338_, _06333_);
  or (_06340_, _06339_, _06006_);
  nor (_06341_, _06009_, _05981_);
  not (_06342_, _05980_);
  and (_06343_, _06255_, _06342_);
  and (_06344_, _06343_, _06260_);
  nor (_06345_, _05980_, _05972_);
  and (_06346_, _06345_, _06260_);
  or (_06347_, _06346_, _06344_);
  nor (_06348_, _06347_, _06341_);
  and (_06349_, _06348_, _06340_);
  and (_06350_, _06336_, _06331_);
  and (_06351_, _06350_, _06260_);
  not (_06352_, _06351_);
  and (_06353_, _06327_, _05852_);
  and (_06354_, _06353_, _06260_);
  nand (_06355_, _06336_, _05850_);
  nor (_06356_, _06355_, _06006_);
  nor (_06357_, _06356_, _06354_);
  and (_06358_, _06357_, _06352_);
  nand (_06359_, _06358_, _06349_);
  nor (_06360_, _06359_, _06330_);
  and (_06361_, _06256_, _05779_);
  and (_06362_, _06280_, _05926_);
  nor (_06363_, _06362_, _06361_);
  not (_06364_, _05958_);
  and (_06365_, _06364_, _05926_);
  nor (_06366_, _05973_, _05965_);
  nor (_06367_, _06366_, _06365_);
  and (_06368_, _06367_, _06363_);
  nor (_06369_, _05973_, _05954_);
  and (_06370_, _06342_, _05852_);
  and (_06371_, _06370_, _06260_);
  nor (_06372_, _06371_, _06369_);
  and (_06373_, _05976_, _05926_);
  not (_06374_, _06373_);
  nor (_06375_, _05973_, _05960_);
  nor (_06376_, _06375_, _06218_);
  and (_06377_, _06376_, _06374_);
  and (_06378_, _06377_, _06372_);
  and (_06379_, _06256_, _05938_);
  nor (_06380_, _06379_, _05927_);
  and (_06381_, _06380_, _06378_);
  and (_06382_, _06381_, _06368_);
  and (_06383_, _06382_, _06360_);
  and (_06384_, _06383_, _05630_);
  nor (_06385_, _06384_, _05597_);
  and (_06386_, _06384_, _05597_);
  nor (_06387_, _06386_, _06385_);
  nor (_06388_, _06383_, _05630_);
  nor (_06389_, _06388_, _06384_);
  and (_06390_, _06389_, _06387_);
  nor (_06391_, _06383_, _06085_);
  and (_06392_, _06383_, _06040_);
  nor (_06393_, _06392_, _06391_);
  nor (_06394_, _06383_, _06033_);
  and (_06395_, _06383_, _06028_);
  nor (_06396_, _06395_, _06394_);
  and (_06397_, _06396_, _06393_);
  and (_06398_, _06397_, _06390_);
  and (_06399_, _06398_, _04719_);
  nor (_06400_, _06389_, _06387_);
  and (_06401_, _06400_, _06397_);
  and (_06402_, _06401_, _04680_);
  nor (_06403_, _06402_, _06399_);
  nor (_06404_, _06396_, _06393_);
  not (_06405_, _06387_);
  nor (_06406_, _06389_, _06405_);
  and (_06407_, _06406_, _06404_);
  and (_06408_, _06407_, _04699_);
  not (_06409_, _06393_);
  nor (_06410_, _06396_, _06409_);
  and (_06411_, _06410_, _06406_);
  and (_06412_, _06411_, _04697_);
  nor (_06413_, _06412_, _06408_);
  and (_06414_, _06413_, _06403_);
  and (_06415_, _06410_, _06390_);
  and (_06416_, _06415_, _04678_);
  and (_06417_, _06410_, _06400_);
  and (_06418_, _06417_, _04717_);
  nor (_06419_, _06418_, _06416_);
  and (_06420_, _06404_, _06400_);
  and (_06421_, _06420_, _04689_);
  and (_06422_, _06389_, _06405_);
  and (_06423_, _06422_, _06404_);
  and (_06424_, _06423_, _04691_);
  nor (_06425_, _06424_, _06421_);
  and (_06426_, _06425_, _06419_);
  and (_06427_, _06426_, _06414_);
  and (_06428_, _06396_, _06409_);
  and (_06429_, _06428_, _06422_);
  and (_06430_, _06429_, _04713_);
  and (_06431_, _06406_, _06397_);
  and (_06432_, _06431_, _04693_);
  nor (_06433_, _06432_, _06430_);
  and (_06434_, _06428_, _06390_);
  and (_06435_, _06434_, _04701_);
  and (_06436_, _06422_, _06397_);
  and (_06437_, _06436_, _04685_);
  nor (_06438_, _06437_, _06435_);
  and (_06439_, _06438_, _06433_);
  and (_06440_, _06404_, _06390_);
  and (_06441_, _06440_, _04704_);
  and (_06442_, _06422_, _06410_);
  and (_06443_, _06442_, _04683_);
  nor (_06444_, _06443_, _06441_);
  and (_06445_, _06428_, _06406_);
  and (_06446_, _06445_, _04706_);
  and (_06447_, _06428_, _06400_);
  and (_06448_, _06447_, _04711_);
  nor (_06449_, _06448_, _06446_);
  and (_06450_, _06449_, _06444_);
  and (_06451_, _06450_, _06439_);
  and (_06452_, _06451_, _06427_);
  nor (_06453_, _06452_, _05982_);
  not (_06454_, _06324_);
  and (_06455_, _06260_, _05926_);
  nor (_06456_, _06455_, _06261_);
  not (_06457_, _06456_);
  and (_06458_, _06457_, _06320_);
  nor (_06459_, _06320_, _06273_);
  not (_06460_, \oc8051_golden_model_1.SP [3]);
  and (_06461_, _06271_, _05926_);
  and (_06462_, _06461_, _06460_);
  nor (_06463_, _06462_, _06459_);
  nor (_06464_, _06012_, _05981_);
  not (_06465_, _06464_);
  nor (_06466_, _06461_, _06272_);
  not (_06467_, _06466_);
  nor (_06468_, _06014_, _05981_);
  nor (_06469_, _06468_, _06341_);
  and (_06470_, _06469_, \oc8051_golden_model_1.PSW [3]);
  or (_06471_, _06470_, _06467_);
  and (_06472_, _06471_, _06465_);
  not (_06473_, _06213_);
  nand (_06474_, _06469_, _06465_);
  and (_06475_, _06474_, _06473_);
  or (_06476_, _06475_, _06472_);
  and (_06477_, _06476_, _06269_);
  and (_06478_, _06477_, _06463_);
  and (_06479_, _06320_, _06268_);
  nor (_06480_, _06006_, _05981_);
  nor (_06481_, _06480_, _06267_);
  not (_06482_, _06481_);
  nor (_06483_, _06482_, _06479_);
  not (_06484_, _06483_);
  nor (_06485_, _06484_, _06478_);
  and (_06486_, _06482_, _06213_);
  nor (_06487_, _06486_, _06457_);
  not (_06488_, _06487_);
  nor (_06489_, _06488_, _06485_);
  nor (_06490_, _06489_, _06458_);
  not (_06491_, _06019_);
  and (_06492_, _06328_, _06491_);
  and (_06493_, _06353_, _06491_);
  nor (_06494_, _06493_, _06492_);
  and (_06495_, _06335_, _06491_);
  and (_06496_, _06332_, _06491_);
  nor (_06497_, _06496_, _06495_);
  and (_06498_, _06336_, _06491_);
  not (_06499_, _06498_);
  and (_06500_, _06499_, _06497_);
  and (_06501_, _06500_, _06494_);
  not (_06502_, _06501_);
  nor (_06503_, _06502_, _06490_);
  and (_06504_, _06491_, _05926_);
  and (_06505_, _06256_, _06491_);
  nor (_06506_, _06505_, _06504_);
  not (_06507_, _06506_);
  nor (_06508_, _06501_, _06213_);
  nor (_06509_, _06508_, _06507_);
  not (_06510_, _06509_);
  nor (_06511_, _06510_, _06503_);
  nor (_06512_, _05981_, _05977_);
  nor (_06513_, _06506_, _06320_);
  nor (_06514_, _06513_, _06512_);
  not (_06515_, _06514_);
  nor (_06516_, _06515_, _06511_);
  not (_06517_, _06512_);
  nor (_06518_, _06517_, _06213_);
  or (_06519_, _06518_, _06516_);
  and (_06520_, _06519_, _06258_);
  and (_06521_, _06320_, _06257_);
  or (_06522_, _06521_, _06520_);
  and (_06523_, _06522_, _05982_);
  or (_06524_, _06523_, _06454_);
  nor (_06525_, _06524_, _06453_);
  or (_06526_, _06525_, _06325_);
  not (_06527_, _05965_);
  and (_06528_, _06256_, _06527_);
  nor (_06529_, _06528_, _06366_);
  nor (_06530_, _05981_, _05965_);
  not (_06531_, _06530_);
  and (_06532_, _06531_, _06529_);
  nor (_06533_, _05981_, _05954_);
  not (_06534_, _06533_);
  not (_06535_, _05954_);
  and (_06536_, _06256_, _06535_);
  nor (_06537_, _06536_, _06369_);
  and (_06538_, _06537_, _06534_);
  and (_06539_, _06538_, _06532_);
  nor (_06540_, _05981_, _05958_);
  not (_06541_, _06540_);
  nor (_06542_, _05981_, _05960_);
  not (_06543_, _06542_);
  not (_06544_, _05960_);
  and (_06545_, _06256_, _06544_);
  nor (_06546_, _06545_, _06375_);
  and (_06547_, _06546_, _06543_);
  and (_06548_, _06547_, _06541_);
  and (_06549_, _06548_, _06539_);
  nand (_06550_, _06549_, _06526_);
  and (_06551_, _06256_, _06364_);
  nor (_06552_, _06549_, _06473_);
  nor (_06553_, _06552_, _06551_);
  and (_06554_, _06553_, _06550_);
  and (_06555_, _06551_, \oc8051_golden_model_1.SP [3]);
  or (_06556_, _06555_, _06365_);
  nor (_06557_, _06556_, _06554_);
  not (_06558_, _06365_);
  nor (_06559_, _06320_, _06558_);
  or (_06560_, _06559_, _06557_);
  and (_06561_, _06560_, _06285_);
  or (_06562_, _06561_, _06284_);
  nand (_06563_, _06562_, _06282_);
  and (_06564_, _06281_, _06460_);
  nor (_06565_, _06564_, _06362_);
  nand (_06566_, _06565_, _06563_);
  not (_06567_, _05779_);
  nor (_06568_, _05981_, _06567_);
  and (_06569_, _06362_, _06320_);
  nor (_06570_, _06569_, _06568_);
  nand (_06571_, _06570_, _06566_);
  and (_06572_, _06568_, _06213_);
  nor (_06573_, _06572_, _05927_);
  and (_06574_, _06573_, _06571_);
  and (_06575_, _06320_, _05927_);
  or (_06576_, _06575_, _06574_);
  nand (_06577_, _06576_, _06279_);
  nor (_06578_, _06279_, _06213_);
  not (_06579_, _06578_);
  and (_06580_, _06579_, _06577_);
  nor (_06581_, _06133_, _00013_);
  nor (_06582_, _06147_, _00054_);
  nor (_06583_, _06582_, _06581_);
  nor (_06584_, _06164_, _00596_);
  nor (_06585_, _06177_, _00249_);
  nor (_06586_, _06585_, _06584_);
  and (_06587_, _06586_, _06583_);
  nor (_06588_, _06137_, _00454_);
  nor (_06589_, _06143_, _00372_);
  nor (_06590_, _06589_, _06588_);
  nor (_06591_, _06153_, _00208_);
  nor (_06592_, _06161_, _43505_);
  nor (_06593_, _06592_, _06591_);
  and (_06594_, _06593_, _06590_);
  and (_06595_, _06594_, _06587_);
  nor (_06596_, _06175_, _00495_);
  nor (_06597_, _06172_, _00331_);
  nor (_06598_, _06597_, _06596_);
  nor (_06599_, _06126_, _00637_);
  nor (_06600_, _06170_, _00536_);
  nor (_06601_, _06600_, _06599_);
  and (_06602_, _06601_, _06598_);
  nor (_06603_, _06166_, _00413_);
  nor (_06604_, _06139_, _00095_);
  nor (_06605_, _06604_, _06603_);
  nor (_06606_, _06151_, _00290_);
  nor (_06607_, _06159_, _00144_);
  nor (_06608_, _06607_, _06606_);
  and (_06609_, _06608_, _06605_);
  and (_06610_, _06609_, _06602_);
  and (_06611_, _06610_, _06595_);
  nor (_06612_, _06611_, _06182_);
  not (_06613_, _06612_);
  nor (_06614_, _06362_, _06257_);
  and (_06615_, _06614_, _06558_);
  and (_06616_, _06506_, _06456_);
  nor (_06617_, _06268_, _05927_);
  and (_06618_, _06617_, _06324_);
  and (_06619_, _06618_, _06616_);
  and (_06620_, _06619_, _06615_);
  nor (_06621_, _06620_, _06613_);
  not (_06622_, _06621_);
  and (_06623_, _06612_, _06272_);
  not (_06624_, _06623_);
  nor (_06625_, _06151_, _00275_);
  nor (_06627_, _06139_, _00080_);
  nor (_06628_, _06627_, _06625_);
  nor (_06629_, _06175_, _00480_);
  nor (_06630_, _06143_, _00357_);
  nor (_06631_, _06630_, _06629_);
  and (_06632_, _06631_, _06628_);
  nor (_06633_, _06177_, _00234_);
  nor (_06634_, _06153_, _00193_);
  nor (_06635_, _06634_, _06633_);
  nor (_06636_, _06161_, _43490_);
  nor (_06637_, _06147_, _00039_);
  nor (_06638_, _06637_, _06636_);
  and (_06639_, _06638_, _06635_);
  and (_06640_, _06639_, _06632_);
  nor (_06641_, _06126_, _00622_);
  nor (_06642_, _06164_, _00574_);
  nor (_06643_, _06642_, _06641_);
  nor (_06644_, _06170_, _00521_);
  nor (_06645_, _06137_, _00439_);
  nor (_06646_, _06645_, _06644_);
  and (_06647_, _06646_, _06643_);
  nor (_06648_, _06159_, _00121_);
  nor (_06649_, _06133_, _43531_);
  nor (_06650_, _06649_, _06648_);
  nor (_06651_, _06166_, _00398_);
  nor (_06652_, _06172_, _00316_);
  nor (_06653_, _06652_, _06651_);
  and (_06654_, _06653_, _06650_);
  and (_06655_, _06654_, _06647_);
  and (_06656_, _06655_, _06640_);
  not (_06657_, _06656_);
  nand (_06658_, _06517_, _06481_);
  nor (_06659_, _06658_, _06474_);
  nand (_06660_, _06659_, _06501_);
  nor (_06661_, _06568_, _06278_);
  and (_06662_, _06661_, _06285_);
  nand (_06663_, _06662_, _06549_);
  or (_06664_, _06663_, _06660_);
  and (_06665_, _06664_, _06657_);
  not (_06666_, _06665_);
  and (_06667_, _06440_, _04653_);
  and (_06668_, _06420_, _04645_);
  nor (_06669_, _06668_, _06667_);
  and (_06670_, _06429_, _04643_);
  and (_06671_, _06431_, _04647_);
  nor (_06672_, _06671_, _06670_);
  and (_06673_, _06672_, _06669_);
  and (_06674_, _06434_, _04660_);
  and (_06675_, _06447_, _04667_);
  nor (_06676_, _06675_, _06674_);
  and (_06677_, _06398_, _04673_);
  and (_06678_, _06401_, _04634_);
  nor (_06679_, _06678_, _06677_);
  and (_06680_, _06679_, _06676_);
  and (_06681_, _06680_, _06673_);
  and (_06682_, _06415_, _04671_);
  and (_06683_, _06442_, _04632_);
  nor (_06684_, _06683_, _06682_);
  and (_06685_, _06407_, _04658_);
  and (_06686_, _06423_, _04665_);
  nor (_06687_, _06686_, _06685_);
  and (_06688_, _06687_, _06684_);
  and (_06689_, _06445_, _04655_);
  and (_06690_, _06436_, _04639_);
  nor (_06691_, _06690_, _06689_);
  and (_06692_, _06411_, _04651_);
  and (_06693_, _06417_, _04637_);
  nor (_06694_, _06693_, _06692_);
  and (_06695_, _06694_, _06691_);
  and (_06696_, _06695_, _06688_);
  and (_06697_, _06696_, _06681_);
  nor (_06698_, _06697_, _05982_);
  nor (_06699_, _06335_, _06328_);
  nor (_06700_, _06699_, _06012_);
  nor (_06701_, _06699_, _06567_);
  nor (_06702_, _06701_, _06700_);
  and (_06703_, _06353_, _06535_);
  not (_06704_, _06703_);
  and (_06705_, _06353_, _05976_);
  not (_06706_, _06014_);
  and (_06707_, _06353_, _06706_);
  nor (_06708_, _06707_, _06705_);
  and (_06709_, _06708_, _06704_);
  and (_06710_, _06709_, _06702_);
  nor (_06711_, _06699_, _05965_);
  nor (_06712_, _06699_, _05960_);
  nor (_06713_, _06712_, _06711_);
  not (_06714_, _06713_);
  not (_06715_, \oc8051_golden_model_1.SP [2]);
  not (_06716_, _06551_);
  nor (_06717_, _06461_, _06281_);
  and (_06718_, _06717_, _06716_);
  nor (_06719_, _06718_, _06715_);
  nor (_06720_, _06719_, _06714_);
  and (_06721_, _06720_, _06710_);
  or (_06722_, _05777_, _05942_);
  nor (_06723_, _06722_, _06699_);
  and (_06724_, _05945_, _05954_);
  nor (_06725_, _05936_, _05699_);
  not (_06726_, _06725_);
  and (_06727_, _06726_, _06724_);
  nor (_06728_, _06727_, _06699_);
  nor (_06729_, _06728_, _06723_);
  not (_06730_, _06699_);
  nand (_06731_, _06006_, _05958_);
  or (_06732_, _06731_, _06706_);
  and (_06733_, _06732_, _06730_);
  and (_06734_, _06327_, _05851_);
  not (_06735_, _06734_);
  and (_06736_, _06006_, _05960_);
  and (_06737_, _06736_, _05963_);
  nor (_06738_, _06737_, _06735_);
  nor (_06739_, _06738_, _06733_);
  and (_06740_, _06739_, _06729_);
  and (_06741_, _06734_, _06266_);
  and (_06742_, _06734_, _06271_);
  nor (_06743_, _06742_, _06741_);
  and (_06744_, _06332_, _06535_);
  not (_06745_, _06744_);
  and (_06746_, _06745_, _06743_);
  and (_06747_, _06734_, _05938_);
  or (_06748_, _05976_, _05944_);
  and (_06749_, _06748_, _06332_);
  nor (_06750_, _06749_, _06747_);
  and (_06751_, _06750_, _06746_);
  and (_06752_, _06734_, _06364_);
  not (_06753_, _06752_);
  and (_06754_, _06734_, _05779_);
  and (_06755_, _06734_, _06527_);
  nor (_06756_, _06755_, _06754_);
  and (_06757_, _06756_, _06753_);
  and (_06758_, _06332_, _06706_);
  and (_06759_, _06353_, _05944_);
  nor (_06760_, _06759_, _06758_);
  and (_06761_, _06760_, _06757_);
  and (_06762_, _06761_, _06751_);
  and (_06763_, _06762_, _06740_);
  and (_06764_, _06763_, _06721_);
  not (_06765_, _06764_);
  nor (_06766_, _06765_, _06698_);
  and (_06767_, _06766_, _06666_);
  and (_06768_, _06767_, _06624_);
  and (_06769_, _06768_, _06622_);
  not (_06770_, \oc8051_golden_model_1.IRAM[0] [0]);
  nor (_06771_, _06279_, _06251_);
  not (_06772_, _06771_);
  nor (_06773_, _06506_, _06214_);
  not (_06774_, _06480_);
  nor (_06775_, _06774_, _06251_);
  or (_06776_, _06465_, _06251_);
  nor (_06777_, _06469_, _06251_);
  not (_06778_, _06017_);
  and (_06779_, _06343_, _06778_);
  nor (_06780_, _06779_, _06707_);
  and (_06781_, _06328_, _06706_);
  not (_06782_, _06781_);
  and (_06783_, _06343_, _06706_);
  nor (_06784_, _06783_, _06468_);
  and (_06785_, _06336_, _05814_);
  nand (_06786_, _06785_, _06706_);
  and (_06787_, _06786_, _06784_);
  and (_06788_, _06787_, _06782_);
  and (_06789_, _06788_, _06780_);
  and (_06790_, _06327_, _05814_);
  not (_06791_, _06790_);
  nor (_06792_, _06343_, _06785_);
  and (_06793_, _06792_, _06791_);
  nor (_06794_, _06793_, _06009_);
  nor (_06795_, _06794_, _06341_);
  and (_06796_, _06795_, _06789_);
  or (_06797_, _06796_, _06777_);
  nand (_06798_, _06797_, _06273_);
  nand (_06799_, _06274_, _06798_);
  not (_06800_, \oc8051_golden_model_1.SP [0]);
  and (_06801_, _06461_, _06800_);
  nor (_06802_, _06801_, _06464_);
  nor (_06803_, _06792_, _06012_);
  and (_06804_, _06790_, _06266_);
  nor (_06805_, _06804_, _06803_);
  and (_06806_, _06805_, _06802_);
  nand (_06807_, _06806_, _06799_);
  nand (_06808_, _06807_, _06776_);
  and (_06809_, _06808_, _06269_);
  or (_06810_, _06270_, _06809_);
  and (_06811_, _06267_, _06251_);
  nor (_06812_, _06792_, _06006_);
  not (_06813_, _06812_);
  nor (_06814_, _06354_, _06330_);
  and (_06815_, _06814_, _06813_);
  not (_06816_, _06815_);
  nor (_06817_, _06816_, _06811_);
  and (_06818_, _06817_, _06810_);
  or (_06819_, _06818_, _06775_);
  nand (_06820_, _06819_, _06456_);
  nor (_06821_, _06456_, _06214_);
  nor (_06822_, _06821_, _06502_);
  nand (_06823_, _06822_, _06820_);
  and (_06824_, _06502_, _06251_);
  and (_06825_, _06343_, _06491_);
  nor (_06826_, _06825_, _06507_);
  not (_06827_, _06826_);
  nor (_06828_, _06827_, _06824_);
  and (_06829_, _06828_, _06823_);
  nor (_06830_, _06829_, _06773_);
  not (_06831_, _06353_);
  and (_06832_, _06329_, _06831_);
  and (_06833_, _06832_, _06792_);
  nor (_06834_, _06833_, _05977_);
  nor (_06835_, _06834_, _06830_);
  nor (_06836_, _06517_, _06251_);
  or (_06837_, _06836_, _06835_);
  and (_06838_, _06837_, _06258_);
  nor (_06839_, _06838_, _06259_);
  nor (_06840_, _06833_, _05945_);
  nor (_06841_, _06840_, _06839_);
  and (_06842_, _06401_, _04578_);
  and (_06843_, _06398_, _04539_);
  nor (_06844_, _06843_, _06842_);
  and (_06845_, _06440_, _04572_);
  and (_06846_, _06434_, _04570_);
  nor (_06847_, _06846_, _06845_);
  and (_06848_, _06847_, _06844_);
  and (_06849_, _06411_, _04563_);
  and (_06850_, _06417_, _04580_);
  nor (_06851_, _06850_, _06849_);
  and (_06852_, _06447_, _04552_);
  and (_06853_, _06436_, _04544_);
  nor (_06854_, _06853_, _06852_);
  and (_06855_, _06854_, _06851_);
  and (_06856_, _06855_, _06848_);
  and (_06857_, _06423_, _04550_);
  and (_06858_, _06442_, _04546_);
  nor (_06859_, _06858_, _06857_);
  and (_06860_, _06407_, _04565_);
  and (_06861_, _06420_, _04554_);
  nor (_06862_, _06861_, _06860_);
  and (_06863_, _06862_, _06859_);
  and (_06864_, _06415_, _04541_);
  and (_06865_, _06431_, _04558_);
  nor (_06866_, _06865_, _06864_);
  and (_06867_, _06445_, _04567_);
  and (_06868_, _06429_, _04560_);
  nor (_06869_, _06868_, _06867_);
  and (_06870_, _06869_, _06866_);
  and (_06871_, _06870_, _06863_);
  and (_06872_, _06871_, _06856_);
  nor (_06873_, _06872_, _05982_);
  or (_06874_, _06873_, _06841_);
  and (_06875_, _06323_, _06214_);
  and (_06876_, _06343_, _06321_);
  nor (_06877_, _06876_, _06322_);
  not (_06878_, _06877_);
  nor (_06879_, _06878_, _06875_);
  and (_06880_, _06879_, _06874_);
  not (_06881_, _06322_);
  nor (_06882_, _06881_, _06214_);
  or (_06883_, _06882_, _06880_);
  and (_06884_, _06343_, _06535_);
  not (_06885_, _06884_);
  and (_06886_, _06336_, _06255_);
  and (_06887_, _06886_, _06535_);
  and (_06888_, _06337_, _06535_);
  nor (_06889_, _06888_, _06887_);
  and (_06890_, _06889_, _06885_);
  and (_06891_, _06328_, _06535_);
  nor (_06892_, _06891_, _06703_);
  and (_06893_, _06892_, _06890_);
  and (_06894_, _06893_, _06883_);
  nor (_06895_, _06538_, _06252_);
  nor (_06896_, _06793_, _05960_);
  nor (_06897_, _06896_, _06895_);
  and (_06898_, _06897_, _06894_);
  nor (_06899_, _06547_, _06252_);
  nor (_06900_, _06793_, _05965_);
  nor (_06901_, _06900_, _06899_);
  and (_06902_, _06901_, _06898_);
  nor (_06903_, _06532_, _06252_);
  nor (_06904_, _06833_, _05958_);
  nor (_06905_, _06904_, _06903_);
  and (_06906_, _06905_, _06902_);
  nor (_06907_, _06541_, _06251_);
  or (_06908_, _06907_, _06906_);
  and (_06909_, _06551_, _06800_);
  nor (_06910_, _06909_, _06365_);
  and (_06911_, _06910_, _06908_);
  nor (_06912_, _06558_, _06214_);
  nor (_06913_, _06912_, _06911_);
  nor (_06914_, _06833_, _05963_);
  nor (_06915_, _06914_, _06913_);
  nor (_06916_, _06285_, _06251_);
  or (_06917_, _06916_, _06915_);
  and (_06918_, _06281_, _06800_);
  nor (_06919_, _06918_, _06362_);
  and (_06920_, _06919_, _06917_);
  not (_06921_, _06362_);
  nor (_06922_, _06921_, _06214_);
  nor (_06923_, _06922_, _06920_);
  nor (_06924_, _06833_, _06567_);
  nor (_06925_, _06924_, _06923_);
  not (_06926_, _06568_);
  nor (_06927_, _06926_, _06251_);
  or (_06928_, _06927_, _06925_);
  and (_06929_, _06928_, _05928_);
  or (_06930_, _06929_, _06215_);
  and (_06931_, _06353_, _05938_);
  and (_06932_, _06792_, _06329_);
  nor (_06933_, _06932_, _06277_);
  nor (_06934_, _06933_, _06931_);
  nand (_06935_, _06934_, _06930_);
  nand (_06936_, _06935_, _06772_);
  or (_06937_, _06936_, _06770_);
  nor (_06938_, _06126_, _00632_);
  nor (_06939_, _06133_, _00008_);
  nor (_06940_, _06939_, _06938_);
  nor (_06941_, _06137_, _00449_);
  nor (_06942_, _06161_, _43500_);
  nor (_06943_, _06942_, _06941_);
  and (_06944_, _06943_, _06940_);
  nor (_06945_, _06143_, _00367_);
  nor (_06946_, _06147_, _00049_);
  nor (_06947_, _06946_, _06945_);
  nor (_06948_, _06177_, _00244_);
  nor (_06949_, _06159_, _00133_);
  nor (_06950_, _06949_, _06948_);
  and (_06951_, _06950_, _06947_);
  and (_06952_, _06951_, _06944_);
  nor (_06953_, _06153_, _00203_);
  nor (_06954_, _06139_, _00090_);
  nor (_06955_, _06954_, _06953_);
  nor (_06956_, _06170_, _00531_);
  nor (_06957_, _06166_, _00408_);
  nor (_06958_, _06957_, _06956_);
  and (_06959_, _06958_, _06955_);
  nor (_06960_, _06164_, _00590_);
  nor (_06961_, _06172_, _00326_);
  nor (_06962_, _06961_, _06960_);
  nor (_06963_, _06175_, _00490_);
  nor (_06964_, _06151_, _00285_);
  nor (_06965_, _06964_, _06963_);
  and (_06966_, _06965_, _06962_);
  and (_06967_, _06966_, _06959_);
  and (_06968_, _06967_, _06952_);
  nor (_06969_, _06968_, _06182_);
  and (_06970_, _06620_, _06273_);
  not (_06971_, _06970_);
  and (_06972_, _06971_, _06969_);
  not (_06973_, _06972_);
  nor (_06974_, _06137_, _00434_);
  nor (_06975_, _06166_, _00393_);
  nor (_06976_, _06975_, _06974_);
  nor (_06977_, _06175_, _00475_);
  nor (_06978_, _06143_, _00352_);
  nor (_06979_, _06978_, _06977_);
  and (_06980_, _06979_, _06976_);
  nor (_06981_, _06159_, _00116_);
  nor (_06982_, _06147_, _00034_);
  nor (_06983_, _06982_, _06981_);
  nor (_06984_, _06151_, _00270_);
  nor (_06985_, _06153_, _00188_);
  nor (_06986_, _06985_, _06984_);
  and (_06987_, _06986_, _06983_);
  and (_06988_, _06987_, _06980_);
  nor (_06989_, _06170_, _00516_);
  nor (_06990_, _06161_, _43485_);
  nor (_06991_, _06990_, _06989_);
  nor (_06992_, _06172_, _00311_);
  nor (_06993_, _06139_, _00075_);
  nor (_06994_, _06993_, _06992_);
  and (_06995_, _06994_, _06991_);
  nor (_06996_, _06126_, _00617_);
  nor (_06997_, _06133_, _43526_);
  nor (_06998_, _06997_, _06996_);
  nor (_06999_, _06164_, _00566_);
  nor (_07000_, _06177_, _00229_);
  nor (_07001_, _07000_, _06999_);
  and (_07002_, _07001_, _06998_);
  and (_07003_, _07002_, _06995_);
  and (_07004_, _07003_, _06988_);
  not (_07005_, _07004_);
  and (_07006_, _07005_, _06664_);
  not (_07007_, _07006_);
  and (_07008_, _06407_, _04612_);
  and (_07009_, _06440_, _04619_);
  nor (_07010_, _07009_, _07008_);
  and (_07011_, _06420_, _04596_);
  and (_07012_, _06411_, _04609_);
  nor (_07013_, _07012_, _07011_);
  and (_07014_, _07013_, _07010_);
  and (_07015_, _06429_, _04626_);
  and (_07016_, _06398_, _04606_);
  nor (_07017_, _07016_, _07015_);
  and (_07018_, _06445_, _04614_);
  and (_07019_, _06447_, _04624_);
  nor (_07020_, _07019_, _07018_);
  and (_07021_, _07020_, _07017_);
  and (_07022_, _07021_, _07014_);
  and (_07023_, _06442_, _04587_);
  and (_07024_, _06436_, _04590_);
  nor (_07025_, _07024_, _07023_);
  and (_07026_, _06417_, _04585_);
  and (_07027_, _06431_, _04598_);
  nor (_07028_, _07027_, _07026_);
  and (_07029_, _07028_, _07025_);
  and (_07030_, _06423_, _04600_);
  and (_07031_, _06401_, _04604_);
  nor (_07032_, _07031_, _07030_);
  and (_07033_, _06415_, _04592_);
  and (_07034_, _06434_, _04617_);
  nor (_07035_, _07034_, _07033_);
  and (_07036_, _07035_, _07032_);
  and (_07037_, _07036_, _07029_);
  and (_07038_, _07037_, _07022_);
  nor (_07039_, _07038_, _05982_);
  and (_07040_, _06886_, _06527_);
  and (_07041_, _06336_, _06334_);
  and (_07042_, _07041_, _06527_);
  nor (_07043_, _07042_, _07040_);
  and (_07044_, _06551_, \oc8051_golden_model_1.SP [1]);
  nor (_07045_, _06355_, _05963_);
  nor (_07046_, _07045_, _07044_);
  nand (_07047_, _07046_, _07043_);
  and (_07048_, _06012_, _06009_);
  nor (_07049_, _07048_, _06355_);
  nor (_07050_, _06355_, _05960_);
  or (_07051_, _07050_, _06356_);
  or (_07052_, _07051_, _07049_);
  or (_07053_, _07052_, _06728_);
  or (_07054_, _07053_, _07047_);
  or (_07055_, _05976_, _06364_);
  nor (_07056_, _07055_, _06706_);
  and (_07057_, _07056_, _06724_);
  nor (_07058_, _07057_, _06355_);
  or (_07059_, _07058_, _06714_);
  nor (_07060_, _07059_, _07054_);
  nor (_07061_, _06355_, _06567_);
  not (_07062_, _07061_);
  or (_07063_, _06355_, _06277_);
  and (_07064_, _07063_, _07062_);
  and (_07065_, _07064_, _06702_);
  nor (_07066_, _06733_, _06723_);
  not (_07067_, \oc8051_golden_model_1.SP [1]);
  nor (_07068_, _06717_, _07067_);
  not (_07069_, _07068_);
  and (_07070_, _07069_, _07066_);
  and (_07071_, _07070_, _07065_);
  and (_07072_, _07071_, _07060_);
  not (_07073_, _07072_);
  nor (_07074_, _07073_, _07039_);
  and (_07075_, _07074_, _07007_);
  and (_07076_, _07075_, _06973_);
  not (_07077_, \oc8051_golden_model_1.IRAM[1] [0]);
  and (_07078_, _06935_, _06772_);
  or (_07079_, _07078_, _07077_);
  and (_07080_, _07079_, _07076_);
  nand (_07081_, _07080_, _06937_);
  not (_07082_, \oc8051_golden_model_1.IRAM[3] [0]);
  or (_07083_, _07078_, _07082_);
  not (_07084_, _07076_);
  not (_07085_, \oc8051_golden_model_1.IRAM[2] [0]);
  or (_07086_, _06936_, _07085_);
  and (_07087_, _07086_, _07084_);
  nand (_07088_, _07087_, _07083_);
  nand (_07089_, _07088_, _07081_);
  nand (_07090_, _07089_, _06769_);
  not (_07091_, _06769_);
  not (_07092_, \oc8051_golden_model_1.IRAM[7] [0]);
  or (_07093_, _07078_, _07092_);
  not (_07094_, \oc8051_golden_model_1.IRAM[6] [0]);
  or (_07095_, _06936_, _07094_);
  and (_07096_, _07095_, _07084_);
  nand (_07097_, _07096_, _07093_);
  not (_07098_, \oc8051_golden_model_1.IRAM[4] [0]);
  or (_07099_, _06936_, _07098_);
  not (_07100_, \oc8051_golden_model_1.IRAM[5] [0]);
  or (_07101_, _07078_, _07100_);
  and (_07102_, _07101_, _07076_);
  nand (_07103_, _07102_, _07099_);
  nand (_07104_, _07103_, _07097_);
  nand (_07105_, _07104_, _07091_);
  nand (_07106_, _07105_, _07090_);
  nand (_07107_, _07106_, _06580_);
  not (_07108_, _06580_);
  nand (_07109_, _06936_, \oc8051_golden_model_1.IRAM[11] [0]);
  nand (_07110_, _07078_, \oc8051_golden_model_1.IRAM[10] [0]);
  and (_07111_, _07110_, _07084_);
  nand (_07112_, _07111_, _07109_);
  nand (_07113_, _07078_, \oc8051_golden_model_1.IRAM[8] [0]);
  nand (_07114_, _06936_, \oc8051_golden_model_1.IRAM[9] [0]);
  and (_07115_, _07114_, _07076_);
  nand (_07116_, _07115_, _07113_);
  nand (_07117_, _07116_, _07112_);
  nand (_07118_, _07117_, _06769_);
  not (_07119_, \oc8051_golden_model_1.IRAM[15] [0]);
  or (_07120_, _07078_, _07119_);
  nand (_07121_, _07078_, \oc8051_golden_model_1.IRAM[14] [0]);
  and (_07122_, _07121_, _07084_);
  nand (_07123_, _07122_, _07120_);
  not (_07124_, \oc8051_golden_model_1.IRAM[12] [0]);
  or (_07125_, _06936_, _07124_);
  nand (_07126_, _06936_, \oc8051_golden_model_1.IRAM[13] [0]);
  and (_07127_, _07126_, _07076_);
  nand (_07128_, _07127_, _07125_);
  nand (_07129_, _07128_, _07123_);
  nand (_07130_, _07129_, _07091_);
  nand (_07131_, _07130_, _07118_);
  nand (_07132_, _07131_, _07108_);
  and (_07133_, _07132_, _07107_);
  and (_07134_, _07133_, _06276_);
  nor (_07135_, _06343_, _06337_);
  nor (_07136_, _06370_, _05935_);
  and (_07137_, _07136_, _07135_);
  nor (_07138_, _07137_, _06017_);
  not (_07139_, _07138_);
  nor (_07140_, _07139_, _07134_);
  and (_07141_, _06335_, _06706_);
  not (_07142_, _07141_);
  nor (_07143_, _07142_, _06182_);
  and (_07144_, _07143_, _06251_);
  nor (_07145_, _07144_, _07140_);
  and (_07146_, _06758_, \oc8051_golden_model_1.SP [0]);
  and (_07147_, _05923_, _05814_);
  and (_07148_, _07147_, _06271_);
  nor (_07149_, _07148_, _07146_);
  and (_07150_, _07149_, _07145_);
  not (_07151_, _06341_);
  nor (_07152_, _07151_, _06182_);
  nor (_07153_, _06343_, _06345_);
  nor (_07154_, _07153_, _06009_);
  not (_07155_, _07154_);
  nor (_07156_, _07155_, _07133_);
  nor (_07157_, _07156_, _07152_);
  and (_07158_, _07157_, _07150_);
  and (_07159_, _07152_, _06252_);
  nor (_07160_, _07159_, _07158_);
  nor (_07161_, _07160_, _06275_);
  not (_07162_, _07161_);
  and (_07163_, _07162_, _06274_);
  nor (_07164_, _06010_, _06800_);
  nor (_07165_, _07164_, _07163_);
  not (_07166_, _06461_);
  nor (_07167_, _07166_, _06182_);
  and (_07168_, _07167_, _06251_);
  and (_07169_, _06785_, _06266_);
  nor (_07170_, _07169_, _06804_);
  not (_07171_, _07170_);
  nor (_07172_, _07171_, _07168_);
  and (_07173_, _07172_, _07165_);
  nor (_07174_, _07153_, _06012_);
  not (_07175_, _07174_);
  nor (_07176_, _07175_, _07133_);
  not (_07177_, _07176_);
  and (_07178_, _07177_, _07173_);
  nor (_07179_, _06269_, _06182_);
  nor (_07180_, _06465_, _06182_);
  and (_07181_, _07180_, _06251_);
  nor (_07182_, _07181_, _07179_);
  and (_07183_, _07182_, _07178_);
  nor (_07184_, _07183_, _06270_);
  or (_07185_, _07184_, _06267_);
  nand (_07186_, _06267_, _06800_);
  nand (_07187_, _07186_, _07185_);
  and (_07188_, _07187_, _06265_);
  nor (_07189_, _07188_, _06263_);
  and (_07190_, _06785_, _06491_);
  nor (_07191_, _06007_, _06800_);
  nor (_07192_, _07191_, _07190_);
  and (_07193_, _07192_, _06494_);
  not (_07194_, _07193_);
  nor (_07195_, _07194_, _07189_);
  nor (_07196_, _06258_, _06182_);
  nor (_07197_, _07153_, _06019_);
  not (_07198_, _07197_);
  nor (_07199_, _07198_, _07133_);
  nor (_07200_, _07199_, _07196_);
  and (_07201_, _07200_, _07195_);
  nor (_07202_, _07201_, _06259_);
  nor (_07203_, _07202_, _06254_);
  nor (_07204_, _05978_, \oc8051_golden_model_1.SP [0]);
  nor (_07205_, _07204_, _07203_);
  and (_07206_, _06343_, _05944_);
  and (_07207_, _06345_, _05944_);
  nor (_07208_, _07207_, _07206_);
  and (_07209_, _06336_, _05851_);
  and (_07210_, _07209_, _05944_);
  and (_07211_, _06699_, _06333_);
  and (_07212_, _06355_, _06831_);
  and (_07213_, _07212_, _07211_);
  nor (_07214_, _07213_, _05945_);
  nor (_07215_, _07214_, _07210_);
  and (_07216_, _07215_, _07208_);
  and (_07217_, _07216_, _05982_);
  nor (_07218_, _07217_, _06182_);
  and (_07219_, _07218_, _06251_);
  and (_07220_, _07147_, _06321_);
  nor (_07221_, _07220_, _07219_);
  not (_07222_, _07221_);
  nor (_07223_, _07222_, _07205_);
  nor (_07224_, _07153_, _05951_);
  not (_07225_, _07224_);
  nor (_07226_, _07225_, _07133_);
  nor (_07227_, _07226_, _06220_);
  and (_07228_, _07227_, _07223_);
  nor (_07229_, _07228_, _06253_);
  nor (_07230_, _07229_, _06217_);
  nor (_07231_, _05952_, \oc8051_golden_model_1.SP [0]);
  nor (_07232_, _07231_, _07230_);
  not (_07233_, _05961_);
  not (_07234_, _06545_);
  nor (_07235_, _07234_, _06182_);
  not (_07236_, _07235_);
  not (_07237_, _06369_);
  nor (_07238_, _07237_, _06182_);
  not (_07239_, _07238_);
  not (_07240_, _06536_);
  nor (_07241_, _07240_, _06182_);
  not (_07242_, _06375_);
  nor (_07243_, _07242_, _06182_);
  nor (_07244_, _07243_, _07241_);
  and (_07245_, _07244_, _07239_);
  and (_07246_, _07245_, _07236_);
  nor (_07247_, _07246_, _06252_);
  nor (_07248_, _07247_, _07233_);
  not (_07249_, _07248_);
  nor (_07250_, _07249_, _07232_);
  nor (_07251_, _05961_, \oc8051_golden_model_1.SP [0]);
  nor (_07252_, _07251_, _07250_);
  not (_07253_, _05959_);
  nor (_07254_, _06529_, _06182_);
  and (_07255_, _07254_, _06251_);
  or (_07256_, _07255_, _07253_);
  nor (_07257_, _07256_, _07252_);
  nor (_07258_, _07257_, _06216_);
  and (_07259_, _07147_, _05779_);
  nor (_07260_, _07259_, _07258_);
  nor (_07261_, _06926_, _06182_);
  and (_07262_, _06343_, _05779_);
  and (_07263_, _06345_, _05779_);
  nor (_07264_, _07263_, _07262_);
  nor (_07265_, _07264_, _07133_);
  nor (_07266_, _07265_, _07261_);
  and (_07267_, _07266_, _07260_);
  and (_07268_, _07261_, _06252_);
  nor (_07269_, _07268_, _07267_);
  nor (_07270_, _06182_, _05928_);
  nor (_07271_, _06361_, _05940_);
  nor (_07272_, _07271_, _06800_);
  nor (_07273_, _07272_, _07270_);
  not (_07274_, _07273_);
  nor (_07275_, _07274_, _07269_);
  nor (_07276_, _07275_, _06215_);
  and (_07277_, _07147_, _05938_);
  nor (_07278_, _07277_, _07276_);
  and (_07279_, _06343_, _05938_);
  and (_07280_, _06345_, _05938_);
  or (_07281_, _07280_, _07279_);
  not (_07282_, _07281_);
  nor (_07283_, _07282_, _07133_);
  not (_07284_, _07283_);
  and (_07285_, _07284_, _07278_);
  nor (_07286_, _06279_, _06182_);
  and (_07287_, _07286_, _06251_);
  not (_07288_, _07287_);
  and (_07289_, _07288_, _07285_);
  and (_07290_, _07286_, _07005_);
  and (_07291_, _06969_, _05927_);
  and (_07292_, _07209_, _05779_);
  nor (_07293_, _07292_, _06754_);
  not (_07294_, _07293_);
  and (_07295_, _07067_, \oc8051_golden_model_1.SP [0]);
  and (_07296_, \oc8051_golden_model_1.SP [1], _06800_);
  nor (_07297_, _07296_, _07295_);
  nor (_07298_, _07297_, _05959_);
  and (_07299_, _07005_, _06220_);
  and (_07300_, _06969_, _06257_);
  not (_07301_, _07297_);
  and (_07302_, _07301_, _06267_);
  not (_07303_, _06267_);
  nor (_07304_, _07153_, _06017_);
  not (_07305_, \oc8051_golden_model_1.IRAM[0] [1]);
  or (_07306_, _06936_, _07305_);
  not (_07307_, \oc8051_golden_model_1.IRAM[1] [1]);
  or (_07308_, _07078_, _07307_);
  and (_07309_, _07308_, _07076_);
  nand (_07310_, _07309_, _07306_);
  not (_07311_, \oc8051_golden_model_1.IRAM[3] [1]);
  or (_07312_, _07078_, _07311_);
  not (_07313_, \oc8051_golden_model_1.IRAM[2] [1]);
  or (_07314_, _06936_, _07313_);
  and (_07315_, _07314_, _07084_);
  nand (_07316_, _07315_, _07312_);
  nand (_07317_, _07316_, _07310_);
  nand (_07318_, _07317_, _06769_);
  not (_07319_, \oc8051_golden_model_1.IRAM[7] [1]);
  or (_07320_, _07078_, _07319_);
  not (_07321_, \oc8051_golden_model_1.IRAM[6] [1]);
  or (_07322_, _06936_, _07321_);
  and (_07323_, _07322_, _07084_);
  nand (_07324_, _07323_, _07320_);
  not (_07325_, \oc8051_golden_model_1.IRAM[4] [1]);
  or (_07326_, _06936_, _07325_);
  not (_07327_, \oc8051_golden_model_1.IRAM[5] [1]);
  or (_07328_, _07078_, _07327_);
  and (_07329_, _07328_, _07076_);
  nand (_07330_, _07329_, _07326_);
  nand (_07331_, _07330_, _07324_);
  nand (_07332_, _07331_, _07091_);
  nand (_07333_, _07332_, _07318_);
  nand (_07334_, _07333_, _06580_);
  nand (_07335_, _06936_, \oc8051_golden_model_1.IRAM[11] [1]);
  nand (_07336_, _07078_, \oc8051_golden_model_1.IRAM[10] [1]);
  and (_07337_, _07336_, _07084_);
  nand (_07338_, _07337_, _07335_);
  nand (_07339_, _07078_, \oc8051_golden_model_1.IRAM[8] [1]);
  nand (_07340_, _06936_, \oc8051_golden_model_1.IRAM[9] [1]);
  and (_07341_, _07340_, _07076_);
  nand (_07342_, _07341_, _07339_);
  nand (_07343_, _07342_, _07338_);
  nand (_07344_, _07343_, _06769_);
  nand (_07345_, _06936_, \oc8051_golden_model_1.IRAM[15] [1]);
  nand (_07346_, _07078_, \oc8051_golden_model_1.IRAM[14] [1]);
  and (_07347_, _07346_, _07084_);
  nand (_07348_, _07347_, _07345_);
  nand (_07349_, _07078_, \oc8051_golden_model_1.IRAM[12] [1]);
  nand (_07350_, _06936_, \oc8051_golden_model_1.IRAM[13] [1]);
  and (_07351_, _07350_, _07076_);
  nand (_07352_, _07351_, _07349_);
  nand (_07353_, _07352_, _07348_);
  nand (_07354_, _07353_, _07091_);
  nand (_07355_, _07354_, _07344_);
  nand (_07356_, _07355_, _07108_);
  nand (_07357_, _07356_, _07334_);
  and (_07358_, _07357_, _06276_);
  or (_07359_, _07358_, _07304_);
  and (_07360_, _07143_, _07004_);
  or (_07361_, _07360_, _07359_);
  and (_07362_, _07297_, _06758_);
  not (_07363_, _07362_);
  and (_07364_, _07209_, _06271_);
  nor (_07365_, _07364_, _06742_);
  and (_07366_, _07365_, _07363_);
  not (_07367_, _07366_);
  nor (_07368_, _07367_, _07361_);
  and (_07369_, _07357_, _07154_);
  nor (_07370_, _07369_, _07152_);
  and (_07371_, _07370_, _07368_);
  and (_07372_, _07152_, _07005_);
  nor (_07373_, _07372_, _07371_);
  and (_07374_, _06968_, _06275_);
  nor (_07375_, _07374_, _07373_);
  or (_07376_, _07301_, _06010_);
  nand (_07377_, _07376_, _07375_);
  and (_07378_, _07167_, _07004_);
  and (_07379_, _07209_, _06266_);
  nor (_07380_, _07379_, _06741_);
  not (_07381_, _07380_);
  nor (_07382_, _07381_, _07378_);
  not (_07383_, _07382_);
  nor (_07384_, _07383_, _07377_);
  and (_07385_, _07357_, _07174_);
  nor (_07386_, _07385_, _07180_);
  and (_07387_, _07386_, _07384_);
  and (_07388_, _07180_, _07005_);
  nor (_07389_, _07388_, _07387_);
  and (_07390_, _06968_, _07179_);
  nor (_07391_, _07390_, _07389_);
  and (_07392_, _07391_, _07303_);
  nor (_07393_, _07392_, _07302_);
  and (_07394_, _06968_, _06264_);
  or (_07395_, _07394_, _07393_);
  nor (_07396_, _07301_, _06007_);
  not (_07397_, _07396_);
  and (_07398_, _07209_, _06491_);
  and (_07399_, _06734_, _06491_);
  nor (_07400_, _07399_, _07398_);
  and (_07401_, _07400_, _07397_);
  not (_07402_, _07401_);
  nor (_07403_, _07402_, _07395_);
  and (_07404_, _07357_, _07197_);
  nor (_07405_, _07404_, _07196_);
  and (_07406_, _07405_, _07403_);
  nor (_07407_, _07406_, _07300_);
  nor (_07408_, _07407_, _06254_);
  nor (_07409_, _07297_, _05978_);
  nor (_07410_, _07409_, _07408_);
  and (_07411_, _07218_, _07004_);
  nor (_07412_, _05951_, _05850_);
  and (_07413_, _07412_, _05923_);
  nor (_07414_, _07413_, _07411_);
  not (_07415_, _07414_);
  nor (_07416_, _07415_, _07410_);
  and (_07417_, _07357_, _07224_);
  nor (_07418_, _07417_, _06220_);
  and (_07419_, _07418_, _07416_);
  nor (_07420_, _07419_, _07299_);
  nor (_07421_, _07420_, _06217_);
  nor (_07422_, _07297_, _05952_);
  nor (_07423_, _07422_, _07421_);
  nor (_07424_, _07246_, _07005_);
  nor (_07425_, _07424_, _07233_);
  not (_07426_, _07425_);
  nor (_07427_, _07426_, _07423_);
  nor (_07428_, _07297_, _05961_);
  nor (_07429_, _07428_, _07427_);
  and (_07430_, _07254_, _07004_);
  or (_07431_, _07430_, _07253_);
  nor (_07432_, _07431_, _07429_);
  nor (_07433_, _07432_, _07298_);
  nor (_07434_, _07433_, _07294_);
  not (_07435_, _07264_);
  and (_07436_, _07357_, _07435_);
  nor (_07437_, _07436_, _07261_);
  and (_07438_, _07437_, _07434_);
  and (_07439_, _07261_, _07005_);
  nor (_07440_, _07439_, _07438_);
  nor (_07441_, _07301_, _07271_);
  nor (_07442_, _07441_, _07270_);
  not (_07443_, _07442_);
  nor (_07444_, _07443_, _07440_);
  nor (_07445_, _07444_, _07291_);
  and (_07446_, _07209_, _05938_);
  nor (_07447_, _07446_, _06747_);
  not (_07448_, _07447_);
  nor (_07449_, _07448_, _07445_);
  and (_07450_, _07357_, _07281_);
  nor (_07451_, _07450_, _07286_);
  and (_07452_, _07451_, _07449_);
  nor (_07453_, _07452_, _07290_);
  not (_07454_, _01354_);
  nor (_07455_, _07211_, _05945_);
  not (_07456_, _07455_);
  not (_07457_, _06759_);
  nor (_07458_, _07210_, _07141_);
  and (_07459_, _07458_, _07457_);
  not (_07460_, _07208_);
  nor (_07461_, _06355_, _05945_);
  nor (_07462_, _07461_, _07460_);
  and (_07463_, _07462_, _07459_);
  and (_07464_, _07463_, _07456_);
  nor (_07465_, _07464_, _06182_);
  nor (_07466_, _07465_, _07235_);
  nor (_07467_, _07167_, _06264_);
  and (_07468_, _07467_, _07466_);
  nor (_07469_, _07180_, _07179_);
  nor (_07470_, _06182_, _05982_);
  not (_07471_, _07470_);
  and (_07472_, _07412_, _06785_);
  nor (_07473_, _07472_, _06492_);
  and (_07474_, _07264_, _07175_);
  and (_07475_, _07474_, _07473_);
  not (_07476_, _07049_);
  and (_07477_, _07476_, _06743_);
  nor (_07478_, _07281_, _07154_);
  and (_07479_, _07478_, _07477_);
  and (_07480_, _07479_, _07475_);
  not (_07481_, _07209_);
  and (_07482_, _07153_, _07481_);
  nor (_07483_, _07482_, _06017_);
  nand (_07484_, _07136_, _05981_);
  and (_07485_, _07484_, _06778_);
  or (_07486_, _07485_, _07483_);
  not (_07487_, _07486_);
  nor (_07488_, _07197_, _06493_);
  and (_07489_, _07488_, _07225_);
  and (_07490_, _07489_, _07487_);
  and (_07491_, _07490_, _07480_);
  and (_07492_, _06350_, _06321_);
  not (_07493_, _07492_);
  and (_07494_, _06007_, _05978_);
  and (_07495_, _06010_, _05952_);
  and (_07496_, _07495_, _07494_);
  and (_07497_, _07496_, _07493_);
  nor (_07498_, _06699_, _06009_);
  not (_07499_, _07498_);
  and (_07500_, _07499_, _06497_);
  and (_07501_, _07500_, _07497_);
  nor (_07502_, _07364_, _07398_);
  and (_07503_, _07502_, _07293_);
  not (_07504_, _06758_);
  and (_07505_, _07041_, _06491_);
  nor (_07506_, _07446_, _07505_);
  and (_07507_, _07506_, _07504_);
  and (_07508_, _07507_, _07503_);
  and (_07509_, _07271_, _05962_);
  and (_07510_, _06327_, _05938_);
  nor (_07511_, _07510_, _06267_);
  and (_07512_, _06886_, _06491_);
  nor (_07513_, _07379_, _07512_);
  and (_07514_, _07513_, _07511_);
  and (_07515_, _07514_, _07509_);
  and (_07516_, _07515_, _07508_);
  and (_07517_, _07516_, _07501_);
  nor (_07518_, _07213_, _05951_);
  not (_07519_, _07518_);
  and (_07520_, _07519_, _07065_);
  and (_07521_, _07520_, _07517_);
  and (_07522_, _07521_, _07491_);
  and (_07523_, _07522_, _07471_);
  and (_07524_, _07523_, _07469_);
  and (_07525_, _07524_, _07468_);
  nor (_07526_, _07261_, _06220_);
  nor (_07527_, _07254_, _07196_);
  and (_07528_, _07527_, _07526_);
  nor (_07529_, _07286_, _07270_);
  nor (_07530_, _07152_, _06275_);
  and (_07531_, _07530_, _07529_);
  and (_07532_, _07531_, _07528_);
  and (_07533_, _07532_, _07245_);
  and (_07534_, _07533_, _07525_);
  nor (_07535_, _07534_, _07454_);
  not (_07536_, _07535_);
  nor (_07537_, _07536_, _07453_);
  and (_07538_, _07537_, _07289_);
  not (_07539_, _07270_);
  or (_07540_, _07539_, _06318_);
  or (_07541_, _07153_, _06567_);
  not (_07542_, \oc8051_golden_model_1.IRAM[0] [3]);
  or (_07543_, _06936_, _07542_);
  not (_07544_, \oc8051_golden_model_1.IRAM[1] [3]);
  or (_07545_, _07078_, _07544_);
  and (_07546_, _07545_, _07076_);
  nand (_07547_, _07546_, _07543_);
  not (_07548_, \oc8051_golden_model_1.IRAM[3] [3]);
  or (_07549_, _07078_, _07548_);
  not (_07550_, \oc8051_golden_model_1.IRAM[2] [3]);
  or (_07551_, _06936_, _07550_);
  and (_07552_, _07551_, _07084_);
  nand (_07553_, _07552_, _07549_);
  nand (_07554_, _07553_, _07547_);
  nand (_07555_, _07554_, _06769_);
  not (_07556_, \oc8051_golden_model_1.IRAM[7] [3]);
  or (_07557_, _07078_, _07556_);
  not (_07558_, \oc8051_golden_model_1.IRAM[6] [3]);
  or (_07559_, _06936_, _07558_);
  and (_07560_, _07559_, _07084_);
  nand (_07561_, _07560_, _07557_);
  not (_07562_, \oc8051_golden_model_1.IRAM[4] [3]);
  or (_07563_, _06936_, _07562_);
  not (_07564_, \oc8051_golden_model_1.IRAM[5] [3]);
  or (_07565_, _07078_, _07564_);
  and (_07566_, _07565_, _07076_);
  nand (_07567_, _07566_, _07563_);
  nand (_07568_, _07567_, _07561_);
  nand (_07569_, _07568_, _07091_);
  nand (_07570_, _07569_, _07555_);
  nand (_07571_, _07570_, _06580_);
  nand (_07572_, _06936_, \oc8051_golden_model_1.IRAM[11] [3]);
  nand (_07573_, _07078_, \oc8051_golden_model_1.IRAM[10] [3]);
  and (_07574_, _07573_, _07084_);
  nand (_07575_, _07574_, _07572_);
  nand (_07576_, _07078_, \oc8051_golden_model_1.IRAM[8] [3]);
  nand (_07577_, _06936_, \oc8051_golden_model_1.IRAM[9] [3]);
  and (_07578_, _07577_, _07076_);
  nand (_07579_, _07578_, _07576_);
  nand (_07580_, _07579_, _07575_);
  nand (_07581_, _07580_, _06769_);
  nand (_07582_, _06936_, \oc8051_golden_model_1.IRAM[15] [3]);
  nand (_07583_, _07078_, \oc8051_golden_model_1.IRAM[14] [3]);
  and (_07584_, _07583_, _07084_);
  nand (_07585_, _07584_, _07582_);
  nand (_07586_, _07078_, \oc8051_golden_model_1.IRAM[12] [3]);
  nand (_07587_, _06936_, \oc8051_golden_model_1.IRAM[13] [3]);
  and (_07588_, _07587_, _07076_);
  nand (_07589_, _07588_, _07586_);
  nand (_07590_, _07589_, _07585_);
  nand (_07591_, _07590_, _07091_);
  nand (_07592_, _07591_, _07581_);
  nand (_07593_, _07592_, _07108_);
  nand (_07594_, _07593_, _07571_);
  not (_07595_, _07594_);
  or (_07596_, _07595_, _07541_);
  and (_07597_, _07594_, _07224_);
  and (_07598_, \oc8051_golden_model_1.SP [1], \oc8051_golden_model_1.SP [0]);
  and (_07599_, _07598_, \oc8051_golden_model_1.SP [2]);
  nor (_07600_, _07599_, \oc8051_golden_model_1.SP [3]);
  and (_07601_, \oc8051_golden_model_1.SP [2], \oc8051_golden_model_1.SP [1]);
  and (_07602_, _07601_, \oc8051_golden_model_1.SP [3]);
  and (_07603_, _07602_, \oc8051_golden_model_1.SP [0]);
  nor (_07604_, _07603_, _07600_);
  not (_07605_, _07604_);
  nor (_07606_, _07605_, _05978_);
  not (_07607_, _06317_);
  and (_07608_, _07607_, _07196_);
  and (_07609_, _07594_, _07197_);
  nor (_07610_, _07605_, _06007_);
  not (_07611_, _06010_);
  and (_07612_, _07594_, _07154_);
  and (_07613_, _07604_, _06758_);
  and (_07614_, _07594_, _06276_);
  not (_07615_, \oc8051_golden_model_1.PSW [3]);
  and (_07616_, _06018_, _07615_);
  nor (_07617_, _07616_, _07614_);
  nor (_07618_, _07617_, _07143_);
  and (_07619_, _07143_, _06213_);
  nor (_07620_, _07619_, _06758_);
  not (_07621_, _07620_);
  nor (_07622_, _07621_, _07618_);
  or (_07623_, _07622_, _07154_);
  nor (_07624_, _07623_, _07613_);
  or (_07625_, _07624_, _07152_);
  nor (_07626_, _07625_, _07612_);
  and (_07627_, _07152_, _06473_);
  or (_07628_, _07627_, _06275_);
  nor (_07629_, _07628_, _07626_);
  and (_07630_, _06318_, _06272_);
  nor (_07631_, _07630_, _07629_);
  nor (_07632_, _07631_, _07611_);
  nor (_07633_, _07604_, _06010_);
  nor (_07634_, _07633_, _07167_);
  not (_07635_, _07634_);
  nor (_07636_, _07635_, _07632_);
  and (_07637_, _07167_, _06473_);
  nor (_07638_, _07637_, _07174_);
  not (_07639_, _07638_);
  nor (_07640_, _07639_, _07636_);
  and (_07641_, _07594_, _07174_);
  nor (_07642_, _07641_, _07180_);
  not (_07643_, _07642_);
  nor (_07644_, _07643_, _07640_);
  and (_07645_, _07180_, _06473_);
  nor (_07646_, _07645_, _07179_);
  not (_07647_, _07646_);
  nor (_07648_, _07647_, _07644_);
  and (_07649_, _06318_, _07179_);
  nor (_07650_, _07649_, _07648_);
  and (_07651_, _07650_, _07303_);
  and (_07652_, _07604_, _06267_);
  nor (_07653_, _07652_, _07651_);
  nor (_07654_, _07653_, _06264_);
  and (_07655_, _06264_, _06320_);
  or (_07656_, _07655_, _07654_);
  and (_07657_, _07656_, _06007_);
  or (_07658_, _07657_, _07197_);
  nor (_07659_, _07658_, _07610_);
  or (_07660_, _07659_, _07196_);
  nor (_07661_, _07660_, _07609_);
  nor (_07662_, _07661_, _07608_);
  nor (_07663_, _07662_, _06254_);
  nor (_07664_, _07663_, _07606_);
  or (_07665_, _07664_, _07218_);
  nand (_07666_, _07218_, _06473_);
  and (_07667_, _07666_, _07225_);
  and (_07668_, _07667_, _07665_);
  or (_07669_, _07668_, _06220_);
  nor (_07670_, _07669_, _07597_);
  nor (_07671_, _06219_, _06214_);
  nor (_07672_, _07671_, _07670_);
  nor (_07673_, _07672_, _06217_);
  nor (_07674_, _07605_, _05952_);
  not (_07675_, _07674_);
  and (_07676_, _07675_, _07246_);
  not (_07677_, _07676_);
  nor (_07678_, _07677_, _07673_);
  nor (_07679_, _07246_, _06473_);
  nor (_07680_, _07679_, _07233_);
  not (_07681_, _07680_);
  nor (_07682_, _07681_, _07678_);
  nor (_07683_, _07605_, _05961_);
  or (_07684_, _07683_, _07254_);
  nor (_07685_, _07684_, _07682_);
  and (_07686_, _07254_, _06213_);
  or (_07687_, _07686_, _07253_);
  nor (_07688_, _07687_, _07685_);
  nor (_07689_, _07605_, _05959_);
  nor (_07690_, _07689_, _07435_);
  not (_07691_, _07690_);
  nor (_07692_, _07691_, _07688_);
  nor (_07693_, _07692_, _07261_);
  and (_07694_, _07693_, _07596_);
  not (_07695_, _07271_);
  and (_07696_, _07261_, _06473_);
  nor (_07697_, _07696_, _07695_);
  not (_07698_, _07697_);
  nor (_07699_, _07698_, _07694_);
  nor (_07700_, _07604_, _07271_);
  nor (_07701_, _07700_, _07270_);
  not (_07702_, _07701_);
  nor (_07703_, _07702_, _07699_);
  nor (_07704_, _07703_, _07281_);
  and (_07705_, _07704_, _07540_);
  and (_07706_, _07594_, _07281_);
  nor (_07707_, _07706_, _07286_);
  not (_07708_, _07707_);
  nor (_07709_, _07708_, _07705_);
  nor (_07710_, _06279_, _06214_);
  nor (_07711_, _07710_, _07709_);
  and (_07712_, _07286_, _06657_);
  and (_07713_, _06612_, _05927_);
  nor (_07714_, _07598_, \oc8051_golden_model_1.SP [2]);
  nor (_07715_, _07714_, _07599_);
  not (_07716_, _07715_);
  nor (_07717_, _07716_, _05959_);
  and (_07718_, _06657_, _06220_);
  and (_07719_, _06612_, _06257_);
  and (_07720_, _07715_, _06267_);
  and (_07721_, _07152_, _06657_);
  not (_07722_, \oc8051_golden_model_1.IRAM[0] [2]);
  or (_07723_, _06936_, _07722_);
  not (_07724_, \oc8051_golden_model_1.IRAM[1] [2]);
  or (_07725_, _07078_, _07724_);
  and (_07726_, _07725_, _07076_);
  nand (_07727_, _07726_, _07723_);
  not (_07728_, \oc8051_golden_model_1.IRAM[3] [2]);
  or (_07729_, _07078_, _07728_);
  not (_07730_, \oc8051_golden_model_1.IRAM[2] [2]);
  or (_07731_, _06936_, _07730_);
  and (_07732_, _07731_, _07084_);
  nand (_07733_, _07732_, _07729_);
  nand (_07734_, _07733_, _07727_);
  nand (_07735_, _07734_, _06769_);
  not (_07736_, \oc8051_golden_model_1.IRAM[7] [2]);
  or (_07737_, _07078_, _07736_);
  not (_07738_, \oc8051_golden_model_1.IRAM[6] [2]);
  or (_07739_, _06936_, _07738_);
  and (_07740_, _07739_, _07084_);
  nand (_07741_, _07740_, _07737_);
  not (_07742_, \oc8051_golden_model_1.IRAM[4] [2]);
  or (_07743_, _06936_, _07742_);
  not (_07744_, \oc8051_golden_model_1.IRAM[5] [2]);
  or (_07745_, _07078_, _07744_);
  and (_07746_, _07745_, _07076_);
  nand (_07747_, _07746_, _07743_);
  nand (_07748_, _07747_, _07741_);
  nand (_07749_, _07748_, _07091_);
  nand (_07750_, _07749_, _07735_);
  nand (_07751_, _07750_, _06580_);
  nand (_07752_, _06936_, \oc8051_golden_model_1.IRAM[11] [2]);
  nand (_07753_, _07078_, \oc8051_golden_model_1.IRAM[10] [2]);
  and (_07754_, _07753_, _07084_);
  nand (_07755_, _07754_, _07752_);
  nand (_07756_, _07078_, \oc8051_golden_model_1.IRAM[8] [2]);
  nand (_07757_, _06936_, \oc8051_golden_model_1.IRAM[9] [2]);
  and (_07758_, _07757_, _07076_);
  nand (_07759_, _07758_, _07756_);
  nand (_07760_, _07759_, _07755_);
  nand (_07761_, _07760_, _06769_);
  not (_07762_, \oc8051_golden_model_1.IRAM[15] [2]);
  or (_07763_, _07078_, _07762_);
  not (_07764_, \oc8051_golden_model_1.IRAM[14] [2]);
  or (_07765_, _06936_, _07764_);
  and (_07766_, _07765_, _07084_);
  nand (_07767_, _07766_, _07763_);
  nand (_07768_, _07078_, \oc8051_golden_model_1.IRAM[12] [2]);
  nand (_07769_, _06936_, \oc8051_golden_model_1.IRAM[13] [2]);
  and (_07770_, _07769_, _07076_);
  nand (_07771_, _07770_, _07768_);
  nand (_07772_, _07771_, _07767_);
  nand (_07773_, _07772_, _07091_);
  nand (_07774_, _07773_, _07761_);
  nand (_07775_, _07774_, _07108_);
  nand (_07776_, _07775_, _07751_);
  or (_07777_, _07776_, _05934_);
  and (_07778_, _07777_, _07485_);
  and (_07779_, _07143_, _06656_);
  nor (_07780_, _07779_, _07778_);
  and (_07781_, _07716_, _06758_);
  and (_07782_, _06336_, _06271_);
  nor (_07783_, _07782_, _07781_);
  and (_07784_, _07783_, _07780_);
  and (_07785_, _07776_, _07154_);
  nor (_07786_, _07785_, _07152_);
  and (_07787_, _07786_, _07784_);
  nor (_07788_, _07787_, _07721_);
  nor (_07789_, _07788_, _06275_);
  nor (_07790_, _07789_, _06623_);
  nor (_07791_, _07715_, _06010_);
  nor (_07792_, _07791_, _07790_);
  and (_07793_, _07167_, _06656_);
  and (_07794_, _06336_, _06266_);
  nor (_07795_, _07794_, _07793_);
  and (_07796_, _07795_, _07792_);
  and (_07797_, _07776_, _07174_);
  nor (_07798_, _07797_, _07180_);
  and (_07799_, _07798_, _07796_);
  and (_07800_, _07180_, _06657_);
  nor (_07801_, _07800_, _07799_);
  and (_07802_, _06611_, _07179_);
  nor (_07803_, _07802_, _07801_);
  and (_07804_, _07803_, _07303_);
  nor (_07805_, _07804_, _07720_);
  and (_07806_, _06264_, _06611_);
  or (_07807_, _07806_, _07805_);
  nor (_07808_, _07715_, _06007_);
  nor (_07809_, _07808_, _06498_);
  not (_07810_, _07809_);
  nor (_07811_, _07810_, _07807_);
  and (_07812_, _07776_, _07197_);
  nor (_07813_, _07812_, _07196_);
  and (_07814_, _07813_, _07811_);
  nor (_07815_, _07814_, _07719_);
  nor (_07816_, _07815_, _06254_);
  nor (_07817_, _07716_, _05978_);
  nor (_07818_, _07817_, _07816_);
  and (_07819_, _07218_, _06656_);
  and (_07820_, _06336_, _06321_);
  nor (_07821_, _07820_, _07819_);
  not (_07822_, _07821_);
  nor (_07823_, _07822_, _07818_);
  and (_07824_, _07776_, _07224_);
  nor (_07825_, _07824_, _06220_);
  and (_07826_, _07825_, _07823_);
  nor (_07827_, _07826_, _07718_);
  nor (_07828_, _07827_, _06217_);
  nor (_07829_, _07716_, _05952_);
  nor (_07830_, _07829_, _07828_);
  nor (_07831_, _07246_, _06657_);
  nor (_07832_, _07831_, _07233_);
  not (_07833_, _07832_);
  nor (_07834_, _07833_, _07830_);
  nor (_07835_, _07716_, _05961_);
  nor (_07836_, _07835_, _07834_);
  and (_07837_, _07254_, _06656_);
  or (_07838_, _07837_, _07253_);
  nor (_07839_, _07838_, _07836_);
  nor (_07840_, _07839_, _07717_);
  and (_07841_, _06336_, _05779_);
  nor (_07842_, _07841_, _07840_);
  and (_07843_, _07776_, _07435_);
  nor (_07844_, _07843_, _07261_);
  and (_07845_, _07844_, _07842_);
  and (_07846_, _07261_, _06657_);
  nor (_07847_, _07846_, _07845_);
  nor (_07848_, _07715_, _07271_);
  nor (_07849_, _07848_, _07270_);
  not (_07850_, _07849_);
  nor (_07851_, _07850_, _07847_);
  nor (_07852_, _07851_, _07713_);
  and (_07853_, _06336_, _05938_);
  nor (_07854_, _07853_, _07852_);
  and (_07855_, _07776_, _07281_);
  nor (_07856_, _07855_, _07286_);
  and (_07857_, _07856_, _07854_);
  nor (_07858_, _07857_, _07712_);
  nor (_07859_, _07858_, _07536_);
  not (_07860_, _07859_);
  nor (_07861_, _07860_, _07711_);
  and (_07862_, _07861_, _07538_);
  or (_07863_, _07862_, \oc8051_golden_model_1.IRAM[15] [7]);
  nand (_07864_, _07601_, _06800_);
  or (_07865_, _07715_, _07296_);
  and (_07866_, _07865_, _07864_);
  and (_07867_, _07602_, _06800_);
  and (_07868_, _07864_, _07605_);
  nor (_07869_, _07868_, _07867_);
  and (_07870_, _07509_, _07504_);
  and (_07871_, _07870_, _07496_);
  nor (_07872_, _07871_, _07454_);
  and (_07873_, _07872_, _07869_);
  and (_07874_, _07873_, _07866_);
  and (_07875_, _07874_, _07295_);
  not (_07876_, _07875_);
  and (_07877_, _07876_, _07863_);
  not (_07878_, _07862_);
  and (_07879_, _06656_, _06473_);
  and (_07880_, _07004_, _06252_);
  and (_07881_, _07880_, _07879_);
  and (_07882_, _06317_, _06182_);
  not (_07883_, _06968_);
  and (_07884_, _07883_, _06611_);
  and (_07885_, _07884_, _07882_);
  and (_07886_, _07885_, _07881_);
  and (_07887_, _07886_, \oc8051_golden_model_1.SBUF [7]);
  not (_07888_, _07887_);
  and (_07889_, _07004_, _06251_);
  and (_07890_, _06656_, _06213_);
  and (_07891_, _07890_, _07889_);
  nor (_07892_, _06968_, _06611_);
  and (_07893_, _07892_, _07882_);
  and (_07894_, _07893_, _07891_);
  and (_07895_, _07894_, \oc8051_golden_model_1.P3 [7]);
  not (_07896_, _06611_);
  and (_07897_, _06968_, _07896_);
  and (_07898_, _07897_, _07882_);
  and (_07899_, _07889_, _07879_);
  and (_07900_, _07899_, _07898_);
  and (_07901_, _07900_, \oc8051_golden_model_1.IE [7]);
  nor (_07902_, _07901_, _07895_);
  and (_07903_, _07902_, _07888_);
  and (_07904_, _07898_, _07891_);
  and (_07905_, _07904_, \oc8051_golden_model_1.P2 [7]);
  and (_07906_, _06968_, _06611_);
  and (_07907_, _07906_, _07882_);
  nor (_07908_, _06656_, _06213_);
  and (_07909_, _07880_, _07908_);
  and (_07910_, _07909_, _07907_);
  and (_07911_, _07910_, \oc8051_golden_model_1.TH1 [7]);
  nor (_07912_, _07911_, _07905_);
  and (_07913_, _07912_, _07903_);
  and (_07914_, _07881_, _07907_);
  and (_07915_, _07914_, \oc8051_golden_model_1.TMOD [7]);
  not (_07916_, _07915_);
  nor (_07917_, _07004_, _06252_);
  and (_07918_, _07879_, _07917_);
  and (_07919_, _07918_, _07907_);
  and (_07920_, _07919_, \oc8051_golden_model_1.TL0 [7]);
  and (_07921_, _07908_, _07889_);
  and (_07922_, _07921_, _07907_);
  and (_07923_, _07922_, \oc8051_golden_model_1.TH0 [7]);
  nor (_07924_, _07923_, _07920_);
  and (_07925_, _07924_, _07916_);
  and (_07926_, _07891_, _07907_);
  and (_07927_, _07926_, \oc8051_golden_model_1.P0 [7]);
  and (_07928_, _07899_, _07907_);
  and (_07929_, _07928_, \oc8051_golden_model_1.TCON [7]);
  nor (_07930_, _07929_, _07927_);
  and (_07931_, _07930_, _07925_);
  and (_07932_, _07931_, _07913_);
  nor (_07933_, _06317_, _06286_);
  and (_07934_, _07933_, _07884_);
  and (_07935_, _07934_, _07891_);
  and (_07936_, _07935_, \oc8051_golden_model_1.PSW [7]);
  not (_07937_, _07936_);
  and (_07938_, _07933_, _07897_);
  and (_07939_, _07938_, _07891_);
  and (_07940_, _07939_, \oc8051_golden_model_1.ACC [7]);
  and (_07941_, _07933_, _07892_);
  and (_07942_, _07941_, _07891_);
  and (_07943_, _07942_, \oc8051_golden_model_1.B [7]);
  nor (_07944_, _07943_, _07940_);
  and (_07945_, _07944_, _07937_);
  and (_07946_, _07899_, _07893_);
  and (_07947_, _07946_, \oc8051_golden_model_1.IP [7]);
  and (_07948_, _07907_, _06213_);
  nor (_07949_, _07004_, _06251_);
  and (_07950_, _07949_, _06657_);
  and (_07951_, _07950_, _07948_);
  and (_07952_, _07951_, \oc8051_golden_model_1.PCON [7]);
  nor (_07953_, _07952_, _07947_);
  and (_07954_, _07953_, _07945_);
  and (_07955_, _07880_, _07890_);
  and (_07956_, _07955_, _07907_);
  and (_07957_, _07956_, \oc8051_golden_model_1.SP [7]);
  not (_07958_, _07957_);
  and (_07959_, _07917_, _06656_);
  and (_07960_, _07959_, _07948_);
  and (_07961_, _07960_, \oc8051_golden_model_1.DPL [7]);
  and (_07962_, _07949_, _07890_);
  and (_07963_, _07962_, _07907_);
  and (_07964_, _07963_, \oc8051_golden_model_1.DPH [7]);
  nor (_07965_, _07964_, _07961_);
  and (_07966_, _07965_, _07958_);
  and (_07967_, _07949_, _07879_);
  and (_07968_, _07967_, _07907_);
  and (_07969_, _07968_, \oc8051_golden_model_1.TL1 [7]);
  not (_07970_, _07969_);
  and (_07971_, _07885_, _07891_);
  and (_07972_, _07971_, \oc8051_golden_model_1.P1 [7]);
  and (_07973_, _07899_, _07885_);
  and (_07974_, _07973_, \oc8051_golden_model_1.SCON [7]);
  nor (_07975_, _07974_, _07972_);
  and (_07976_, _07975_, _07970_);
  and (_07977_, _07976_, _07966_);
  and (_07978_, _07977_, _07954_);
  and (_07979_, _07978_, _07932_);
  not (_07980_, \oc8051_golden_model_1.IRAM[0] [7]);
  or (_07981_, _06936_, _07980_);
  not (_07982_, \oc8051_golden_model_1.IRAM[1] [7]);
  or (_07983_, _07078_, _07982_);
  and (_07984_, _07983_, _07076_);
  nand (_07985_, _07984_, _07981_);
  not (_07986_, \oc8051_golden_model_1.IRAM[3] [7]);
  or (_07987_, _07078_, _07986_);
  not (_07988_, \oc8051_golden_model_1.IRAM[2] [7]);
  or (_07989_, _06936_, _07988_);
  and (_07990_, _07989_, _07084_);
  nand (_07991_, _07990_, _07987_);
  nand (_07992_, _07991_, _07985_);
  nand (_07993_, _07992_, _06769_);
  not (_07994_, \oc8051_golden_model_1.IRAM[7] [7]);
  or (_07995_, _07078_, _07994_);
  not (_07996_, \oc8051_golden_model_1.IRAM[6] [7]);
  or (_07997_, _06936_, _07996_);
  and (_07998_, _07997_, _07084_);
  nand (_07999_, _07998_, _07995_);
  not (_08000_, \oc8051_golden_model_1.IRAM[4] [7]);
  or (_08001_, _06936_, _08000_);
  not (_08002_, \oc8051_golden_model_1.IRAM[5] [7]);
  or (_08003_, _07078_, _08002_);
  and (_08004_, _08003_, _07076_);
  nand (_08005_, _08004_, _08001_);
  nand (_08006_, _08005_, _07999_);
  nand (_08007_, _08006_, _07091_);
  nand (_08008_, _08007_, _07993_);
  nand (_08009_, _08008_, _06580_);
  not (_08010_, \oc8051_golden_model_1.IRAM[11] [7]);
  or (_08011_, _07078_, _08010_);
  not (_08012_, \oc8051_golden_model_1.IRAM[10] [7]);
  or (_08013_, _06936_, _08012_);
  and (_08014_, _08013_, _07084_);
  nand (_08015_, _08014_, _08011_);
  not (_08016_, \oc8051_golden_model_1.IRAM[8] [7]);
  or (_08017_, _06936_, _08016_);
  not (_08018_, \oc8051_golden_model_1.IRAM[9] [7]);
  or (_08019_, _07078_, _08018_);
  and (_08020_, _08019_, _07076_);
  nand (_08021_, _08020_, _08017_);
  nand (_08022_, _08021_, _08015_);
  nand (_08023_, _08022_, _06769_);
  not (_08024_, \oc8051_golden_model_1.IRAM[15] [7]);
  or (_08025_, _07078_, _08024_);
  not (_08026_, \oc8051_golden_model_1.IRAM[14] [7]);
  or (_08027_, _06936_, _08026_);
  and (_08028_, _08027_, _07084_);
  nand (_08029_, _08028_, _08025_);
  not (_08030_, \oc8051_golden_model_1.IRAM[12] [7]);
  or (_08031_, _06936_, _08030_);
  not (_08032_, \oc8051_golden_model_1.IRAM[13] [7]);
  or (_08033_, _07078_, _08032_);
  and (_08034_, _08033_, _07076_);
  nand (_08035_, _08034_, _08031_);
  nand (_08036_, _08035_, _08029_);
  nand (_08037_, _08036_, _07091_);
  nand (_08038_, _08037_, _08023_);
  nand (_08039_, _08038_, _07108_);
  nand (_08040_, _08039_, _08009_);
  or (_08041_, _08040_, _06182_);
  and (_08042_, _08041_, _07979_);
  not (_08043_, _08042_);
  and (_08044_, _07904_, \oc8051_golden_model_1.P2 [6]);
  not (_08045_, _08044_);
  and (_08046_, _07886_, \oc8051_golden_model_1.SBUF [6]);
  not (_08047_, _08046_);
  and (_08048_, _07894_, \oc8051_golden_model_1.P3 [6]);
  and (_08049_, _07900_, \oc8051_golden_model_1.IE [6]);
  nor (_08050_, _08049_, _08048_);
  and (_08051_, _08050_, _08047_);
  and (_08052_, _08051_, _08045_);
  and (_08053_, _07926_, \oc8051_golden_model_1.P0 [6]);
  not (_08054_, _08053_);
  and (_08055_, _07960_, \oc8051_golden_model_1.DPL [6]);
  and (_08056_, _07963_, \oc8051_golden_model_1.DPH [6]);
  nor (_08057_, _08056_, _08055_);
  and (_08058_, _08057_, _08054_);
  and (_08059_, _07971_, \oc8051_golden_model_1.P1 [6]);
  and (_08060_, _07973_, \oc8051_golden_model_1.SCON [6]);
  nor (_08061_, _08060_, _08059_);
  and (_08062_, _07968_, \oc8051_golden_model_1.TL1 [6]);
  and (_08063_, _07910_, \oc8051_golden_model_1.TH1 [6]);
  nor (_08064_, _08063_, _08062_);
  and (_08065_, _08064_, _08061_);
  and (_08066_, _08065_, _08058_);
  and (_08067_, _08066_, _08052_);
  and (_08068_, _07935_, \oc8051_golden_model_1.PSW [6]);
  not (_08069_, _08068_);
  and (_08070_, _07942_, \oc8051_golden_model_1.B [6]);
  and (_08071_, _07939_, \oc8051_golden_model_1.ACC [6]);
  nor (_08072_, _08071_, _08070_);
  and (_08073_, _08072_, _08069_);
  and (_08074_, _07946_, \oc8051_golden_model_1.IP [6]);
  and (_08075_, _07951_, \oc8051_golden_model_1.PCON [6]);
  nor (_08076_, _08075_, _08074_);
  and (_08077_, _08076_, _08073_);
  and (_08078_, _07928_, \oc8051_golden_model_1.TCON [6]);
  not (_08079_, _08078_);
  and (_08080_, _07922_, \oc8051_golden_model_1.TH0 [6]);
  and (_08081_, _07919_, \oc8051_golden_model_1.TL0 [6]);
  nor (_08082_, _08081_, _08080_);
  and (_08083_, _08082_, _08079_);
  and (_08084_, _07914_, \oc8051_golden_model_1.TMOD [6]);
  and (_08085_, _07956_, \oc8051_golden_model_1.SP [6]);
  nor (_08086_, _08085_, _08084_);
  and (_08087_, _08086_, _08083_);
  and (_08088_, _08087_, _08077_);
  and (_08089_, _08088_, _08067_);
  not (_08090_, \oc8051_golden_model_1.IRAM[0] [6]);
  or (_08091_, _06936_, _08090_);
  not (_08092_, \oc8051_golden_model_1.IRAM[1] [6]);
  or (_08093_, _07078_, _08092_);
  and (_08094_, _08093_, _07076_);
  nand (_08095_, _08094_, _08091_);
  not (_08096_, \oc8051_golden_model_1.IRAM[3] [6]);
  or (_08097_, _07078_, _08096_);
  not (_08098_, \oc8051_golden_model_1.IRAM[2] [6]);
  or (_08099_, _06936_, _08098_);
  and (_08100_, _08099_, _07084_);
  nand (_08101_, _08100_, _08097_);
  nand (_08102_, _08101_, _08095_);
  nand (_08103_, _08102_, _06769_);
  not (_08104_, \oc8051_golden_model_1.IRAM[7] [6]);
  or (_08105_, _07078_, _08104_);
  not (_08106_, \oc8051_golden_model_1.IRAM[6] [6]);
  or (_08107_, _06936_, _08106_);
  and (_08108_, _08107_, _07084_);
  nand (_08109_, _08108_, _08105_);
  not (_08110_, \oc8051_golden_model_1.IRAM[4] [6]);
  or (_08111_, _06936_, _08110_);
  not (_08112_, \oc8051_golden_model_1.IRAM[5] [6]);
  or (_08113_, _07078_, _08112_);
  and (_08114_, _08113_, _07076_);
  nand (_08115_, _08114_, _08111_);
  nand (_08116_, _08115_, _08109_);
  nand (_08117_, _08116_, _07091_);
  nand (_08118_, _08117_, _08103_);
  nand (_08119_, _08118_, _06580_);
  nand (_08120_, _06936_, \oc8051_golden_model_1.IRAM[11] [6]);
  nand (_08121_, _07078_, \oc8051_golden_model_1.IRAM[10] [6]);
  and (_08122_, _08121_, _07084_);
  nand (_08123_, _08122_, _08120_);
  nand (_08124_, _07078_, \oc8051_golden_model_1.IRAM[8] [6]);
  nand (_08125_, _06936_, \oc8051_golden_model_1.IRAM[9] [6]);
  and (_08126_, _08125_, _07076_);
  nand (_08127_, _08126_, _08124_);
  nand (_08128_, _08127_, _08123_);
  nand (_08129_, _08128_, _06769_);
  nand (_08130_, _06936_, \oc8051_golden_model_1.IRAM[15] [6]);
  nand (_08131_, _07078_, \oc8051_golden_model_1.IRAM[14] [6]);
  and (_08132_, _08131_, _07084_);
  nand (_08133_, _08132_, _08130_);
  nand (_08134_, _07078_, \oc8051_golden_model_1.IRAM[12] [6]);
  nand (_08135_, _06936_, \oc8051_golden_model_1.IRAM[13] [6]);
  and (_08136_, _08135_, _07076_);
  nand (_08137_, _08136_, _08134_);
  nand (_08138_, _08137_, _08133_);
  nand (_08139_, _08138_, _07091_);
  nand (_08140_, _08139_, _08129_);
  nand (_08141_, _08140_, _07108_);
  nand (_08142_, _08141_, _08119_);
  or (_08143_, _08142_, _06182_);
  and (_08144_, _08143_, _08089_);
  not (_08145_, _08144_);
  and (_08146_, _07935_, \oc8051_golden_model_1.PSW [5]);
  and (_08147_, _07942_, \oc8051_golden_model_1.B [5]);
  nor (_08148_, _08147_, _08146_);
  and (_08149_, _07973_, \oc8051_golden_model_1.SCON [5]);
  and (_08150_, _07894_, \oc8051_golden_model_1.P3 [5]);
  nor (_08151_, _08150_, _08149_);
  and (_08152_, _08151_, _08148_);
  and (_08153_, _07919_, \oc8051_golden_model_1.TL0 [5]);
  and (_08154_, _07939_, \oc8051_golden_model_1.ACC [5]);
  nor (_08155_, _08154_, _08153_);
  and (_08156_, _07922_, \oc8051_golden_model_1.TH0 [5]);
  and (_08157_, _07904_, \oc8051_golden_model_1.P2 [5]);
  nor (_08158_, _08157_, _08156_);
  and (_08159_, _08158_, _08155_);
  and (_08160_, _07971_, \oc8051_golden_model_1.P1 [5]);
  and (_08161_, _07900_, \oc8051_golden_model_1.IE [5]);
  nor (_08162_, _08161_, _08160_);
  and (_08163_, _07886_, \oc8051_golden_model_1.SBUF [5]);
  and (_08164_, _07946_, \oc8051_golden_model_1.IP [5]);
  nor (_08165_, _08164_, _08163_);
  and (_08166_, _08165_, _08162_);
  and (_08167_, _08166_, _08159_);
  and (_08168_, _08167_, _08152_);
  and (_08169_, _07926_, \oc8051_golden_model_1.P0 [5]);
  not (_08170_, _08169_);
  and (_08171_, _07960_, \oc8051_golden_model_1.DPL [5]);
  and (_08172_, _07880_, _06656_);
  and (_08173_, _07948_, _08172_);
  and (_08174_, _08173_, \oc8051_golden_model_1.SP [5]);
  nor (_08175_, _08174_, _08171_);
  and (_08176_, _08175_, _08170_);
  and (_08177_, _07928_, \oc8051_golden_model_1.TCON [5]);
  and (_08178_, _07914_, \oc8051_golden_model_1.TMOD [5]);
  nor (_08179_, _08178_, _08177_);
  and (_08180_, _07968_, \oc8051_golden_model_1.TL1 [5]);
  and (_08181_, _07910_, \oc8051_golden_model_1.TH1 [5]);
  nor (_08182_, _08181_, _08180_);
  and (_08183_, _08182_, _08179_);
  and (_08184_, _07951_, \oc8051_golden_model_1.PCON [5]);
  and (_08185_, _07949_, _06656_);
  and (_08186_, _08185_, _07948_);
  and (_08187_, _08186_, \oc8051_golden_model_1.DPH [5]);
  nor (_08188_, _08187_, _08184_);
  and (_08189_, _08188_, _08183_);
  and (_08190_, _08189_, _08176_);
  and (_08191_, _08190_, _08168_);
  not (_08192_, \oc8051_golden_model_1.IRAM[0] [5]);
  or (_08193_, _06936_, _08192_);
  not (_08194_, \oc8051_golden_model_1.IRAM[1] [5]);
  or (_08195_, _07078_, _08194_);
  and (_08196_, _08195_, _07076_);
  nand (_08197_, _08196_, _08193_);
  not (_08198_, \oc8051_golden_model_1.IRAM[3] [5]);
  or (_08199_, _07078_, _08198_);
  not (_08200_, \oc8051_golden_model_1.IRAM[2] [5]);
  or (_08201_, _06936_, _08200_);
  and (_08202_, _08201_, _07084_);
  nand (_08203_, _08202_, _08199_);
  nand (_08204_, _08203_, _08197_);
  nand (_08205_, _08204_, _06769_);
  not (_08206_, \oc8051_golden_model_1.IRAM[7] [5]);
  or (_08207_, _07078_, _08206_);
  not (_08208_, \oc8051_golden_model_1.IRAM[6] [5]);
  or (_08209_, _06936_, _08208_);
  and (_08210_, _08209_, _07084_);
  nand (_08211_, _08210_, _08207_);
  not (_08212_, \oc8051_golden_model_1.IRAM[4] [5]);
  or (_08213_, _06936_, _08212_);
  not (_08214_, \oc8051_golden_model_1.IRAM[5] [5]);
  or (_08215_, _07078_, _08214_);
  and (_08216_, _08215_, _07076_);
  nand (_08217_, _08216_, _08213_);
  nand (_08218_, _08217_, _08211_);
  nand (_08219_, _08218_, _07091_);
  nand (_08220_, _08219_, _08205_);
  nand (_08221_, _08220_, _06580_);
  nand (_08222_, _06936_, \oc8051_golden_model_1.IRAM[11] [5]);
  nand (_08223_, _07078_, \oc8051_golden_model_1.IRAM[10] [5]);
  and (_08224_, _08223_, _07084_);
  nand (_08225_, _08224_, _08222_);
  nand (_08226_, _07078_, \oc8051_golden_model_1.IRAM[8] [5]);
  nand (_08227_, _06936_, \oc8051_golden_model_1.IRAM[9] [5]);
  and (_08228_, _08227_, _07076_);
  nand (_08229_, _08228_, _08226_);
  nand (_08230_, _08229_, _08225_);
  nand (_08231_, _08230_, _06769_);
  nand (_08232_, _06936_, \oc8051_golden_model_1.IRAM[15] [5]);
  nand (_08233_, _07078_, \oc8051_golden_model_1.IRAM[14] [5]);
  and (_08234_, _08233_, _07084_);
  nand (_08235_, _08234_, _08232_);
  nand (_08236_, _07078_, \oc8051_golden_model_1.IRAM[12] [5]);
  nand (_08237_, _06936_, \oc8051_golden_model_1.IRAM[13] [5]);
  and (_08238_, _08237_, _07076_);
  nand (_08239_, _08238_, _08236_);
  nand (_08240_, _08239_, _08235_);
  nand (_08241_, _08240_, _07091_);
  nand (_08242_, _08241_, _08231_);
  nand (_08243_, _08242_, _07108_);
  nand (_08244_, _08243_, _08221_);
  or (_08245_, _08244_, _06182_);
  and (_08246_, _08245_, _08191_);
  not (_08247_, _08246_);
  and (_08248_, _07900_, \oc8051_golden_model_1.IE [3]);
  and (_08249_, _07946_, \oc8051_golden_model_1.IP [3]);
  nor (_08250_, _08249_, _08248_);
  and (_08251_, _07886_, \oc8051_golden_model_1.SBUF [3]);
  and (_08252_, _07904_, \oc8051_golden_model_1.P2 [3]);
  nor (_08253_, _08252_, _08251_);
  and (_08254_, _08253_, _08250_);
  and (_08255_, _07894_, \oc8051_golden_model_1.P3 [3]);
  and (_08256_, _07939_, \oc8051_golden_model_1.ACC [3]);
  nor (_08257_, _08256_, _08255_);
  and (_08258_, _07935_, \oc8051_golden_model_1.PSW [3]);
  and (_08259_, _07942_, \oc8051_golden_model_1.B [3]);
  nor (_08260_, _08259_, _08258_);
  and (_08261_, _08260_, _08257_);
  and (_08262_, _07971_, \oc8051_golden_model_1.P1 [3]);
  and (_08263_, _07973_, \oc8051_golden_model_1.SCON [3]);
  nor (_08264_, _08263_, _08262_);
  and (_08265_, _07919_, \oc8051_golden_model_1.TL0 [3]);
  and (_08266_, _07922_, \oc8051_golden_model_1.TH0 [3]);
  nor (_08267_, _08266_, _08265_);
  and (_08268_, _08267_, _08264_);
  and (_08269_, _08268_, _08261_);
  and (_08270_, _08269_, _08254_);
  and (_08271_, _07926_, \oc8051_golden_model_1.P0 [3]);
  not (_08272_, _08271_);
  and (_08273_, _07960_, \oc8051_golden_model_1.DPL [3]);
  and (_08274_, _08173_, \oc8051_golden_model_1.SP [3]);
  nor (_08275_, _08274_, _08273_);
  and (_08276_, _08275_, _08272_);
  and (_08277_, _07928_, \oc8051_golden_model_1.TCON [3]);
  and (_08278_, _07914_, \oc8051_golden_model_1.TMOD [3]);
  nor (_08279_, _08278_, _08277_);
  and (_08280_, _07968_, \oc8051_golden_model_1.TL1 [3]);
  and (_08281_, _07910_, \oc8051_golden_model_1.TH1 [3]);
  nor (_08282_, _08281_, _08280_);
  and (_08283_, _08282_, _08279_);
  and (_08284_, _07951_, \oc8051_golden_model_1.PCON [3]);
  and (_08285_, _08186_, \oc8051_golden_model_1.DPH [3]);
  nor (_08286_, _08285_, _08284_);
  and (_08287_, _08286_, _08283_);
  and (_08288_, _08287_, _08276_);
  and (_08289_, _08288_, _08270_);
  or (_08290_, _07594_, _06182_);
  and (_08291_, _08290_, _08289_);
  not (_08292_, _08291_);
  and (_08293_, _07886_, \oc8051_golden_model_1.SBUF [1]);
  not (_08294_, _08293_);
  and (_08295_, _07900_, \oc8051_golden_model_1.IE [1]);
  and (_08296_, _07894_, \oc8051_golden_model_1.P3 [1]);
  nor (_08297_, _08296_, _08295_);
  and (_08298_, _08297_, _08294_);
  and (_08299_, _07904_, \oc8051_golden_model_1.P2 [1]);
  and (_08300_, _07968_, \oc8051_golden_model_1.TL1 [1]);
  nor (_08301_, _08300_, _08299_);
  and (_08302_, _08301_, _08298_);
  and (_08303_, _07914_, \oc8051_golden_model_1.TMOD [1]);
  not (_08304_, _08303_);
  and (_08305_, _07919_, \oc8051_golden_model_1.TL0 [1]);
  and (_08306_, _07922_, \oc8051_golden_model_1.TH0 [1]);
  nor (_08307_, _08306_, _08305_);
  and (_08308_, _08307_, _08304_);
  and (_08309_, _07928_, \oc8051_golden_model_1.TCON [1]);
  and (_08310_, _07956_, \oc8051_golden_model_1.SP [1]);
  nor (_08311_, _08310_, _08309_);
  and (_08312_, _08311_, _08308_);
  and (_08313_, _08312_, _08302_);
  and (_08314_, _07939_, \oc8051_golden_model_1.ACC [1]);
  and (_08315_, _07942_, \oc8051_golden_model_1.B [1]);
  nor (_08316_, _08315_, _08314_);
  and (_08317_, _07935_, \oc8051_golden_model_1.PSW [1]);
  not (_08318_, _08317_);
  and (_08319_, _08318_, _08316_);
  and (_08320_, _07946_, \oc8051_golden_model_1.IP [1]);
  and (_08321_, _07951_, \oc8051_golden_model_1.PCON [1]);
  nor (_08322_, _08321_, _08320_);
  and (_08323_, _08322_, _08319_);
  and (_08324_, _07926_, \oc8051_golden_model_1.P0 [1]);
  not (_08325_, _08324_);
  and (_08326_, _07960_, \oc8051_golden_model_1.DPL [1]);
  and (_08327_, _07963_, \oc8051_golden_model_1.DPH [1]);
  nor (_08328_, _08327_, _08326_);
  and (_08329_, _08328_, _08325_);
  and (_08330_, _07910_, \oc8051_golden_model_1.TH1 [1]);
  not (_08331_, _08330_);
  and (_08332_, _07973_, \oc8051_golden_model_1.SCON [1]);
  and (_08333_, _07971_, \oc8051_golden_model_1.P1 [1]);
  nor (_08334_, _08333_, _08332_);
  and (_08335_, _08334_, _08331_);
  and (_08336_, _08335_, _08329_);
  and (_08337_, _08336_, _08323_);
  and (_08338_, _08337_, _08313_);
  or (_08339_, _07357_, _06182_);
  and (_08340_, _08339_, _08338_);
  not (_08341_, _08340_);
  and (_08342_, _07904_, \oc8051_golden_model_1.P2 [0]);
  not (_08343_, _08342_);
  and (_08344_, _07886_, \oc8051_golden_model_1.SBUF [0]);
  not (_08345_, _08344_);
  and (_08346_, _07900_, \oc8051_golden_model_1.IE [0]);
  and (_08347_, _07894_, \oc8051_golden_model_1.P3 [0]);
  nor (_08348_, _08347_, _08346_);
  and (_08349_, _08348_, _08345_);
  and (_08350_, _08349_, _08343_);
  and (_08351_, _07960_, \oc8051_golden_model_1.DPL [0]);
  and (_08352_, _07963_, \oc8051_golden_model_1.DPH [0]);
  nor (_08353_, _08352_, _08351_);
  and (_08354_, _07926_, \oc8051_golden_model_1.P0 [0]);
  not (_08355_, _08354_);
  and (_08356_, _08355_, _08353_);
  and (_08357_, _07968_, \oc8051_golden_model_1.TL1 [0]);
  and (_08358_, _07910_, \oc8051_golden_model_1.TH1 [0]);
  nor (_08359_, _08358_, _08357_);
  and (_08360_, _07973_, \oc8051_golden_model_1.SCON [0]);
  and (_08361_, _07971_, \oc8051_golden_model_1.P1 [0]);
  nor (_08362_, _08361_, _08360_);
  and (_08363_, _08362_, _08359_);
  and (_08364_, _08363_, _08356_);
  and (_08365_, _08364_, _08350_);
  and (_08366_, _07935_, \oc8051_golden_model_1.PSW [0]);
  not (_08367_, _08366_);
  and (_08368_, _07939_, \oc8051_golden_model_1.ACC [0]);
  and (_08369_, _07942_, \oc8051_golden_model_1.B [0]);
  nor (_08370_, _08369_, _08368_);
  and (_08371_, _08370_, _08367_);
  and (_08372_, _07946_, \oc8051_golden_model_1.IP [0]);
  and (_08373_, _07951_, \oc8051_golden_model_1.PCON [0]);
  nor (_08374_, _08373_, _08372_);
  and (_08375_, _08374_, _08371_);
  and (_08376_, _07914_, \oc8051_golden_model_1.TMOD [0]);
  not (_08377_, _08376_);
  and (_08378_, _07919_, \oc8051_golden_model_1.TL0 [0]);
  and (_08379_, _07922_, \oc8051_golden_model_1.TH0 [0]);
  nor (_08380_, _08379_, _08378_);
  and (_08381_, _08380_, _08377_);
  and (_08382_, _07928_, \oc8051_golden_model_1.TCON [0]);
  and (_08383_, _07956_, \oc8051_golden_model_1.SP [0]);
  nor (_08384_, _08383_, _08382_);
  and (_08385_, _08384_, _08381_);
  and (_08386_, _08385_, _08375_);
  and (_08387_, _08386_, _08365_);
  not (_08388_, _08387_);
  and (_08389_, _07133_, _06286_);
  or (_08390_, _08389_, _08388_);
  and (_08391_, _08390_, _08341_);
  and (_08392_, _07886_, \oc8051_golden_model_1.SBUF [2]);
  not (_08393_, _08392_);
  and (_08394_, _07900_, \oc8051_golden_model_1.IE [2]);
  and (_08395_, _07894_, \oc8051_golden_model_1.P3 [2]);
  nor (_08396_, _08395_, _08394_);
  and (_08397_, _08396_, _08393_);
  and (_08398_, _07904_, \oc8051_golden_model_1.P2 [2]);
  and (_08399_, _07968_, \oc8051_golden_model_1.TL1 [2]);
  nor (_08400_, _08399_, _08398_);
  and (_08401_, _08400_, _08397_);
  and (_08402_, _07928_, \oc8051_golden_model_1.TCON [2]);
  not (_08403_, _08402_);
  and (_08404_, _07922_, \oc8051_golden_model_1.TH0 [2]);
  and (_08405_, _07919_, \oc8051_golden_model_1.TL0 [2]);
  nor (_08406_, _08405_, _08404_);
  and (_08407_, _08406_, _08403_);
  and (_08408_, _07914_, \oc8051_golden_model_1.TMOD [2]);
  and (_08409_, _07926_, \oc8051_golden_model_1.P0 [2]);
  nor (_08410_, _08409_, _08408_);
  and (_08411_, _08410_, _08407_);
  and (_08412_, _08411_, _08401_);
  and (_08413_, _07935_, \oc8051_golden_model_1.PSW [2]);
  not (_08414_, _08413_);
  and (_08415_, _07939_, \oc8051_golden_model_1.ACC [2]);
  and (_08416_, _07942_, \oc8051_golden_model_1.B [2]);
  nor (_08417_, _08416_, _08415_);
  and (_08418_, _08417_, _08414_);
  and (_08419_, _07946_, \oc8051_golden_model_1.IP [2]);
  and (_08420_, _07951_, \oc8051_golden_model_1.PCON [2]);
  nor (_08421_, _08420_, _08419_);
  and (_08422_, _08421_, _08418_);
  and (_08423_, _07956_, \oc8051_golden_model_1.SP [2]);
  not (_08424_, _08423_);
  and (_08425_, _07960_, \oc8051_golden_model_1.DPL [2]);
  and (_08426_, _07963_, \oc8051_golden_model_1.DPH [2]);
  nor (_08427_, _08426_, _08425_);
  and (_08428_, _08427_, _08424_);
  and (_08429_, _07910_, \oc8051_golden_model_1.TH1 [2]);
  not (_08430_, _08429_);
  and (_08431_, _07973_, \oc8051_golden_model_1.SCON [2]);
  and (_08432_, _07971_, \oc8051_golden_model_1.P1 [2]);
  nor (_08433_, _08432_, _08431_);
  and (_08434_, _08433_, _08430_);
  and (_08435_, _08434_, _08428_);
  and (_08436_, _08435_, _08422_);
  and (_08437_, _08436_, _08412_);
  or (_08438_, _07776_, _06182_);
  and (_08439_, _08438_, _08437_);
  not (_08440_, _08439_);
  and (_08441_, _08440_, _08391_);
  and (_08442_, _08441_, _08292_);
  and (_08443_, _07904_, \oc8051_golden_model_1.P2 [4]);
  not (_08444_, _08443_);
  and (_08445_, _07886_, \oc8051_golden_model_1.SBUF [4]);
  not (_08446_, _08445_);
  and (_08447_, _07894_, \oc8051_golden_model_1.P3 [4]);
  and (_08448_, _07900_, \oc8051_golden_model_1.IE [4]);
  nor (_08449_, _08448_, _08447_);
  and (_08450_, _08449_, _08446_);
  and (_08451_, _08450_, _08444_);
  and (_08452_, _07956_, \oc8051_golden_model_1.SP [4]);
  not (_08453_, _08452_);
  and (_08454_, _07960_, \oc8051_golden_model_1.DPL [4]);
  and (_08455_, _07963_, \oc8051_golden_model_1.DPH [4]);
  nor (_08456_, _08455_, _08454_);
  and (_08457_, _08456_, _08453_);
  and (_08458_, _07971_, \oc8051_golden_model_1.P1 [4]);
  and (_08459_, _07973_, \oc8051_golden_model_1.SCON [4]);
  nor (_08460_, _08459_, _08458_);
  and (_08461_, _07910_, \oc8051_golden_model_1.TH1 [4]);
  and (_08462_, _07968_, \oc8051_golden_model_1.TL1 [4]);
  nor (_08463_, _08462_, _08461_);
  and (_08464_, _08463_, _08460_);
  and (_08465_, _08464_, _08457_);
  and (_08466_, _08465_, _08451_);
  and (_08467_, _07935_, \oc8051_golden_model_1.PSW [4]);
  not (_08468_, _08467_);
  and (_08469_, _07939_, \oc8051_golden_model_1.ACC [4]);
  and (_08470_, _07942_, \oc8051_golden_model_1.B [4]);
  nor (_08471_, _08470_, _08469_);
  and (_08472_, _08471_, _08468_);
  and (_08473_, _07946_, \oc8051_golden_model_1.IP [4]);
  and (_08474_, _07951_, \oc8051_golden_model_1.PCON [4]);
  nor (_08475_, _08474_, _08473_);
  and (_08476_, _08475_, _08472_);
  and (_08477_, _07928_, \oc8051_golden_model_1.TCON [4]);
  not (_08478_, _08477_);
  and (_08479_, _07919_, \oc8051_golden_model_1.TL0 [4]);
  and (_08480_, _07922_, \oc8051_golden_model_1.TH0 [4]);
  nor (_08481_, _08480_, _08479_);
  and (_08482_, _08481_, _08478_);
  and (_08483_, _07914_, \oc8051_golden_model_1.TMOD [4]);
  and (_08484_, _07926_, \oc8051_golden_model_1.P0 [4]);
  nor (_08485_, _08484_, _08483_);
  and (_08486_, _08485_, _08482_);
  and (_08487_, _08486_, _08476_);
  and (_08488_, _08487_, _08466_);
  not (_08489_, \oc8051_golden_model_1.IRAM[0] [4]);
  or (_08490_, _06936_, _08489_);
  not (_08491_, \oc8051_golden_model_1.IRAM[1] [4]);
  or (_08492_, _07078_, _08491_);
  and (_08493_, _08492_, _07076_);
  nand (_08494_, _08493_, _08490_);
  not (_08495_, \oc8051_golden_model_1.IRAM[3] [4]);
  or (_08496_, _07078_, _08495_);
  not (_08497_, \oc8051_golden_model_1.IRAM[2] [4]);
  or (_08498_, _06936_, _08497_);
  and (_08499_, _08498_, _07084_);
  nand (_08500_, _08499_, _08496_);
  nand (_08501_, _08500_, _08494_);
  nand (_08502_, _08501_, _06769_);
  not (_08503_, \oc8051_golden_model_1.IRAM[7] [4]);
  or (_08504_, _07078_, _08503_);
  not (_08505_, \oc8051_golden_model_1.IRAM[6] [4]);
  or (_08506_, _06936_, _08505_);
  and (_08507_, _08506_, _07084_);
  nand (_08508_, _08507_, _08504_);
  not (_08509_, \oc8051_golden_model_1.IRAM[4] [4]);
  or (_08510_, _06936_, _08509_);
  not (_08511_, \oc8051_golden_model_1.IRAM[5] [4]);
  or (_08512_, _07078_, _08511_);
  and (_08513_, _08512_, _07076_);
  nand (_08514_, _08513_, _08510_);
  nand (_08515_, _08514_, _08508_);
  nand (_08516_, _08515_, _07091_);
  nand (_08517_, _08516_, _08502_);
  nand (_08518_, _08517_, _06580_);
  nand (_08519_, _06936_, \oc8051_golden_model_1.IRAM[11] [4]);
  nand (_08520_, _07078_, \oc8051_golden_model_1.IRAM[10] [4]);
  and (_08521_, _08520_, _07084_);
  nand (_08522_, _08521_, _08519_);
  nand (_08523_, _07078_, \oc8051_golden_model_1.IRAM[8] [4]);
  nand (_08524_, _06936_, \oc8051_golden_model_1.IRAM[9] [4]);
  and (_08525_, _08524_, _07076_);
  nand (_08526_, _08525_, _08523_);
  nand (_08527_, _08526_, _08522_);
  nand (_08528_, _08527_, _06769_);
  nand (_08529_, _06936_, \oc8051_golden_model_1.IRAM[15] [4]);
  nand (_08530_, _07078_, \oc8051_golden_model_1.IRAM[14] [4]);
  and (_08531_, _08530_, _07084_);
  nand (_08532_, _08531_, _08529_);
  nand (_08533_, _07078_, \oc8051_golden_model_1.IRAM[12] [4]);
  nand (_08534_, _06936_, \oc8051_golden_model_1.IRAM[13] [4]);
  and (_08535_, _08534_, _07076_);
  nand (_08536_, _08535_, _08533_);
  nand (_08537_, _08536_, _08532_);
  nand (_08538_, _08537_, _07091_);
  nand (_08539_, _08538_, _08528_);
  nand (_08540_, _08539_, _07108_);
  nand (_08541_, _08540_, _08518_);
  or (_08542_, _08541_, _06182_);
  and (_08543_, _08542_, _08488_);
  not (_08544_, _08543_);
  and (_08545_, _08544_, _08442_);
  and (_08546_, _08545_, _08247_);
  and (_08547_, _08546_, _08145_);
  or (_08548_, _08547_, _08043_);
  nand (_08549_, _08547_, _08043_);
  and (_08550_, _08549_, _08548_);
  and (_08551_, _08550_, _07286_);
  not (_08552_, _08040_);
  and (_08553_, _08541_, _08244_);
  and (_08554_, _07776_, _07594_);
  not (_08555_, _07133_);
  and (_08556_, _07357_, _08555_);
  and (_08557_, _08556_, _08554_);
  and (_08558_, _08557_, _08553_);
  and (_08559_, _08558_, _08142_);
  or (_08560_, _08559_, _08552_);
  nand (_08561_, _08559_, _08552_);
  and (_08562_, _08561_, _08560_);
  and (_08563_, _06337_, _05779_);
  and (_08564_, _06350_, _05779_);
  nor (_08565_, _08564_, _08563_);
  nor (_08566_, _07211_, _06567_);
  nor (_08567_, _07212_, _06567_);
  nor (_08568_, _08567_, _08566_);
  and (_08569_, _08568_, _08565_);
  or (_08570_, _08569_, _08562_);
  not (_08571_, _07243_);
  not (_08572_, \oc8051_golden_model_1.ACC [7]);
  and (_08573_, _08042_, _08572_);
  nor (_08574_, _08042_, _08572_);
  nor (_08575_, _08574_, _08573_);
  and (_08576_, _08575_, _07241_);
  not (_08577_, _07241_);
  and (_08578_, _06420_, _04431_);
  and (_08579_, _06445_, _04415_);
  nor (_08580_, _08579_, _08578_);
  and (_08581_, _06434_, _04434_);
  and (_08582_, _06436_, _04419_);
  nor (_08583_, _08582_, _08581_);
  and (_08584_, _08583_, _08580_);
  and (_08585_, _06417_, _04355_);
  and (_08586_, _06415_, _04439_);
  nor (_08587_, _08586_, _08585_);
  and (_08588_, _06411_, _04387_);
  and (_08589_, _06431_, _04392_);
  nor (_08590_, _08589_, _08588_);
  and (_08591_, _08590_, _08587_);
  and (_08592_, _08591_, _08584_);
  and (_08593_, _06447_, _04397_);
  and (_08594_, _06429_, _04406_);
  nor (_08595_, _08594_, _08593_);
  and (_08596_, _06440_, _04401_);
  and (_08597_, _06401_, _04381_);
  nor (_08598_, _08597_, _08596_);
  and (_08599_, _08598_, _08595_);
  and (_08600_, _06407_, _04423_);
  and (_08601_, _06398_, _04442_);
  nor (_08602_, _08601_, _08600_);
  and (_08603_, _06423_, _04411_);
  and (_08604_, _06442_, _04426_);
  nor (_08605_, _08604_, _08603_);
  and (_08606_, _08605_, _08602_);
  and (_08607_, _08606_, _08599_);
  and (_08608_, _08607_, _08592_);
  nand (_08609_, _08608_, _06220_);
  not (_08610_, _07179_);
  and (_08611_, _07948_, \oc8051_golden_model_1.P0 [7]);
  not (_08612_, _06214_);
  nor (_08613_, _06969_, _08612_);
  and (_08614_, _06613_, _06320_);
  and (_08615_, _08614_, _08613_);
  and (_08616_, _08615_, _07907_);
  and (_08617_, _08616_, \oc8051_golden_model_1.TCON [7]);
  nor (_08618_, _06612_, _06320_);
  and (_08619_, _08618_, _08613_);
  and (_08620_, _08619_, _07885_);
  and (_08621_, _08620_, \oc8051_golden_model_1.P1 [7]);
  and (_08622_, _08615_, _07885_);
  and (_08623_, _08622_, \oc8051_golden_model_1.SCON [7]);
  and (_08624_, _08619_, _07898_);
  and (_08625_, _08624_, \oc8051_golden_model_1.P2 [7]);
  and (_08626_, _08615_, _07898_);
  and (_08627_, _08626_, \oc8051_golden_model_1.IE [7]);
  and (_08628_, _08619_, _07893_);
  and (_08629_, _08628_, \oc8051_golden_model_1.P3 [7]);
  and (_08630_, _08619_, _07934_);
  and (_08631_, _08630_, \oc8051_golden_model_1.PSW [7]);
  and (_08632_, _08615_, _07893_);
  and (_08633_, _08632_, \oc8051_golden_model_1.IP [7]);
  and (_08634_, _07941_, _08619_);
  and (_08635_, _08634_, \oc8051_golden_model_1.B [7]);
  and (_08636_, _08619_, _07938_);
  and (_08637_, _08636_, \oc8051_golden_model_1.ACC [7]);
  or (_08638_, _08637_, _08635_);
  or (_08639_, _08638_, _08633_);
  or (_08640_, _08639_, _08631_);
  or (_08641_, _08640_, _08629_);
  or (_08642_, _08641_, _08627_);
  or (_08643_, _08642_, _08625_);
  or (_08644_, _08643_, _08623_);
  or (_08645_, _08644_, _08621_);
  or (_08646_, _08645_, _08617_);
  nor (_08647_, _08646_, _08611_);
  and (_08648_, _08647_, _08041_);
  nor (_08649_, _08648_, _07950_);
  or (_08650_, _08649_, _08610_);
  not (_08651_, _06275_);
  not (_08652_, _07152_);
  nor (_08653_, _07213_, _06009_);
  nor (_08654_, _08653_, _07364_);
  or (_08655_, _08654_, _08562_);
  and (_08656_, \oc8051_golden_model_1.PC [5], \oc8051_golden_model_1.PC [4]);
  and (_08657_, _08656_, \oc8051_golden_model_1.PC [6]);
  and (_08658_, _08657_, _05929_);
  and (_08659_, _08658_, \oc8051_golden_model_1.PC [7]);
  nor (_08660_, _08658_, \oc8051_golden_model_1.PC [7]);
  nor (_08661_, _08660_, _08659_);
  and (_08662_, _08661_, _06758_);
  nor (_08663_, _06758_, _08572_);
  nor (_08664_, _08663_, _08662_);
  nand (_08665_, _08664_, _08654_);
  and (_08666_, _08665_, _08655_);
  or (_08667_, _08666_, _07154_);
  nor (_08668_, \oc8051_golden_model_1.SP [1], \oc8051_golden_model_1.SP [0]);
  and (_08669_, _08668_, _06715_);
  nor (_08670_, _08669_, _06460_);
  nor (_08671_, \oc8051_golden_model_1.SP [2], \oc8051_golden_model_1.SP [1]);
  and (_08672_, _08671_, _06460_);
  and (_08673_, _08672_, _06800_);
  nor (_08674_, _08673_, _08670_);
  nor (_08675_, _06551_, _06281_);
  nor (_08676_, _08675_, _08674_);
  and (_08677_, _07594_, _07198_);
  and (_08678_, _07197_, _06213_);
  not (_08679_, _08678_);
  nand (_08680_, _08679_, _08675_);
  nor (_08681_, _08680_, _08677_);
  nor (_08682_, _08681_, _08676_);
  nor (_08683_, _08668_, _06715_);
  nor (_08684_, _08683_, _08669_);
  nor (_08685_, _08684_, _08675_);
  not (_08686_, _08685_);
  nand (_08687_, _07776_, _07198_);
  and (_08688_, _07197_, _06656_);
  not (_08689_, _08688_);
  and (_08690_, _08689_, _08675_);
  nand (_08691_, _08690_, _08687_);
  and (_08692_, _08691_, _08686_);
  or (_08693_, _07197_, _07133_);
  and (_08694_, _07197_, _06251_);
  not (_08695_, _08694_);
  and (_08696_, _08695_, _08675_);
  nand (_08697_, _08696_, _08693_);
  nor (_08698_, _08675_, \oc8051_golden_model_1.SP [0]);
  not (_08699_, _08698_);
  and (_08700_, _08699_, _08697_);
  nand (_08701_, _08700_, \oc8051_golden_model_1.IRAM[0] [7]);
  nor (_08702_, _08675_, _07297_);
  not (_08703_, _08702_);
  or (_08704_, _07357_, _07197_);
  or (_08705_, _07198_, _07004_);
  and (_08706_, _08705_, _08675_);
  nand (_08707_, _08706_, _08704_);
  and (_08708_, _08707_, _08703_);
  not (_08709_, _08708_);
  or (_08710_, _08700_, _07982_);
  and (_08711_, _08710_, _08709_);
  nand (_08712_, _08711_, _08701_);
  nand (_08713_, _08700_, \oc8051_golden_model_1.IRAM[2] [7]);
  or (_08714_, _08700_, _07986_);
  and (_08715_, _08714_, _08708_);
  nand (_08716_, _08715_, _08713_);
  nand (_08717_, _08716_, _08712_);
  nand (_08718_, _08717_, _08692_);
  not (_08719_, _08692_);
  nand (_08720_, _08700_, \oc8051_golden_model_1.IRAM[4] [7]);
  or (_08721_, _08700_, _08002_);
  and (_08722_, _08721_, _08709_);
  nand (_08723_, _08722_, _08720_);
  nand (_08724_, _08700_, \oc8051_golden_model_1.IRAM[6] [7]);
  or (_08725_, _08700_, _07994_);
  and (_08726_, _08725_, _08708_);
  nand (_08727_, _08726_, _08724_);
  nand (_08728_, _08727_, _08723_);
  nand (_08729_, _08728_, _08719_);
  nand (_08730_, _08729_, _08718_);
  nand (_08731_, _08730_, _08682_);
  not (_08732_, _08682_);
  nand (_08733_, _08700_, \oc8051_golden_model_1.IRAM[10] [7]);
  or (_08734_, _08700_, _08010_);
  and (_08735_, _08734_, _08708_);
  nand (_08736_, _08735_, _08733_);
  nand (_08737_, _08700_, \oc8051_golden_model_1.IRAM[8] [7]);
  or (_08738_, _08700_, _08018_);
  and (_08739_, _08738_, _08709_);
  nand (_08740_, _08739_, _08737_);
  nand (_08741_, _08740_, _08736_);
  nand (_08742_, _08741_, _08692_);
  nand (_08743_, _08700_, \oc8051_golden_model_1.IRAM[12] [7]);
  or (_08744_, _08700_, _08032_);
  and (_08745_, _08744_, _08709_);
  nand (_08746_, _08745_, _08743_);
  nand (_08747_, _08700_, \oc8051_golden_model_1.IRAM[14] [7]);
  or (_08748_, _08700_, _08024_);
  and (_08749_, _08748_, _08708_);
  nand (_08750_, _08749_, _08747_);
  nand (_08751_, _08750_, _08746_);
  nand (_08752_, _08751_, _08719_);
  nand (_08753_, _08752_, _08742_);
  nand (_08754_, _08753_, _08732_);
  and (_08755_, _08754_, _08731_);
  or (_08756_, _08755_, _07155_);
  and (_08757_, _08756_, _08667_);
  and (_08758_, _08757_, _08652_);
  and (_08759_, _08543_, _08246_);
  not (_08760_, _08390_);
  and (_08761_, _08760_, _08340_);
  and (_08762_, _08439_, _08291_);
  and (_08763_, _08762_, _08761_);
  and (_08764_, _08763_, _08759_);
  and (_08765_, _08764_, _08144_);
  or (_08766_, _08765_, _08043_);
  nand (_08767_, _08765_, _08043_);
  and (_08768_, _08767_, _08766_);
  and (_08769_, _08768_, _07152_);
  or (_08770_, _08769_, _08758_);
  and (_08771_, _08770_, _08651_);
  not (_08772_, _07950_);
  nand (_08773_, _08648_, _08772_);
  and (_08774_, _08773_, _06275_);
  or (_08775_, _08774_, _07611_);
  or (_08776_, _08775_, _08771_);
  nor (_08777_, _08661_, _06010_);
  nor (_08778_, _08777_, _07167_);
  and (_08779_, _08778_, _08776_);
  and (_08780_, _08552_, _07167_);
  or (_08781_, _08780_, _07179_);
  or (_08782_, _08781_, _08779_);
  and (_08783_, _08782_, _08650_);
  or (_08784_, _08783_, _06267_);
  nand (_08785_, _08042_, _06267_);
  and (_08786_, _08785_, _06265_);
  and (_08787_, _08786_, _08784_);
  nor (_08788_, _08648_, _08772_);
  not (_08789_, _08788_);
  and (_08790_, _08789_, _08773_);
  and (_08791_, _08790_, _06264_);
  or (_08792_, _08791_, _08787_);
  and (_08793_, _08792_, _06007_);
  not (_08794_, _08661_);
  or (_08795_, _08794_, _06007_);
  nand (_08796_, _08795_, _06501_);
  or (_08797_, _08796_, _08793_);
  nand (_08798_, _08042_, _06502_);
  and (_08799_, _08798_, _08797_);
  or (_08800_, _08799_, _07197_);
  not (_08801_, _07196_);
  and (_08802_, _08755_, _06286_);
  nand (_08803_, _07979_, _07197_);
  or (_08804_, _08803_, _08802_);
  and (_08805_, _08804_, _08801_);
  and (_08806_, _08805_, _08800_);
  and (_08807_, _07950_, \oc8051_golden_model_1.PSW [7]);
  or (_08808_, _08807_, _08649_);
  and (_08809_, _08808_, _07196_);
  or (_08810_, _08809_, _06254_);
  or (_08811_, _08810_, _08806_);
  nor (_08812_, _07215_, _06182_);
  nor (_08813_, _08661_, _05978_);
  nor (_08814_, _08813_, _08812_);
  and (_08815_, _08814_, _08811_);
  nor (_08816_, _07208_, _06182_);
  not (_08817_, _08812_);
  nor (_08818_, _08040_, _08817_);
  or (_08819_, _08818_, _08816_);
  or (_08820_, _08819_, _08815_);
  not (_08821_, _08816_);
  or (_08822_, _08755_, _08821_);
  and (_08823_, _08822_, _07471_);
  and (_08824_, _08823_, _08820_);
  not (_08825_, _08608_);
  nor (_08826_, _08825_, _08040_);
  and (_08827_, _06423_, _04849_);
  and (_08828_, _06445_, _04839_);
  nor (_08829_, _08828_, _08827_);
  and (_08830_, _06447_, _04851_);
  and (_08831_, _06436_, _04823_);
  nor (_08832_, _08831_, _08830_);
  and (_08833_, _08832_, _08829_);
  and (_08834_, _06411_, _04835_);
  and (_08835_, _06431_, _04831_);
  nor (_08836_, _08835_, _08834_);
  and (_08837_, _06415_, _04855_);
  and (_08838_, _06442_, _04816_);
  nor (_08839_, _08838_, _08837_);
  and (_08840_, _08839_, _08836_);
  and (_08841_, _08840_, _08833_);
  and (_08842_, _06434_, _04844_);
  and (_08843_, _06429_, _04827_);
  nor (_08844_, _08843_, _08842_);
  and (_08845_, _06440_, _04837_);
  and (_08846_, _06401_, _04818_);
  nor (_08847_, _08846_, _08845_);
  and (_08848_, _08847_, _08844_);
  and (_08849_, _06407_, _04842_);
  and (_08850_, _06398_, _04857_);
  nor (_08851_, _08850_, _08849_);
  and (_08852_, _06420_, _04829_);
  and (_08853_, _06417_, _04821_);
  nor (_08854_, _08853_, _08852_);
  and (_08855_, _08854_, _08851_);
  and (_08856_, _08855_, _08848_);
  and (_08857_, _08856_, _08841_);
  and (_08858_, _08857_, _08825_);
  and (_08859_, _06407_, _04750_);
  and (_08860_, _06442_, _04724_);
  nor (_08861_, _08860_, _08859_);
  and (_08862_, _06411_, _04743_);
  and (_08863_, _06431_, _04739_);
  nor (_08864_, _08863_, _08862_);
  and (_08865_, _08864_, _08861_);
  and (_08866_, _06445_, _04747_);
  and (_08868_, _06429_, _04735_);
  nor (_08869_, _08868_, _08866_);
  and (_08870_, _06440_, _04745_);
  and (_08871_, _06423_, _04757_);
  nor (_08872_, _08871_, _08870_);
  and (_08873_, _08872_, _08869_);
  and (_08874_, _08873_, _08865_);
  and (_08875_, _06447_, _04759_);
  and (_08876_, _06398_, _04765_);
  nor (_08877_, _08876_, _08875_);
  and (_08879_, _06436_, _04731_);
  and (_08880_, _06401_, _04726_);
  nor (_08881_, _08880_, _08879_);
  and (_08882_, _08881_, _08877_);
  and (_08883_, _06417_, _04729_);
  and (_08884_, _06415_, _04763_);
  nor (_08885_, _08884_, _08883_);
  and (_08886_, _06420_, _04737_);
  and (_08887_, _06434_, _04752_);
  nor (_08888_, _08887_, _08886_);
  and (_08890_, _08888_, _08885_);
  and (_08891_, _08890_, _08882_);
  and (_08892_, _08891_, _08874_);
  and (_08893_, _06445_, _04793_);
  and (_08894_, _06401_, _04772_);
  nor (_08895_, _08894_, _08893_);
  and (_08896_, _06440_, _04791_);
  and (_08897_, _06431_, _04781_);
  nor (_08898_, _08897_, _08896_);
  and (_08899_, _08898_, _08895_);
  and (_08901_, _06420_, _04783_);
  and (_08902_, _06423_, _04785_);
  nor (_08903_, _08902_, _08901_);
  and (_08904_, _06434_, _04798_);
  and (_08905_, _06429_, _04805_);
  nor (_08906_, _08905_, _08904_);
  and (_08907_, _08906_, _08903_);
  and (_08908_, _08907_, _08899_);
  and (_08909_, _06415_, _04809_);
  and (_08910_, _06442_, _04770_);
  nor (_08912_, _08910_, _08909_);
  and (_08913_, _06436_, _04777_);
  and (_08914_, _06398_, _04811_);
  nor (_08915_, _08914_, _08913_);
  and (_08916_, _08915_, _08912_);
  and (_08917_, _06407_, _04796_);
  and (_08918_, _06447_, _04803_);
  nor (_08919_, _08918_, _08917_);
  and (_08920_, _06411_, _04789_);
  and (_08921_, _06417_, _04775_);
  nor (_08923_, _08921_, _08920_);
  and (_08924_, _08923_, _08919_);
  and (_08925_, _08924_, _08916_);
  and (_08926_, _08925_, _08908_);
  and (_08927_, _08926_, _08892_);
  and (_08928_, _08927_, _08858_);
  and (_08929_, _07038_, _06872_);
  not (_08930_, _06452_);
  and (_08931_, _06697_, _08930_);
  and (_08932_, _08931_, _08929_);
  and (_08934_, _08932_, _08928_);
  and (_08935_, _08934_, \oc8051_golden_model_1.TCON [7]);
  not (_08936_, _07038_);
  and (_08937_, _08936_, _06872_);
  and (_08938_, _08937_, _08931_);
  and (_08939_, _08938_, _08928_);
  and (_08940_, _08939_, \oc8051_golden_model_1.TL0 [7]);
  or (_08941_, _08940_, _08935_);
  and (_08942_, _06697_, _06452_);
  and (_08943_, _08942_, _08929_);
  and (_08944_, _08943_, _08928_);
  and (_08945_, _08944_, \oc8051_golden_model_1.P0 [7]);
  not (_08946_, _08926_);
  and (_08947_, _08946_, _08892_);
  nor (_08948_, _08857_, _08608_);
  and (_08949_, _08948_, _08943_);
  and (_08950_, _08949_, _08947_);
  and (_08951_, _08950_, \oc8051_golden_model_1.ACC [7]);
  or (_08952_, _08951_, _08945_);
  or (_08953_, _08952_, _08941_);
  not (_08954_, _06872_);
  and (_08955_, _07038_, _08954_);
  and (_08956_, _08955_, _08931_);
  and (_08957_, _08956_, _08928_);
  and (_08958_, _08957_, \oc8051_golden_model_1.TMOD [7]);
  not (_08959_, _08892_);
  and (_08960_, _08926_, _08959_);
  and (_08961_, _08960_, _08858_);
  and (_08962_, _08961_, _08943_);
  and (_08963_, _08962_, \oc8051_golden_model_1.P1 [7]);
  or (_08964_, _08963_, _08958_);
  and (_08965_, _08961_, _08932_);
  and (_08966_, _08965_, \oc8051_golden_model_1.SCON [7]);
  nor (_08967_, _08926_, _08892_);
  and (_08968_, _08967_, _08949_);
  and (_08969_, _08968_, \oc8051_golden_model_1.B [7]);
  or (_08970_, _08969_, _08966_);
  or (_08971_, _08970_, _08964_);
  or (_08972_, _08971_, _08953_);
  not (_08973_, _06697_);
  nor (_08974_, _07038_, _06872_);
  and (_08975_, _08974_, _08928_);
  and (_08976_, _08975_, _06452_);
  and (_08977_, _08976_, _08973_);
  and (_08978_, _08977_, \oc8051_golden_model_1.PCON [7]);
  and (_08979_, _08976_, _06697_);
  and (_08980_, _08979_, \oc8051_golden_model_1.DPH [7]);
  or (_08981_, _08980_, _08978_);
  or (_08982_, _08981_, _08972_);
  and (_08983_, _08942_, _08928_);
  and (_08984_, _08983_, _08937_);
  and (_08985_, _08984_, \oc8051_golden_model_1.DPL [7]);
  and (_08986_, _08975_, _08931_);
  and (_08987_, _08986_, \oc8051_golden_model_1.TL1 [7]);
  and (_08988_, _08955_, _08983_);
  and (_08989_, _08988_, \oc8051_golden_model_1.SP [7]);
  or (_08990_, _08989_, _08987_);
  or (_08991_, _08990_, _08985_);
  and (_08992_, _08947_, _08858_);
  and (_08993_, _08992_, _08932_);
  and (_08994_, _08993_, \oc8051_golden_model_1.IE [7]);
  and (_08995_, _08967_, _08858_);
  and (_08996_, _08995_, _08932_);
  and (_08997_, _08996_, \oc8051_golden_model_1.IP [7]);
  or (_08998_, _08997_, _08994_);
  and (_08999_, _08992_, _08943_);
  and (_09000_, _08999_, \oc8051_golden_model_1.P2 [7]);
  and (_09001_, _08995_, _08943_);
  and (_09002_, _09001_, \oc8051_golden_model_1.P3 [7]);
  or (_09003_, _09002_, _09000_);
  or (_09004_, _09003_, _08998_);
  and (_09005_, _08961_, _08956_);
  and (_09006_, _09005_, \oc8051_golden_model_1.SBUF [7]);
  and (_09007_, _08960_, _08949_);
  and (_09008_, _09007_, \oc8051_golden_model_1.PSW [7]);
  or (_09009_, _09008_, _09006_);
  or (_09010_, _09009_, _09004_);
  nor (_09011_, _06697_, _06452_);
  and (_09012_, _09011_, _08928_);
  and (_09013_, _09012_, _08929_);
  and (_09014_, _09013_, \oc8051_golden_model_1.TH0 [7]);
  and (_09015_, _09012_, _08955_);
  and (_09016_, _09015_, \oc8051_golden_model_1.TH1 [7]);
  or (_09017_, _09016_, _09014_);
  or (_09018_, _09017_, _09010_);
  or (_09019_, _09018_, _08991_);
  or (_09020_, _09019_, _08982_);
  or (_09021_, _09020_, _08826_);
  and (_09022_, _09021_, _07470_);
  nor (_09023_, _07211_, _05951_);
  not (_09024_, _09023_);
  nor (_09025_, _07212_, _05951_);
  not (_09026_, _09025_);
  and (_09027_, _07209_, _06321_);
  nor (_09028_, _09027_, _07224_);
  and (_09029_, _09028_, _09026_);
  and (_09030_, _09029_, _09024_);
  not (_09031_, _09030_);
  or (_09032_, _09031_, _09022_);
  or (_09033_, _09032_, _08824_);
  or (_09034_, _09030_, _06182_);
  and (_09035_, _09034_, _09033_);
  or (_09036_, _09035_, _06220_);
  and (_09037_, _09036_, _08609_);
  or (_09038_, _09037_, _06217_);
  nor (_09039_, _08661_, _05952_);
  nor (_09040_, _09039_, _07238_);
  and (_09041_, _09040_, _09038_);
  nor (_09042_, _08608_, _08042_);
  and (_09043_, _08608_, _08042_);
  nor (_09044_, _09043_, _09042_);
  and (_09045_, _09044_, _07238_);
  or (_09046_, _09045_, _09041_);
  and (_09047_, _09046_, _08577_);
  or (_09048_, _09047_, _08576_);
  and (_09049_, _09048_, _08571_);
  and (_09050_, _09042_, _07243_);
  or (_09051_, _09050_, _09049_);
  and (_09052_, _09051_, _07236_);
  and (_09053_, _08574_, _07235_);
  or (_09054_, _09053_, _07233_);
  or (_09055_, _09054_, _09052_);
  not (_09056_, _06366_);
  nor (_09057_, _09056_, _06182_);
  nor (_09058_, _08661_, _05961_);
  nor (_09059_, _09058_, _09057_);
  and (_09060_, _09059_, _09055_);
  not (_09061_, _06528_);
  nor (_09062_, _09061_, _06182_);
  not (_09063_, _09043_);
  and (_09064_, _09063_, _09057_);
  or (_09065_, _09064_, _09062_);
  or (_09066_, _09065_, _09060_);
  nand (_09067_, _08573_, _09062_);
  and (_09068_, _09067_, _05959_);
  and (_09069_, _09068_, _09066_);
  or (_09070_, _08794_, _05959_);
  nand (_09071_, _09070_, _08569_);
  or (_09072_, _09071_, _09069_);
  and (_09073_, _09072_, _08570_);
  or (_09074_, _09073_, _07435_);
  not (_09075_, _07261_);
  not (_09076_, _08755_);
  nand (_09077_, _08700_, \oc8051_golden_model_1.IRAM[0] [6]);
  or (_09078_, _08700_, _08092_);
  and (_09079_, _09078_, _08709_);
  nand (_09080_, _09079_, _09077_);
  nand (_09081_, _08700_, \oc8051_golden_model_1.IRAM[2] [6]);
  or (_09082_, _08700_, _08096_);
  and (_09083_, _09082_, _08708_);
  nand (_09084_, _09083_, _09081_);
  nand (_09085_, _09084_, _09080_);
  nand (_09086_, _09085_, _08692_);
  nand (_09087_, _08700_, \oc8051_golden_model_1.IRAM[4] [6]);
  or (_09088_, _08700_, _08112_);
  and (_09089_, _09088_, _08709_);
  nand (_09090_, _09089_, _09087_);
  nand (_09091_, _08700_, \oc8051_golden_model_1.IRAM[6] [6]);
  or (_09092_, _08700_, _08104_);
  and (_09093_, _09092_, _08708_);
  nand (_09094_, _09093_, _09091_);
  nand (_09095_, _09094_, _09090_);
  nand (_09096_, _09095_, _08719_);
  and (_09097_, _09096_, _08682_);
  and (_09098_, _09097_, _09086_);
  not (_09099_, _08700_);
  or (_09100_, _09099_, \oc8051_golden_model_1.IRAM[10] [6]);
  or (_09101_, _08700_, \oc8051_golden_model_1.IRAM[11] [6]);
  nand (_09102_, _09101_, _09100_);
  nand (_09103_, _09102_, _08708_);
  or (_09104_, _09099_, \oc8051_golden_model_1.IRAM[8] [6]);
  or (_09105_, _08700_, \oc8051_golden_model_1.IRAM[9] [6]);
  nand (_09106_, _09105_, _09104_);
  nand (_09107_, _09106_, _08709_);
  nand (_09108_, _09107_, _09103_);
  nand (_09109_, _09108_, _08692_);
  or (_09110_, _09099_, \oc8051_golden_model_1.IRAM[14] [6]);
  or (_09111_, _08700_, \oc8051_golden_model_1.IRAM[15] [6]);
  nand (_09112_, _09111_, _09110_);
  nand (_09113_, _09112_, _08708_);
  or (_09114_, _09099_, \oc8051_golden_model_1.IRAM[12] [6]);
  or (_09115_, _08700_, \oc8051_golden_model_1.IRAM[13] [6]);
  nand (_09116_, _09115_, _09114_);
  nand (_09117_, _09116_, _08709_);
  nand (_09118_, _09117_, _09113_);
  nand (_09119_, _09118_, _08719_);
  and (_09120_, _09119_, _08732_);
  and (_09121_, _09120_, _09109_);
  nor (_09122_, _09121_, _09098_);
  nand (_09123_, _08700_, \oc8051_golden_model_1.IRAM[0] [5]);
  or (_09124_, _08700_, _08194_);
  and (_09125_, _09124_, _08709_);
  nand (_09126_, _09125_, _09123_);
  nand (_09127_, _08700_, \oc8051_golden_model_1.IRAM[2] [5]);
  or (_09128_, _08700_, _08198_);
  and (_09129_, _09128_, _08708_);
  nand (_09130_, _09129_, _09127_);
  nand (_09131_, _09130_, _09126_);
  nand (_09132_, _09131_, _08692_);
  nand (_09133_, _08700_, \oc8051_golden_model_1.IRAM[4] [5]);
  or (_09134_, _08700_, _08214_);
  and (_09135_, _09134_, _08709_);
  nand (_09136_, _09135_, _09133_);
  nand (_09137_, _08700_, \oc8051_golden_model_1.IRAM[6] [5]);
  or (_09138_, _08700_, _08206_);
  and (_09139_, _09138_, _08708_);
  nand (_09140_, _09139_, _09137_);
  nand (_09141_, _09140_, _09136_);
  nand (_09142_, _09141_, _08719_);
  and (_09143_, _09142_, _08682_);
  and (_09144_, _09143_, _09132_);
  or (_09145_, _09099_, \oc8051_golden_model_1.IRAM[10] [5]);
  or (_09146_, _08700_, \oc8051_golden_model_1.IRAM[11] [5]);
  nand (_09147_, _09146_, _09145_);
  nand (_09148_, _09147_, _08708_);
  or (_09149_, _09099_, \oc8051_golden_model_1.IRAM[8] [5]);
  or (_09150_, _08700_, \oc8051_golden_model_1.IRAM[9] [5]);
  nand (_09151_, _09150_, _09149_);
  nand (_09152_, _09151_, _08709_);
  nand (_09153_, _09152_, _09148_);
  nand (_09154_, _09153_, _08692_);
  or (_09155_, _09099_, \oc8051_golden_model_1.IRAM[14] [5]);
  or (_09156_, _08700_, \oc8051_golden_model_1.IRAM[15] [5]);
  nand (_09157_, _09156_, _09155_);
  nand (_09158_, _09157_, _08708_);
  or (_09159_, _09099_, \oc8051_golden_model_1.IRAM[12] [5]);
  or (_09160_, _08700_, \oc8051_golden_model_1.IRAM[13] [5]);
  nand (_09161_, _09160_, _09159_);
  nand (_09162_, _09161_, _08709_);
  nand (_09163_, _09162_, _09158_);
  nand (_09164_, _09163_, _08719_);
  and (_09165_, _09164_, _08732_);
  and (_09166_, _09165_, _09154_);
  nor (_09167_, _09166_, _09144_);
  nand (_09168_, _08700_, \oc8051_golden_model_1.IRAM[0] [4]);
  or (_09169_, _08700_, _08491_);
  and (_09170_, _09169_, _08709_);
  nand (_09171_, _09170_, _09168_);
  nand (_09172_, _08700_, \oc8051_golden_model_1.IRAM[2] [4]);
  or (_09173_, _08700_, _08495_);
  and (_09174_, _09173_, _08708_);
  nand (_09175_, _09174_, _09172_);
  nand (_09176_, _09175_, _09171_);
  nand (_09177_, _09176_, _08692_);
  nand (_09178_, _08700_, \oc8051_golden_model_1.IRAM[4] [4]);
  or (_09179_, _08700_, _08511_);
  and (_09180_, _09179_, _08709_);
  nand (_09181_, _09180_, _09178_);
  nand (_09182_, _08700_, \oc8051_golden_model_1.IRAM[6] [4]);
  or (_09183_, _08700_, _08503_);
  and (_09184_, _09183_, _08708_);
  nand (_09185_, _09184_, _09182_);
  nand (_09186_, _09185_, _09181_);
  nand (_09187_, _09186_, _08719_);
  and (_09188_, _09187_, _08682_);
  and (_09189_, _09188_, _09177_);
  or (_09190_, _09099_, \oc8051_golden_model_1.IRAM[10] [4]);
  or (_09191_, _08700_, \oc8051_golden_model_1.IRAM[11] [4]);
  nand (_09192_, _09191_, _09190_);
  nand (_09193_, _09192_, _08708_);
  or (_09194_, _09099_, \oc8051_golden_model_1.IRAM[8] [4]);
  or (_09195_, _08700_, \oc8051_golden_model_1.IRAM[9] [4]);
  nand (_09196_, _09195_, _09194_);
  nand (_09197_, _09196_, _08709_);
  nand (_09198_, _09197_, _09193_);
  nand (_09199_, _09198_, _08692_);
  or (_09200_, _09099_, \oc8051_golden_model_1.IRAM[14] [4]);
  or (_09201_, _08700_, \oc8051_golden_model_1.IRAM[15] [4]);
  nand (_09202_, _09201_, _09200_);
  nand (_09203_, _09202_, _08708_);
  or (_09204_, _09099_, \oc8051_golden_model_1.IRAM[12] [4]);
  or (_09205_, _08700_, \oc8051_golden_model_1.IRAM[13] [4]);
  nand (_09206_, _09205_, _09204_);
  nand (_09207_, _09206_, _08709_);
  nand (_09208_, _09207_, _09203_);
  nand (_09209_, _09208_, _08719_);
  and (_09210_, _09209_, _08732_);
  and (_09211_, _09210_, _09199_);
  nor (_09212_, _09211_, _09189_);
  nand (_09213_, _08700_, \oc8051_golden_model_1.IRAM[0] [3]);
  or (_09214_, _08700_, _07544_);
  and (_09215_, _09214_, _08709_);
  nand (_09216_, _09215_, _09213_);
  nand (_09217_, _08700_, \oc8051_golden_model_1.IRAM[2] [3]);
  or (_09218_, _08700_, _07548_);
  and (_09219_, _09218_, _08708_);
  nand (_09220_, _09219_, _09217_);
  nand (_09221_, _09220_, _09216_);
  nand (_09222_, _09221_, _08692_);
  nand (_09223_, _08700_, \oc8051_golden_model_1.IRAM[4] [3]);
  or (_09224_, _08700_, _07564_);
  and (_09225_, _09224_, _08709_);
  nand (_09226_, _09225_, _09223_);
  nand (_09227_, _08700_, \oc8051_golden_model_1.IRAM[6] [3]);
  or (_09228_, _08700_, _07556_);
  and (_09229_, _09228_, _08708_);
  nand (_09230_, _09229_, _09227_);
  nand (_09231_, _09230_, _09226_);
  nand (_09232_, _09231_, _08719_);
  and (_09233_, _09232_, _08682_);
  and (_09234_, _09233_, _09222_);
  or (_09235_, _09099_, \oc8051_golden_model_1.IRAM[10] [3]);
  or (_09236_, _08700_, \oc8051_golden_model_1.IRAM[11] [3]);
  nand (_09237_, _09236_, _09235_);
  nand (_09238_, _09237_, _08708_);
  or (_09239_, _09099_, \oc8051_golden_model_1.IRAM[8] [3]);
  or (_09240_, _08700_, \oc8051_golden_model_1.IRAM[9] [3]);
  nand (_09241_, _09240_, _09239_);
  nand (_09242_, _09241_, _08709_);
  nand (_09243_, _09242_, _09238_);
  nand (_09244_, _09243_, _08692_);
  or (_09245_, _09099_, \oc8051_golden_model_1.IRAM[14] [3]);
  or (_09246_, _08700_, \oc8051_golden_model_1.IRAM[15] [3]);
  nand (_09247_, _09246_, _09245_);
  nand (_09248_, _09247_, _08708_);
  or (_09249_, _09099_, \oc8051_golden_model_1.IRAM[12] [3]);
  or (_09250_, _08700_, \oc8051_golden_model_1.IRAM[13] [3]);
  nand (_09251_, _09250_, _09249_);
  nand (_09252_, _09251_, _08709_);
  nand (_09253_, _09252_, _09248_);
  nand (_09254_, _09253_, _08719_);
  and (_09255_, _09254_, _08732_);
  and (_09256_, _09255_, _09244_);
  nor (_09257_, _09256_, _09234_);
  nand (_09258_, _08700_, \oc8051_golden_model_1.IRAM[0] [2]);
  or (_09259_, _08700_, _07724_);
  and (_09260_, _09259_, _08709_);
  nand (_09261_, _09260_, _09258_);
  nand (_09262_, _08700_, \oc8051_golden_model_1.IRAM[2] [2]);
  or (_09263_, _08700_, _07728_);
  and (_09264_, _09263_, _08708_);
  nand (_09265_, _09264_, _09262_);
  nand (_09266_, _09265_, _09261_);
  nand (_09267_, _09266_, _08692_);
  nand (_09268_, _08700_, \oc8051_golden_model_1.IRAM[4] [2]);
  or (_09269_, _08700_, _07744_);
  and (_09270_, _09269_, _08709_);
  nand (_09271_, _09270_, _09268_);
  nand (_09272_, _08700_, \oc8051_golden_model_1.IRAM[6] [2]);
  or (_09273_, _08700_, _07736_);
  and (_09274_, _09273_, _08708_);
  nand (_09275_, _09274_, _09272_);
  nand (_09276_, _09275_, _09271_);
  nand (_09277_, _09276_, _08719_);
  and (_09278_, _09277_, _08682_);
  and (_09279_, _09278_, _09267_);
  or (_09280_, _09099_, \oc8051_golden_model_1.IRAM[10] [2]);
  or (_09281_, _08700_, \oc8051_golden_model_1.IRAM[11] [2]);
  nand (_09282_, _09281_, _09280_);
  nand (_09283_, _09282_, _08708_);
  or (_09284_, _09099_, \oc8051_golden_model_1.IRAM[8] [2]);
  or (_09285_, _08700_, \oc8051_golden_model_1.IRAM[9] [2]);
  nand (_09286_, _09285_, _09284_);
  nand (_09287_, _09286_, _08709_);
  nand (_09288_, _09287_, _09283_);
  nand (_09289_, _09288_, _08692_);
  nand (_09290_, _08700_, _07764_);
  or (_09291_, _08700_, \oc8051_golden_model_1.IRAM[15] [2]);
  nand (_09292_, _09291_, _09290_);
  nand (_09293_, _09292_, _08708_);
  or (_09294_, _09099_, \oc8051_golden_model_1.IRAM[12] [2]);
  or (_09295_, _08700_, \oc8051_golden_model_1.IRAM[13] [2]);
  nand (_09296_, _09295_, _09294_);
  nand (_09297_, _09296_, _08709_);
  nand (_09298_, _09297_, _09293_);
  nand (_09299_, _09298_, _08719_);
  and (_09300_, _09299_, _08732_);
  and (_09301_, _09300_, _09289_);
  nor (_09302_, _09301_, _09279_);
  nand (_09303_, _08700_, \oc8051_golden_model_1.IRAM[0] [1]);
  or (_09304_, _08700_, _07307_);
  and (_09305_, _09304_, _08709_);
  nand (_09306_, _09305_, _09303_);
  nand (_09307_, _08700_, \oc8051_golden_model_1.IRAM[2] [1]);
  or (_09308_, _08700_, _07311_);
  and (_09309_, _09308_, _08708_);
  nand (_09310_, _09309_, _09307_);
  nand (_09311_, _09310_, _09306_);
  nand (_09312_, _09311_, _08692_);
  nand (_09313_, _08700_, \oc8051_golden_model_1.IRAM[4] [1]);
  or (_09314_, _08700_, _07327_);
  and (_09315_, _09314_, _08709_);
  nand (_09316_, _09315_, _09313_);
  nand (_09317_, _08700_, \oc8051_golden_model_1.IRAM[6] [1]);
  or (_09318_, _08700_, _07319_);
  and (_09319_, _09318_, _08708_);
  nand (_09320_, _09319_, _09317_);
  nand (_09321_, _09320_, _09316_);
  nand (_09322_, _09321_, _08719_);
  and (_09323_, _09322_, _08682_);
  and (_09324_, _09323_, _09312_);
  or (_09325_, _09099_, \oc8051_golden_model_1.IRAM[10] [1]);
  or (_09326_, _08700_, \oc8051_golden_model_1.IRAM[11] [1]);
  nand (_09327_, _09326_, _09325_);
  nand (_09328_, _09327_, _08708_);
  or (_09329_, _09099_, \oc8051_golden_model_1.IRAM[8] [1]);
  or (_09330_, _08700_, \oc8051_golden_model_1.IRAM[9] [1]);
  nand (_09331_, _09330_, _09329_);
  nand (_09332_, _09331_, _08709_);
  nand (_09333_, _09332_, _09328_);
  nand (_09334_, _09333_, _08692_);
  or (_09335_, _09099_, \oc8051_golden_model_1.IRAM[14] [1]);
  or (_09336_, _08700_, \oc8051_golden_model_1.IRAM[15] [1]);
  nand (_09337_, _09336_, _09335_);
  nand (_09338_, _09337_, _08708_);
  or (_09339_, _09099_, \oc8051_golden_model_1.IRAM[12] [1]);
  or (_09340_, _08700_, \oc8051_golden_model_1.IRAM[13] [1]);
  nand (_09341_, _09340_, _09339_);
  nand (_09342_, _09341_, _08709_);
  nand (_09343_, _09342_, _09338_);
  nand (_09344_, _09343_, _08719_);
  and (_09345_, _09344_, _08732_);
  and (_09346_, _09345_, _09334_);
  nor (_09347_, _09346_, _09324_);
  nand (_09348_, _08700_, \oc8051_golden_model_1.IRAM[0] [0]);
  or (_09349_, _08700_, _07077_);
  and (_09350_, _09349_, _08709_);
  nand (_09351_, _09350_, _09348_);
  nand (_09352_, _08700_, \oc8051_golden_model_1.IRAM[2] [0]);
  or (_09353_, _08700_, _07082_);
  and (_09354_, _09353_, _08708_);
  nand (_09355_, _09354_, _09352_);
  nand (_09356_, _09355_, _09351_);
  nand (_09357_, _09356_, _08692_);
  nand (_09358_, _08700_, \oc8051_golden_model_1.IRAM[4] [0]);
  or (_09359_, _08700_, _07100_);
  and (_09360_, _09359_, _08709_);
  nand (_09361_, _09360_, _09358_);
  nand (_09362_, _08700_, \oc8051_golden_model_1.IRAM[6] [0]);
  or (_09363_, _08700_, _07092_);
  and (_09364_, _09363_, _08708_);
  nand (_09365_, _09364_, _09362_);
  nand (_09366_, _09365_, _09361_);
  nand (_09367_, _09366_, _08719_);
  and (_09368_, _09367_, _08682_);
  and (_09369_, _09368_, _09357_);
  or (_09370_, _09099_, \oc8051_golden_model_1.IRAM[10] [0]);
  or (_09371_, _08700_, \oc8051_golden_model_1.IRAM[11] [0]);
  nand (_09372_, _09371_, _09370_);
  nand (_09373_, _09372_, _08708_);
  or (_09374_, _09099_, \oc8051_golden_model_1.IRAM[8] [0]);
  or (_09375_, _08700_, \oc8051_golden_model_1.IRAM[9] [0]);
  nand (_09376_, _09375_, _09374_);
  nand (_09377_, _09376_, _08709_);
  nand (_09378_, _09377_, _09373_);
  nand (_09379_, _09378_, _08692_);
  nand (_09380_, _08700_, \oc8051_golden_model_1.IRAM[14] [0]);
  or (_09381_, _08700_, _07119_);
  and (_09382_, _09381_, _09380_);
  nand (_09383_, _09382_, _08708_);
  nand (_09384_, _08700_, _07124_);
  or (_09385_, _08700_, \oc8051_golden_model_1.IRAM[13] [0]);
  nand (_09386_, _09385_, _09384_);
  nand (_09387_, _09386_, _08709_);
  nand (_09388_, _09387_, _09383_);
  nand (_09389_, _09388_, _08719_);
  and (_09390_, _09389_, _08732_);
  and (_09391_, _09390_, _09379_);
  or (_09392_, _09391_, _09369_);
  not (_09393_, _09392_);
  and (_09394_, _09393_, _09347_);
  and (_09395_, _09394_, _09302_);
  and (_09396_, _09395_, _09257_);
  and (_09397_, _09396_, _09212_);
  and (_09398_, _09397_, _09167_);
  and (_09399_, _09398_, _09122_);
  nor (_09400_, _09399_, _09076_);
  and (_09401_, _09399_, _09076_);
  or (_09402_, _09401_, _09400_);
  or (_09403_, _09402_, _07541_);
  and (_09404_, _09403_, _09075_);
  and (_09405_, _09404_, _09074_);
  and (_09406_, _08768_, _07261_);
  or (_09407_, _09406_, _06361_);
  or (_09408_, _09407_, _09405_);
  and (_09409_, _08657_, \oc8051_golden_model_1.PC [7]);
  and (_09410_, _05634_, \oc8051_golden_model_1.PC [2]);
  and (_09411_, _09410_, \oc8051_golden_model_1.PC [3]);
  and (_09412_, _09411_, _09409_);
  and (_09413_, _09411_, _08657_);
  nor (_09414_, _09413_, \oc8051_golden_model_1.PC [7]);
  nor (_09415_, _09414_, _09412_);
  not (_09416_, _09415_);
  nand (_09417_, _09416_, _06361_);
  and (_09418_, _09417_, _09408_);
  or (_09419_, _09418_, _05940_);
  and (_09420_, _08794_, _05940_);
  nor (_09421_, _09420_, _07270_);
  and (_09422_, _09421_, _09419_);
  and (_09423_, _08649_, _07270_);
  and (_09424_, _05938_, _05923_);
  or (_09425_, _09424_, _09423_);
  or (_09426_, _09425_, _09422_);
  not (_09427_, _09424_);
  not (_09428_, _08142_);
  not (_09429_, _08244_);
  not (_09430_, _08541_);
  not (_09431_, _07776_);
  not (_09432_, _07357_);
  and (_09433_, _09432_, _07133_);
  and (_09434_, _09433_, _09431_);
  and (_09435_, _09434_, _07595_);
  and (_09436_, _09435_, _09430_);
  and (_09437_, _09436_, _09429_);
  and (_09438_, _09437_, _09428_);
  nand (_09439_, _09438_, _08552_);
  or (_09440_, _09438_, _08552_);
  and (_09441_, _09440_, _09439_);
  or (_09442_, _09441_, _09427_);
  and (_09443_, _09442_, _09426_);
  or (_09444_, _09443_, _07281_);
  not (_09445_, _07286_);
  or (_09446_, _09121_, _09098_);
  or (_09447_, _09166_, _09144_);
  or (_09448_, _09211_, _09189_);
  or (_09449_, _09256_, _09234_);
  or (_09450_, _09301_, _09279_);
  or (_09451_, _09346_, _09324_);
  and (_09452_, _09392_, _09451_);
  and (_09453_, _09452_, _09450_);
  and (_09454_, _09453_, _09449_);
  and (_09455_, _09454_, _09448_);
  and (_09456_, _09455_, _09447_);
  and (_09457_, _09456_, _09446_);
  nor (_09458_, _09457_, _09076_);
  and (_09459_, _09457_, _09076_);
  or (_09460_, _09459_, _09458_);
  or (_09461_, _09460_, _07282_);
  and (_09462_, _09461_, _09445_);
  and (_09463_, _09462_, _09444_);
  or (_09464_, _09463_, _08551_);
  and (_09465_, _09464_, _07535_);
  or (_09466_, _09465_, _07878_);
  and (_09467_, _09466_, _07877_);
  not (_09468_, \oc8051_golden_model_1.PC [15]);
  and (_09469_, \oc8051_golden_model_1.PC [12], \oc8051_golden_model_1.PC [13]);
  and (_09470_, \oc8051_golden_model_1.PC [11], \oc8051_golden_model_1.PC [10]);
  and (_09471_, \oc8051_golden_model_1.PC [9], \oc8051_golden_model_1.PC [8]);
  and (_09472_, _09471_, _09470_);
  and (_09473_, _09472_, _09412_);
  and (_09474_, _09473_, _09469_);
  and (_09475_, _09474_, \oc8051_golden_model_1.PC [14]);
  and (_09476_, _09475_, _09468_);
  nor (_09477_, _09475_, _09468_);
  or (_09478_, _09477_, _09476_);
  not (_09479_, _09478_);
  nand (_09480_, _09479_, _06361_);
  and (_09481_, _09472_, _08659_);
  and (_09482_, _09481_, _09469_);
  and (_09483_, _09482_, \oc8051_golden_model_1.PC [14]);
  and (_09485_, _09483_, _09468_);
  nor (_09486_, _09483_, _09468_);
  or (_09487_, _09486_, _09485_);
  or (_09488_, _09487_, _06361_);
  and (_09489_, _09488_, _09480_);
  and (_09490_, _09489_, _07872_);
  and (_09491_, _09490_, _07875_);
  or (_40572_, _09491_, _09467_);
  not (_09492_, \oc8051_golden_model_1.B [7]);
  nor (_09493_, _01347_, _09492_);
  nor (_09494_, _07942_, _09492_);
  and (_09495_, _08575_, _07942_);
  or (_09496_, _09495_, _09494_);
  and (_09497_, _09496_, _06536_);
  not (_09498_, _07942_);
  nor (_09499_, _08040_, _09498_);
  or (_09500_, _09499_, _09494_);
  or (_09501_, _09500_, _07215_);
  nor (_09502_, _08634_, _09492_);
  and (_09503_, _08649_, _08634_);
  or (_09505_, _09503_, _09502_);
  and (_09506_, _09505_, _06268_);
  and (_09507_, _08768_, _07942_);
  or (_09508_, _09507_, _09494_);
  or (_09509_, _09508_, _07151_);
  and (_09510_, _07942_, \oc8051_golden_model_1.ACC [7]);
  or (_09511_, _09510_, _09494_);
  and (_09512_, _09511_, _07141_);
  nor (_09513_, _07141_, _09492_);
  or (_09514_, _09513_, _06341_);
  or (_09515_, _09514_, _09512_);
  and (_09516_, _09515_, _06273_);
  and (_09517_, _09516_, _09509_);
  and (_09518_, _08773_, _08634_);
  or (_09519_, _09518_, _09502_);
  and (_09520_, _09519_, _06272_);
  or (_09521_, _09520_, _06461_);
  or (_09522_, _09521_, _09517_);
  or (_09523_, _09500_, _07166_);
  and (_09524_, _09523_, _09522_);
  or (_09525_, _09524_, _06464_);
  or (_09526_, _09511_, _06465_);
  and (_09527_, _09526_, _06269_);
  and (_09528_, _09527_, _09525_);
  or (_09529_, _09528_, _09506_);
  and (_09530_, _09529_, _06262_);
  and (_09531_, _06370_, _06491_);
  or (_09532_, _09502_, _08789_);
  and (_09533_, _09532_, _06261_);
  and (_09534_, _09533_, _09519_);
  or (_09535_, _09534_, _09531_);
  or (_09536_, _09535_, _09530_);
  not (_09537_, _09531_);
  and (_09538_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [7]);
  and (_09539_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [6]);
  and (_09540_, _09539_, _09538_);
  and (_09541_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [7]);
  and (_09542_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [6]);
  nor (_09543_, _09542_, _09541_);
  nor (_09544_, _09543_, _09540_);
  and (_09545_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [6]);
  and (_09546_, \oc8051_golden_model_1.ACC [3], \oc8051_golden_model_1.B [7]);
  and (_09547_, _09546_, _09545_);
  and (_09548_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [7]);
  and (_09549_, _09548_, _09539_);
  and (_09550_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [5]);
  nor (_09551_, _09548_, _09539_);
  nor (_09552_, _09551_, _09549_);
  and (_09553_, _09552_, _09550_);
  nor (_09554_, _09553_, _09549_);
  and (_09555_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [7]);
  and (_09556_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [6]);
  and (_09557_, _09556_, _09555_);
  nor (_09558_, _09556_, _09555_);
  nor (_09559_, _09558_, _09557_);
  not (_09560_, _09559_);
  nor (_09561_, _09560_, _09554_);
  and (_09562_, _09560_, _09554_);
  nor (_09563_, _09562_, _09561_);
  and (_09564_, _09563_, _09547_);
  nor (_09565_, _09563_, _09547_);
  nor (_09566_, _09565_, _09564_);
  and (_09567_, _09566_, _09544_);
  and (_09568_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [7]);
  and (_09569_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [6]);
  and (_09570_, _09569_, _09568_);
  nor (_09571_, _09569_, _09568_);
  nor (_09572_, _09571_, _09570_);
  and (_09573_, _09572_, _09540_);
  nor (_09574_, _09572_, _09540_);
  nor (_09575_, _09574_, _09573_);
  and (_09576_, _09575_, _09557_);
  nor (_09577_, _09575_, _09557_);
  nor (_09578_, _09577_, _09576_);
  and (_09579_, _09578_, _09538_);
  nor (_09580_, _09578_, _09538_);
  nor (_09581_, _09580_, _09579_);
  and (_09582_, _09581_, _09567_);
  nor (_09583_, _09564_, _09561_);
  not (_09584_, _09583_);
  nor (_09585_, _09581_, _09567_);
  nor (_09586_, _09585_, _09582_);
  and (_09587_, _09586_, _09584_);
  nor (_09588_, _09587_, _09582_);
  nor (_09589_, _09576_, _09573_);
  not (_09590_, _09589_);
  and (_09591_, \oc8051_golden_model_1.ACC [6], \oc8051_golden_model_1.B [7]);
  and (_09592_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [7]);
  and (_09593_, _09592_, _09591_);
  nor (_09594_, _09592_, _09591_);
  nor (_09595_, _09594_, _09593_);
  and (_09596_, _09595_, _09570_);
  nor (_09597_, _09595_, _09570_);
  nor (_09598_, _09597_, _09596_);
  and (_09599_, _09598_, _09579_);
  nor (_09600_, _09598_, _09579_);
  nor (_09601_, _09600_, _09599_);
  and (_09602_, _09601_, _09590_);
  nor (_09603_, _09601_, _09590_);
  nor (_09604_, _09603_, _09602_);
  not (_09605_, _09604_);
  nor (_09606_, _09605_, _09588_);
  and (_09607_, \oc8051_golden_model_1.ACC [7], \oc8051_golden_model_1.B [7]);
  not (_09608_, _09607_);
  nor (_09609_, _09608_, _09569_);
  nor (_09610_, _09609_, _09596_);
  nor (_09611_, _09602_, _09599_);
  nor (_09612_, _09611_, _09610_);
  and (_09613_, _09611_, _09610_);
  nor (_09614_, _09613_, _09612_);
  and (_09615_, _09614_, _09606_);
  or (_09616_, _09612_, _09593_);
  or (_09617_, _09616_, _09615_);
  and (_09618_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [6]);
  and (_09619_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [7]);
  and (_09620_, _09619_, _09618_);
  not (_09621_, _09618_);
  and (_09622_, _09619_, _09621_);
  and (_09623_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [5]);
  and (_09624_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [3]);
  and (_09625_, _09624_, _09539_);
  and (_09626_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [6]);
  and (_09627_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [4]);
  nor (_09628_, _09627_, _09626_);
  nor (_09629_, _09628_, _09625_);
  and (_09630_, _09629_, _09623_);
  nor (_09631_, _09629_, _09623_);
  nor (_09632_, _09631_, _09630_);
  and (_09633_, _09632_, _09622_);
  nor (_09634_, _09633_, _09620_);
  nor (_09635_, _09552_, _09550_);
  nor (_09636_, _09635_, _09553_);
  not (_09637_, _09636_);
  nor (_09638_, _09637_, _09634_);
  and (_09639_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [3]);
  and (_09640_, \oc8051_golden_model_1.ACC [2], \oc8051_golden_model_1.B [7]);
  and (_09641_, _09640_, _09639_);
  nor (_09642_, _09630_, _09625_);
  nor (_09643_, _09546_, _09545_);
  nor (_09644_, _09643_, _09547_);
  not (_09645_, _09644_);
  nor (_09646_, _09645_, _09642_);
  and (_09647_, _09645_, _09642_);
  nor (_09648_, _09647_, _09646_);
  and (_09649_, _09648_, _09641_);
  nor (_09650_, _09648_, _09641_);
  nor (_09651_, _09650_, _09649_);
  and (_09652_, _09637_, _09634_);
  nor (_09653_, _09652_, _09638_);
  and (_09654_, _09653_, _09651_);
  nor (_09655_, _09654_, _09638_);
  not (_09656_, _09655_);
  nor (_09657_, _09566_, _09544_);
  nor (_09658_, _09657_, _09567_);
  and (_09660_, _09658_, _09656_);
  nor (_09661_, _09649_, _09646_);
  not (_09663_, _09661_);
  nor (_09664_, _09658_, _09656_);
  nor (_09666_, _09664_, _09660_);
  and (_09667_, _09666_, _09663_);
  nor (_09669_, _09667_, _09660_);
  nor (_09670_, _09586_, _09584_);
  nor (_09672_, _09670_, _09587_);
  not (_09673_, _09672_);
  nor (_09675_, _09673_, _09669_);
  and (_09676_, _09605_, _09588_);
  nor (_09678_, _09676_, _09606_);
  and (_09679_, _09678_, _09675_);
  and (_09681_, _09679_, _09614_);
  and (_09682_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [7]);
  and (_09684_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [6]);
  and (_09685_, _09684_, _09682_);
  and (_09687_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [2]);
  and (_09688_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [7]);
  nor (_09690_, _09688_, _09618_);
  nor (_09691_, _09690_, _09685_);
  and (_09693_, _09691_, _09687_);
  nor (_09694_, _09693_, _09685_);
  and (_09696_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [6]);
  nor (_09697_, _09696_, _09682_);
  nor (_09698_, _09697_, _09620_);
  not (_09699_, _09698_);
  nor (_09700_, _09699_, _09694_);
  and (_09701_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [3]);
  and (_09702_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [4]);
  and (_09703_, _09702_, _09624_);
  nor (_09704_, _09702_, _09624_);
  nor (_09705_, _09704_, _09703_);
  and (_09706_, _09705_, _09701_);
  nor (_09707_, _09705_, _09701_);
  nor (_09708_, _09707_, _09706_);
  and (_09709_, _09699_, _09694_);
  nor (_09710_, _09709_, _09700_);
  and (_09711_, _09710_, _09708_);
  nor (_09712_, _09711_, _09700_);
  nor (_09713_, _09632_, _09622_);
  nor (_09714_, _09713_, _09633_);
  not (_09715_, _09714_);
  nor (_09716_, _09715_, _09712_);
  and (_09717_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [2]);
  and (_09718_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [7]);
  and (_09719_, _09718_, _09717_);
  nor (_09720_, _09706_, _09703_);
  nor (_09721_, _09640_, _09639_);
  nor (_09722_, _09721_, _09641_);
  not (_09723_, _09722_);
  nor (_09724_, _09723_, _09720_);
  and (_09725_, _09723_, _09720_);
  nor (_09726_, _09725_, _09724_);
  and (_09727_, _09726_, _09719_);
  nor (_09728_, _09726_, _09719_);
  nor (_09729_, _09728_, _09727_);
  and (_09730_, _09715_, _09712_);
  nor (_09731_, _09730_, _09716_);
  and (_09732_, _09731_, _09729_);
  nor (_09733_, _09732_, _09716_);
  nor (_09734_, _09653_, _09651_);
  nor (_09735_, _09734_, _09654_);
  not (_09736_, _09735_);
  nor (_09737_, _09736_, _09733_);
  nor (_09738_, _09727_, _09724_);
  not (_09739_, _09738_);
  and (_09740_, _09736_, _09733_);
  nor (_09741_, _09740_, _09737_);
  and (_09742_, _09741_, _09739_);
  nor (_09743_, _09742_, _09737_);
  nor (_09744_, _09666_, _09663_);
  nor (_09745_, _09744_, _09667_);
  not (_09746_, _09745_);
  nor (_09747_, _09746_, _09743_);
  and (_09748_, _09673_, _09669_);
  nor (_09749_, _09748_, _09675_);
  and (_09750_, _09749_, _09747_);
  nor (_09751_, _09678_, _09675_);
  nor (_09752_, _09751_, _09679_);
  and (_09753_, _09752_, _09750_);
  nor (_09755_, _09752_, _09750_);
  nor (_09757_, _09755_, _09753_);
  and (_09758_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [0]);
  and (_09760_, _09758_, _09618_);
  and (_09761_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [2]);
  and (_09763_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [1]);
  nor (_09764_, _09763_, _09684_);
  nor (_09766_, _09764_, _09760_);
  and (_09767_, _09766_, _09761_);
  nor (_09769_, _09767_, _09760_);
  not (_09770_, _09769_);
  nor (_09772_, _09691_, _09687_);
  nor (_09773_, _09772_, _09693_);
  and (_09775_, _09773_, _09770_);
  and (_09776_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [2]);
  and (_09778_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [3]);
  and (_09779_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [3]);
  and (_09781_, _09779_, _09778_);
  nor (_09782_, _09779_, _09778_);
  nor (_09784_, _09782_, _09781_);
  and (_09785_, _09784_, _09776_);
  nor (_09787_, _09784_, _09776_);
  nor (_09788_, _09787_, _09785_);
  nor (_09790_, _09773_, _09770_);
  nor (_09791_, _09790_, _09775_);
  and (_09792_, _09791_, _09788_);
  nor (_09793_, _09792_, _09775_);
  nor (_09794_, _09710_, _09708_);
  nor (_09795_, _09794_, _09711_);
  not (_09796_, _09795_);
  nor (_09797_, _09796_, _09793_);
  and (_09798_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [0]);
  and (_09799_, _09798_, _09718_);
  nor (_09800_, _09785_, _09781_);
  nor (_09801_, _09718_, _09717_);
  nor (_09802_, _09801_, _09719_);
  not (_09803_, _09802_);
  nor (_09804_, _09803_, _09800_);
  and (_09805_, _09803_, _09800_);
  nor (_09806_, _09805_, _09804_);
  and (_09807_, _09806_, _09799_);
  nor (_09808_, _09806_, _09799_);
  nor (_09809_, _09808_, _09807_);
  and (_09810_, _09796_, _09793_);
  nor (_09811_, _09810_, _09797_);
  and (_09812_, _09811_, _09809_);
  nor (_09813_, _09812_, _09797_);
  nor (_09814_, _09731_, _09729_);
  nor (_09815_, _09814_, _09732_);
  not (_09816_, _09815_);
  nor (_09817_, _09816_, _09813_);
  nor (_09818_, _09807_, _09804_);
  not (_09819_, _09818_);
  and (_09820_, _09816_, _09813_);
  nor (_09821_, _09820_, _09817_);
  and (_09822_, _09821_, _09819_);
  nor (_09823_, _09822_, _09817_);
  nor (_09824_, _09741_, _09739_);
  nor (_09825_, _09824_, _09742_);
  not (_09826_, _09825_);
  nor (_09827_, _09826_, _09823_);
  and (_09828_, _09746_, _09743_);
  nor (_09829_, _09828_, _09747_);
  and (_09830_, _09829_, _09827_);
  nor (_09831_, _09749_, _09747_);
  nor (_09832_, _09831_, _09750_);
  nand (_09833_, _09832_, _09830_);
  and (_09834_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [1]);
  and (_09835_, _09834_, _09758_);
  and (_09836_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [3]);
  nor (_09837_, _09834_, _09758_);
  nor (_09838_, _09837_, _09835_);
  and (_09839_, _09838_, _09836_);
  nor (_09840_, _09839_, _09835_);
  not (_09841_, _09840_);
  nor (_09842_, _09766_, _09761_);
  nor (_09843_, _09842_, _09767_);
  and (_09844_, _09843_, _09841_);
  and (_09845_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [5]);
  and (_09846_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [3]);
  and (_09847_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [2]);
  and (_09848_, _09847_, _09846_);
  nor (_09849_, _09847_, _09846_);
  nor (_09850_, _09849_, _09848_);
  and (_09851_, _09850_, _09845_);
  nor (_09852_, _09850_, _09845_);
  nor (_09853_, _09852_, _09851_);
  nor (_09854_, _09843_, _09841_);
  nor (_09855_, _09854_, _09844_);
  and (_09856_, _09855_, _09853_);
  nor (_09857_, _09856_, _09844_);
  not (_09858_, _09857_);
  nor (_09859_, _09791_, _09788_);
  nor (_09860_, _09859_, _09792_);
  and (_09861_, _09860_, _09858_);
  nor (_09862_, _09851_, _09848_);
  and (_09863_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [6]);
  and (_09864_, \oc8051_golden_model_1.ACC [0], \oc8051_golden_model_1.B [7]);
  nor (_09865_, _09864_, _09863_);
  nor (_09866_, _09865_, _09799_);
  not (_09867_, _09866_);
  nor (_09868_, _09867_, _09862_);
  and (_09869_, _09867_, _09862_);
  nor (_09870_, _09869_, _09868_);
  nor (_09871_, _09860_, _09858_);
  nor (_09872_, _09871_, _09861_);
  and (_09873_, _09872_, _09870_);
  nor (_09874_, _09873_, _09861_);
  nor (_09875_, _09811_, _09809_);
  nor (_09876_, _09875_, _09812_);
  not (_09877_, _09876_);
  nor (_09878_, _09877_, _09874_);
  and (_09879_, _09877_, _09874_);
  nor (_09880_, _09879_, _09878_);
  and (_09881_, _09880_, _09868_);
  nor (_09882_, _09881_, _09878_);
  nor (_09883_, _09821_, _09819_);
  nor (_09884_, _09883_, _09822_);
  not (_09885_, _09884_);
  nor (_09886_, _09885_, _09882_);
  and (_09887_, _09826_, _09823_);
  nor (_09888_, _09887_, _09827_);
  and (_09889_, _09888_, _09886_);
  nor (_09890_, _09829_, _09827_);
  nor (_09891_, _09890_, _09830_);
  and (_09892_, _09891_, _09889_);
  nor (_09893_, _09891_, _09889_);
  nor (_09894_, _09893_, _09892_);
  and (_09895_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [0]);
  and (_09896_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [3]);
  and (_09897_, _09896_, _09895_);
  and (_09898_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [2]);
  nor (_09899_, _09896_, _09895_);
  nor (_09900_, _09899_, _09897_);
  and (_09901_, _09900_, _09898_);
  nor (_09902_, _09901_, _09897_);
  not (_09903_, _09902_);
  nor (_09904_, _09838_, _09836_);
  nor (_09905_, _09904_, _09839_);
  and (_09906_, _09905_, _09903_);
  and (_09907_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [0]);
  and (_09908_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [2]);
  and (_09909_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [4]);
  and (_09910_, _09909_, _09908_);
  nor (_09911_, _09909_, _09908_);
  nor (_09912_, _09911_, _09910_);
  and (_09913_, _09912_, _09907_);
  nor (_09914_, _09912_, _09907_);
  nor (_09915_, _09914_, _09913_);
  nor (_09916_, _09905_, _09903_);
  nor (_09917_, _09916_, _09906_);
  and (_09918_, _09917_, _09915_);
  nor (_09919_, _09918_, _09906_);
  not (_09920_, _09919_);
  nor (_09921_, _09855_, _09853_);
  nor (_09922_, _09921_, _09856_);
  and (_09923_, _09922_, _09920_);
  not (_09924_, _09798_);
  nor (_09925_, _09913_, _09910_);
  nor (_09926_, _09925_, _09924_);
  and (_09927_, _09925_, _09924_);
  nor (_09928_, _09927_, _09926_);
  nor (_09929_, _09922_, _09920_);
  nor (_09930_, _09929_, _09923_);
  and (_09931_, _09930_, _09928_);
  nor (_09932_, _09931_, _09923_);
  not (_09933_, _09932_);
  nor (_09934_, _09872_, _09870_);
  nor (_09935_, _09934_, _09873_);
  and (_09936_, _09935_, _09933_);
  nor (_09937_, _09935_, _09933_);
  nor (_09938_, _09937_, _09936_);
  and (_09939_, _09938_, _09926_);
  nor (_09940_, _09939_, _09936_);
  nor (_09941_, _09880_, _09868_);
  nor (_09942_, _09941_, _09881_);
  not (_09943_, _09942_);
  nor (_09944_, _09943_, _09940_);
  and (_09945_, _09885_, _09882_);
  nor (_09946_, _09945_, _09886_);
  and (_09947_, _09946_, _09944_);
  nor (_09948_, _09888_, _09886_);
  nor (_09949_, _09948_, _09889_);
  nand (_09950_, _09949_, _09947_);
  or (_09951_, _09949_, _09947_);
  and (_09952_, _09951_, _09950_);
  and (_09953_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [3]);
  and (_09954_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [2]);
  and (_09955_, _09954_, _09953_);
  and (_09956_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [2]);
  nor (_09957_, _09954_, _09953_);
  nor (_09958_, _09957_, _09955_);
  and (_09959_, _09958_, _09956_);
  nor (_09960_, _09959_, _09955_);
  not (_09961_, _09960_);
  nor (_09962_, _09900_, _09898_);
  nor (_09963_, _09962_, _09901_);
  and (_09964_, _09963_, _09961_);
  and (_09965_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [0]);
  and (_09966_, _09965_, _09909_);
  and (_09967_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [3]);
  and (_09968_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [0]);
  nor (_09969_, _09968_, _09967_);
  nor (_09970_, _09969_, _09966_);
  nor (_09971_, _09963_, _09961_);
  nor (_09972_, _09971_, _09964_);
  and (_09973_, _09972_, _09970_);
  nor (_09974_, _09973_, _09964_);
  not (_09975_, _09974_);
  nor (_09976_, _09917_, _09915_);
  nor (_09977_, _09976_, _09918_);
  and (_09978_, _09977_, _09975_);
  nor (_09979_, _09977_, _09975_);
  nor (_09980_, _09979_, _09978_);
  and (_09981_, _09980_, _09966_);
  nor (_09982_, _09981_, _09978_);
  not (_09983_, _09982_);
  nor (_09984_, _09930_, _09928_);
  nor (_09985_, _09984_, _09931_);
  and (_09986_, _09985_, _09983_);
  nor (_09987_, _09938_, _09926_);
  nor (_09988_, _09987_, _09939_);
  and (_09989_, _09988_, _09986_);
  and (_09990_, _09943_, _09940_);
  nor (_09991_, _09990_, _09944_);
  and (_09992_, _09991_, _09989_);
  nor (_09993_, _09946_, _09944_);
  nor (_09994_, _09993_, _09947_);
  and (_09995_, _09994_, _09992_);
  nor (_09996_, _09994_, _09992_);
  nor (_09997_, _09996_, _09995_);
  and (_09998_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [2]);
  and (_09999_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [1]);
  and (_10000_, _09999_, _09998_);
  and (_10001_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [0]);
  nor (_10002_, _09999_, _09998_);
  nor (_10003_, _10002_, _10000_);
  and (_10004_, _10003_, _10001_);
  nor (_10005_, _10004_, _10000_);
  not (_10006_, _10005_);
  nor (_10007_, _09958_, _09956_);
  nor (_10008_, _10007_, _09959_);
  and (_10009_, _10008_, _10006_);
  nor (_10010_, _10008_, _10006_);
  nor (_10011_, _10010_, _10009_);
  and (_10012_, _10011_, _09965_);
  nor (_10013_, _10012_, _10009_);
  not (_10014_, _10013_);
  nor (_10015_, _09972_, _09970_);
  nor (_10016_, _10015_, _09973_);
  and (_10017_, _10016_, _10014_);
  nor (_10018_, _09980_, _09966_);
  nor (_10019_, _10018_, _09981_);
  and (_10020_, _10019_, _10017_);
  nor (_10021_, _09985_, _09983_);
  nor (_10022_, _10021_, _09986_);
  and (_10023_, _10022_, _10020_);
  nor (_10024_, _09988_, _09986_);
  nor (_10025_, _10024_, _09989_);
  and (_10026_, _10025_, _10023_);
  nor (_10027_, _09991_, _09989_);
  nor (_10028_, _10027_, _09992_);
  and (_10029_, _10028_, _10026_);
  and (_10030_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [0]);
  and (_10031_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [0]);
  and (_10032_, _10031_, _10030_);
  nor (_10033_, _10003_, _10001_);
  nor (_10034_, _10033_, _10004_);
  and (_10035_, _10034_, _10032_);
  nor (_10036_, _10011_, _09965_);
  nor (_10037_, _10036_, _10012_);
  and (_10038_, _10037_, _10035_);
  nor (_10039_, _10016_, _10014_);
  nor (_10040_, _10039_, _10017_);
  and (_10041_, _10040_, _10038_);
  nor (_10042_, _10019_, _10017_);
  nor (_10043_, _10042_, _10020_);
  and (_10044_, _10043_, _10041_);
  nor (_10045_, _10022_, _10020_);
  nor (_10046_, _10045_, _10023_);
  and (_10047_, _10046_, _10044_);
  nor (_10048_, _10025_, _10023_);
  nor (_10049_, _10048_, _10026_);
  and (_10050_, _10049_, _10047_);
  nor (_10051_, _10028_, _10026_);
  nor (_10052_, _10051_, _10029_);
  and (_10053_, _10052_, _10050_);
  nor (_10054_, _10053_, _10029_);
  not (_10055_, _10054_);
  and (_10056_, _10055_, _09997_);
  or (_10057_, _10056_, _09995_);
  nand (_10058_, _10057_, _09952_);
  and (_10059_, _10058_, _09950_);
  not (_10060_, _10059_);
  and (_10061_, _10060_, _09894_);
  or (_10062_, _10061_, _09892_);
  or (_10063_, _09832_, _09830_);
  and (_10064_, _10063_, _09833_);
  nand (_10065_, _10064_, _10062_);
  and (_10066_, _10065_, _09833_);
  not (_10067_, _10066_);
  and (_10068_, _10067_, _09757_);
  or (_10069_, _10068_, _09753_);
  nor (_10070_, _09679_, _09606_);
  and (_10071_, _10070_, _09614_);
  nor (_10072_, _10070_, _09614_);
  or (_10073_, _10072_, _10071_);
  and (_10074_, _10073_, _10069_);
  or (_10075_, _10074_, _09681_);
  or (_10076_, _10075_, _09617_);
  or (_10077_, _10076_, _09537_);
  and (_10078_, _10077_, _06258_);
  and (_10079_, _10078_, _09536_);
  not (_10080_, _07215_);
  and (_10081_, _08808_, _08634_);
  or (_10082_, _10081_, _09502_);
  and (_10083_, _10082_, _06257_);
  or (_10084_, _10083_, _10080_);
  or (_10085_, _10084_, _10079_);
  and (_10086_, _10085_, _09501_);
  or (_10087_, _10086_, _07460_);
  and (_10088_, _08755_, _07942_);
  or (_10089_, _09494_, _07208_);
  or (_10090_, _10089_, _10088_);
  and (_10091_, _10090_, _05982_);
  and (_10092_, _10091_, _10087_);
  and (_10093_, _06370_, _05944_);
  not (_10094_, _05982_);
  and (_10095_, _09021_, _07942_);
  or (_10096_, _10095_, _09494_);
  and (_10097_, _10096_, _10094_);
  or (_10098_, _10097_, _10093_);
  or (_10099_, _10098_, _10092_);
  not (_10100_, _10093_);
  not (_10101_, \oc8051_golden_model_1.B [1]);
  nor (_10102_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.B [4]);
  nor (_10103_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.B [3]);
  and (_10104_, _10103_, _10102_);
  and (_10105_, _10104_, _10101_);
  not (_10106_, \oc8051_golden_model_1.B [0]);
  and (_10107_, _10106_, \oc8051_golden_model_1.ACC [7]);
  nor (_10108_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.B [7]);
  and (_10109_, _10108_, _10107_);
  and (_10110_, _10109_, _10105_);
  and (_10111_, \oc8051_golden_model_1.B [0], _08572_);
  not (_10112_, _10111_);
  and (_10113_, _10108_, _10105_);
  and (_10114_, _10113_, _10112_);
  or (_10115_, _10114_, _08572_);
  not (_10116_, \oc8051_golden_model_1.ACC [6]);
  and (_10117_, \oc8051_golden_model_1.B [0], _10116_);
  nor (_10118_, _10117_, _08572_);
  nor (_10119_, _10118_, _10101_);
  not (_10120_, _10119_);
  and (_10121_, _10108_, _10104_);
  and (_10122_, _10121_, _10120_);
  nor (_10123_, _10122_, _10115_);
  nor (_10124_, _10123_, _10110_);
  and (_10125_, _10122_, \oc8051_golden_model_1.B [0]);
  nor (_10126_, _10125_, _10116_);
  and (_10127_, _10126_, _10101_);
  nor (_10128_, _10126_, _10101_);
  nor (_10129_, _10128_, _10127_);
  nor (_10130_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [0]);
  nor (_10131_, _10130_, _09758_);
  nor (_10132_, _10131_, \oc8051_golden_model_1.ACC [4]);
  and (_10133_, \oc8051_golden_model_1.ACC [4], _10106_);
  nor (_10134_, _10133_, \oc8051_golden_model_1.ACC [5]);
  not (_10135_, \oc8051_golden_model_1.ACC [4]);
  and (_10136_, _10135_, \oc8051_golden_model_1.B [0]);
  nor (_10137_, _10136_, _10134_);
  nor (_10138_, _10137_, _10132_);
  not (_10139_, _10138_);
  and (_10140_, _10139_, _10129_);
  nor (_10141_, _10124_, \oc8051_golden_model_1.B [2]);
  nor (_10142_, _10141_, _10127_);
  not (_10143_, _10142_);
  nor (_10144_, _10143_, _10140_);
  not (_10145_, \oc8051_golden_model_1.B [3]);
  nor (_10146_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.B [7]);
  and (_10147_, _10146_, _10102_);
  and (_10148_, _10147_, _10145_);
  and (_10149_, \oc8051_golden_model_1.B [2], _08572_);
  not (_10150_, _10149_);
  and (_10151_, _10150_, _10148_);
  not (_10152_, _10151_);
  nor (_10153_, _10152_, _10144_);
  nor (_10154_, _10153_, _10124_);
  nor (_10155_, _10154_, _10110_);
  and (_10156_, _10147_, \oc8051_golden_model_1.ACC [7]);
  nor (_10157_, _10156_, _10148_);
  nor (_10158_, _10155_, \oc8051_golden_model_1.B [3]);
  not (_10159_, \oc8051_golden_model_1.B [2]);
  nor (_10160_, _10139_, _10129_);
  nor (_10161_, _10160_, _10140_);
  not (_10162_, _10161_);
  and (_10163_, _10162_, _10153_);
  nor (_10164_, _10153_, _10126_);
  nor (_10165_, _10164_, _10163_);
  and (_10166_, _10165_, _10159_);
  nor (_10167_, _10165_, _10159_);
  nor (_10168_, _10167_, _10166_);
  not (_10169_, _10168_);
  not (_10170_, \oc8051_golden_model_1.ACC [5]);
  nor (_10171_, _10153_, _10170_);
  and (_10172_, _10153_, _10131_);
  or (_10173_, _10172_, _10171_);
  and (_10174_, _10173_, _10101_);
  nor (_10175_, _10173_, _10101_);
  nor (_10176_, _10175_, _10136_);
  nor (_10177_, _10176_, _10174_);
  nor (_10178_, _10177_, _10169_);
  or (_10179_, _10178_, _10166_);
  nor (_10180_, _10179_, _10158_);
  nor (_10181_, _10180_, _10157_);
  nor (_10182_, _10181_, _10155_);
  nor (_10183_, _10182_, _10110_);
  not (_10184_, _10181_);
  and (_10185_, _10177_, _10169_);
  nor (_10186_, _10185_, _10178_);
  nor (_10187_, _10186_, _10184_);
  nor (_10188_, _10181_, _10165_);
  nor (_10189_, _10188_, _10187_);
  and (_10190_, _10189_, _10145_);
  nor (_10191_, _10189_, _10145_);
  nor (_10192_, _10191_, _10190_);
  not (_10193_, _10192_);
  nor (_10194_, _10181_, _10173_);
  nor (_10195_, _10175_, _10174_);
  and (_10196_, _10195_, _10136_);
  nor (_10197_, _10195_, _10136_);
  nor (_10198_, _10197_, _10196_);
  and (_10199_, _10198_, _10181_);
  or (_10200_, _10199_, _10194_);
  nor (_10201_, _10200_, \oc8051_golden_model_1.B [2]);
  and (_10202_, _10200_, \oc8051_golden_model_1.B [2]);
  nor (_10203_, _10136_, _10133_);
  and (_10204_, _10181_, _10203_);
  nor (_10205_, _10181_, \oc8051_golden_model_1.ACC [4]);
  nor (_10206_, _10205_, _10204_);
  and (_10207_, _10206_, _10101_);
  nor (_10208_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [3]);
  nor (_10209_, _10208_, _09953_);
  nor (_10210_, _10209_, \oc8051_golden_model_1.ACC [2]);
  and (_10211_, _10106_, \oc8051_golden_model_1.ACC [2]);
  nor (_10212_, _10211_, \oc8051_golden_model_1.ACC [3]);
  not (_10213_, \oc8051_golden_model_1.ACC [2]);
  and (_10214_, \oc8051_golden_model_1.B [0], _10213_);
  nor (_10215_, _10214_, _10212_);
  nor (_10216_, _10215_, _10210_);
  not (_10217_, _10216_);
  nor (_10218_, _10206_, _10101_);
  nor (_10219_, _10218_, _10207_);
  and (_10220_, _10219_, _10217_);
  nor (_10221_, _10220_, _10207_);
  nor (_10222_, _10221_, _10202_);
  nor (_10223_, _10222_, _10201_);
  nor (_10224_, _10223_, _10193_);
  nor (_10225_, _10183_, \oc8051_golden_model_1.B [4]);
  nor (_10226_, _10225_, _10190_);
  not (_10227_, _10226_);
  nor (_10228_, _10227_, _10224_);
  not (_10229_, \oc8051_golden_model_1.B [5]);
  and (_10230_, _10146_, _10229_);
  not (_10231_, _10230_);
  and (_10232_, \oc8051_golden_model_1.B [4], _08572_);
  nor (_10233_, _10232_, _10231_);
  not (_10234_, _10233_);
  nor (_10235_, _10234_, _10228_);
  nor (_10236_, _10235_, _10183_);
  nor (_10237_, _10236_, _10110_);
  and (_10238_, _10146_, \oc8051_golden_model_1.ACC [7]);
  nor (_10239_, _10238_, _10230_);
  nor (_10240_, _10237_, \oc8051_golden_model_1.B [5]);
  not (_10241_, \oc8051_golden_model_1.B [4]);
  and (_10242_, _10223_, _10193_);
  nor (_10243_, _10242_, _10224_);
  not (_10244_, _10243_);
  and (_10245_, _10244_, _10235_);
  nor (_10246_, _10235_, _10189_);
  nor (_10247_, _10246_, _10245_);
  and (_10248_, _10247_, _10241_);
  nor (_10249_, _10247_, _10241_);
  nor (_10250_, _10249_, _10248_);
  not (_10251_, _10250_);
  nor (_10252_, _10235_, _10200_);
  nor (_10253_, _10202_, _10201_);
  and (_10254_, _10253_, _10221_);
  nor (_10255_, _10253_, _10221_);
  nor (_10256_, _10255_, _10254_);
  not (_10257_, _10256_);
  and (_10258_, _10257_, _10235_);
  nor (_10259_, _10258_, _10252_);
  nor (_10260_, _10259_, \oc8051_golden_model_1.B [3]);
  and (_10261_, _10259_, \oc8051_golden_model_1.B [3]);
  nor (_10262_, _10219_, _10217_);
  nor (_10263_, _10262_, _10220_);
  not (_10264_, _10263_);
  and (_10265_, _10264_, _10235_);
  nor (_10266_, _10235_, _10206_);
  nor (_10267_, _10266_, _10265_);
  and (_10268_, _10267_, _10159_);
  nor (_10269_, _10235_, _06055_);
  and (_10270_, _10235_, _10209_);
  or (_10271_, _10270_, _10269_);
  and (_10272_, _10271_, _10101_);
  nor (_10273_, _10271_, _10101_);
  nor (_10274_, _10273_, _10214_);
  nor (_10275_, _10274_, _10272_);
  nor (_10276_, _10267_, _10159_);
  nor (_10277_, _10276_, _10268_);
  not (_10278_, _10277_);
  nor (_10279_, _10278_, _10275_);
  nor (_10280_, _10279_, _10268_);
  nor (_10281_, _10280_, _10261_);
  nor (_10282_, _10281_, _10260_);
  nor (_10283_, _10282_, _10251_);
  or (_10284_, _10283_, _10248_);
  nor (_10285_, _10284_, _10240_);
  nor (_10286_, _10285_, _10239_);
  nor (_10287_, _10286_, _10237_);
  not (_10288_, _10286_);
  and (_10289_, _10282_, _10251_);
  nor (_10290_, _10289_, _10283_);
  nor (_10291_, _10290_, _10288_);
  nor (_10292_, _10286_, _10247_);
  nor (_10293_, _10292_, _10291_);
  and (_10294_, _10293_, _10229_);
  nor (_10295_, _10293_, _10229_);
  nor (_10296_, _10295_, _10294_);
  not (_10297_, _10296_);
  nor (_10298_, _10286_, _10259_);
  nor (_10299_, _10261_, _10260_);
  nor (_10300_, _10299_, _10280_);
  and (_10301_, _10299_, _10280_);
  or (_10302_, _10301_, _10300_);
  and (_10303_, _10302_, _10286_);
  or (_10304_, _10303_, _10298_);
  and (_10305_, _10304_, _10241_);
  nor (_10306_, _10304_, _10241_);
  and (_10307_, _10278_, _10275_);
  nor (_10308_, _10307_, _10279_);
  nor (_10309_, _10308_, _10288_);
  nor (_10310_, _10286_, _10267_);
  nor (_10311_, _10310_, _10309_);
  and (_10312_, _10311_, _10145_);
  nor (_10313_, _10273_, _10272_);
  nor (_10314_, _10313_, _10214_);
  and (_10315_, _10313_, _10214_);
  or (_10316_, _10315_, _10314_);
  nor (_10317_, _10316_, _10288_);
  nor (_10318_, _10286_, _10271_);
  nor (_10319_, _10318_, _10317_);
  and (_10320_, _10319_, _10159_);
  nor (_10321_, _10319_, _10159_);
  nor (_10322_, _10214_, _10211_);
  and (_10323_, _10286_, _10322_);
  nor (_10324_, _10286_, \oc8051_golden_model_1.ACC [2]);
  nor (_10325_, _10324_, _10323_);
  and (_10326_, _10325_, _10101_);
  and (_10327_, _06042_, \oc8051_golden_model_1.B [0]);
  not (_10328_, _10327_);
  nor (_10329_, _10325_, _10101_);
  nor (_10330_, _10329_, _10326_);
  and (_10331_, _10330_, _10328_);
  nor (_10332_, _10331_, _10326_);
  nor (_10333_, _10332_, _10321_);
  nor (_10334_, _10333_, _10320_);
  nor (_10335_, _10311_, _10145_);
  nor (_10336_, _10335_, _10312_);
  not (_10337_, _10336_);
  nor (_10338_, _10337_, _10334_);
  nor (_10339_, _10338_, _10312_);
  nor (_10340_, _10339_, _10306_);
  nor (_10341_, _10340_, _10305_);
  nor (_10342_, _10341_, _10297_);
  nor (_10343_, _10342_, _10294_);
  and (_10344_, \oc8051_golden_model_1.ACC [7], _09492_);
  nor (_10345_, _10344_, _10146_);
  nor (_10346_, _10345_, _10343_);
  not (_10347_, _10146_);
  nor (_10348_, _10287_, _10110_);
  nor (_10349_, _10348_, _10347_);
  nor (_10350_, _10349_, _10346_);
  and (_10351_, _10350_, _10287_);
  or (_10352_, _10351_, _10110_);
  nor (_10353_, _10352_, _09492_);
  nor (_10354_, _10352_, \oc8051_golden_model_1.B [7]);
  nor (_10355_, _10354_, _09607_);
  not (_10356_, _10355_);
  not (_10357_, \oc8051_golden_model_1.B [6]);
  and (_10358_, _10341_, _10297_);
  nor (_10359_, _10358_, _10342_);
  nor (_10360_, _10359_, _10350_);
  not (_10361_, _10350_);
  nor (_10362_, _10361_, _10293_);
  nor (_10363_, _10362_, _10360_);
  nor (_10364_, _10363_, _10357_);
  and (_10365_, _10363_, _10357_);
  nor (_10366_, _10306_, _10305_);
  nor (_10367_, _10366_, _10339_);
  and (_10368_, _10366_, _10339_);
  or (_10369_, _10368_, _10367_);
  nor (_10370_, _10369_, _10350_);
  nor (_10371_, _10361_, _10304_);
  nor (_10372_, _10371_, _10370_);
  nor (_10373_, _10372_, _10229_);
  and (_10374_, _10372_, _10229_);
  not (_10375_, _10374_);
  and (_10376_, _10337_, _10334_);
  nor (_10377_, _10376_, _10338_);
  nor (_10378_, _10377_, _10350_);
  nor (_10379_, _10361_, _10311_);
  nor (_10380_, _10379_, _10378_);
  nor (_10381_, _10380_, _10241_);
  and (_10382_, _10350_, _10319_);
  nor (_10383_, _10321_, _10320_);
  and (_10384_, _10383_, _10332_);
  nor (_10385_, _10383_, _10332_);
  nor (_10386_, _10385_, _10384_);
  nor (_10387_, _10386_, _10350_);
  or (_10388_, _10387_, _10382_);
  and (_10389_, _10388_, _10145_);
  nor (_10390_, _10388_, _10145_);
  nor (_10391_, _10390_, _10389_);
  nor (_10392_, _10330_, _10328_);
  nor (_10393_, _10392_, _10331_);
  nor (_10394_, _10393_, _10350_);
  nor (_10395_, _10361_, _10325_);
  nor (_10396_, _10395_, _10394_);
  nor (_10397_, _10396_, _10159_);
  and (_10398_, _10396_, _10159_);
  nor (_10399_, _10398_, _10397_);
  and (_10400_, _10399_, _10391_);
  and (_10401_, _10350_, _06042_);
  nor (_10402_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [0]);
  nor (_10403_, _10402_, _10030_);
  nor (_10404_, _10350_, _10403_);
  nor (_10405_, _10404_, _10401_);
  and (_10406_, _10405_, _10101_);
  nor (_10407_, _10405_, _10101_);
  and (_10408_, _10106_, \oc8051_golden_model_1.ACC [0]);
  not (_10409_, _10408_);
  nor (_10410_, _10409_, _10407_);
  nor (_10411_, _10410_, _10406_);
  and (_10412_, _10411_, _10400_);
  and (_10413_, _10397_, _10391_);
  nor (_10414_, _10413_, _10390_);
  not (_10415_, _10414_);
  nor (_10416_, _10415_, _10412_);
  and (_10417_, _10380_, _10241_);
  nor (_10418_, _10417_, _10416_);
  or (_10419_, _10418_, _10381_);
  and (_10420_, _10419_, _10375_);
  nor (_10421_, _10420_, _10373_);
  nor (_10422_, _10421_, _10365_);
  or (_10423_, _10422_, _10364_);
  and (_10424_, _10423_, _10356_);
  nor (_10425_, _10424_, _10353_);
  nor (_10426_, _10417_, _10381_);
  nor (_10427_, _10374_, _10373_);
  and (_10428_, _10427_, _10426_);
  nor (_10429_, _10365_, _10364_);
  and (_10430_, _10429_, _10356_);
  and (_10431_, _10430_, _10428_);
  nor (_10432_, _10407_, _10406_);
  and (_10433_, \oc8051_golden_model_1.B [0], _06097_);
  not (_10434_, _10433_);
  and (_10435_, _10434_, _10432_);
  and (_10436_, _10435_, _10409_);
  and (_10437_, _10436_, _10400_);
  and (_10438_, _10437_, _10431_);
  nor (_10439_, _10438_, _10425_);
  or (_10440_, _10439_, _10110_);
  and (_10441_, _10440_, _10352_);
  or (_10442_, _10441_, _10100_);
  and (_10443_, _10442_, _10099_);
  and (_10444_, _10443_, _06219_);
  and (_10445_, _08825_, _07942_);
  or (_10446_, _10445_, _09494_);
  and (_10447_, _10446_, _06218_);
  or (_10448_, _10447_, _06369_);
  or (_10449_, _10448_, _10444_);
  and (_10450_, _09044_, _07942_);
  or (_10451_, _10450_, _09494_);
  or (_10452_, _10451_, _07237_);
  and (_10453_, _10452_, _07240_);
  and (_10454_, _10453_, _10449_);
  or (_10455_, _10454_, _09497_);
  and (_10456_, _10455_, _07242_);
  or (_10457_, _09494_, _08043_);
  and (_10458_, _10446_, _06375_);
  and (_10459_, _10458_, _10457_);
  or (_10460_, _10459_, _10456_);
  and (_10461_, _10460_, _07234_);
  and (_10462_, _09511_, _06545_);
  and (_10463_, _10462_, _10457_);
  or (_10464_, _10463_, _06366_);
  or (_10465_, _10464_, _10461_);
  nor (_10466_, _09043_, _09498_);
  or (_10467_, _09494_, _09056_);
  or (_10468_, _10467_, _10466_);
  and (_10469_, _10468_, _09061_);
  and (_10470_, _10469_, _10465_);
  nor (_10471_, _08573_, _09498_);
  or (_10472_, _10471_, _09494_);
  and (_10473_, _10472_, _06528_);
  or (_10474_, _10473_, _06568_);
  or (_10475_, _10474_, _10470_);
  or (_10476_, _09508_, _06926_);
  and (_10477_, _10476_, _05928_);
  and (_10478_, _10477_, _10475_);
  and (_10479_, _09505_, _05927_);
  or (_10480_, _10479_, _06278_);
  or (_10481_, _10480_, _10478_);
  and (_10482_, _08550_, _07942_);
  or (_10483_, _09494_, _06279_);
  or (_10484_, _10483_, _10482_);
  and (_10485_, _10484_, _01347_);
  and (_10486_, _10485_, _10481_);
  or (_10487_, _10486_, _09493_);
  and (_40573_, _10487_, _42618_);
  nor (_10488_, _01347_, _08572_);
  nor (_10489_, _07939_, _08572_);
  not (_10490_, _07939_);
  nor (_10491_, _09043_, _10490_);
  or (_10492_, _10491_, _10489_);
  and (_10493_, _10492_, _06366_);
  and (_10494_, _08040_, _08572_);
  nor (_10495_, _10494_, _07043_);
  and (_10496_, _06370_, _06544_);
  not (_10497_, _10496_);
  nor (_10498_, _08755_, \oc8051_golden_model_1.ACC [7]);
  and (_10499_, _08755_, \oc8051_golden_model_1.ACC [7]);
  nor (_10500_, _10499_, _10498_);
  and (_10501_, _06345_, _06535_);
  nor (_10502_, _10501_, _06884_);
  or (_10503_, _10502_, _10500_);
  nor (_10504_, _08040_, _08572_);
  nor (_10505_, _10504_, _10494_);
  and (_10506_, _07041_, _06535_);
  or (_10507_, _10506_, _06703_);
  nor (_10508_, _10507_, _06887_);
  not (_10509_, _10508_);
  and (_10510_, _10509_, _10505_);
  or (_10511_, _06182_, _05975_);
  nor (_10512_, _08040_, _10490_);
  or (_10513_, _10512_, _10489_);
  or (_10514_, _10513_, _07215_);
  not (_10515_, _05984_);
  and (_10516_, _06370_, _05976_);
  not (_10517_, _10516_);
  and (_10518_, _07949_, \oc8051_golden_model_1.PSW [7]);
  and (_10519_, _10518_, _07908_);
  and (_10520_, _10519_, _07892_);
  and (_10521_, _10520_, _07607_);
  and (_10522_, _10521_, _06286_);
  nor (_10523_, _10521_, _06286_);
  or (_10524_, _10523_, _10522_);
  nor (_10525_, _10524_, _08572_);
  and (_10526_, _10524_, _08572_);
  nor (_10527_, _10526_, _10525_);
  not (_10528_, _10527_);
  nor (_10529_, _10520_, _07607_);
  nor (_10530_, _10529_, _10521_);
  nor (_10531_, _10530_, _10116_);
  and (_10532_, _10519_, _07883_);
  nor (_10533_, _10532_, _07896_);
  nor (_10534_, _10533_, _10520_);
  and (_10535_, _10534_, _10170_);
  nor (_10536_, _10534_, _10170_);
  nor (_10537_, _10519_, _07883_);
  nor (_10538_, _10537_, _10532_);
  nor (_10539_, _10538_, _10135_);
  nor (_10540_, _10539_, _10536_);
  nor (_10541_, _10540_, _10535_);
  nor (_10542_, _10536_, _10535_);
  not (_10543_, _10542_);
  and (_10544_, _10538_, _10135_);
  or (_10545_, _10544_, _10539_);
  or (_10546_, _10545_, _10543_);
  nor (_10547_, _08807_, _06473_);
  nor (_10548_, _10547_, _10519_);
  nor (_10549_, _10548_, _06055_);
  and (_10550_, _10548_, _06055_);
  nor (_10551_, _10550_, _10549_);
  nor (_10552_, _10518_, _06657_);
  nor (_10553_, _10552_, _08807_);
  nor (_10554_, _10553_, _10213_);
  and (_10555_, _10553_, _10213_);
  nor (_10556_, _10555_, _10554_);
  and (_10557_, _10556_, _10551_);
  not (_10558_, \oc8051_golden_model_1.PSW [7]);
  nor (_10559_, _06251_, _10558_);
  nor (_10560_, _10559_, _07005_);
  nor (_10561_, _10560_, _10518_);
  nor (_10562_, _10561_, _06042_);
  and (_10563_, _06251_, _10558_);
  nor (_10564_, _10563_, _10559_);
  and (_10565_, _10564_, _06097_);
  and (_10566_, _10561_, _06042_);
  nor (_10567_, _10562_, _10566_);
  not (_10568_, _10567_);
  nor (_10569_, _10568_, _10565_);
  or (_10570_, _10569_, _10562_);
  and (_10571_, _10570_, _10557_);
  and (_10572_, _10554_, _10551_);
  or (_10573_, _10572_, _10549_);
  nor (_10574_, _10573_, _10571_);
  nor (_10575_, _10574_, _10546_);
  nor (_10576_, _10575_, _10541_);
  and (_10577_, _10530_, _10116_);
  nor (_10578_, _10531_, _10577_);
  not (_10579_, _10578_);
  nor (_10580_, _10579_, _10576_);
  or (_10581_, _10580_, _10531_);
  and (_10582_, _10581_, _10528_);
  nor (_10583_, _10581_, _10528_);
  or (_10584_, _10583_, _10582_);
  or (_10585_, _10584_, _10517_);
  and (_10586_, _06343_, _05976_);
  and (_10587_, _06345_, _05976_);
  nor (_10588_, _10587_, _10586_);
  and (_10589_, _09392_, \oc8051_golden_model_1.PSW [7]);
  and (_10590_, _10589_, _09451_);
  and (_10591_, _10590_, _09450_);
  and (_10592_, _10591_, _09449_);
  and (_10593_, _10592_, _09448_);
  and (_10594_, _10593_, _09447_);
  and (_10595_, _10594_, _09446_);
  nor (_10596_, _10595_, _09076_);
  and (_10597_, _10595_, _09076_);
  nor (_10598_, _10597_, _10596_);
  and (_10599_, _10598_, \oc8051_golden_model_1.ACC [7]);
  nor (_10600_, _10598_, \oc8051_golden_model_1.ACC [7]);
  nor (_10601_, _10600_, _10599_);
  not (_10602_, _10601_);
  nor (_10603_, _10594_, _09446_);
  nor (_10604_, _10603_, _10595_);
  nor (_10605_, _10604_, _10116_);
  nor (_10606_, _10593_, _09447_);
  nor (_10607_, _10606_, _10594_);
  and (_10608_, _10607_, _10170_);
  nor (_10609_, _10607_, _10170_);
  nor (_10610_, _10609_, _10608_);
  not (_10611_, _10610_);
  nor (_10612_, _10592_, _09448_);
  nor (_10613_, _10612_, _10593_);
  nor (_10614_, _10613_, _10135_);
  and (_10615_, _10613_, _10135_);
  or (_10616_, _10615_, _10614_);
  or (_10617_, _10616_, _10611_);
  nor (_10618_, _10591_, _09449_);
  nor (_10619_, _10618_, _10592_);
  nor (_10620_, _10619_, _06055_);
  and (_10621_, _10619_, _06055_);
  nor (_10622_, _10621_, _10620_);
  nor (_10623_, _10590_, _09450_);
  nor (_10624_, _10623_, _10591_);
  nor (_10625_, _10624_, _10213_);
  and (_10626_, _10624_, _10213_);
  nor (_10627_, _10626_, _10625_);
  and (_10628_, _10627_, _10622_);
  nor (_10629_, _10589_, _09451_);
  nor (_10630_, _10629_, _10590_);
  nor (_10631_, _10630_, _06042_);
  and (_10632_, _10630_, _06042_);
  nor (_10633_, _09392_, \oc8051_golden_model_1.PSW [7]);
  nor (_10634_, _10633_, _10589_);
  and (_10635_, _10634_, _06097_);
  nor (_10636_, _10635_, _10632_);
  or (_10637_, _10636_, _10631_);
  and (_10638_, _10637_, _10628_);
  and (_10639_, _10625_, _10622_);
  or (_10640_, _10639_, _10620_);
  nor (_10641_, _10640_, _10638_);
  nor (_10642_, _10641_, _10617_);
  and (_10643_, _10614_, _10610_);
  nor (_10644_, _10643_, _10609_);
  not (_10645_, _10644_);
  nor (_10646_, _10645_, _10642_);
  and (_10647_, _10604_, _10116_);
  nor (_10648_, _10605_, _10647_);
  not (_10649_, _10648_);
  nor (_10650_, _10649_, _10646_);
  or (_10651_, _10650_, _10605_);
  and (_10652_, _10651_, _10602_);
  nor (_10653_, _10651_, _10602_);
  or (_10654_, _10653_, _10652_);
  or (_10655_, _10654_, _10588_);
  not (_10656_, _10588_);
  and (_10657_, _07133_, \oc8051_golden_model_1.PSW [7]);
  and (_10658_, _10657_, _09432_);
  and (_10659_, _10658_, _09431_);
  and (_10661_, _10659_, _07595_);
  and (_10662_, _10661_, _09430_);
  and (_10663_, _10662_, _09429_);
  and (_10664_, _10663_, _09428_);
  and (_10665_, _10664_, _08040_);
  nor (_10666_, _10664_, _08040_);
  or (_10667_, _10666_, _10665_);
  nor (_10668_, _10667_, _08572_);
  and (_10669_, _10667_, _08572_);
  nor (_10670_, _10669_, _10668_);
  not (_10672_, _10670_);
  nor (_10673_, _10663_, _09428_);
  nor (_10674_, _10673_, _10664_);
  nor (_10675_, _10674_, _10116_);
  nor (_10676_, _10662_, _09429_);
  nor (_10677_, _10676_, _10663_);
  and (_10678_, _10677_, _10170_);
  nor (_10679_, _10677_, _10170_);
  nor (_10680_, _10661_, _09430_);
  nor (_10681_, _10680_, _10662_);
  nor (_10683_, _10681_, _10135_);
  nor (_10684_, _10683_, _10679_);
  nor (_10685_, _10684_, _10678_);
  nor (_10686_, _10679_, _10678_);
  not (_10687_, _10686_);
  and (_10688_, _10681_, _10135_);
  or (_10689_, _10688_, _10683_);
  or (_10690_, _10689_, _10687_);
  nor (_10691_, _10659_, _07595_);
  nor (_10692_, _10691_, _10661_);
  nor (_10694_, _10692_, _06055_);
  and (_10695_, _10692_, _06055_);
  nor (_10696_, _10695_, _10694_);
  nor (_10697_, _10658_, _09431_);
  nor (_10698_, _10697_, _10659_);
  nor (_10699_, _10698_, _10213_);
  and (_10700_, _10698_, _10213_);
  nor (_10701_, _10700_, _10699_);
  and (_10702_, _10701_, _10696_);
  nor (_10703_, _10657_, _09432_);
  nor (_10705_, _10703_, _10658_);
  nor (_10706_, _10705_, _06042_);
  and (_10707_, _10705_, _06042_);
  nor (_10708_, _07133_, \oc8051_golden_model_1.PSW [7]);
  nor (_10709_, _10708_, _10657_);
  and (_10710_, _10709_, _06097_);
  nor (_10711_, _10710_, _10707_);
  or (_10712_, _10711_, _10706_);
  nand (_10713_, _10712_, _10702_);
  and (_10714_, _10699_, _10696_);
  nor (_10716_, _10714_, _10694_);
  and (_10717_, _10716_, _10713_);
  nor (_10718_, _10717_, _10690_);
  nor (_10719_, _10718_, _10685_);
  and (_10720_, _10674_, _10116_);
  nor (_10721_, _10675_, _10720_);
  not (_10722_, _10721_);
  nor (_10723_, _10722_, _10719_);
  or (_10724_, _10723_, _10675_);
  and (_10725_, _10724_, _10672_);
  nor (_10727_, _10724_, _10672_);
  or (_10728_, _10727_, _10725_);
  and (_10729_, _07041_, _05976_);
  and (_10730_, _06327_, _05976_);
  nor (_10731_, _10730_, _10729_);
  and (_10732_, _06336_, _05972_);
  and (_10733_, _10732_, _05976_);
  not (_10734_, _10733_);
  and (_10735_, _10734_, _10731_);
  or (_10736_, _10735_, _10728_);
  not (_10737_, _10735_);
  nor (_10738_, _10049_, _10047_);
  nor (_10739_, _10738_, _10050_);
  or (_10740_, _10739_, _09537_);
  not (_10741_, _06700_);
  nor (_10742_, _07794_, _06741_);
  and (_10743_, _10742_, _10741_);
  not (_10744_, _10743_);
  nand (_10745_, _10744_, _08040_);
  nor (_10746_, _08636_, _08572_);
  and (_10747_, _08773_, _08636_);
  or (_10748_, _10747_, _10746_);
  or (_10749_, _10748_, _06273_);
  and (_10750_, _10749_, _07166_);
  not (_10751_, _06784_);
  nor (_10752_, _06345_, _07209_);
  and (_10753_, _10752_, _07212_);
  nor (_10754_, _10753_, _06014_);
  nor (_10755_, _10754_, _10751_);
  not (_10756_, _10755_);
  nand (_10757_, _10756_, _08040_);
  and (_10758_, _06370_, _06706_);
  not (_10759_, _10758_);
  nor (_10760_, _06781_, _08572_);
  and (_10761_, _06781_, _08572_);
  nor (_10762_, _10761_, _10760_);
  nand (_10763_, _10762_, _10755_);
  and (_10764_, _10763_, _10759_);
  and (_10765_, _10764_, _10757_);
  and (_10766_, _10758_, _08755_);
  or (_10767_, _10766_, _10765_);
  not (_10768_, _06015_);
  nor (_10769_, _06341_, _10768_);
  and (_10770_, _10769_, _10767_);
  and (_10771_, _08768_, _07939_);
  or (_10772_, _10771_, _10489_);
  and (_10773_, _10772_, _06341_);
  or (_10774_, _10773_, _10770_);
  and (_10775_, _06370_, _06271_);
  not (_10776_, _10775_);
  and (_10777_, _10776_, _10774_);
  nor (_10778_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.ACC [2]);
  nor (_10779_, _10778_, _06055_);
  and (_10780_, _10779_, \oc8051_golden_model_1.ACC [4]);
  and (_10781_, _10780_, \oc8051_golden_model_1.ACC [5]);
  and (_10782_, _10781_, \oc8051_golden_model_1.ACC [6]);
  and (_10783_, _10782_, \oc8051_golden_model_1.ACC [7]);
  nor (_10784_, _10782_, \oc8051_golden_model_1.ACC [7]);
  nor (_10785_, _10784_, _10783_);
  nor (_10786_, _10780_, \oc8051_golden_model_1.ACC [5]);
  nor (_10787_, _10786_, _10781_);
  nor (_10788_, _10781_, \oc8051_golden_model_1.ACC [6]);
  nor (_10789_, _10788_, _10782_);
  nor (_10790_, _10789_, _10787_);
  not (_10791_, _10790_);
  and (_10792_, _10791_, _10785_);
  not (_10793_, _10792_);
  nor (_10794_, _10783_, \oc8051_golden_model_1.PSW [7]);
  and (_10795_, _10794_, _10793_);
  nor (_10796_, _10795_, _10790_);
  or (_10797_, _10796_, _10785_);
  and (_10798_, _10793_, _10775_);
  and (_10799_, _10798_, _10797_);
  or (_10800_, _10799_, _06272_);
  or (_10801_, _10800_, _10777_);
  and (_10802_, _10801_, _10750_);
  and (_10803_, _10513_, _06461_);
  or (_10804_, _10803_, _10744_);
  or (_10805_, _10804_, _10802_);
  and (_10806_, _10805_, _10745_);
  or (_10807_, _10806_, _07174_);
  or (_10808_, _08755_, _07175_);
  and (_10809_, _10808_, _06465_);
  and (_10810_, _10809_, _10807_);
  and (_10811_, _06370_, _06266_);
  nor (_10812_, _08042_, _06465_);
  or (_10813_, _10812_, _10811_);
  or (_10814_, _10813_, _10810_);
  nand (_10815_, _10811_, _06055_);
  and (_10816_, _10815_, _10814_);
  or (_10817_, _10816_, _06268_);
  and (_10818_, _08649_, _08636_);
  or (_10819_, _10818_, _10746_);
  or (_10820_, _10819_, _06269_);
  and (_10821_, _10820_, _06262_);
  and (_10822_, _10821_, _10817_);
  or (_10823_, _10746_, _08789_);
  and (_10824_, _10823_, _06261_);
  and (_10825_, _10824_, _10748_);
  or (_10826_, _10825_, _09531_);
  or (_10827_, _10826_, _10822_);
  and (_10828_, _10827_, _10740_);
  or (_10829_, _10828_, _10737_);
  and (_10830_, _10829_, _10736_);
  or (_10831_, _10830_, _10656_);
  and (_10832_, _10831_, _06517_);
  and (_10833_, _10832_, _10655_);
  and (_10834_, _08390_, \oc8051_golden_model_1.PSW [7]);
  and (_10835_, _10834_, _08341_);
  and (_10836_, _10835_, _08440_);
  and (_10837_, _10836_, _08292_);
  and (_10838_, _10837_, _08544_);
  and (_10839_, _10838_, _08247_);
  and (_10840_, _10839_, _08145_);
  nor (_10841_, _10840_, _08042_);
  and (_10842_, _10840_, _08042_);
  nor (_10843_, _10842_, _10841_);
  and (_10844_, _10843_, \oc8051_golden_model_1.ACC [7]);
  nor (_10845_, _10843_, \oc8051_golden_model_1.ACC [7]);
  nor (_10846_, _10845_, _10844_);
  not (_10847_, _10846_);
  nor (_10848_, _10839_, _08145_);
  nor (_10849_, _10848_, _10840_);
  nor (_10850_, _10849_, _10116_);
  nor (_10851_, _10838_, _08247_);
  nor (_10852_, _10851_, _10839_);
  and (_10853_, _10852_, _10170_);
  nor (_10854_, _10852_, _10170_);
  nor (_10855_, _10837_, _08544_);
  nor (_10856_, _10855_, _10838_);
  nor (_10857_, _10856_, _10135_);
  nor (_10858_, _10857_, _10854_);
  nor (_10859_, _10858_, _10853_);
  nor (_10860_, _10854_, _10853_);
  not (_10861_, _10860_);
  and (_10862_, _10856_, _10135_);
  or (_10863_, _10862_, _10857_);
  or (_10864_, _10863_, _10861_);
  nor (_10865_, _10836_, _08292_);
  nor (_10866_, _10865_, _10837_);
  nor (_10867_, _10866_, _06055_);
  and (_10868_, _10866_, _06055_);
  nor (_10869_, _10868_, _10867_);
  nor (_10870_, _10835_, _08440_);
  nor (_10871_, _10870_, _10836_);
  nor (_10872_, _10871_, _10213_);
  and (_10873_, _10871_, _10213_);
  nor (_10874_, _10873_, _10872_);
  and (_10875_, _10874_, _10869_);
  nor (_10876_, _10834_, _08341_);
  nor (_10877_, _10876_, _10835_);
  nor (_10878_, _10877_, _06042_);
  and (_10879_, _10877_, _06042_);
  nor (_10880_, _08390_, \oc8051_golden_model_1.PSW [7]);
  nor (_10881_, _10880_, _10834_);
  and (_10882_, _10881_, _06097_);
  nor (_10883_, _10882_, _10879_);
  or (_10884_, _10883_, _10878_);
  nand (_10885_, _10884_, _10875_);
  and (_10886_, _10872_, _10869_);
  nor (_10887_, _10886_, _10867_);
  and (_10888_, _10887_, _10885_);
  nor (_10889_, _10888_, _10864_);
  nor (_10890_, _10889_, _10859_);
  and (_10891_, _10849_, _10116_);
  nor (_10892_, _10850_, _10891_);
  not (_10893_, _10892_);
  nor (_10894_, _10893_, _10890_);
  or (_10895_, _10894_, _10850_);
  and (_10896_, _10895_, _10847_);
  nor (_10897_, _10895_, _10847_);
  or (_10898_, _10897_, _10896_);
  and (_10899_, _10898_, _06512_);
  or (_10900_, _10899_, _10516_);
  or (_10901_, _10900_, _10833_);
  and (_10902_, _10901_, _10585_);
  or (_10903_, _10902_, _10515_);
  or (_10904_, _06182_, _05984_);
  and (_10905_, _10904_, _06258_);
  and (_10906_, _10905_, _10903_);
  and (_10907_, _08808_, _08636_);
  or (_10908_, _10907_, _10746_);
  and (_10909_, _10908_, _06257_);
  or (_10910_, _10909_, _10080_);
  or (_10911_, _10910_, _10906_);
  and (_10912_, _10911_, _10514_);
  or (_10913_, _10912_, _07460_);
  and (_10914_, _08755_, _07939_);
  or (_10915_, _10489_, _07208_);
  or (_10916_, _10915_, _10914_);
  and (_10917_, _10916_, _05982_);
  and (_10918_, _10917_, _10913_);
  and (_10919_, _09021_, _07939_);
  or (_10920_, _10919_, _10489_);
  and (_10921_, _10920_, _10094_);
  or (_10922_, _10921_, _10093_);
  or (_10923_, _10922_, _10918_);
  or (_10924_, _10114_, _10100_);
  and (_10925_, _10924_, _10923_);
  or (_10926_, _10925_, _05974_);
  and (_10927_, _10926_, _10511_);
  or (_10928_, _10927_, _06218_);
  and (_10929_, _06370_, _06321_);
  not (_10930_, _10929_);
  and (_10931_, _08825_, _07939_);
  nor (_10932_, _10931_, _10489_);
  nand (_10933_, _10932_, _06218_);
  and (_10934_, _10933_, _10930_);
  and (_10935_, _10934_, _10928_);
  and (_10936_, _10929_, _06182_);
  nor (_10937_, _07211_, _05954_);
  or (_10938_, _10937_, _10936_);
  or (_10939_, _10938_, _10935_);
  not (_10940_, _10937_);
  or (_10941_, _10940_, _10505_);
  and (_10942_, _10941_, _10508_);
  and (_10943_, _10942_, _10939_);
  or (_10944_, _10943_, _10510_);
  and (_10945_, _07209_, _06535_);
  not (_10946_, _10945_);
  and (_10947_, _10946_, _10944_);
  not (_10948_, _10502_);
  and (_10949_, _10945_, _10505_);
  or (_10950_, _10949_, _10948_);
  or (_10951_, _10950_, _10947_);
  and (_10952_, _10951_, _10503_);
  or (_10953_, _10952_, _06533_);
  and (_10954_, _06370_, _06535_);
  not (_10955_, _10954_);
  or (_10956_, _08575_, _06534_);
  and (_10957_, _10956_, _10955_);
  nand (_10958_, _10957_, _10953_);
  nor (_10959_, _06182_, \oc8051_golden_model_1.ACC [7]);
  and (_10960_, _06182_, \oc8051_golden_model_1.ACC [7]);
  nor (_10961_, _10960_, _10959_);
  nand (_10962_, _10954_, _10961_);
  and (_10963_, _10962_, _07237_);
  and (_10964_, _10963_, _10958_);
  and (_10965_, _09044_, _07939_);
  nor (_10966_, _10965_, _10489_);
  and (_10967_, _10966_, _06369_);
  or (_10968_, _10967_, _10964_);
  and (_10969_, _10968_, _07240_);
  nor (_10970_, _10489_, _07240_);
  nor (_10971_, _07482_, _05960_);
  not (_10972_, _10971_);
  and (_10973_, _06886_, _06544_);
  and (_10974_, _07041_, _06544_);
  nor (_10975_, _10974_, _10973_);
  and (_10976_, _06327_, _06544_);
  not (_10977_, _10976_);
  and (_10978_, _10977_, _10975_);
  and (_10979_, _10978_, _10972_);
  not (_10980_, _10979_);
  or (_10981_, _10980_, _10970_);
  or (_10982_, _10981_, _10969_);
  nor (_10983_, _07153_, _05960_);
  nand (_10984_, _10983_, _10499_);
  and (_10985_, _06336_, _06544_);
  nor (_10986_, _10985_, _10976_);
  not (_10987_, _10986_);
  nand (_10988_, _10987_, _10504_);
  and (_10989_, _10988_, _06543_);
  and (_10990_, _10989_, _10984_);
  and (_10991_, _10990_, _10982_);
  nor (_10992_, _08574_, _06543_);
  or (_10993_, _10992_, _10991_);
  and (_10994_, _10993_, _10497_);
  nor (_10995_, _10960_, _10497_);
  or (_10996_, _10995_, _06375_);
  nor (_10997_, _10996_, _10994_);
  nor (_10998_, _06755_, _06711_);
  not (_10999_, _10998_);
  or (_11000_, _10932_, _07242_);
  nor (_11001_, _11000_, _08573_);
  or (_11002_, _11001_, _10999_);
  or (_11003_, _11002_, _10997_);
  nand (_11004_, _10999_, _10494_);
  and (_11005_, _11004_, _07043_);
  and (_11006_, _11005_, _11003_);
  or (_11007_, _11006_, _10495_);
  and (_11008_, _07209_, _06527_);
  not (_11009_, _11008_);
  and (_11010_, _11009_, _11007_);
  and (_11011_, _06343_, _06527_);
  and (_11012_, _06345_, _06527_);
  nor (_11013_, _11012_, _11011_);
  not (_11014_, _11013_);
  nor (_11015_, _11009_, _10494_);
  or (_11016_, _11015_, _11014_);
  or (_11017_, _11016_, _11010_);
  nand (_11018_, _11014_, _10498_);
  and (_11019_, _11018_, _06531_);
  and (_11020_, _11019_, _11017_);
  and (_11021_, _06370_, _06527_);
  nor (_11022_, _11021_, _06530_);
  not (_11023_, _11022_);
  not (_11024_, _11021_);
  nand (_11025_, _11024_, _08573_);
  and (_11026_, _11025_, _11023_);
  or (_11027_, _11026_, _11020_);
  nand (_11028_, _11021_, _10959_);
  and (_11029_, _11028_, _09056_);
  and (_11030_, _11029_, _11027_);
  or (_11031_, _11030_, _10493_);
  nor (_11032_, _07041_, _06353_);
  nor (_11033_, _11032_, _05958_);
  nor (_11034_, _07211_, _05958_);
  or (_11035_, _11034_, _11033_);
  and (_11036_, _10732_, _06364_);
  nor (_11037_, _11036_, _11035_);
  and (_11038_, _11037_, _11031_);
  and (_11039_, _06343_, _06364_);
  and (_11040_, _06345_, _06364_);
  or (_11041_, _11040_, _11039_);
  and (_11042_, _10674_, \oc8051_golden_model_1.ACC [6]);
  and (_11043_, _10677_, \oc8051_golden_model_1.ACC [5]);
  nand (_11044_, _10681_, \oc8051_golden_model_1.ACC [4]);
  and (_11045_, _10692_, \oc8051_golden_model_1.ACC [3]);
  and (_11046_, _10698_, \oc8051_golden_model_1.ACC [2]);
  and (_11047_, _10705_, \oc8051_golden_model_1.ACC [1]);
  nor (_11048_, _10707_, _10706_);
  not (_11049_, _11048_);
  and (_11050_, _10709_, \oc8051_golden_model_1.ACC [0]);
  and (_11051_, _11050_, _11049_);
  nor (_11052_, _11051_, _11047_);
  nor (_11053_, _11052_, _10701_);
  nor (_11054_, _11053_, _11046_);
  nor (_11055_, _11054_, _10696_);
  or (_11056_, _11055_, _11045_);
  nand (_11057_, _11056_, _10689_);
  and (_11058_, _11057_, _11044_);
  nor (_11059_, _11058_, _10686_);
  or (_11060_, _11059_, _11043_);
  and (_11061_, _11060_, _10722_);
  nor (_11062_, _11061_, _11042_);
  and (_11063_, _11062_, _10670_);
  nor (_11064_, _11062_, _10670_);
  or (_11065_, _11064_, _11037_);
  nor (_11066_, _11065_, _11063_);
  or (_11067_, _11066_, _11041_);
  or (_11068_, _11067_, _11038_);
  not (_11069_, _11041_);
  nand (_11070_, _10604_, \oc8051_golden_model_1.ACC [6]);
  and (_11071_, _10607_, \oc8051_golden_model_1.ACC [5]);
  nand (_11072_, _10613_, \oc8051_golden_model_1.ACC [4]);
  and (_11073_, _10619_, \oc8051_golden_model_1.ACC [3]);
  and (_11074_, _10624_, \oc8051_golden_model_1.ACC [2]);
  and (_11075_, _10630_, \oc8051_golden_model_1.ACC [1]);
  nor (_11076_, _10632_, _10631_);
  not (_11077_, _11076_);
  and (_11078_, _10634_, \oc8051_golden_model_1.ACC [0]);
  and (_11079_, _11078_, _11077_);
  nor (_11080_, _11079_, _11075_);
  nor (_11081_, _11080_, _10627_);
  nor (_11082_, _11081_, _11074_);
  nor (_11083_, _11082_, _10622_);
  or (_11084_, _11083_, _11073_);
  nand (_11085_, _11084_, _10616_);
  and (_11086_, _11085_, _11072_);
  nor (_11087_, _11086_, _10610_);
  or (_11088_, _11087_, _11071_);
  nand (_11089_, _11088_, _10649_);
  and (_11090_, _11089_, _11070_);
  nor (_11091_, _11090_, _10601_);
  and (_11092_, _11090_, _10601_);
  nor (_11093_, _11092_, _11091_);
  or (_11094_, _11093_, _11069_);
  and (_11095_, _11094_, _06541_);
  and (_11096_, _11095_, _11068_);
  and (_11097_, _06370_, _06364_);
  nand (_11098_, _10849_, \oc8051_golden_model_1.ACC [6]);
  and (_11099_, _10852_, \oc8051_golden_model_1.ACC [5]);
  nand (_11100_, _10856_, \oc8051_golden_model_1.ACC [4]);
  and (_11101_, _10866_, \oc8051_golden_model_1.ACC [3]);
  and (_11102_, _10871_, \oc8051_golden_model_1.ACC [2]);
  and (_11103_, _10877_, \oc8051_golden_model_1.ACC [1]);
  nor (_11104_, _10879_, _10878_);
  not (_11105_, _11104_);
  and (_11106_, _10881_, \oc8051_golden_model_1.ACC [0]);
  and (_11107_, _11106_, _11105_);
  nor (_11108_, _11107_, _11103_);
  nor (_11109_, _11108_, _10874_);
  nor (_11110_, _11109_, _11102_);
  nor (_11111_, _11110_, _10869_);
  or (_11112_, _11111_, _11101_);
  nand (_11113_, _11112_, _10863_);
  and (_11114_, _11113_, _11100_);
  nor (_11115_, _11114_, _10860_);
  or (_11116_, _11115_, _11099_);
  nand (_11117_, _11116_, _10893_);
  and (_11118_, _11117_, _11098_);
  nor (_11119_, _11118_, _10846_);
  and (_11120_, _11118_, _10846_);
  nor (_11121_, _11120_, _11119_);
  and (_11122_, _11121_, _06540_);
  or (_11123_, _11122_, _11097_);
  or (_11124_, _11123_, _11096_);
  nor (_11125_, _05973_, _05958_);
  not (_11126_, _11125_);
  not (_11127_, _11097_);
  and (_11128_, _10530_, \oc8051_golden_model_1.ACC [6]);
  and (_11129_, _10534_, \oc8051_golden_model_1.ACC [5]);
  nand (_11130_, _10538_, \oc8051_golden_model_1.ACC [4]);
  and (_11131_, _10548_, \oc8051_golden_model_1.ACC [3]);
  and (_11132_, _10553_, \oc8051_golden_model_1.ACC [2]);
  and (_11133_, _10561_, \oc8051_golden_model_1.ACC [1]);
  and (_11134_, _10564_, \oc8051_golden_model_1.ACC [0]);
  and (_11135_, _11134_, _10568_);
  nor (_11136_, _11135_, _11133_);
  nor (_11137_, _11136_, _10556_);
  nor (_11138_, _11137_, _11132_);
  nor (_11139_, _11138_, _10551_);
  or (_11140_, _11139_, _11131_);
  nand (_11141_, _11140_, _10545_);
  and (_11142_, _11141_, _11130_);
  nor (_11143_, _11142_, _10542_);
  or (_11144_, _11143_, _11129_);
  and (_11145_, _11144_, _10579_);
  nor (_11146_, _11145_, _11128_);
  nor (_11147_, _11146_, _10527_);
  and (_11148_, _11146_, _10527_);
  nor (_11149_, _11148_, _11147_);
  or (_11150_, _11149_, _11127_);
  and (_11151_, _11150_, _11126_);
  and (_11152_, _11151_, _11124_);
  nand (_11153_, _11125_, \oc8051_golden_model_1.ACC [6]);
  and (_11154_, _07209_, _06280_);
  and (_11155_, _06327_, _06280_);
  or (_11156_, _11155_, _07045_);
  nor (_11157_, _11156_, _11154_);
  nand (_11158_, _11157_, _11153_);
  or (_11159_, _11158_, _11152_);
  nor (_11160_, _08142_, _10116_);
  not (_11161_, _11160_);
  nand (_11162_, _08142_, _10116_);
  and (_11163_, _11162_, _11161_);
  nor (_11164_, _08244_, _10170_);
  and (_11165_, _08244_, _10170_);
  nor (_11166_, _11165_, _11164_);
  nor (_11167_, _08541_, _10135_);
  not (_11168_, _11167_);
  nand (_11169_, _08541_, _10135_);
  and (_11170_, _11169_, _11168_);
  nor (_11171_, _07594_, _06055_);
  and (_11172_, _07594_, _06055_);
  nor (_11173_, _07776_, _10213_);
  and (_11174_, _07776_, _10213_);
  nor (_11175_, _11174_, _11173_);
  nor (_11176_, _07357_, _06042_);
  and (_11177_, _07357_, _06042_);
  nor (_11178_, _11177_, _11176_);
  and (_11179_, _07133_, \oc8051_golden_model_1.ACC [0]);
  and (_11180_, _11179_, _11178_);
  nor (_11181_, _11180_, _11176_);
  not (_11182_, _11181_);
  and (_11183_, _11182_, _11175_);
  nor (_11184_, _11183_, _11173_);
  nor (_11185_, _11184_, _11172_);
  or (_11186_, _11185_, _11171_);
  and (_11187_, _11186_, _11170_);
  nor (_11188_, _11187_, _11167_);
  not (_11189_, _11188_);
  and (_11190_, _11189_, _11166_);
  or (_11191_, _11190_, _11164_);
  and (_11192_, _11191_, _11163_);
  nor (_11193_, _11192_, _11160_);
  and (_11194_, _11193_, _10505_);
  nor (_11195_, _11193_, _10505_);
  or (_11196_, _11195_, _11194_);
  or (_11197_, _11196_, _11157_);
  and (_11198_, _11197_, _11159_);
  and (_11199_, _06343_, _06280_);
  and (_11200_, _06345_, _06280_);
  or (_11201_, _11200_, _11199_);
  or (_11202_, _11201_, _11198_);
  not (_11203_, _11201_);
  and (_11204_, _09446_, \oc8051_golden_model_1.ACC [6]);
  or (_11205_, _09446_, \oc8051_golden_model_1.ACC [6]);
  not (_11206_, _11204_);
  and (_11207_, _11206_, _11205_);
  and (_11208_, _09447_, \oc8051_golden_model_1.ACC [5]);
  and (_11209_, _09167_, _10170_);
  or (_11210_, _11209_, _11208_);
  and (_11211_, _09448_, \oc8051_golden_model_1.ACC [4]);
  not (_11212_, _11211_);
  or (_11213_, _09448_, \oc8051_golden_model_1.ACC [4]);
  and (_11214_, _11212_, _11213_);
  and (_11215_, _09449_, \oc8051_golden_model_1.ACC [3]);
  and (_11216_, _09257_, _06055_);
  and (_11217_, _09450_, \oc8051_golden_model_1.ACC [2]);
  and (_11218_, _09302_, _10213_);
  nor (_11219_, _11217_, _11218_);
  and (_11220_, _09451_, \oc8051_golden_model_1.ACC [1]);
  and (_11221_, _09347_, _06042_);
  nor (_11222_, _11220_, _11221_);
  and (_11223_, _09392_, \oc8051_golden_model_1.ACC [0]);
  and (_11224_, _11223_, _11222_);
  nor (_11225_, _11224_, _11220_);
  not (_11226_, _11225_);
  and (_11227_, _11226_, _11219_);
  nor (_11228_, _11227_, _11217_);
  nor (_11229_, _11228_, _11216_);
  or (_11230_, _11229_, _11215_);
  nand (_11231_, _11230_, _11214_);
  and (_11232_, _11231_, _11212_);
  nor (_11233_, _11232_, _11210_);
  or (_11234_, _11233_, _11208_);
  and (_11235_, _11234_, _11207_);
  nor (_11236_, _11235_, _11204_);
  and (_11237_, _11236_, _10500_);
  nor (_11238_, _11236_, _10500_);
  or (_11239_, _11238_, _11237_);
  or (_11240_, _11239_, _11203_);
  and (_11241_, _11240_, _06285_);
  and (_11242_, _11241_, _11202_);
  and (_11243_, _06370_, _06280_);
  nor (_11244_, _08144_, _10116_);
  not (_11245_, _11244_);
  and (_11246_, _08144_, _10116_);
  nor (_11247_, _11246_, _11244_);
  nor (_11248_, _08246_, _10170_);
  and (_11249_, _08246_, _10170_);
  nor (_11250_, _11249_, _11248_);
  nor (_11251_, _08543_, _10135_);
  not (_11252_, _11251_);
  and (_11253_, _08543_, _10135_);
  nor (_11254_, _11253_, _11251_);
  nor (_11255_, _08291_, _06055_);
  and (_11256_, _08291_, _06055_);
  nor (_11257_, _08439_, _10213_);
  and (_11258_, _08439_, _10213_);
  nor (_11259_, _11258_, _11257_);
  nor (_11260_, _08340_, _06042_);
  and (_11261_, _08340_, _06042_);
  nor (_11262_, _11261_, _11260_);
  and (_11263_, _08390_, \oc8051_golden_model_1.ACC [0]);
  and (_11264_, _11263_, _11262_);
  nor (_11265_, _11264_, _11260_);
  not (_11266_, _11265_);
  and (_11267_, _11266_, _11259_);
  nor (_11268_, _11267_, _11257_);
  nor (_11269_, _11268_, _11256_);
  or (_11270_, _11269_, _11255_);
  nand (_11271_, _11270_, _11254_);
  and (_11272_, _11271_, _11252_);
  not (_11273_, _11272_);
  and (_11274_, _11273_, _11250_);
  or (_11275_, _11274_, _11248_);
  nand (_11276_, _11275_, _11247_);
  and (_11277_, _11276_, _11245_);
  nor (_11278_, _11277_, _08575_);
  and (_11279_, _11277_, _08575_);
  or (_11280_, _11279_, _11278_);
  and (_11281_, _11280_, _06283_);
  or (_11282_, _11281_, _11243_);
  or (_11283_, _11282_, _11242_);
  nor (_11284_, _05973_, _05963_);
  not (_11285_, _11284_);
  nor (_11286_, _06317_, _10116_);
  not (_11287_, _11286_);
  and (_11288_, _06317_, _10116_);
  nor (_11289_, _11286_, _11288_);
  nor (_11290_, _06611_, _10170_);
  and (_11291_, _06611_, _10170_);
  nor (_11292_, _06968_, _10135_);
  not (_11293_, _11292_);
  and (_11294_, _06968_, _10135_);
  nor (_11295_, _11292_, _11294_);
  nor (_11296_, _06213_, _06055_);
  and (_11297_, _06213_, _06055_);
  nor (_11298_, _06656_, _10213_);
  and (_11299_, _06656_, _10213_);
  nor (_11300_, _11298_, _11299_);
  nor (_11301_, _07004_, _06042_);
  nor (_11302_, _06251_, _06097_);
  and (_11303_, _07004_, \oc8051_golden_model_1.ACC [1]);
  nor (_11304_, _07004_, \oc8051_golden_model_1.ACC [1]);
  nor (_11305_, _11304_, _11303_);
  not (_11306_, _11305_);
  and (_11307_, _11306_, _11302_);
  nor (_11308_, _11307_, _11301_);
  not (_11309_, _11308_);
  and (_11310_, _11309_, _11300_);
  nor (_11311_, _11310_, _11298_);
  nor (_11312_, _11311_, _11297_);
  or (_11313_, _11312_, _11296_);
  nand (_11314_, _11313_, _11295_);
  and (_11315_, _11314_, _11293_);
  nor (_11316_, _11315_, _11291_);
  or (_11317_, _11316_, _11290_);
  nand (_11318_, _11317_, _11289_);
  and (_11319_, _11318_, _11287_);
  and (_11320_, _11319_, _10961_);
  not (_11321_, _11243_);
  nor (_11322_, _11319_, _10961_);
  or (_11323_, _11322_, _11321_);
  or (_11324_, _11323_, _11320_);
  and (_11325_, _11324_, _11285_);
  and (_11326_, _11325_, _11283_);
  and (_11327_, _11284_, \oc8051_golden_model_1.ACC [6]);
  or (_11328_, _11327_, _06568_);
  or (_11329_, _11328_, _11326_);
  and (_11330_, _06370_, _05779_);
  not (_11331_, _11330_);
  or (_11332_, _10772_, _06926_);
  and (_11333_, _11332_, _11331_);
  and (_11334_, _11333_, _11329_);
  nor (_11335_, _05973_, _06567_);
  and (_11336_, _10778_, _06097_);
  and (_11337_, _11336_, _06055_);
  and (_11338_, _11337_, _10135_);
  and (_11339_, _11338_, _10170_);
  and (_11340_, _11339_, _10116_);
  nor (_11341_, _11340_, _08572_);
  and (_11342_, _11340_, _08572_);
  or (_11343_, _11342_, _11341_);
  and (_11344_, _11343_, _11330_);
  or (_11345_, _11344_, _11335_);
  or (_11346_, _11345_, _11334_);
  nand (_11347_, _11335_, _10558_);
  and (_11348_, _11347_, _05928_);
  and (_11349_, _11348_, _11346_);
  and (_11350_, _10819_, _05927_);
  or (_11351_, _11350_, _06278_);
  or (_11352_, _11351_, _11349_);
  and (_11353_, _06370_, _05938_);
  not (_11354_, _11353_);
  and (_11355_, _08550_, _07939_);
  or (_11356_, _11355_, _10489_);
  or (_11357_, _11356_, _06279_);
  and (_11358_, _11357_, _11354_);
  and (_11359_, _11358_, _11352_);
  nor (_11360_, _05973_, _06277_);
  and (_11361_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.ACC [0]);
  and (_11362_, _11361_, \oc8051_golden_model_1.ACC [2]);
  and (_11363_, _11362_, \oc8051_golden_model_1.ACC [3]);
  and (_11364_, _11363_, \oc8051_golden_model_1.ACC [4]);
  and (_11365_, _11364_, \oc8051_golden_model_1.ACC [5]);
  and (_11366_, _11365_, \oc8051_golden_model_1.ACC [6]);
  nor (_11367_, _11366_, _08572_);
  and (_11368_, _11366_, _08572_);
  or (_11369_, _11368_, _11367_);
  and (_11370_, _11369_, _11353_);
  or (_11371_, _11370_, _11360_);
  or (_11372_, _11371_, _11359_);
  nand (_11373_, _11360_, _06097_);
  and (_11374_, _11373_, _01347_);
  and (_11375_, _11374_, _11372_);
  or (_11376_, _11375_, _10488_);
  and (_40574_, _11376_, _42618_);
  not (_11377_, \oc8051_golden_model_1.PCON [7]);
  nor (_11378_, _01347_, _11377_);
  nor (_11379_, _07951_, _11377_);
  not (_11380_, _07951_);
  nor (_11381_, _08573_, _11380_);
  or (_11382_, _11381_, _11379_);
  and (_11383_, _11382_, _06528_);
  and (_11384_, _08575_, _07951_);
  or (_11385_, _11384_, _11379_);
  and (_11386_, _11385_, _06536_);
  and (_11387_, _08768_, _07951_);
  or (_11388_, _11387_, _11379_);
  or (_11389_, _11388_, _07151_);
  and (_11390_, _07951_, \oc8051_golden_model_1.ACC [7]);
  or (_11391_, _11390_, _11379_);
  and (_11392_, _11391_, _07141_);
  nor (_11393_, _07141_, _11377_);
  or (_11394_, _11393_, _06341_);
  or (_11395_, _11394_, _11392_);
  and (_11396_, _11395_, _07166_);
  and (_11397_, _11396_, _11389_);
  nor (_11398_, _08040_, _11380_);
  or (_11399_, _11398_, _11379_);
  and (_11400_, _11399_, _06461_);
  or (_11401_, _11400_, _11397_);
  and (_11402_, _11401_, _06465_);
  and (_11403_, _11391_, _06464_);
  or (_11404_, _11403_, _10080_);
  or (_11405_, _11404_, _11402_);
  or (_11406_, _11399_, _07215_);
  and (_11407_, _11406_, _11405_);
  or (_11408_, _11407_, _07460_);
  and (_11409_, _08755_, _07951_);
  or (_11410_, _11379_, _07208_);
  or (_11411_, _11410_, _11409_);
  and (_11412_, _11411_, _05982_);
  and (_11413_, _11412_, _11408_);
  and (_11414_, _09021_, _07951_);
  or (_11415_, _11414_, _11379_);
  and (_11416_, _11415_, _10094_);
  or (_11417_, _11416_, _06218_);
  or (_11418_, _11417_, _11413_);
  and (_11419_, _08825_, _07951_);
  or (_11420_, _11419_, _11379_);
  or (_11421_, _11420_, _06219_);
  and (_11422_, _11421_, _11418_);
  or (_11423_, _11422_, _06369_);
  and (_11424_, _09044_, _07951_);
  or (_11425_, _11424_, _11379_);
  or (_11426_, _11425_, _07237_);
  and (_11427_, _11426_, _07240_);
  and (_11428_, _11427_, _11423_);
  or (_11429_, _11428_, _11386_);
  and (_11430_, _11429_, _07242_);
  or (_11431_, _11379_, _08043_);
  and (_11432_, _11420_, _06375_);
  and (_11433_, _11432_, _11431_);
  or (_11434_, _11433_, _11430_);
  and (_11435_, _11434_, _07234_);
  and (_11436_, _11391_, _06545_);
  and (_11437_, _11436_, _11431_);
  or (_11438_, _11437_, _06366_);
  or (_11439_, _11438_, _11435_);
  nor (_11440_, _09043_, _11380_);
  or (_11441_, _11379_, _09056_);
  or (_11442_, _11441_, _11440_);
  and (_11443_, _11442_, _09061_);
  and (_11444_, _11443_, _11439_);
  or (_11445_, _11444_, _11383_);
  and (_11446_, _11445_, _06926_);
  and (_11447_, _11388_, _06568_);
  or (_11448_, _11447_, _06278_);
  or (_11449_, _11448_, _11446_);
  and (_11450_, _08550_, _07951_);
  or (_11451_, _11379_, _06279_);
  or (_11452_, _11451_, _11450_);
  and (_11453_, _11452_, _01347_);
  and (_11454_, _11453_, _11449_);
  or (_11455_, _11454_, _11378_);
  and (_40575_, _11455_, _42618_);
  and (_11456_, _01351_, \oc8051_golden_model_1.TMOD [7]);
  not (_11457_, _07914_);
  and (_11458_, _11457_, \oc8051_golden_model_1.TMOD [7]);
  nor (_11459_, _08573_, _11457_);
  or (_11460_, _11459_, _11458_);
  and (_11461_, _11460_, _06528_);
  and (_11462_, _08575_, _07914_);
  or (_11463_, _11462_, _11458_);
  and (_11464_, _11463_, _06536_);
  and (_11465_, _08768_, _07914_);
  or (_11466_, _11465_, _11458_);
  or (_11467_, _11466_, _07151_);
  and (_11468_, _07914_, \oc8051_golden_model_1.ACC [7]);
  or (_11469_, _11468_, _11458_);
  and (_11470_, _11469_, _07141_);
  and (_11471_, _07142_, \oc8051_golden_model_1.TMOD [7]);
  or (_11472_, _11471_, _06341_);
  or (_11473_, _11472_, _11470_);
  and (_11474_, _11473_, _07166_);
  and (_11475_, _11474_, _11467_);
  nor (_11476_, _08040_, _11457_);
  or (_11477_, _11476_, _11458_);
  and (_11478_, _11477_, _06461_);
  or (_11479_, _11478_, _11475_);
  and (_11480_, _11479_, _06465_);
  and (_11481_, _11469_, _06464_);
  or (_11482_, _11481_, _10080_);
  or (_11483_, _11482_, _11480_);
  or (_11484_, _11477_, _07215_);
  and (_11485_, _11484_, _11483_);
  or (_11486_, _11485_, _07460_);
  and (_11487_, _08755_, _07914_);
  or (_11488_, _11458_, _07208_);
  or (_11489_, _11488_, _11487_);
  and (_11490_, _11489_, _05982_);
  and (_11491_, _11490_, _11486_);
  and (_11492_, _09021_, _07914_);
  or (_11493_, _11492_, _11458_);
  and (_11494_, _11493_, _10094_);
  or (_11495_, _11494_, _06218_);
  or (_11496_, _11495_, _11491_);
  and (_11497_, _08825_, _07914_);
  or (_11498_, _11497_, _11458_);
  or (_11499_, _11498_, _06219_);
  and (_11500_, _11499_, _11496_);
  or (_11501_, _11500_, _06369_);
  and (_11502_, _09044_, _07914_);
  or (_11503_, _11502_, _11458_);
  or (_11504_, _11503_, _07237_);
  and (_11505_, _11504_, _07240_);
  and (_11506_, _11505_, _11501_);
  or (_11507_, _11506_, _11464_);
  and (_11508_, _11507_, _07242_);
  or (_11509_, _11458_, _08043_);
  and (_11510_, _11498_, _06375_);
  and (_11511_, _11510_, _11509_);
  or (_11512_, _11511_, _11508_);
  and (_11513_, _11512_, _07234_);
  and (_11514_, _11469_, _06545_);
  and (_11515_, _11514_, _11509_);
  or (_11516_, _11515_, _06366_);
  or (_11517_, _11516_, _11513_);
  nor (_11518_, _09043_, _11457_);
  or (_11519_, _11458_, _09056_);
  or (_11520_, _11519_, _11518_);
  and (_11521_, _11520_, _09061_);
  and (_11522_, _11521_, _11517_);
  or (_11523_, _11522_, _11461_);
  and (_11524_, _11523_, _06926_);
  and (_11525_, _11466_, _06568_);
  or (_11526_, _11525_, _06278_);
  or (_11527_, _11526_, _11524_);
  and (_11528_, _08550_, _07914_);
  or (_11529_, _11458_, _06279_);
  or (_11530_, _11529_, _11528_);
  and (_11531_, _11530_, _01347_);
  and (_11532_, _11531_, _11527_);
  or (_11533_, _11532_, _11456_);
  and (_40576_, _11533_, _42618_);
  not (_11534_, \oc8051_golden_model_1.DPL [7]);
  nor (_11535_, _01347_, _11534_);
  nor (_11536_, _07960_, _11534_);
  not (_11537_, _07960_);
  nor (_11538_, _08573_, _11537_);
  or (_11539_, _11538_, _11536_);
  and (_11540_, _11539_, _06528_);
  and (_11541_, _08575_, _07960_);
  or (_11542_, _11541_, _11536_);
  and (_11543_, _11542_, _06536_);
  nor (_11544_, _08040_, _11537_);
  or (_11545_, _11544_, _11536_);
  or (_11546_, _11545_, _07215_);
  and (_11547_, _08768_, _07960_);
  or (_11548_, _11547_, _11536_);
  or (_11549_, _11548_, _07151_);
  and (_11550_, _07960_, \oc8051_golden_model_1.ACC [7]);
  or (_11551_, _11550_, _11536_);
  and (_11552_, _11551_, _07141_);
  nor (_11553_, _07141_, _11534_);
  or (_11554_, _11553_, _06341_);
  or (_11555_, _11554_, _11552_);
  and (_11556_, _11555_, _07166_);
  and (_11557_, _11556_, _11549_);
  and (_11558_, _11545_, _06461_);
  or (_11559_, _11558_, _06464_);
  or (_11560_, _11559_, _11557_);
  nor (_11561_, _06019_, _05973_);
  not (_11562_, _11561_);
  or (_11563_, _11551_, _06465_);
  and (_11564_, _11563_, _11562_);
  and (_11565_, _11564_, _11560_);
  and (_11566_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.DPL [0]);
  and (_11567_, _11566_, \oc8051_golden_model_1.DPL [2]);
  and (_11568_, _11567_, \oc8051_golden_model_1.DPL [3]);
  and (_11569_, _11568_, \oc8051_golden_model_1.DPL [4]);
  and (_11570_, _11569_, \oc8051_golden_model_1.DPL [5]);
  and (_11571_, _11570_, \oc8051_golden_model_1.DPL [6]);
  nor (_11572_, _11571_, \oc8051_golden_model_1.DPL [7]);
  and (_11573_, _11571_, \oc8051_golden_model_1.DPL [7]);
  nor (_11574_, _11573_, _11572_);
  and (_11575_, _11574_, _11561_);
  or (_11576_, _11575_, _11565_);
  and (_11577_, _11576_, _06374_);
  nor (_11578_, _08608_, _06374_);
  or (_11579_, _11578_, _10080_);
  or (_11580_, _11579_, _11577_);
  and (_11581_, _11580_, _11546_);
  or (_11582_, _11581_, _07460_);
  and (_11583_, _08755_, _07960_);
  or (_11584_, _11536_, _07208_);
  or (_11585_, _11584_, _11583_);
  and (_11586_, _11585_, _05982_);
  and (_11587_, _11586_, _11582_);
  and (_11588_, _09021_, _07960_);
  or (_11589_, _11588_, _11536_);
  and (_11590_, _11589_, _10094_);
  or (_11591_, _11590_, _06218_);
  or (_11592_, _11591_, _11587_);
  and (_11593_, _08825_, _07960_);
  or (_11594_, _11593_, _11536_);
  or (_11595_, _11594_, _06219_);
  and (_11596_, _11595_, _11592_);
  or (_11597_, _11596_, _06369_);
  and (_11598_, _09044_, _07960_);
  or (_11599_, _11598_, _11536_);
  or (_11600_, _11599_, _07237_);
  and (_11601_, _11600_, _07240_);
  and (_11602_, _11601_, _11597_);
  or (_11603_, _11602_, _11543_);
  and (_11604_, _11603_, _07242_);
  or (_11605_, _11536_, _08043_);
  and (_11606_, _11594_, _06375_);
  and (_11607_, _11606_, _11605_);
  or (_11608_, _11607_, _11604_);
  and (_11609_, _11608_, _07234_);
  and (_11610_, _11551_, _06545_);
  and (_11611_, _11610_, _11605_);
  or (_11612_, _11611_, _06366_);
  or (_11613_, _11612_, _11609_);
  nor (_11614_, _09043_, _11537_);
  or (_11615_, _11536_, _09056_);
  or (_11616_, _11615_, _11614_);
  and (_11617_, _11616_, _09061_);
  and (_11618_, _11617_, _11613_);
  or (_11619_, _11618_, _11540_);
  and (_11620_, _11619_, _06926_);
  and (_11621_, _11548_, _06568_);
  or (_11622_, _11621_, _06278_);
  or (_11623_, _11622_, _11620_);
  and (_11624_, _08550_, _07960_);
  or (_11625_, _11536_, _06279_);
  or (_11626_, _11625_, _11624_);
  and (_11627_, _11626_, _01347_);
  and (_11628_, _11627_, _11623_);
  or (_11629_, _11628_, _11535_);
  and (_40577_, _11629_, _42618_);
  not (_11630_, \oc8051_golden_model_1.DPH [7]);
  nor (_11631_, _01347_, _11630_);
  nor (_11632_, _07963_, _11630_);
  not (_11633_, _08186_);
  nor (_11634_, _08573_, _11633_);
  or (_11635_, _11634_, _11632_);
  and (_11636_, _11635_, _06528_);
  and (_11637_, _08575_, _08186_);
  or (_11638_, _11637_, _11632_);
  and (_11639_, _11638_, _06536_);
  nor (_11640_, _08040_, _11633_);
  or (_11641_, _11640_, _11632_);
  or (_11642_, _11641_, _07215_);
  and (_11643_, _08768_, _08186_);
  or (_11644_, _11643_, _11632_);
  or (_11645_, _11644_, _07151_);
  and (_11646_, _07963_, \oc8051_golden_model_1.ACC [7]);
  or (_11647_, _11646_, _11632_);
  and (_11648_, _11647_, _07141_);
  nor (_11649_, _07141_, _11630_);
  or (_11650_, _11649_, _06341_);
  or (_11651_, _11650_, _11648_);
  and (_11652_, _11651_, _07166_);
  and (_11653_, _11652_, _11645_);
  and (_11654_, _11641_, _06461_);
  or (_11655_, _11654_, _06464_);
  or (_11656_, _11655_, _11653_);
  or (_11657_, _11647_, _06465_);
  and (_11658_, _11657_, _11562_);
  and (_11659_, _11658_, _11656_);
  and (_11660_, _11573_, \oc8051_golden_model_1.DPH [0]);
  and (_11661_, _11660_, \oc8051_golden_model_1.DPH [1]);
  and (_11662_, _11661_, \oc8051_golden_model_1.DPH [2]);
  and (_11663_, _11662_, \oc8051_golden_model_1.DPH [3]);
  and (_11664_, _11663_, \oc8051_golden_model_1.DPH [4]);
  and (_11665_, _11664_, \oc8051_golden_model_1.DPH [5]);
  and (_11666_, _11665_, \oc8051_golden_model_1.DPH [6]);
  nor (_11667_, _11666_, _11630_);
  and (_11668_, _11666_, _11630_);
  or (_11669_, _11668_, _11667_);
  and (_11670_, _11669_, _11561_);
  or (_11671_, _11670_, _11659_);
  and (_11672_, _11671_, _06374_);
  and (_11673_, _06373_, _06182_);
  or (_11674_, _11673_, _10080_);
  or (_11675_, _11674_, _11672_);
  and (_11676_, _11675_, _11642_);
  or (_11677_, _11676_, _07460_);
  or (_11678_, _11632_, _07208_);
  and (_11679_, _08755_, _07963_);
  or (_11680_, _11679_, _11678_);
  and (_11681_, _11680_, _05982_);
  and (_11682_, _11681_, _11677_);
  and (_11683_, _09021_, _07963_);
  or (_11684_, _11683_, _11632_);
  and (_11685_, _11684_, _10094_);
  or (_11686_, _11685_, _06218_);
  or (_11687_, _11686_, _11682_);
  and (_11688_, _08825_, _07963_);
  or (_11689_, _11688_, _11632_);
  or (_11690_, _11689_, _06219_);
  and (_11691_, _11690_, _11687_);
  or (_11692_, _11691_, _06369_);
  and (_11693_, _09044_, _07963_);
  or (_11694_, _11693_, _11632_);
  or (_11695_, _11694_, _07237_);
  and (_11696_, _11695_, _07240_);
  and (_11697_, _11696_, _11692_);
  or (_11698_, _11697_, _11639_);
  and (_11699_, _11698_, _07242_);
  or (_11700_, _11632_, _08043_);
  and (_11701_, _11689_, _06375_);
  and (_11702_, _11701_, _11700_);
  or (_11703_, _11702_, _11699_);
  and (_11704_, _11703_, _07234_);
  and (_11705_, _11647_, _06545_);
  and (_11706_, _11705_, _11700_);
  or (_11707_, _11706_, _06366_);
  or (_11708_, _11707_, _11704_);
  nor (_11709_, _09043_, _11633_);
  or (_11710_, _11632_, _09056_);
  or (_11711_, _11710_, _11709_);
  and (_11712_, _11711_, _09061_);
  and (_11713_, _11712_, _11708_);
  or (_11714_, _11713_, _11636_);
  and (_11715_, _11714_, _06926_);
  and (_11716_, _11644_, _06568_);
  or (_11717_, _11716_, _06278_);
  or (_11718_, _11717_, _11715_);
  and (_11719_, _08550_, _08186_);
  or (_11720_, _11632_, _06279_);
  or (_11721_, _11720_, _11719_);
  and (_11722_, _11721_, _01347_);
  and (_11723_, _11722_, _11718_);
  or (_11724_, _11723_, _11631_);
  and (_40580_, _11724_, _42618_);
  and (_11725_, _01351_, \oc8051_golden_model_1.TL1 [7]);
  not (_11726_, _07968_);
  and (_11727_, _11726_, \oc8051_golden_model_1.TL1 [7]);
  nor (_11728_, _08573_, _11726_);
  or (_11729_, _11728_, _11727_);
  and (_11730_, _11729_, _06528_);
  and (_11731_, _08575_, _07968_);
  or (_11732_, _11731_, _11727_);
  and (_11733_, _11732_, _06536_);
  and (_11734_, _08768_, _07968_);
  or (_11735_, _11734_, _11727_);
  or (_11736_, _11735_, _07151_);
  and (_11737_, _07968_, \oc8051_golden_model_1.ACC [7]);
  or (_11738_, _11737_, _11727_);
  and (_11739_, _11738_, _07141_);
  and (_11740_, _07142_, \oc8051_golden_model_1.TL1 [7]);
  or (_11741_, _11740_, _06341_);
  or (_11742_, _11741_, _11739_);
  and (_11743_, _11742_, _07166_);
  and (_11744_, _11743_, _11736_);
  nor (_11745_, _08040_, _11726_);
  or (_11746_, _11745_, _11727_);
  and (_11747_, _11746_, _06461_);
  or (_11748_, _11747_, _11744_);
  and (_11749_, _11748_, _06465_);
  and (_11750_, _11738_, _06464_);
  or (_11751_, _11750_, _10080_);
  or (_11752_, _11751_, _11749_);
  or (_11753_, _11746_, _07215_);
  and (_11754_, _11753_, _11752_);
  or (_11755_, _11754_, _07460_);
  and (_11756_, _08755_, _07968_);
  or (_11757_, _11727_, _07208_);
  or (_11758_, _11757_, _11756_);
  and (_11759_, _11758_, _05982_);
  and (_11760_, _11759_, _11755_);
  and (_11761_, _09021_, _07968_);
  or (_11762_, _11761_, _11727_);
  and (_11763_, _11762_, _10094_);
  or (_11764_, _11763_, _06218_);
  or (_11765_, _11764_, _11760_);
  and (_11766_, _08825_, _07968_);
  or (_11767_, _11766_, _11727_);
  or (_11768_, _11767_, _06219_);
  and (_11769_, _11768_, _11765_);
  or (_11770_, _11769_, _06369_);
  and (_11771_, _09044_, _07968_);
  or (_11772_, _11771_, _11727_);
  or (_11773_, _11772_, _07237_);
  and (_11774_, _11773_, _07240_);
  and (_11775_, _11774_, _11770_);
  or (_11776_, _11775_, _11733_);
  and (_11777_, _11776_, _07242_);
  or (_11778_, _11727_, _08043_);
  and (_11779_, _11767_, _06375_);
  and (_11780_, _11779_, _11778_);
  or (_11781_, _11780_, _11777_);
  and (_11782_, _11781_, _07234_);
  and (_11783_, _11738_, _06545_);
  and (_11784_, _11783_, _11778_);
  or (_11785_, _11784_, _06366_);
  or (_11786_, _11785_, _11782_);
  nor (_11787_, _09043_, _11726_);
  or (_11788_, _11727_, _09056_);
  or (_11789_, _11788_, _11787_);
  and (_11790_, _11789_, _09061_);
  and (_11791_, _11790_, _11786_);
  or (_11792_, _11791_, _11730_);
  and (_11793_, _11792_, _06926_);
  and (_11794_, _11735_, _06568_);
  or (_11795_, _11794_, _06278_);
  or (_11796_, _11795_, _11793_);
  and (_11797_, _08550_, _07968_);
  or (_11798_, _11727_, _06279_);
  or (_11799_, _11798_, _11797_);
  and (_11800_, _11799_, _01347_);
  and (_11801_, _11800_, _11796_);
  or (_11802_, _11801_, _11725_);
  and (_40581_, _11802_, _42618_);
  and (_11803_, _01351_, \oc8051_golden_model_1.TL0 [7]);
  not (_11804_, _07919_);
  and (_11805_, _11804_, \oc8051_golden_model_1.TL0 [7]);
  nor (_11806_, _08573_, _11804_);
  or (_11807_, _11806_, _11805_);
  and (_11808_, _11807_, _06528_);
  and (_11809_, _08575_, _07919_);
  or (_11810_, _11809_, _11805_);
  and (_11811_, _11810_, _06536_);
  nor (_11812_, _08040_, _11804_);
  or (_11813_, _11812_, _11805_);
  or (_11814_, _11813_, _07215_);
  and (_11815_, _08768_, _07919_);
  or (_11816_, _11815_, _11805_);
  or (_11817_, _11816_, _07151_);
  and (_11818_, _07919_, \oc8051_golden_model_1.ACC [7]);
  or (_11819_, _11818_, _11805_);
  and (_11820_, _11819_, _07141_);
  and (_11821_, _07142_, \oc8051_golden_model_1.TL0 [7]);
  or (_11822_, _11821_, _06341_);
  or (_11823_, _11822_, _11820_);
  and (_11824_, _11823_, _07166_);
  and (_11825_, _11824_, _11817_);
  and (_11826_, _11813_, _06461_);
  or (_11827_, _11826_, _11825_);
  and (_11828_, _11827_, _06465_);
  and (_11829_, _11819_, _06464_);
  or (_11830_, _11829_, _10080_);
  or (_11831_, _11830_, _11828_);
  and (_11832_, _11831_, _11814_);
  or (_11833_, _11832_, _07460_);
  and (_11834_, _08755_, _07919_);
  or (_11835_, _11805_, _07208_);
  or (_11836_, _11835_, _11834_);
  and (_11837_, _11836_, _05982_);
  and (_11838_, _11837_, _11833_);
  and (_11839_, _09021_, _07919_);
  or (_11840_, _11839_, _11805_);
  and (_11841_, _11840_, _10094_);
  or (_11842_, _11841_, _06218_);
  or (_11843_, _11842_, _11838_);
  and (_11844_, _08825_, _07919_);
  or (_11845_, _11844_, _11805_);
  or (_11846_, _11845_, _06219_);
  and (_11847_, _11846_, _11843_);
  or (_11848_, _11847_, _06369_);
  and (_11849_, _09044_, _07919_);
  or (_11850_, _11849_, _11805_);
  or (_11851_, _11850_, _07237_);
  and (_11852_, _11851_, _07240_);
  and (_11853_, _11852_, _11848_);
  or (_11854_, _11853_, _11811_);
  and (_11855_, _11854_, _07242_);
  or (_11856_, _11805_, _08043_);
  and (_11857_, _11845_, _06375_);
  and (_11858_, _11857_, _11856_);
  or (_11859_, _11858_, _11855_);
  and (_11860_, _11859_, _07234_);
  and (_11861_, _11819_, _06545_);
  and (_11862_, _11861_, _11856_);
  or (_11863_, _11862_, _06366_);
  or (_11864_, _11863_, _11860_);
  nor (_11865_, _09043_, _11804_);
  or (_11866_, _11805_, _09056_);
  or (_11867_, _11866_, _11865_);
  and (_11868_, _11867_, _09061_);
  and (_11869_, _11868_, _11864_);
  or (_11870_, _11869_, _11808_);
  and (_11871_, _11870_, _06926_);
  and (_11872_, _11816_, _06568_);
  or (_11873_, _11872_, _06278_);
  or (_11874_, _11873_, _11871_);
  and (_11875_, _08550_, _07919_);
  or (_11876_, _11805_, _06279_);
  or (_11877_, _11876_, _11875_);
  and (_11878_, _11877_, _01347_);
  and (_11879_, _11878_, _11874_);
  or (_11880_, _11879_, _11803_);
  and (_40582_, _11880_, _42618_);
  and (_11881_, _01351_, \oc8051_golden_model_1.TCON [7]);
  not (_11882_, _07928_);
  and (_11883_, _11882_, \oc8051_golden_model_1.TCON [7]);
  and (_11884_, _08575_, _07928_);
  or (_11885_, _11884_, _11883_);
  and (_11886_, _11885_, _06536_);
  nor (_11887_, _08040_, _11882_);
  or (_11888_, _11887_, _11883_);
  or (_11889_, _11888_, _07215_);
  not (_11890_, _08616_);
  and (_11891_, _11890_, \oc8051_golden_model_1.TCON [7]);
  and (_11892_, _08649_, _08616_);
  or (_11893_, _11892_, _11891_);
  and (_11894_, _11893_, _06268_);
  and (_11895_, _08768_, _07928_);
  or (_11896_, _11895_, _11883_);
  or (_11897_, _11896_, _07151_);
  and (_11898_, _07928_, \oc8051_golden_model_1.ACC [7]);
  or (_11899_, _11898_, _11883_);
  and (_11900_, _11899_, _07141_);
  and (_11901_, _07142_, \oc8051_golden_model_1.TCON [7]);
  or (_11902_, _11901_, _06341_);
  or (_11903_, _11902_, _11900_);
  and (_11904_, _11903_, _06273_);
  and (_11905_, _11904_, _11897_);
  and (_11906_, _08773_, _08616_);
  or (_11907_, _11906_, _11891_);
  and (_11908_, _11907_, _06272_);
  or (_11909_, _11908_, _06461_);
  or (_11910_, _11909_, _11905_);
  or (_11911_, _11888_, _07166_);
  and (_11912_, _11911_, _11910_);
  or (_11913_, _11912_, _06464_);
  or (_11914_, _11899_, _06465_);
  and (_11915_, _11914_, _06269_);
  and (_11916_, _11915_, _11913_);
  or (_11917_, _11916_, _11894_);
  and (_11918_, _11917_, _06262_);
  and (_11919_, _08790_, _08616_);
  or (_11920_, _11919_, _11891_);
  and (_11921_, _11920_, _06261_);
  or (_11922_, _11921_, _11918_);
  and (_11923_, _11922_, _06258_);
  and (_11924_, _08808_, _08616_);
  or (_11925_, _11924_, _11891_);
  and (_11926_, _11925_, _06257_);
  or (_11927_, _11926_, _10080_);
  or (_11928_, _11927_, _11923_);
  and (_11929_, _11928_, _11889_);
  or (_11930_, _11929_, _07460_);
  and (_11931_, _08755_, _07928_);
  or (_11932_, _11883_, _07208_);
  or (_11933_, _11932_, _11931_);
  and (_11934_, _11933_, _05982_);
  and (_11935_, _11934_, _11930_);
  and (_11936_, _09021_, _07928_);
  or (_11937_, _11936_, _11883_);
  and (_11938_, _11937_, _10094_);
  or (_11939_, _11938_, _06218_);
  or (_11940_, _11939_, _11935_);
  and (_11941_, _08825_, _07928_);
  or (_11942_, _11941_, _11883_);
  or (_11943_, _11942_, _06219_);
  and (_11944_, _11943_, _11940_);
  or (_11945_, _11944_, _06369_);
  and (_11946_, _09044_, _07928_);
  or (_11947_, _11946_, _11883_);
  or (_11948_, _11947_, _07237_);
  and (_11949_, _11948_, _07240_);
  and (_11950_, _11949_, _11945_);
  or (_11951_, _11950_, _11886_);
  and (_11952_, _11951_, _07242_);
  or (_11953_, _11883_, _08043_);
  and (_11954_, _11942_, _06375_);
  and (_11955_, _11954_, _11953_);
  or (_11956_, _11955_, _11952_);
  and (_11957_, _11956_, _07234_);
  and (_11958_, _11899_, _06545_);
  and (_11959_, _11958_, _11953_);
  or (_11960_, _11959_, _06366_);
  or (_11961_, _11960_, _11957_);
  nor (_11962_, _09043_, _11882_);
  or (_11963_, _11883_, _09056_);
  or (_11964_, _11963_, _11962_);
  and (_11965_, _11964_, _09061_);
  and (_11966_, _11965_, _11961_);
  nor (_11967_, _08573_, _11882_);
  or (_11968_, _11967_, _11883_);
  and (_11969_, _11968_, _06528_);
  or (_11970_, _11969_, _06568_);
  or (_11971_, _11970_, _11966_);
  or (_11972_, _11896_, _06926_);
  and (_11973_, _11972_, _05928_);
  and (_11974_, _11973_, _11971_);
  and (_11975_, _11893_, _05927_);
  or (_11976_, _11975_, _06278_);
  or (_11977_, _11976_, _11974_);
  and (_11978_, _08550_, _07928_);
  or (_11979_, _11883_, _06279_);
  or (_11980_, _11979_, _11978_);
  and (_11981_, _11980_, _01347_);
  and (_11982_, _11981_, _11977_);
  or (_11983_, _11982_, _11881_);
  and (_40583_, _11983_, _42618_);
  and (_11984_, _01351_, \oc8051_golden_model_1.TH1 [7]);
  not (_11985_, _07910_);
  and (_11986_, _11985_, \oc8051_golden_model_1.TH1 [7]);
  nor (_11987_, _08573_, _11985_);
  or (_11988_, _11987_, _11986_);
  and (_11989_, _11988_, _06528_);
  and (_11990_, _08575_, _07910_);
  or (_11991_, _11990_, _11986_);
  and (_11992_, _11991_, _06536_);
  nor (_11993_, _08040_, _11985_);
  or (_11994_, _11993_, _11986_);
  or (_11995_, _11994_, _07215_);
  and (_11996_, _08768_, _07910_);
  or (_11997_, _11996_, _11986_);
  or (_11998_, _11997_, _07151_);
  and (_11999_, _07910_, \oc8051_golden_model_1.ACC [7]);
  or (_12000_, _11999_, _11986_);
  and (_12001_, _12000_, _07141_);
  and (_12002_, _07142_, \oc8051_golden_model_1.TH1 [7]);
  or (_12003_, _12002_, _06341_);
  or (_12004_, _12003_, _12001_);
  and (_12005_, _12004_, _07166_);
  and (_12006_, _12005_, _11998_);
  and (_12007_, _11994_, _06461_);
  or (_12008_, _12007_, _12006_);
  and (_12009_, _12008_, _06465_);
  and (_12010_, _12000_, _06464_);
  or (_12011_, _12010_, _10080_);
  or (_12012_, _12011_, _12009_);
  and (_12013_, _12012_, _11995_);
  or (_12014_, _12013_, _07460_);
  and (_12015_, _08755_, _07910_);
  or (_12016_, _11986_, _07208_);
  or (_12017_, _12016_, _12015_);
  and (_12018_, _12017_, _05982_);
  and (_12019_, _12018_, _12014_);
  and (_12020_, _09021_, _07910_);
  or (_12021_, _12020_, _11986_);
  and (_12022_, _12021_, _10094_);
  or (_12023_, _12022_, _06218_);
  or (_12024_, _12023_, _12019_);
  and (_12025_, _08825_, _07910_);
  or (_12026_, _12025_, _11986_);
  or (_12027_, _12026_, _06219_);
  and (_12028_, _12027_, _12024_);
  or (_12029_, _12028_, _06369_);
  and (_12030_, _09044_, _07910_);
  or (_12031_, _12030_, _11986_);
  or (_12032_, _12031_, _07237_);
  and (_12033_, _12032_, _07240_);
  and (_12034_, _12033_, _12029_);
  or (_12035_, _12034_, _11992_);
  and (_12036_, _12035_, _07242_);
  or (_12037_, _11986_, _08043_);
  and (_12038_, _12026_, _06375_);
  and (_12039_, _12038_, _12037_);
  or (_12040_, _12039_, _12036_);
  and (_12041_, _12040_, _07234_);
  and (_12042_, _12000_, _06545_);
  and (_12043_, _12042_, _12037_);
  or (_12044_, _12043_, _06366_);
  or (_12045_, _12044_, _12041_);
  nor (_12046_, _09043_, _11985_);
  or (_12047_, _11986_, _09056_);
  or (_12048_, _12047_, _12046_);
  and (_12049_, _12048_, _09061_);
  and (_12050_, _12049_, _12045_);
  or (_12051_, _12050_, _11989_);
  and (_12052_, _12051_, _06926_);
  and (_12053_, _11997_, _06568_);
  or (_12054_, _12053_, _06278_);
  or (_12055_, _12054_, _12052_);
  and (_12056_, _08550_, _07910_);
  or (_12057_, _11986_, _06279_);
  or (_12058_, _12057_, _12056_);
  and (_12059_, _12058_, _01347_);
  and (_12060_, _12059_, _12055_);
  or (_12061_, _12060_, _11984_);
  and (_40584_, _12061_, _42618_);
  and (_12062_, _01351_, \oc8051_golden_model_1.TH0 [7]);
  not (_12063_, _07922_);
  and (_12064_, _12063_, \oc8051_golden_model_1.TH0 [7]);
  nor (_12065_, _08573_, _12063_);
  or (_12066_, _12065_, _12064_);
  and (_12067_, _12066_, _06528_);
  and (_12068_, _08575_, _07922_);
  or (_12069_, _12068_, _12064_);
  and (_12070_, _12069_, _06536_);
  nor (_12071_, _08040_, _12063_);
  or (_12072_, _12071_, _12064_);
  or (_12073_, _12072_, _07215_);
  and (_12074_, _08768_, _07922_);
  or (_12075_, _12074_, _12064_);
  or (_12076_, _12075_, _07151_);
  and (_12077_, _07922_, \oc8051_golden_model_1.ACC [7]);
  or (_12078_, _12077_, _12064_);
  and (_12079_, _12078_, _07141_);
  and (_12080_, _07142_, \oc8051_golden_model_1.TH0 [7]);
  or (_12081_, _12080_, _06341_);
  or (_12082_, _12081_, _12079_);
  and (_12083_, _12082_, _07166_);
  and (_12084_, _12083_, _12076_);
  and (_12085_, _12072_, _06461_);
  or (_12086_, _12085_, _12084_);
  and (_12087_, _12086_, _06465_);
  and (_12088_, _12078_, _06464_);
  or (_12089_, _12088_, _10080_);
  or (_12090_, _12089_, _12087_);
  and (_12091_, _12090_, _12073_);
  or (_12092_, _12091_, _07460_);
  and (_12093_, _08755_, _07922_);
  or (_12094_, _12064_, _07208_);
  or (_12095_, _12094_, _12093_);
  and (_12096_, _12095_, _05982_);
  and (_12097_, _12096_, _12092_);
  and (_12098_, _09021_, _07922_);
  or (_12099_, _12098_, _12064_);
  and (_12100_, _12099_, _10094_);
  or (_12101_, _12100_, _06218_);
  or (_12102_, _12101_, _12097_);
  and (_12103_, _08825_, _07922_);
  or (_12104_, _12103_, _12064_);
  or (_12105_, _12104_, _06219_);
  and (_12106_, _12105_, _12102_);
  or (_12107_, _12106_, _06369_);
  and (_12108_, _09044_, _07922_);
  or (_12109_, _12108_, _12064_);
  or (_12110_, _12109_, _07237_);
  and (_12111_, _12110_, _07240_);
  and (_12112_, _12111_, _12107_);
  or (_12113_, _12112_, _12070_);
  and (_12114_, _12113_, _07242_);
  or (_12115_, _12064_, _08043_);
  and (_12116_, _12104_, _06375_);
  and (_12117_, _12116_, _12115_);
  or (_12118_, _12117_, _12114_);
  and (_12119_, _12118_, _07234_);
  and (_12120_, _12078_, _06545_);
  and (_12121_, _12120_, _12115_);
  or (_12122_, _12121_, _06366_);
  or (_12123_, _12122_, _12119_);
  nor (_12124_, _09043_, _12063_);
  or (_12125_, _12064_, _09056_);
  or (_12126_, _12125_, _12124_);
  and (_12127_, _12126_, _09061_);
  and (_12128_, _12127_, _12123_);
  or (_12129_, _12128_, _12067_);
  and (_12130_, _12129_, _06926_);
  and (_12131_, _12075_, _06568_);
  or (_12132_, _12131_, _06278_);
  or (_12133_, _12132_, _12130_);
  and (_12134_, _08550_, _07922_);
  or (_12135_, _12064_, _06279_);
  or (_12136_, _12135_, _12134_);
  and (_12137_, _12136_, _01347_);
  and (_12138_, _12137_, _12133_);
  or (_12139_, _12138_, _12062_);
  and (_40585_, _12139_, _42618_);
  not (_12140_, _06379_);
  nor (_12141_, _11360_, _11353_);
  not (_12142_, _05616_);
  and (_12143_, _09409_, _12142_);
  and (_12144_, _12143_, _09472_);
  and (_12145_, _12144_, _09469_);
  and (_12146_, _12145_, \oc8051_golden_model_1.PC [14]);
  and (_12147_, _12146_, _09468_);
  nor (_12148_, _12146_, _09468_);
  or (_12149_, _12148_, _12147_);
  nor (_12150_, _12149_, _12141_);
  and (_12151_, _11203_, _11157_);
  nor (_12152_, _12151_, _12149_);
  nor (_12153_, _11097_, _06540_);
  and (_12154_, _11069_, _11037_);
  nor (_12155_, _12154_, _12149_);
  not (_12156_, _07042_);
  and (_12157_, _10998_, _12156_);
  nor (_12158_, _11008_, _07040_);
  not (_12159_, _12158_);
  or (_12160_, _12159_, _11012_);
  nor (_12161_, _12160_, _11011_);
  and (_12162_, _12161_, _12157_);
  nor (_12163_, _12162_, _12149_);
  nor (_12164_, _10496_, _06542_);
  nor (_12165_, _12149_, _10979_);
  nor (_12166_, _10954_, _06533_);
  nor (_12167_, _07482_, _05954_);
  nor (_12168_, _12167_, _10509_);
  and (_12169_, _12168_, _10940_);
  nor (_12170_, _12169_, _12149_);
  nor (_12171_, _09487_, _09030_);
  nor (_12172_, _10093_, _05974_);
  nor (_12173_, _09479_, _05982_);
  nor (_12174_, _06006_, _05973_);
  not (_12175_, _12174_);
  not (_12176_, _06371_);
  not (_12177_, _06347_);
  and (_12178_, _09412_, \oc8051_golden_model_1.PC [8]);
  and (_12179_, _12178_, \oc8051_golden_model_1.PC [9]);
  and (_12180_, _12179_, \oc8051_golden_model_1.PC [10]);
  and (_12181_, _12180_, \oc8051_golden_model_1.PC [11]);
  and (_12182_, _12181_, \oc8051_golden_model_1.PC [12]);
  and (_12183_, _12182_, \oc8051_golden_model_1.PC [13]);
  and (_12184_, _12183_, \oc8051_golden_model_1.PC [14]);
  nor (_12185_, _12183_, \oc8051_golden_model_1.PC [14]);
  nor (_12186_, _12185_, _12184_);
  not (_12187_, _12186_);
  nor (_12188_, _12187_, _08608_);
  and (_12189_, _12187_, _08608_);
  nor (_12190_, _12189_, _12188_);
  not (_12191_, _12190_);
  nor (_12192_, _12182_, \oc8051_golden_model_1.PC [13]);
  nor (_12193_, _12192_, _12183_);
  not (_12194_, _12193_);
  nor (_12195_, _12194_, _08608_);
  and (_12196_, _12194_, _08608_);
  nor (_12197_, _12181_, \oc8051_golden_model_1.PC [12]);
  nor (_12198_, _12197_, _12182_);
  not (_12199_, _12198_);
  nor (_12200_, _12199_, _08608_);
  nor (_12201_, _12179_, \oc8051_golden_model_1.PC [10]);
  nor (_12202_, _12201_, _12180_);
  not (_12203_, _12202_);
  nor (_12204_, _12203_, _08608_);
  not (_12205_, _12204_);
  nor (_12206_, _12180_, \oc8051_golden_model_1.PC [11]);
  nor (_12207_, _12206_, _12181_);
  not (_12208_, _12207_);
  nor (_12209_, _12208_, _08608_);
  and (_12210_, _12208_, _08608_);
  nor (_12211_, _12210_, _12209_);
  and (_12212_, _12203_, _08608_);
  nor (_12213_, _12212_, _12204_);
  and (_12214_, _12213_, _12211_);
  nor (_12215_, _12178_, \oc8051_golden_model_1.PC [9]);
  nor (_12216_, _12215_, _12179_);
  not (_12217_, _12216_);
  nor (_12218_, _12217_, _08608_);
  and (_12219_, _12217_, _08608_);
  nor (_12220_, _12219_, _12218_);
  nor (_12221_, _09416_, _08608_);
  and (_12222_, _09416_, _08608_);
  and (_12223_, _09411_, _08656_);
  nor (_12224_, _12223_, \oc8051_golden_model_1.PC [6]);
  nor (_12225_, _12224_, _09413_);
  not (_12226_, _12225_);
  nor (_12227_, _12226_, _08857_);
  and (_12228_, _12226_, _08857_);
  nor (_12229_, _12228_, _12227_);
  not (_12230_, _12229_);
  and (_12231_, _09411_, \oc8051_golden_model_1.PC [4]);
  nor (_12232_, _12231_, \oc8051_golden_model_1.PC [5]);
  nor (_12233_, _12232_, _12223_);
  not (_12234_, _12233_);
  nor (_12235_, _12234_, _08926_);
  and (_12236_, _12234_, _08926_);
  nor (_12237_, _09411_, \oc8051_golden_model_1.PC [4]);
  nor (_12238_, _12237_, _12231_);
  not (_12239_, _12238_);
  nor (_12240_, _12239_, _08892_);
  nor (_12241_, _09410_, \oc8051_golden_model_1.PC [3]);
  nor (_12242_, _12241_, _09411_);
  not (_12243_, _12242_);
  nor (_12244_, _12243_, _06452_);
  and (_12245_, _12243_, _06452_);
  nor (_12246_, _05634_, \oc8051_golden_model_1.PC [2]);
  nor (_12247_, _12246_, _09410_);
  not (_12248_, _12247_);
  nor (_12249_, _12248_, _06697_);
  nor (_12250_, _07038_, _06111_);
  nor (_12251_, _06872_, \oc8051_golden_model_1.PC [0]);
  and (_12252_, _07038_, _06111_);
  nor (_12253_, _12252_, _12250_);
  and (_12254_, _12253_, _12251_);
  nor (_12255_, _12254_, _12250_);
  and (_12256_, _12248_, _06697_);
  nor (_12257_, _12256_, _12249_);
  not (_12258_, _12257_);
  nor (_12259_, _12258_, _12255_);
  nor (_12260_, _12259_, _12249_);
  nor (_12261_, _12260_, _12245_);
  nor (_12262_, _12261_, _12244_);
  and (_12263_, _12239_, _08892_);
  nor (_12264_, _12263_, _12240_);
  not (_12265_, _12264_);
  nor (_12266_, _12265_, _12262_);
  nor (_12267_, _12266_, _12240_);
  nor (_12268_, _12267_, _12236_);
  nor (_12269_, _12268_, _12235_);
  nor (_12270_, _12269_, _12230_);
  nor (_12271_, _12270_, _12227_);
  nor (_12272_, _12271_, _12222_);
  or (_12273_, _12272_, _12221_);
  nor (_12274_, _09412_, \oc8051_golden_model_1.PC [8]);
  nor (_12275_, _12274_, _12178_);
  not (_12276_, _12275_);
  nor (_12277_, _12276_, _08608_);
  and (_12278_, _12276_, _08608_);
  nor (_12279_, _12278_, _12277_);
  and (_12280_, _12279_, _12273_);
  and (_12281_, _12280_, _12220_);
  and (_12282_, _12281_, _12214_);
  nor (_12283_, _12277_, _12218_);
  not (_12284_, _12283_);
  and (_12285_, _12284_, _12214_);
  or (_12286_, _12285_, _12209_);
  nor (_12287_, _12286_, _12282_);
  and (_12288_, _12287_, _12205_);
  and (_12289_, _12199_, _08608_);
  nor (_12290_, _12289_, _12200_);
  not (_12291_, _12290_);
  nor (_12292_, _12291_, _12288_);
  nor (_12293_, _12292_, _12200_);
  nor (_12294_, _12293_, _12196_);
  nor (_12295_, _12294_, _12195_);
  nor (_12296_, _12295_, _12191_);
  nor (_12297_, _12296_, _12188_);
  and (_12298_, _09479_, _08608_);
  nor (_12299_, _09479_, _08608_);
  nor (_12300_, _12299_, _12298_);
  and (_12301_, _12300_, _12297_);
  nor (_12302_, _12300_, _12297_);
  nor (_12303_, _12302_, _12301_);
  nor (_12304_, _08755_, _06286_);
  nor (_12305_, _12304_, _08802_);
  or (_12306_, _09446_, _06317_);
  or (_12307_, _09122_, _07607_);
  and (_12308_, _12307_, _12306_);
  and (_12309_, _12308_, _12305_);
  or (_12310_, _09167_, _07896_);
  or (_12311_, _09447_, _06611_);
  and (_12312_, _12311_, _12310_);
  or (_12313_, _09212_, _07883_);
  or (_12314_, _09448_, _06968_);
  and (_12315_, _12314_, _12313_);
  and (_12316_, _12315_, _12312_);
  and (_12317_, _12316_, _12309_);
  or (_12318_, _09449_, _06213_);
  or (_12319_, _09257_, _06473_);
  and (_12320_, _12319_, _12318_);
  or (_12321_, _09450_, _06656_);
  or (_12322_, _09302_, _06657_);
  and (_12323_, _12322_, _12321_);
  and (_12324_, _12323_, _12320_);
  or (_12325_, _09451_, _07004_);
  or (_12326_, _09347_, _07005_);
  and (_12327_, _12326_, _12325_);
  or (_12328_, _09392_, _06251_);
  nand (_12329_, _09392_, _06251_);
  and (_12330_, _12329_, _12328_);
  and (_12331_, _12330_, _12327_);
  and (_12332_, _12331_, _12324_);
  and (_12333_, _12332_, _12317_);
  or (_12334_, _12333_, _12303_);
  nand (_12335_, _12332_, _12317_);
  or (_12336_, _12335_, _09479_);
  nand (_12337_, _12336_, _12334_);
  nor (_12338_, _12337_, _12177_);
  not (_12339_, _08041_);
  and (_12340_, _08040_, _06182_);
  nor (_12341_, _12340_, _12339_);
  nor (_12342_, _08142_, _07607_);
  and (_12343_, _08142_, _07607_);
  nor (_12344_, _12343_, _12342_);
  and (_12345_, _12344_, _12341_);
  or (_12346_, _08244_, _07896_);
  and (_12347_, _08244_, _07896_);
  not (_12348_, _12347_);
  and (_12349_, _12348_, _12346_);
  and (_12350_, _08541_, _07883_);
  nor (_12351_, _08541_, _07883_);
  nor (_12352_, _12351_, _12350_);
  and (_12353_, _12352_, _12349_);
  and (_12354_, _12353_, _12345_);
  and (_12355_, _07594_, _06473_);
  and (_12356_, _07776_, _06657_);
  nor (_12357_, _12356_, _12355_);
  or (_12358_, _07594_, _06473_);
  or (_12359_, _07776_, _06657_);
  and (_12360_, _12359_, _12358_);
  and (_12361_, _12360_, _12357_);
  or (_12362_, _07357_, _07005_);
  and (_12363_, _07357_, _07005_);
  not (_12364_, _12363_);
  and (_12365_, _12364_, _12362_);
  nand (_12366_, _07133_, _06251_);
  or (_12367_, _07133_, _06251_);
  and (_12368_, _12367_, _12366_);
  and (_12369_, _12368_, _12365_);
  and (_12370_, _12369_, _12361_);
  and (_12371_, _12370_, _12354_);
  nand (_12372_, _12371_, _09479_);
  and (_12373_, _07209_, _06260_);
  not (_12374_, _12373_);
  not (_12375_, _06357_);
  nor (_12376_, _07211_, _06006_);
  nor (_12377_, _12376_, _12375_);
  and (_12378_, _12377_, _12374_);
  not (_12379_, _12378_);
  not (_12380_, _12303_);
  or (_12381_, _12371_, _12380_);
  and (_12382_, _12381_, _12379_);
  and (_12383_, _12382_, _12372_);
  and (_12384_, _09487_, _06464_);
  not (_12385_, _12149_);
  and (_12386_, _12385_, _07154_);
  not (_12387_, _08654_);
  not (_12388_, _09487_);
  and (_12389_, _08142_, _08040_);
  and (_12390_, _12389_, _08553_);
  and (_12391_, _07357_, _07133_);
  and (_12392_, _12391_, _08554_);
  nand (_12393_, _12392_, _12390_);
  or (_12394_, _12393_, _12388_);
  and (_12395_, _08659_, \oc8051_golden_model_1.PC [8]);
  and (_12396_, _12395_, \oc8051_golden_model_1.PC [9]);
  and (_12397_, _12396_, \oc8051_golden_model_1.PC [10]);
  and (_12398_, _12397_, \oc8051_golden_model_1.PC [11]);
  and (_12399_, _12398_, \oc8051_golden_model_1.PC [12]);
  and (_12400_, _12399_, \oc8051_golden_model_1.PC [13]);
  and (_12401_, _12400_, \oc8051_golden_model_1.PC [14]);
  nor (_12402_, _12400_, \oc8051_golden_model_1.PC [14]);
  nor (_12403_, _12402_, _12401_);
  and (_12404_, _12403_, _06182_);
  nor (_12405_, _12403_, _06182_);
  nor (_12406_, _12405_, _12404_);
  not (_12407_, _12406_);
  nor (_12408_, _12399_, \oc8051_golden_model_1.PC [13]);
  nor (_12409_, _12408_, _12400_);
  nor (_12410_, _12409_, _06182_);
  and (_12411_, _12409_, _06182_);
  not (_12412_, _12411_);
  nor (_12413_, _12398_, \oc8051_golden_model_1.PC [12]);
  nor (_12414_, _12413_, _12399_);
  and (_12415_, _12414_, _06182_);
  nor (_12416_, _12397_, \oc8051_golden_model_1.PC [11]);
  nor (_12417_, _12416_, _12398_);
  and (_12418_, _12417_, _06182_);
  nor (_12419_, _12417_, _06182_);
  nor (_12420_, _12396_, \oc8051_golden_model_1.PC [10]);
  nor (_12421_, _12420_, _12397_);
  and (_12422_, _12421_, _06182_);
  nor (_12423_, _12421_, _06182_);
  nor (_12424_, _12423_, _12422_);
  nor (_12425_, _12395_, \oc8051_golden_model_1.PC [9]);
  nor (_12426_, _12425_, _12396_);
  nor (_12427_, _12426_, _06182_);
  and (_12428_, _12426_, _06182_);
  not (_12429_, _12428_);
  nor (_12430_, _08659_, \oc8051_golden_model_1.PC [8]);
  nor (_12431_, _12430_, _12395_);
  and (_12432_, _12431_, _06182_);
  and (_12433_, _08661_, _06182_);
  nor (_12434_, _08661_, _06182_);
  nor (_12435_, _12434_, _12433_);
  not (_12436_, _12435_);
  and (_12437_, _08656_, _05929_);
  nor (_12438_, _12437_, \oc8051_golden_model_1.PC [6]);
  nor (_12439_, _12438_, _08658_);
  not (_12440_, _12439_);
  nor (_12441_, _12440_, _06317_);
  and (_12442_, _12440_, _06317_);
  nor (_12443_, _12442_, _12441_);
  and (_12444_, _05929_, \oc8051_golden_model_1.PC [4]);
  nor (_12445_, _12444_, \oc8051_golden_model_1.PC [5]);
  nor (_12446_, _12445_, _12437_);
  not (_12447_, _12446_);
  nor (_12448_, _12447_, _06611_);
  and (_12449_, _12447_, _06611_);
  nor (_12450_, _05929_, \oc8051_golden_model_1.PC [4]);
  nor (_12451_, _12450_, _12444_);
  not (_12452_, _12451_);
  nor (_12453_, _12452_, _06968_);
  nor (_12454_, _06213_, _06033_);
  and (_12455_, _06213_, _06033_);
  nor (_12456_, _06656_, _06085_);
  nor (_12457_, _07004_, \oc8051_golden_model_1.PC [1]);
  nor (_12458_, _06251_, _05630_);
  and (_12459_, _07004_, \oc8051_golden_model_1.PC [1]);
  nor (_12460_, _12459_, _12457_);
  and (_12461_, _12460_, _12458_);
  nor (_12462_, _12461_, _12457_);
  and (_12463_, _06656_, _06085_);
  nor (_12464_, _12463_, _12456_);
  not (_12465_, _12464_);
  nor (_12466_, _12465_, _12462_);
  nor (_12467_, _12466_, _12456_);
  nor (_12468_, _12467_, _12455_);
  nor (_12469_, _12468_, _12454_);
  and (_12470_, _12452_, _06968_);
  nor (_12471_, _12470_, _12453_);
  not (_12472_, _12471_);
  nor (_12473_, _12472_, _12469_);
  nor (_12474_, _12473_, _12453_);
  nor (_12475_, _12474_, _12449_);
  or (_12476_, _12475_, _12448_);
  and (_12477_, _12476_, _12443_);
  nor (_12478_, _12477_, _12441_);
  nor (_12479_, _12478_, _12436_);
  nor (_12480_, _12479_, _12433_);
  nor (_12481_, _12431_, _06182_);
  nor (_12482_, _12481_, _12432_);
  not (_12483_, _12482_);
  nor (_12484_, _12483_, _12480_);
  nor (_12485_, _12484_, _12432_);
  and (_12486_, _12485_, _12429_);
  or (_12487_, _12486_, _12427_);
  not (_12488_, _12487_);
  and (_12489_, _12488_, _12424_);
  nor (_12490_, _12489_, _12422_);
  nor (_12491_, _12490_, _12419_);
  or (_12492_, _12491_, _12418_);
  nor (_12493_, _12414_, _06182_);
  nor (_12494_, _12493_, _12415_);
  and (_12495_, _12494_, _12492_);
  nor (_12496_, _12495_, _12415_);
  and (_12497_, _12496_, _12412_);
  or (_12498_, _12497_, _12410_);
  nor (_12499_, _12498_, _12407_);
  nor (_12500_, _12499_, _12404_);
  nor (_12501_, _09487_, _06182_);
  and (_12502_, _09487_, _06182_);
  nor (_12503_, _12502_, _12501_);
  and (_12504_, _12503_, _12500_);
  nor (_12505_, _12503_, _12500_);
  nor (_12506_, _12505_, _12504_);
  and (_12507_, _12392_, _12390_);
  or (_12508_, _12507_, _12506_);
  nand (_12509_, _12508_, _12394_);
  nand (_12510_, _12509_, _12387_);
  nor (_12511_, _10758_, _10768_);
  and (_12512_, _12511_, _10755_);
  nor (_12513_, _07486_, _06781_);
  and (_12514_, _12513_, _12512_);
  or (_12515_, _12514_, _12149_);
  not (_12516_, _12512_);
  nor (_12517_, _07141_, _06758_);
  or (_12518_, _12517_, _09487_);
  nor (_12519_, _07141_, \oc8051_golden_model_1.PC [15]);
  and (_12520_, _12519_, _07504_);
  nand (_12521_, _12520_, _12513_);
  and (_12522_, _12521_, _12518_);
  or (_12523_, _12522_, _12516_);
  and (_12524_, _12523_, _08654_);
  and (_12525_, _12524_, _12515_);
  nor (_12526_, _12525_, _07154_);
  and (_12527_, _12526_, _12510_);
  nor (_12528_, _12527_, _12386_);
  and (_12529_, _12528_, _07151_);
  and (_12530_, _08390_, _08340_);
  and (_12531_, _08762_, _12530_);
  and (_12532_, _08144_, _08042_);
  and (_12533_, _12532_, _08759_);
  nand (_12534_, _12533_, _12531_);
  or (_12535_, _12534_, _09478_);
  and (_12536_, _12533_, _12531_);
  or (_12537_, _12536_, _12380_);
  and (_12538_, _12537_, _12535_);
  and (_12539_, _12538_, _06341_);
  nor (_12540_, _06009_, _05973_);
  nor (_12541_, _12540_, _10775_);
  not (_12542_, _12541_);
  or (_12543_, _12542_, _12539_);
  or (_12544_, _12543_, _12529_);
  and (_12545_, _06466_, _06010_);
  not (_12546_, _12545_);
  nor (_12547_, _12541_, _12149_);
  nor (_12548_, _12547_, _12546_);
  nand (_12549_, _12548_, _12544_);
  and (_12550_, _10743_, _07175_);
  not (_12551_, _12550_);
  nor (_12552_, _12545_, _12388_);
  nor (_12553_, _12552_, _12551_);
  nand (_12554_, _12553_, _12549_);
  nor (_12555_, _12550_, _12149_);
  nor (_12556_, _12555_, _06464_);
  and (_12557_, _12556_, _12554_);
  or (_12558_, _12557_, _12384_);
  nor (_12559_, _06012_, _05973_);
  nor (_12560_, _12559_, _10811_);
  nand (_12561_, _12560_, _12558_);
  nor (_12562_, _12560_, _12385_);
  not (_12563_, _06013_);
  nor (_12564_, _06267_, _12563_);
  and (_12565_, _12564_, _06269_);
  not (_12566_, _12565_);
  nor (_12567_, _12566_, _12562_);
  nand (_12568_, _12567_, _12561_);
  nor (_12569_, _12565_, _09487_);
  not (_12570_, _12569_);
  and (_12571_, _12570_, _12378_);
  and (_12572_, _12571_, _12568_);
  or (_12573_, _12572_, _12383_);
  nor (_12574_, _12573_, _06347_);
  or (_12575_, _12574_, _06480_);
  nor (_12576_, _12575_, _12338_);
  nor (_12577_, _11256_, _11255_);
  nor (_12578_, _12577_, _11259_);
  not (_12579_, _11262_);
  nor (_12580_, _08390_, \oc8051_golden_model_1.ACC [0]);
  or (_12581_, _12580_, _11263_);
  and (_12582_, _12581_, _12579_);
  and (_12583_, _12582_, _12578_);
  nor (_12584_, _11250_, _11254_);
  nor (_12585_, _11247_, _08575_);
  and (_12586_, _12585_, _12584_);
  and (_12587_, _12586_, _12583_);
  nor (_12588_, _12587_, _12303_);
  and (_12589_, _12587_, _09478_);
  nor (_12590_, _12589_, _12588_);
  nor (_12591_, _12590_, _06774_);
  or (_12592_, _12591_, _12576_);
  nand (_12593_, _12592_, _12176_);
  nor (_12594_, _11296_, _11297_);
  nor (_12595_, _12594_, _11300_);
  and (_12596_, _06251_, _06097_);
  nor (_12597_, _12596_, _11302_);
  nor (_12598_, _11306_, _12597_);
  and (_12599_, _12598_, _12595_);
  nor (_12600_, _11290_, _11291_);
  nor (_12601_, _12600_, _11295_);
  nor (_12602_, _11289_, _10961_);
  and (_12603_, _12602_, _12601_);
  and (_12604_, _12603_, _12599_);
  nand (_12605_, _12604_, _09478_);
  or (_12606_, _12604_, _12303_);
  and (_12607_, _12606_, _12605_);
  or (_12608_, _12607_, _12176_);
  nand (_12609_, _12608_, _12593_);
  nand (_12610_, _12609_, _12175_);
  and (_12611_, _12174_, _12149_);
  not (_12612_, _12611_);
  not (_12613_, _06007_);
  nor (_12614_, _06261_, _12613_);
  nor (_12615_, _06355_, _06019_);
  nor (_12616_, _07399_, _12615_);
  and (_12617_, _12616_, _12614_);
  not (_12618_, _06492_);
  nor (_12619_, _06495_, _06455_);
  and (_12620_, _12619_, _12618_);
  nor (_12621_, _07197_, _07398_);
  and (_12622_, _12621_, _12620_);
  and (_12623_, _12622_, _12617_);
  and (_12624_, _12623_, _12612_);
  nand (_12625_, _12624_, _12610_);
  nor (_12626_, _12623_, _09487_);
  nor (_12627_, _06019_, _05981_);
  not (_12628_, _12627_);
  nor (_12629_, _11561_, _09531_);
  and (_12630_, _12629_, _12628_);
  not (_12631_, _12630_);
  nor (_12632_, _12631_, _12626_);
  nand (_12633_, _12632_, _12625_);
  nor (_12634_, _12630_, _12385_);
  and (_12635_, _06506_, _06020_);
  not (_12636_, _12635_);
  nor (_12637_, _12636_, _12634_);
  and (_12638_, _12637_, _12633_);
  and (_12639_, _10735_, _10588_);
  or (_12640_, _12635_, _09487_);
  nand (_12641_, _12640_, _12639_);
  or (_12642_, _12641_, _12638_);
  nor (_12643_, _10516_, _06512_);
  not (_12644_, _12643_);
  nor (_12645_, _12639_, _12385_);
  nor (_12646_, _12645_, _12644_);
  nand (_12647_, _12646_, _12642_);
  nor (_12648_, _12643_, _09487_);
  nor (_12649_, _12648_, _10515_);
  nand (_12650_, _12649_, _12647_);
  nor (_12651_, _12385_, _05984_);
  nor (_12652_, _06257_, _06254_);
  not (_12653_, _12652_);
  nor (_12654_, _12653_, _12651_);
  nand (_12655_, _12654_, _12650_);
  nor (_12656_, _12652_, _09487_);
  nor (_12657_, _12656_, _06373_);
  nand (_12658_, _12657_, _12655_);
  not (_12659_, _07216_);
  and (_12660_, _09478_, _06373_);
  nor (_12661_, _12660_, _12659_);
  nand (_12662_, _12661_, _12658_);
  nor (_12663_, _09487_, _07216_);
  nor (_12664_, _12663_, _10094_);
  and (_12665_, _12664_, _12662_);
  or (_12666_, _12665_, _12173_);
  nand (_12667_, _12666_, _12172_);
  not (_12668_, _05946_);
  nor (_12669_, _06323_, _12668_);
  not (_12670_, _12669_);
  nor (_12671_, _12172_, _12385_);
  nor (_12672_, _12671_, _12670_);
  nand (_12673_, _12672_, _12667_);
  and (_12674_, _05944_, _05926_);
  nor (_12675_, _12669_, _09487_);
  nor (_12676_, _12675_, _12674_);
  nand (_12678_, _12676_, _12673_);
  not (_12679_, _12674_);
  nor (_12680_, _12679_, _12506_);
  nor (_12681_, _12680_, _09031_);
  and (_12682_, _12681_, _12678_);
  or (_12683_, _12682_, _12171_);
  nand (_12684_, _12683_, _06219_);
  and (_12685_, _09479_, _06218_);
  nor (_12686_, _12685_, _10929_);
  and (_12687_, _12686_, _12684_);
  and (_12688_, _10929_, _09487_);
  or (_12689_, _12688_, _12687_);
  nor (_12690_, _05973_, _05951_);
  not (_12691_, _12690_);
  nand (_12692_, _12691_, _12689_);
  not (_12693_, \oc8051_golden_model_1.DPH [0]);
  and (_12694_, \oc8051_golden_model_1.DPL [7], \oc8051_golden_model_1.ACC [7]);
  nor (_12695_, \oc8051_golden_model_1.DPL [7], \oc8051_golden_model_1.ACC [7]);
  and (_12696_, \oc8051_golden_model_1.DPL [6], \oc8051_golden_model_1.ACC [6]);
  nor (_12697_, \oc8051_golden_model_1.DPL [6], \oc8051_golden_model_1.ACC [6]);
  nor (_12699_, _12697_, _12696_);
  not (_12700_, _12699_);
  and (_12701_, \oc8051_golden_model_1.DPL [5], \oc8051_golden_model_1.ACC [5]);
  nor (_12702_, \oc8051_golden_model_1.DPL [5], \oc8051_golden_model_1.ACC [5]);
  nor (_12703_, _12702_, _12701_);
  not (_12704_, _12703_);
  and (_12705_, \oc8051_golden_model_1.DPL [4], \oc8051_golden_model_1.ACC [4]);
  nor (_12706_, _06001_, _05997_);
  nor (_12707_, \oc8051_golden_model_1.DPL [4], \oc8051_golden_model_1.ACC [4]);
  nor (_12708_, _12707_, _12705_);
  not (_12709_, _12708_);
  nor (_12710_, _12709_, _12706_);
  nor (_12711_, _12710_, _12705_);
  nor (_12712_, _12711_, _12704_);
  nor (_12713_, _12712_, _12701_);
  nor (_12714_, _12713_, _12700_);
  nor (_12715_, _12714_, _12696_);
  nor (_12716_, _12715_, _12695_);
  nor (_12717_, _12716_, _12694_);
  nor (_12718_, _12717_, _12693_);
  and (_12719_, _12718_, \oc8051_golden_model_1.DPH [1]);
  and (_12720_, _12719_, \oc8051_golden_model_1.DPH [2]);
  and (_12721_, _12720_, \oc8051_golden_model_1.DPH [3]);
  and (_12722_, _12721_, \oc8051_golden_model_1.DPH [4]);
  and (_12723_, _12722_, \oc8051_golden_model_1.DPH [5]);
  and (_12724_, _12723_, \oc8051_golden_model_1.DPH [6]);
  and (_12725_, _12724_, \oc8051_golden_model_1.DPH [7]);
  nor (_12726_, _12724_, \oc8051_golden_model_1.DPH [7]);
  nor (_12727_, _12726_, _12725_);
  and (_12728_, _12727_, _12690_);
  nor (_12729_, _06322_, _06217_);
  not (_12730_, _12729_);
  nor (_12731_, _12730_, _12728_);
  nand (_12732_, _12731_, _12692_);
  and (_12733_, _06321_, _05926_);
  nor (_12734_, _12729_, _09487_);
  nor (_12735_, _12734_, _12733_);
  nand (_12736_, _12735_, _12732_);
  not (_12737_, _12169_);
  and (_12738_, _11342_, _09487_);
  nor (_12739_, _12506_, _11342_);
  or (_12740_, _12739_, _12738_);
  and (_12741_, _12740_, _12733_);
  nor (_12742_, _12741_, _12737_);
  and (_12743_, _12742_, _12736_);
  or (_12744_, _12743_, _12170_);
  nand (_12745_, _12744_, _12166_);
  nor (_12746_, _12166_, _09487_);
  nor (_12747_, _12746_, _06369_);
  nand (_12748_, _12747_, _12745_);
  and (_12749_, _09478_, _06369_);
  not (_12750_, _05955_);
  nor (_12751_, _06536_, _12750_);
  not (_12752_, _12751_);
  nor (_12753_, _12752_, _12749_);
  nand (_12754_, _12753_, _12748_);
  and (_12755_, _06535_, _05926_);
  nor (_12756_, _12751_, _09487_);
  nor (_12757_, _12756_, _12755_);
  nand (_12758_, _12757_, _12754_);
  not (_12759_, _11342_);
  and (_12760_, _12759_, _09487_);
  nor (_12761_, _12506_, _12759_);
  or (_12762_, _12761_, _12760_);
  and (_12763_, _12762_, _12755_);
  nor (_12764_, _12763_, _10980_);
  and (_12765_, _12764_, _12758_);
  or (_12766_, _12765_, _12165_);
  nand (_12767_, _12766_, _12164_);
  nor (_12768_, _12164_, _09487_);
  nor (_12769_, _12768_, _06375_);
  nand (_12770_, _12769_, _12767_);
  and (_12771_, _09478_, _06375_);
  nor (_12772_, _06545_, _07233_);
  not (_12773_, _12772_);
  nor (_12774_, _12773_, _12771_);
  nand (_12775_, _12774_, _12770_);
  and (_12776_, _06544_, _05926_);
  nor (_12777_, _12772_, _09487_);
  nor (_12778_, _12777_, _12776_);
  nand (_12779_, _12778_, _12775_);
  not (_12780_, _12162_);
  and (_12781_, _12506_, _10558_);
  not (_12782_, _12776_);
  nor (_12783_, _09487_, _10558_);
  nor (_12784_, _12783_, _12782_);
  not (_12785_, _12784_);
  nor (_12786_, _12785_, _12781_);
  nor (_12787_, _12786_, _12780_);
  and (_12788_, _12787_, _12779_);
  or (_12789_, _12788_, _12163_);
  nand (_12790_, _12789_, _11022_);
  nor (_12791_, _11022_, _09487_);
  nor (_12792_, _12791_, _06366_);
  nand (_12793_, _12792_, _12790_);
  and (_12794_, _09478_, _06366_);
  not (_12795_, _05966_);
  nor (_12796_, _06528_, _12795_);
  not (_12797_, _12796_);
  nor (_12798_, _12797_, _12794_);
  nand (_12799_, _12798_, _12793_);
  and (_12800_, _06527_, _05926_);
  nor (_12801_, _12796_, _09487_);
  nor (_12802_, _12801_, _12800_);
  nand (_12803_, _12802_, _12799_);
  not (_12804_, _12154_);
  and (_12805_, _09487_, _10558_);
  nor (_12806_, _12506_, _10558_);
  or (_12807_, _12806_, _12805_);
  and (_12808_, _12807_, _12800_);
  nor (_12809_, _12808_, _12804_);
  and (_12810_, _12809_, _12803_);
  or (_12811_, _12810_, _12155_);
  nand (_12812_, _12811_, _12153_);
  nor (_12813_, _12153_, _09487_);
  nor (_12814_, _12813_, _11125_);
  and (_12815_, _12814_, _12812_);
  and (_12816_, _12149_, _11125_);
  or (_12817_, _12816_, _06551_);
  nor (_12818_, _12817_, _12815_);
  and (_12819_, _08040_, _06551_);
  or (_12820_, _12819_, _12818_);
  nand (_12821_, _12820_, _05959_);
  nor (_12822_, _09487_, _05959_);
  nor (_12823_, _12822_, _06365_);
  nand (_12824_, _12823_, _12821_);
  not (_12825_, _07959_);
  and (_12826_, _07948_, \oc8051_golden_model_1.P0 [2]);
  and (_12827_, _08616_, \oc8051_golden_model_1.TCON [2]);
  and (_12828_, _08620_, \oc8051_golden_model_1.P1 [2]);
  and (_12829_, _08622_, \oc8051_golden_model_1.SCON [2]);
  and (_12830_, _08624_, \oc8051_golden_model_1.P2 [2]);
  and (_12831_, _08626_, \oc8051_golden_model_1.IE [2]);
  and (_12832_, _08628_, \oc8051_golden_model_1.P3 [2]);
  and (_12833_, _08632_, \oc8051_golden_model_1.IP [2]);
  and (_12834_, _08630_, \oc8051_golden_model_1.PSW [2]);
  and (_12835_, _08636_, \oc8051_golden_model_1.ACC [2]);
  and (_12836_, _08634_, \oc8051_golden_model_1.B [2]);
  or (_12837_, _12836_, _12835_);
  or (_12838_, _12837_, _12834_);
  or (_12839_, _12838_, _12833_);
  or (_12840_, _12839_, _12832_);
  or (_12841_, _12840_, _12831_);
  or (_12842_, _12841_, _12830_);
  or (_12843_, _12842_, _12829_);
  or (_12844_, _12843_, _12828_);
  or (_12845_, _12844_, _12827_);
  nor (_12846_, _12845_, _12826_);
  and (_12847_, _12846_, _08438_);
  nor (_12848_, _12847_, _12825_);
  not (_12849_, _08172_);
  and (_12850_, _07948_, \oc8051_golden_model_1.P0 [1]);
  and (_12851_, _08616_, \oc8051_golden_model_1.TCON [1]);
  and (_12852_, _08620_, \oc8051_golden_model_1.P1 [1]);
  and (_12853_, _08622_, \oc8051_golden_model_1.SCON [1]);
  and (_12854_, _08624_, \oc8051_golden_model_1.P2 [1]);
  and (_12855_, _08626_, \oc8051_golden_model_1.IE [1]);
  and (_12856_, _08628_, \oc8051_golden_model_1.P3 [1]);
  and (_12857_, _08632_, \oc8051_golden_model_1.IP [1]);
  and (_12858_, _08630_, \oc8051_golden_model_1.PSW [1]);
  and (_12859_, _08636_, \oc8051_golden_model_1.ACC [1]);
  and (_12860_, _08634_, \oc8051_golden_model_1.B [1]);
  or (_12861_, _12860_, _12859_);
  or (_12862_, _12861_, _12858_);
  or (_12863_, _12862_, _12857_);
  or (_12864_, _12863_, _12856_);
  or (_12865_, _12864_, _12855_);
  or (_12866_, _12865_, _12854_);
  or (_12867_, _12866_, _12853_);
  or (_12868_, _12867_, _12852_);
  or (_12869_, _12868_, _12851_);
  nor (_12870_, _12869_, _12850_);
  and (_12871_, _12870_, _08339_);
  nor (_12872_, _12871_, _12849_);
  nor (_12873_, _12872_, _12848_);
  and (_12874_, _08628_, \oc8051_golden_model_1.P3 [4]);
  and (_12875_, _08626_, \oc8051_golden_model_1.IE [4]);
  nor (_12876_, _12875_, _12874_);
  and (_12877_, _08622_, \oc8051_golden_model_1.SCON [4]);
  and (_12878_, _08624_, \oc8051_golden_model_1.P2 [4]);
  nor (_12879_, _12878_, _12877_);
  and (_12880_, _12879_, _12876_);
  and (_12881_, _08630_, \oc8051_golden_model_1.PSW [4]);
  and (_12882_, _08632_, \oc8051_golden_model_1.IP [4]);
  and (_12883_, _08636_, \oc8051_golden_model_1.ACC [4]);
  and (_12884_, _08634_, \oc8051_golden_model_1.B [4]);
  or (_12885_, _12884_, _12883_);
  or (_12886_, _12885_, _12882_);
  nor (_12887_, _12886_, _12881_);
  and (_12888_, _08616_, \oc8051_golden_model_1.TCON [4]);
  and (_12889_, _07948_, \oc8051_golden_model_1.P0 [4]);
  and (_12890_, _08620_, \oc8051_golden_model_1.P1 [4]);
  or (_12891_, _12890_, _12889_);
  nor (_12892_, _12891_, _12888_);
  and (_12893_, _12892_, _12887_);
  and (_12894_, _12893_, _12880_);
  and (_12895_, _12894_, _08542_);
  and (_12896_, _07889_, _06657_);
  not (_12897_, _12896_);
  nor (_12898_, _12897_, _12895_);
  nor (_12899_, _12898_, _08788_);
  and (_12900_, _12899_, _12873_);
  and (_12901_, _07889_, _06656_);
  not (_12902_, _12901_);
  and (_12903_, _07948_, \oc8051_golden_model_1.P0 [0]);
  and (_12904_, _08616_, \oc8051_golden_model_1.TCON [0]);
  and (_12905_, _08620_, \oc8051_golden_model_1.P1 [0]);
  and (_12906_, _08622_, \oc8051_golden_model_1.SCON [0]);
  and (_12907_, _08624_, \oc8051_golden_model_1.P2 [0]);
  and (_12908_, _08626_, \oc8051_golden_model_1.IE [0]);
  and (_12909_, _08628_, \oc8051_golden_model_1.P3 [0]);
  and (_12910_, _08632_, \oc8051_golden_model_1.IP [0]);
  and (_12911_, _08630_, \oc8051_golden_model_1.PSW [0]);
  and (_12912_, _08636_, \oc8051_golden_model_1.ACC [0]);
  and (_12913_, _08634_, \oc8051_golden_model_1.B [0]);
  or (_12914_, _12913_, _12912_);
  or (_12915_, _12914_, _12911_);
  or (_12916_, _12915_, _12910_);
  or (_12917_, _12916_, _12909_);
  or (_12918_, _12917_, _12908_);
  or (_12919_, _12918_, _12907_);
  or (_12920_, _12919_, _12906_);
  or (_12921_, _12920_, _12905_);
  or (_12922_, _12921_, _12904_);
  nor (_12923_, _12922_, _12903_);
  not (_12924_, _12923_);
  nor (_12925_, _12924_, _08389_);
  nor (_12926_, _12925_, _12902_);
  and (_12927_, _08632_, \oc8051_golden_model_1.IP [6]);
  and (_12928_, _08622_, \oc8051_golden_model_1.SCON [6]);
  nor (_12929_, _12928_, _12927_);
  and (_12930_, _08630_, \oc8051_golden_model_1.PSW [6]);
  and (_12931_, _08634_, \oc8051_golden_model_1.B [6]);
  and (_12932_, _08636_, \oc8051_golden_model_1.ACC [6]);
  or (_12933_, _12932_, _12931_);
  nor (_12934_, _12933_, _12930_);
  and (_12935_, _08616_, \oc8051_golden_model_1.TCON [6]);
  and (_12936_, _07948_, \oc8051_golden_model_1.P0 [6]);
  and (_12937_, _08620_, \oc8051_golden_model_1.P1 [6]);
  or (_12938_, _12937_, _12936_);
  nor (_12939_, _12938_, _12935_);
  and (_12940_, _08624_, \oc8051_golden_model_1.P2 [6]);
  and (_12941_, _08628_, \oc8051_golden_model_1.P3 [6]);
  and (_12942_, _08626_, \oc8051_golden_model_1.IE [6]);
  or (_12943_, _12942_, _12941_);
  nor (_12944_, _12943_, _12940_);
  and (_12945_, _12944_, _12939_);
  and (_12946_, _12945_, _12934_);
  and (_12947_, _12946_, _12929_);
  and (_12948_, _12947_, _08143_);
  and (_12949_, _07917_, _06657_);
  not (_12950_, _12949_);
  nor (_12951_, _12950_, _12948_);
  nor (_12952_, _12951_, _12926_);
  not (_12953_, _08185_);
  and (_12954_, _07948_, \oc8051_golden_model_1.P0 [3]);
  and (_12955_, _08616_, \oc8051_golden_model_1.TCON [3]);
  and (_12956_, _08620_, \oc8051_golden_model_1.P1 [3]);
  and (_12957_, _08622_, \oc8051_golden_model_1.SCON [3]);
  and (_12958_, _08624_, \oc8051_golden_model_1.P2 [3]);
  and (_12959_, _08626_, \oc8051_golden_model_1.IE [3]);
  and (_12960_, _08628_, \oc8051_golden_model_1.P3 [3]);
  and (_12961_, _08632_, \oc8051_golden_model_1.IP [3]);
  and (_12962_, _08630_, \oc8051_golden_model_1.PSW [3]);
  and (_12963_, _08634_, \oc8051_golden_model_1.B [3]);
  and (_12964_, _08636_, \oc8051_golden_model_1.ACC [3]);
  or (_12965_, _12964_, _12963_);
  or (_12966_, _12965_, _12962_);
  or (_12967_, _12966_, _12961_);
  or (_12968_, _12967_, _12960_);
  or (_12969_, _12968_, _12959_);
  or (_12970_, _12969_, _12958_);
  or (_12971_, _12970_, _12957_);
  or (_12972_, _12971_, _12956_);
  or (_12973_, _12972_, _12955_);
  nor (_12974_, _12973_, _12954_);
  and (_12975_, _12974_, _08290_);
  nor (_12976_, _12975_, _12953_);
  and (_12977_, _07948_, \oc8051_golden_model_1.P0 [5]);
  and (_12978_, _08616_, \oc8051_golden_model_1.TCON [5]);
  and (_12979_, _08620_, \oc8051_golden_model_1.P1 [5]);
  and (_12980_, _08622_, \oc8051_golden_model_1.SCON [5]);
  and (_12981_, _08624_, \oc8051_golden_model_1.P2 [5]);
  and (_12982_, _08626_, \oc8051_golden_model_1.IE [5]);
  and (_12983_, _08628_, \oc8051_golden_model_1.P3 [5]);
  and (_12984_, _08632_, \oc8051_golden_model_1.IP [5]);
  and (_12985_, _08630_, \oc8051_golden_model_1.PSW [5]);
  and (_12986_, _08636_, \oc8051_golden_model_1.ACC [5]);
  and (_12987_, _08634_, \oc8051_golden_model_1.B [5]);
  or (_12988_, _12987_, _12986_);
  or (_12989_, _12988_, _12985_);
  or (_12990_, _12989_, _12984_);
  or (_12991_, _12990_, _12983_);
  or (_12992_, _12991_, _12982_);
  or (_12993_, _12992_, _12981_);
  or (_12994_, _12993_, _12980_);
  or (_12995_, _12994_, _12979_);
  or (_12996_, _12995_, _12978_);
  nor (_12997_, _12996_, _12977_);
  and (_12998_, _12997_, _08245_);
  and (_12999_, _07880_, _06657_);
  not (_13000_, _12999_);
  nor (_13001_, _13000_, _12998_);
  nor (_13002_, _13001_, _12976_);
  and (_13003_, _13002_, _12952_);
  and (_13004_, _13003_, _12900_);
  nor (_13005_, _09478_, _13004_);
  and (_13006_, _12303_, _13004_);
  or (_13007_, _13006_, _06558_);
  or (_13008_, _13007_, _13005_);
  and (_13009_, _13008_, _12151_);
  and (_13010_, _13009_, _12824_);
  or (_13011_, _13010_, _12152_);
  nor (_13012_, _11243_, _06283_);
  nand (_13013_, _13012_, _13011_);
  nor (_13014_, _13012_, _09487_);
  nor (_13015_, _13014_, _11284_);
  and (_13016_, _13015_, _13013_);
  and (_13017_, _12149_, _11284_);
  or (_13018_, _13017_, _06281_);
  nor (_13019_, _13018_, _13016_);
  and (_13020_, _08040_, _06281_);
  or (_13021_, _13020_, _13019_);
  nand (_13022_, _13021_, _05964_);
  nor (_13023_, _09487_, _05964_);
  nor (_13024_, _13023_, _06362_);
  nand (_13025_, _13024_, _13022_);
  nor (_13026_, _12380_, _13004_);
  and (_13027_, _09479_, _13004_);
  nor (_13028_, _13027_, _13026_);
  and (_13029_, _13028_, _06362_);
  and (_13030_, _08569_, _07264_);
  not (_13031_, _13030_);
  nor (_13032_, _13031_, _13029_);
  nand (_13033_, _13032_, _13025_);
  nor (_13034_, _13030_, _12149_);
  nor (_13035_, _13034_, _06568_);
  nand (_13036_, _13035_, _13033_);
  nor (_13037_, _11335_, _11330_);
  not (_13038_, _13037_);
  and (_13039_, _09487_, _06568_);
  nor (_13040_, _13039_, _13038_);
  nand (_13041_, _13040_, _13036_);
  nor (_13042_, _12149_, _13037_);
  nor (_13043_, _13042_, _06361_);
  nand (_13044_, _13043_, _13041_);
  and (_13045_, _06361_, _06182_);
  nor (_13046_, _13045_, _05940_);
  nand (_13047_, _13046_, _13044_);
  and (_13048_, _12388_, _05940_);
  nor (_13049_, _13048_, _05927_);
  nand (_13050_, _13049_, _13047_);
  and (_13051_, _13028_, _05927_);
  nor (_13052_, _09424_, _07281_);
  not (_13053_, _13052_);
  nor (_13054_, _13053_, _13051_);
  nand (_13055_, _13054_, _13050_);
  nor (_13056_, _13052_, _12149_);
  nor (_13057_, _13056_, _06278_);
  nand (_13058_, _13057_, _13055_);
  not (_13059_, _12141_);
  and (_13060_, _09487_, _06278_);
  nor (_13061_, _13060_, _13059_);
  and (_13062_, _13061_, _13058_);
  or (_13063_, _13062_, _12150_);
  nand (_13064_, _13063_, _12140_);
  nor (_13065_, _12140_, _06182_);
  nor (_13066_, _13065_, _05939_);
  nand (_13067_, _13066_, _13064_);
  and (_13068_, _05938_, _05926_);
  and (_13069_, _09487_, _05939_);
  nor (_13070_, _13069_, _13068_);
  and (_13071_, _13070_, _13067_);
  and (_13072_, _13068_, _12385_);
  nor (_13073_, _13072_, _13071_);
  or (_13074_, _13073_, _01351_);
  or (_13075_, _01347_, \oc8051_golden_model_1.PC [15]);
  and (_13076_, _13075_, _42618_);
  and (_40586_, _13076_, _13074_);
  not (_13077_, _07904_);
  and (_13078_, _13077_, \oc8051_golden_model_1.P2 [7]);
  and (_13079_, _08575_, _07904_);
  or (_13080_, _13079_, _13078_);
  and (_13081_, _13080_, _06536_);
  nor (_13082_, _08040_, _13077_);
  or (_13083_, _13082_, _13078_);
  or (_13084_, _13083_, _07215_);
  not (_13085_, _08624_);
  and (_13086_, _13085_, \oc8051_golden_model_1.P2 [7]);
  and (_13087_, _08649_, _08624_);
  or (_13088_, _13087_, _13086_);
  and (_13089_, _13088_, _06268_);
  and (_13090_, _08768_, _07904_);
  or (_13091_, _13090_, _13078_);
  or (_13092_, _13091_, _07151_);
  and (_13093_, _07904_, \oc8051_golden_model_1.ACC [7]);
  or (_13094_, _13093_, _13078_);
  and (_13095_, _13094_, _07141_);
  and (_13096_, _07142_, \oc8051_golden_model_1.P2 [7]);
  or (_13097_, _13096_, _06341_);
  or (_13098_, _13097_, _13095_);
  and (_13099_, _13098_, _06273_);
  and (_13100_, _13099_, _13092_);
  and (_13101_, _08773_, _08624_);
  or (_13102_, _13101_, _13086_);
  and (_13103_, _13102_, _06272_);
  or (_13104_, _13103_, _06461_);
  or (_13105_, _13104_, _13100_);
  or (_13106_, _13083_, _07166_);
  and (_13107_, _13106_, _13105_);
  or (_13108_, _13107_, _06464_);
  or (_13109_, _13094_, _06465_);
  and (_13110_, _13109_, _06269_);
  and (_13111_, _13110_, _13108_);
  or (_13112_, _13111_, _13089_);
  and (_13113_, _13112_, _06262_);
  or (_13114_, _13086_, _08789_);
  and (_13115_, _13114_, _06261_);
  and (_13116_, _13115_, _13102_);
  or (_13117_, _13116_, _13113_);
  and (_13118_, _13117_, _06258_);
  and (_13119_, _08808_, _08624_);
  or (_13120_, _13119_, _13086_);
  and (_13121_, _13120_, _06257_);
  or (_13122_, _13121_, _10080_);
  or (_13123_, _13122_, _13118_);
  and (_13124_, _13123_, _13084_);
  or (_13125_, _13124_, _07460_);
  and (_13126_, _08755_, _07904_);
  or (_13127_, _13078_, _07208_);
  or (_13128_, _13127_, _13126_);
  and (_13129_, _13128_, _05982_);
  and (_13130_, _13129_, _13125_);
  and (_13131_, _09021_, _07904_);
  or (_13132_, _13131_, _13078_);
  and (_13133_, _13132_, _10094_);
  or (_13134_, _13133_, _06218_);
  or (_13135_, _13134_, _13130_);
  and (_13136_, _08825_, _07904_);
  or (_13137_, _13136_, _13078_);
  or (_13138_, _13137_, _06219_);
  and (_13139_, _13138_, _13135_);
  or (_13140_, _13139_, _06369_);
  and (_13141_, _09044_, _07904_);
  or (_13142_, _13141_, _13078_);
  or (_13143_, _13142_, _07237_);
  and (_13144_, _13143_, _07240_);
  and (_13145_, _13144_, _13140_);
  or (_13146_, _13145_, _13081_);
  and (_13147_, _13146_, _07242_);
  or (_13148_, _13078_, _08043_);
  and (_13149_, _13137_, _06375_);
  and (_13150_, _13149_, _13148_);
  or (_13151_, _13150_, _13147_);
  and (_13152_, _13151_, _07234_);
  and (_13153_, _13094_, _06545_);
  and (_13154_, _13153_, _13148_);
  or (_13155_, _13154_, _06366_);
  or (_13156_, _13155_, _13152_);
  nor (_13157_, _09043_, _13077_);
  or (_13158_, _13078_, _09056_);
  or (_13159_, _13158_, _13157_);
  and (_13160_, _13159_, _09061_);
  and (_13161_, _13160_, _13156_);
  nor (_13162_, _08573_, _13077_);
  or (_13163_, _13162_, _13078_);
  and (_13164_, _13163_, _06528_);
  or (_13165_, _13164_, _06568_);
  or (_13166_, _13165_, _13161_);
  or (_13167_, _13091_, _06926_);
  and (_13168_, _13167_, _05928_);
  and (_13169_, _13168_, _13166_);
  and (_13170_, _13088_, _05927_);
  or (_13171_, _13170_, _06278_);
  or (_13172_, _13171_, _13169_);
  and (_13173_, _08550_, _07904_);
  or (_13174_, _13078_, _06279_);
  or (_13175_, _13174_, _13173_);
  and (_13176_, _13175_, _01347_);
  and (_13177_, _13176_, _13172_);
  nor (_13178_, \oc8051_golden_model_1.P2 [7], rst);
  nor (_13179_, _13178_, _01354_);
  or (_40587_, _13179_, _13177_);
  not (_13180_, _07894_);
  and (_13181_, _13180_, \oc8051_golden_model_1.P3 [7]);
  and (_13182_, _08575_, _07894_);
  or (_13183_, _13182_, _13181_);
  and (_13184_, _13183_, _06536_);
  nor (_13185_, _08040_, _13180_);
  or (_13186_, _13185_, _13181_);
  or (_13187_, _13186_, _07215_);
  not (_13188_, _08628_);
  and (_13189_, _13188_, \oc8051_golden_model_1.P3 [7]);
  and (_13190_, _08649_, _08628_);
  or (_13191_, _13190_, _13189_);
  and (_13192_, _13191_, _06268_);
  and (_13193_, _08768_, _07894_);
  or (_13194_, _13193_, _13181_);
  or (_13195_, _13194_, _07151_);
  and (_13196_, _07894_, \oc8051_golden_model_1.ACC [7]);
  or (_13197_, _13196_, _13181_);
  and (_13198_, _13197_, _07141_);
  and (_13199_, _07142_, \oc8051_golden_model_1.P3 [7]);
  or (_13200_, _13199_, _06341_);
  or (_13201_, _13200_, _13198_);
  and (_13202_, _13201_, _06273_);
  and (_13203_, _13202_, _13195_);
  and (_13204_, _08773_, _08628_);
  or (_13205_, _13204_, _13189_);
  and (_13206_, _13205_, _06272_);
  or (_13207_, _13206_, _06461_);
  or (_13208_, _13207_, _13203_);
  or (_13209_, _13186_, _07166_);
  and (_13210_, _13209_, _13208_);
  or (_13211_, _13210_, _06464_);
  or (_13212_, _13197_, _06465_);
  and (_13213_, _13212_, _06269_);
  and (_13214_, _13213_, _13211_);
  or (_13215_, _13214_, _13192_);
  and (_13216_, _13215_, _06262_);
  and (_13217_, _08790_, _08628_);
  or (_13218_, _13217_, _13189_);
  and (_13219_, _13218_, _06261_);
  or (_13220_, _13219_, _13216_);
  and (_13221_, _13220_, _06258_);
  and (_13222_, _08808_, _08628_);
  or (_13223_, _13222_, _13189_);
  and (_13224_, _13223_, _06257_);
  or (_13225_, _13224_, _10080_);
  or (_13226_, _13225_, _13221_);
  and (_13227_, _13226_, _13187_);
  or (_13228_, _13227_, _07460_);
  and (_13229_, _08755_, _07894_);
  or (_13230_, _13181_, _07208_);
  or (_13231_, _13230_, _13229_);
  and (_13232_, _13231_, _05982_);
  and (_13233_, _13232_, _13228_);
  and (_13234_, _09021_, _07894_);
  or (_13235_, _13234_, _13181_);
  and (_13236_, _13235_, _10094_);
  or (_13237_, _13236_, _06218_);
  or (_13238_, _13237_, _13233_);
  and (_13239_, _08825_, _07894_);
  or (_13240_, _13239_, _13181_);
  or (_13241_, _13240_, _06219_);
  and (_13242_, _13241_, _13238_);
  or (_13243_, _13242_, _06369_);
  and (_13244_, _09044_, _07894_);
  or (_13245_, _13244_, _13181_);
  or (_13246_, _13245_, _07237_);
  and (_13247_, _13246_, _07240_);
  and (_13248_, _13247_, _13243_);
  or (_13249_, _13248_, _13184_);
  and (_13250_, _13249_, _07242_);
  or (_13251_, _13181_, _08043_);
  and (_13252_, _13240_, _06375_);
  and (_13253_, _13252_, _13251_);
  or (_13254_, _13253_, _13250_);
  and (_13255_, _13254_, _07234_);
  and (_13256_, _13197_, _06545_);
  and (_13257_, _13256_, _13251_);
  or (_13258_, _13257_, _06366_);
  or (_13259_, _13258_, _13255_);
  nor (_13260_, _09043_, _13180_);
  or (_13261_, _13181_, _09056_);
  or (_13262_, _13261_, _13260_);
  and (_13263_, _13262_, _09061_);
  and (_13264_, _13263_, _13259_);
  nor (_13265_, _08573_, _13180_);
  or (_13266_, _13265_, _13181_);
  and (_13267_, _13266_, _06528_);
  or (_13268_, _13267_, _06568_);
  or (_13269_, _13268_, _13264_);
  or (_13270_, _13194_, _06926_);
  and (_13271_, _13270_, _05928_);
  and (_13272_, _13271_, _13269_);
  and (_13273_, _13191_, _05927_);
  or (_13274_, _13273_, _06278_);
  or (_13275_, _13274_, _13272_);
  and (_13276_, _08550_, _07894_);
  or (_13277_, _13181_, _06279_);
  or (_13278_, _13277_, _13276_);
  and (_13279_, _13278_, _01347_);
  and (_13280_, _13279_, _13275_);
  nor (_13281_, \oc8051_golden_model_1.P3 [7], rst);
  nor (_13282_, _13281_, _01354_);
  or (_40588_, _13282_, _13280_);
  not (_13283_, _07926_);
  and (_13284_, _13283_, \oc8051_golden_model_1.P0 [7]);
  and (_13285_, _08575_, _07926_);
  or (_13286_, _13285_, _13284_);
  and (_13287_, _13286_, _06536_);
  nor (_13288_, _08040_, _13283_);
  or (_13289_, _13288_, _13284_);
  or (_13290_, _13289_, _07215_);
  not (_13291_, _07948_);
  and (_13292_, _13291_, \oc8051_golden_model_1.P0 [7]);
  and (_13293_, _08649_, _07948_);
  or (_13294_, _13293_, _13292_);
  and (_13295_, _13294_, _06268_);
  and (_13296_, _08768_, _07926_);
  or (_13297_, _13296_, _13284_);
  or (_13298_, _13297_, _07151_);
  and (_13299_, _07926_, \oc8051_golden_model_1.ACC [7]);
  or (_13300_, _13299_, _13284_);
  and (_13301_, _13300_, _07141_);
  and (_13302_, _07142_, \oc8051_golden_model_1.P0 [7]);
  or (_13303_, _13302_, _06341_);
  or (_13304_, _13303_, _13301_);
  and (_13305_, _13304_, _06273_);
  and (_13306_, _13305_, _13298_);
  and (_13307_, _08773_, _07948_);
  or (_13308_, _13307_, _13292_);
  and (_13309_, _13308_, _06272_);
  or (_13310_, _13309_, _06461_);
  or (_13311_, _13310_, _13306_);
  or (_13312_, _13289_, _07166_);
  and (_13313_, _13312_, _13311_);
  or (_13314_, _13313_, _06464_);
  or (_13315_, _13300_, _06465_);
  and (_13316_, _13315_, _06269_);
  and (_13317_, _13316_, _13314_);
  or (_13318_, _13317_, _13295_);
  and (_13319_, _13318_, _06262_);
  and (_13320_, _08790_, _07948_);
  or (_13321_, _13320_, _13292_);
  and (_13322_, _13321_, _06261_);
  or (_13323_, _13322_, _13319_);
  and (_13324_, _13323_, _06258_);
  and (_13325_, _08808_, _07948_);
  or (_13326_, _13325_, _13292_);
  and (_13327_, _13326_, _06257_);
  or (_13328_, _13327_, _10080_);
  or (_13329_, _13328_, _13324_);
  and (_13330_, _13329_, _13290_);
  or (_13331_, _13330_, _07460_);
  and (_13332_, _08755_, _07926_);
  or (_13333_, _13284_, _07208_);
  or (_13334_, _13333_, _13332_);
  and (_13335_, _13334_, _05982_);
  and (_13336_, _13335_, _13331_);
  and (_13337_, _09021_, _07926_);
  or (_13338_, _13337_, _13284_);
  and (_13339_, _13338_, _10094_);
  or (_13340_, _13339_, _06218_);
  or (_13341_, _13340_, _13336_);
  and (_13342_, _08825_, _07926_);
  or (_13343_, _13342_, _13284_);
  or (_13344_, _13343_, _06219_);
  and (_13345_, _13344_, _13341_);
  or (_13346_, _13345_, _06369_);
  and (_13347_, _09044_, _07926_);
  or (_13348_, _13347_, _13284_);
  or (_13349_, _13348_, _07237_);
  and (_13350_, _13349_, _07240_);
  and (_13351_, _13350_, _13346_);
  or (_13352_, _13351_, _13287_);
  and (_13353_, _13352_, _07242_);
  or (_13354_, _13284_, _08043_);
  and (_13355_, _13343_, _06375_);
  and (_13356_, _13355_, _13354_);
  or (_13357_, _13356_, _13353_);
  and (_13358_, _13357_, _07234_);
  and (_13359_, _13300_, _06545_);
  and (_13360_, _13359_, _13354_);
  or (_13361_, _13360_, _06366_);
  or (_13362_, _13361_, _13358_);
  nor (_13363_, _09043_, _13283_);
  or (_13364_, _13284_, _09056_);
  or (_13365_, _13364_, _13363_);
  and (_13366_, _13365_, _09061_);
  and (_13367_, _13366_, _13362_);
  nor (_13368_, _08573_, _13283_);
  or (_13369_, _13368_, _13284_);
  and (_13370_, _13369_, _06528_);
  or (_13371_, _13370_, _06568_);
  or (_13372_, _13371_, _13367_);
  or (_13373_, _13297_, _06926_);
  and (_13374_, _13373_, _05928_);
  and (_13375_, _13374_, _13372_);
  and (_13376_, _13294_, _05927_);
  or (_13377_, _13376_, _06278_);
  or (_13378_, _13377_, _13375_);
  and (_13379_, _08550_, _07926_);
  or (_13380_, _13284_, _06279_);
  or (_13381_, _13380_, _13379_);
  and (_13382_, _13381_, _01347_);
  and (_13383_, _13382_, _13378_);
  nor (_13384_, \oc8051_golden_model_1.P0 [7], rst);
  nor (_13385_, _13384_, _01354_);
  or (_40589_, _13385_, _13383_);
  nor (_13386_, \oc8051_golden_model_1.P1 [7], rst);
  nor (_13387_, _13386_, _01354_);
  not (_13388_, _07971_);
  and (_13389_, _13388_, \oc8051_golden_model_1.P1 [7]);
  and (_13390_, _08575_, _07971_);
  or (_13391_, _13390_, _13389_);
  and (_13392_, _13391_, _06536_);
  nor (_13393_, _08040_, _13388_);
  or (_13394_, _13393_, _13389_);
  or (_13395_, _13394_, _07215_);
  not (_13396_, _08620_);
  and (_13397_, _13396_, \oc8051_golden_model_1.P1 [7]);
  and (_13398_, _08649_, _08620_);
  or (_13399_, _13398_, _13397_);
  and (_13400_, _13399_, _06268_);
  and (_13401_, _08768_, _07971_);
  or (_13402_, _13401_, _13389_);
  or (_13403_, _13402_, _07151_);
  and (_13404_, _07971_, \oc8051_golden_model_1.ACC [7]);
  or (_13405_, _13404_, _13389_);
  and (_13406_, _13405_, _07141_);
  and (_13407_, _07142_, \oc8051_golden_model_1.P1 [7]);
  or (_13408_, _13407_, _06341_);
  or (_13409_, _13408_, _13406_);
  and (_13410_, _13409_, _06273_);
  and (_13411_, _13410_, _13403_);
  and (_13412_, _08773_, _08620_);
  or (_13413_, _13412_, _13397_);
  and (_13414_, _13413_, _06272_);
  or (_13415_, _13414_, _06461_);
  or (_13416_, _13415_, _13411_);
  or (_13417_, _13394_, _07166_);
  and (_13418_, _13417_, _13416_);
  or (_13419_, _13418_, _06464_);
  or (_13420_, _13405_, _06465_);
  and (_13421_, _13420_, _06269_);
  and (_13422_, _13421_, _13419_);
  or (_13423_, _13422_, _13400_);
  and (_13424_, _13423_, _06262_);
  or (_13425_, _13397_, _08789_);
  and (_13426_, _13425_, _06261_);
  and (_13427_, _13426_, _13413_);
  or (_13428_, _13427_, _13424_);
  and (_13429_, _13428_, _06258_);
  and (_13430_, _08808_, _08620_);
  or (_13431_, _13430_, _13397_);
  and (_13432_, _13431_, _06257_);
  or (_13433_, _13432_, _10080_);
  or (_13434_, _13433_, _13429_);
  and (_13435_, _13434_, _13395_);
  or (_13436_, _13435_, _07460_);
  and (_13437_, _08755_, _07971_);
  or (_13438_, _13389_, _07208_);
  or (_13439_, _13438_, _13437_);
  and (_13440_, _13439_, _05982_);
  and (_13441_, _13440_, _13436_);
  and (_13442_, _09021_, _07971_);
  or (_13443_, _13442_, _13389_);
  and (_13444_, _13443_, _10094_);
  or (_13445_, _13444_, _06218_);
  or (_13446_, _13445_, _13441_);
  and (_13447_, _08825_, _07971_);
  or (_13448_, _13447_, _13389_);
  or (_13449_, _13448_, _06219_);
  and (_13450_, _13449_, _13446_);
  or (_13451_, _13450_, _06369_);
  and (_13452_, _09044_, _07971_);
  or (_13453_, _13452_, _13389_);
  or (_13454_, _13453_, _07237_);
  and (_13455_, _13454_, _07240_);
  and (_13456_, _13455_, _13451_);
  or (_13457_, _13456_, _13392_);
  and (_13458_, _13457_, _07242_);
  or (_13459_, _13389_, _08043_);
  and (_13460_, _13448_, _06375_);
  and (_13461_, _13460_, _13459_);
  or (_13462_, _13461_, _13458_);
  and (_13463_, _13462_, _07234_);
  and (_13464_, _13405_, _06545_);
  and (_13465_, _13464_, _13459_);
  or (_13466_, _13465_, _06366_);
  or (_13467_, _13466_, _13463_);
  nor (_13468_, _09043_, _13388_);
  or (_13469_, _13389_, _09056_);
  or (_13470_, _13469_, _13468_);
  and (_13471_, _13470_, _09061_);
  and (_13472_, _13471_, _13467_);
  nor (_13473_, _08573_, _13388_);
  or (_13474_, _13473_, _13389_);
  and (_13475_, _13474_, _06528_);
  or (_13476_, _13475_, _06568_);
  or (_13477_, _13476_, _13472_);
  or (_13478_, _13402_, _06926_);
  and (_13479_, _13478_, _05928_);
  and (_13480_, _13479_, _13477_);
  and (_13481_, _13399_, _05927_);
  or (_13482_, _13481_, _06278_);
  or (_13483_, _13482_, _13480_);
  and (_13484_, _08550_, _07971_);
  or (_13485_, _13389_, _06279_);
  or (_13486_, _13485_, _13484_);
  and (_13487_, _13486_, _01347_);
  and (_13488_, _13487_, _13483_);
  or (_40591_, _13488_, _13387_);
  and (_13489_, _01351_, \oc8051_golden_model_1.IP [7]);
  not (_13490_, _07946_);
  and (_13491_, _13490_, \oc8051_golden_model_1.IP [7]);
  and (_13492_, _08575_, _07946_);
  or (_13493_, _13492_, _13491_);
  and (_13494_, _13493_, _06536_);
  nor (_13495_, _08040_, _13490_);
  or (_13496_, _13495_, _13491_);
  or (_13497_, _13496_, _07215_);
  not (_13498_, _08632_);
  and (_13499_, _13498_, \oc8051_golden_model_1.IP [7]);
  and (_13500_, _08649_, _08632_);
  or (_13501_, _13500_, _13499_);
  and (_13502_, _13501_, _06268_);
  and (_13503_, _08768_, _07946_);
  or (_13504_, _13503_, _13491_);
  or (_13505_, _13504_, _07151_);
  and (_13506_, _07946_, \oc8051_golden_model_1.ACC [7]);
  or (_13507_, _13506_, _13491_);
  and (_13508_, _13507_, _07141_);
  and (_13509_, _07142_, \oc8051_golden_model_1.IP [7]);
  or (_13510_, _13509_, _06341_);
  or (_13511_, _13510_, _13508_);
  and (_13512_, _13511_, _06273_);
  and (_13513_, _13512_, _13505_);
  and (_13514_, _08773_, _08632_);
  or (_13515_, _13514_, _13499_);
  and (_13516_, _13515_, _06272_);
  or (_13517_, _13516_, _06461_);
  or (_13518_, _13517_, _13513_);
  or (_13519_, _13496_, _07166_);
  and (_13520_, _13519_, _13518_);
  or (_13521_, _13520_, _06464_);
  or (_13522_, _13507_, _06465_);
  and (_13523_, _13522_, _06269_);
  and (_13524_, _13523_, _13521_);
  or (_13525_, _13524_, _13502_);
  and (_13526_, _13525_, _06262_);
  and (_13527_, _08790_, _08632_);
  or (_13528_, _13527_, _13499_);
  and (_13529_, _13528_, _06261_);
  or (_13530_, _13529_, _13526_);
  and (_13531_, _13530_, _06258_);
  and (_13532_, _08808_, _08632_);
  or (_13533_, _13532_, _13499_);
  and (_13534_, _13533_, _06257_);
  or (_13535_, _13534_, _10080_);
  or (_13536_, _13535_, _13531_);
  and (_13537_, _13536_, _13497_);
  or (_13538_, _13537_, _07460_);
  and (_13539_, _08755_, _07946_);
  or (_13540_, _13491_, _07208_);
  or (_13541_, _13540_, _13539_);
  and (_13542_, _13541_, _05982_);
  and (_13543_, _13542_, _13538_);
  and (_13544_, _09021_, _07946_);
  or (_13545_, _13544_, _13491_);
  and (_13546_, _13545_, _10094_);
  or (_13547_, _13546_, _06218_);
  or (_13548_, _13547_, _13543_);
  and (_13549_, _08825_, _07946_);
  or (_13550_, _13549_, _13491_);
  or (_13551_, _13550_, _06219_);
  and (_13552_, _13551_, _13548_);
  or (_13553_, _13552_, _06369_);
  and (_13554_, _09044_, _07946_);
  or (_13555_, _13554_, _13491_);
  or (_13556_, _13555_, _07237_);
  and (_13557_, _13556_, _07240_);
  and (_13558_, _13557_, _13553_);
  or (_13559_, _13558_, _13494_);
  and (_13560_, _13559_, _07242_);
  or (_13561_, _13491_, _08043_);
  and (_13562_, _13550_, _06375_);
  and (_13563_, _13562_, _13561_);
  or (_13564_, _13563_, _13560_);
  and (_13565_, _13564_, _07234_);
  and (_13566_, _13507_, _06545_);
  and (_13567_, _13566_, _13561_);
  or (_13568_, _13567_, _06366_);
  or (_13569_, _13568_, _13565_);
  nor (_13570_, _09043_, _13490_);
  or (_13571_, _13491_, _09056_);
  or (_13572_, _13571_, _13570_);
  and (_13573_, _13572_, _09061_);
  and (_13574_, _13573_, _13569_);
  nor (_13575_, _08573_, _13490_);
  or (_13576_, _13575_, _13491_);
  and (_13577_, _13576_, _06528_);
  or (_13578_, _13577_, _06568_);
  or (_13579_, _13578_, _13574_);
  or (_13580_, _13504_, _06926_);
  and (_13581_, _13580_, _05928_);
  and (_13582_, _13581_, _13579_);
  and (_13583_, _13501_, _05927_);
  or (_13584_, _13583_, _06278_);
  or (_13585_, _13584_, _13582_);
  and (_13586_, _08550_, _07946_);
  or (_13587_, _13491_, _06279_);
  or (_13588_, _13587_, _13586_);
  and (_13589_, _13588_, _01347_);
  and (_13590_, _13589_, _13585_);
  or (_13591_, _13590_, _13489_);
  and (_40592_, _13591_, _42618_);
  and (_13592_, _01351_, \oc8051_golden_model_1.IE [7]);
  not (_13593_, _07900_);
  and (_13594_, _13593_, \oc8051_golden_model_1.IE [7]);
  and (_13595_, _08575_, _07900_);
  or (_13596_, _13595_, _13594_);
  and (_13597_, _13596_, _06536_);
  nor (_13598_, _08040_, _13593_);
  or (_13599_, _13598_, _13594_);
  or (_13600_, _13599_, _07215_);
  not (_13601_, _08626_);
  and (_13602_, _13601_, \oc8051_golden_model_1.IE [7]);
  and (_13603_, _08649_, _08626_);
  or (_13604_, _13603_, _13602_);
  and (_13605_, _13604_, _06268_);
  and (_13606_, _08768_, _07900_);
  or (_13607_, _13606_, _13594_);
  or (_13608_, _13607_, _07151_);
  and (_13609_, _07900_, \oc8051_golden_model_1.ACC [7]);
  or (_13610_, _13609_, _13594_);
  and (_13611_, _13610_, _07141_);
  and (_13612_, _07142_, \oc8051_golden_model_1.IE [7]);
  or (_13614_, _13612_, _06341_);
  or (_13615_, _13614_, _13611_);
  and (_13616_, _13615_, _06273_);
  and (_13617_, _13616_, _13608_);
  and (_13618_, _08773_, _08626_);
  or (_13619_, _13618_, _13602_);
  and (_13620_, _13619_, _06272_);
  or (_13621_, _13620_, _06461_);
  or (_13622_, _13621_, _13617_);
  or (_13623_, _13599_, _07166_);
  and (_13625_, _13623_, _13622_);
  or (_13626_, _13625_, _06464_);
  or (_13627_, _13610_, _06465_);
  and (_13628_, _13627_, _06269_);
  and (_13629_, _13628_, _13626_);
  or (_13630_, _13629_, _13605_);
  and (_13631_, _13630_, _06262_);
  and (_13632_, _08790_, _08626_);
  or (_13633_, _13632_, _13602_);
  and (_13634_, _13633_, _06261_);
  or (_13636_, _13634_, _13631_);
  and (_13637_, _13636_, _06258_);
  and (_13638_, _08808_, _08626_);
  or (_13639_, _13638_, _13602_);
  and (_13640_, _13639_, _06257_);
  or (_13641_, _13640_, _10080_);
  or (_13642_, _13641_, _13637_);
  and (_13643_, _13642_, _13600_);
  or (_13644_, _13643_, _07460_);
  and (_13645_, _08755_, _07900_);
  or (_13647_, _13594_, _07208_);
  or (_13648_, _13647_, _13645_);
  and (_13649_, _13648_, _05982_);
  and (_13650_, _13649_, _13644_);
  and (_13651_, _09021_, _07900_);
  or (_13652_, _13651_, _13594_);
  and (_13653_, _13652_, _10094_);
  or (_13654_, _13653_, _06218_);
  or (_13655_, _13654_, _13650_);
  and (_13656_, _08825_, _07900_);
  or (_13658_, _13656_, _13594_);
  or (_13659_, _13658_, _06219_);
  and (_13660_, _13659_, _13655_);
  or (_13661_, _13660_, _06369_);
  and (_13662_, _09044_, _07900_);
  or (_13663_, _13662_, _13594_);
  or (_13664_, _13663_, _07237_);
  and (_13665_, _13664_, _07240_);
  and (_13666_, _13665_, _13661_);
  or (_13667_, _13666_, _13597_);
  and (_13669_, _13667_, _07242_);
  or (_13670_, _13594_, _08043_);
  and (_13671_, _13658_, _06375_);
  and (_13672_, _13671_, _13670_);
  or (_13673_, _13672_, _13669_);
  and (_13674_, _13673_, _07234_);
  and (_13675_, _13610_, _06545_);
  and (_13676_, _13675_, _13670_);
  or (_13677_, _13676_, _06366_);
  or (_13678_, _13677_, _13674_);
  nor (_13680_, _09043_, _13593_);
  or (_13681_, _13594_, _09056_);
  or (_13682_, _13681_, _13680_);
  and (_13683_, _13682_, _09061_);
  and (_13684_, _13683_, _13678_);
  nor (_13685_, _08573_, _13593_);
  or (_13686_, _13685_, _13594_);
  and (_13687_, _13686_, _06528_);
  or (_13688_, _13687_, _06568_);
  or (_13689_, _13688_, _13684_);
  or (_13691_, _13607_, _06926_);
  and (_13692_, _13691_, _05928_);
  and (_13693_, _13692_, _13689_);
  and (_13694_, _13604_, _05927_);
  or (_13695_, _13694_, _06278_);
  or (_13696_, _13695_, _13693_);
  and (_13697_, _08550_, _07900_);
  or (_13698_, _13594_, _06279_);
  or (_13699_, _13698_, _13697_);
  and (_13700_, _13699_, _01347_);
  and (_13702_, _13700_, _13696_);
  or (_13703_, _13702_, _13592_);
  and (_40593_, _13703_, _42618_);
  and (_13704_, _01351_, \oc8051_golden_model_1.SCON [7]);
  not (_13705_, _07973_);
  and (_13706_, _13705_, \oc8051_golden_model_1.SCON [7]);
  and (_13707_, _08575_, _07973_);
  or (_13708_, _13707_, _13706_);
  and (_13709_, _13708_, _06536_);
  nor (_13710_, _08040_, _13705_);
  or (_13712_, _13710_, _13706_);
  or (_13713_, _13712_, _07215_);
  not (_13714_, _08622_);
  and (_13715_, _13714_, \oc8051_golden_model_1.SCON [7]);
  and (_13716_, _08649_, _08622_);
  or (_13717_, _13716_, _13715_);
  and (_13718_, _13717_, _06268_);
  and (_13719_, _08768_, _07973_);
  or (_13720_, _13719_, _13706_);
  or (_13721_, _13720_, _07151_);
  and (_13723_, _07973_, \oc8051_golden_model_1.ACC [7]);
  or (_13724_, _13723_, _13706_);
  and (_13725_, _13724_, _07141_);
  and (_13726_, _07142_, \oc8051_golden_model_1.SCON [7]);
  or (_13727_, _13726_, _06341_);
  or (_13728_, _13727_, _13725_);
  and (_13729_, _13728_, _06273_);
  and (_13730_, _13729_, _13721_);
  and (_13731_, _08773_, _08622_);
  or (_13732_, _13731_, _13715_);
  and (_13734_, _13732_, _06272_);
  or (_13735_, _13734_, _06461_);
  or (_13736_, _13735_, _13730_);
  or (_13737_, _13712_, _07166_);
  and (_13738_, _13737_, _13736_);
  or (_13739_, _13738_, _06464_);
  or (_13740_, _13724_, _06465_);
  and (_13741_, _13740_, _06269_);
  and (_13742_, _13741_, _13739_);
  or (_13743_, _13742_, _13718_);
  and (_13745_, _13743_, _06262_);
  and (_13746_, _08790_, _08622_);
  or (_13747_, _13746_, _13715_);
  and (_13748_, _13747_, _06261_);
  or (_13749_, _13748_, _13745_);
  and (_13750_, _13749_, _06258_);
  and (_13751_, _08808_, _08622_);
  or (_13752_, _13751_, _13715_);
  and (_13753_, _13752_, _06257_);
  or (_13754_, _13753_, _10080_);
  or (_13756_, _13754_, _13750_);
  and (_13757_, _13756_, _13713_);
  or (_13758_, _13757_, _07460_);
  and (_13759_, _08755_, _07973_);
  or (_13760_, _13706_, _07208_);
  or (_13761_, _13760_, _13759_);
  and (_13762_, _13761_, _05982_);
  and (_13763_, _13762_, _13758_);
  and (_13764_, _09021_, _07973_);
  or (_13765_, _13764_, _13706_);
  and (_13766_, _13765_, _10094_);
  or (_13767_, _13766_, _06218_);
  or (_13768_, _13767_, _13763_);
  and (_13769_, _08825_, _07973_);
  or (_13770_, _13769_, _13706_);
  or (_13771_, _13770_, _06219_);
  and (_13772_, _13771_, _13768_);
  or (_13773_, _13772_, _06369_);
  and (_13774_, _09044_, _07973_);
  or (_13775_, _13774_, _13706_);
  or (_13776_, _13775_, _07237_);
  and (_13777_, _13776_, _07240_);
  and (_13778_, _13777_, _13773_);
  or (_13779_, _13778_, _13709_);
  and (_13780_, _13779_, _07242_);
  or (_13781_, _13706_, _08043_);
  and (_13782_, _13770_, _06375_);
  and (_13783_, _13782_, _13781_);
  or (_13784_, _13783_, _13780_);
  and (_13785_, _13784_, _07234_);
  and (_13786_, _13724_, _06545_);
  and (_13787_, _13786_, _13781_);
  or (_13788_, _13787_, _06366_);
  or (_13789_, _13788_, _13785_);
  nor (_13790_, _09043_, _13705_);
  or (_13791_, _13706_, _09056_);
  or (_13792_, _13791_, _13790_);
  and (_13793_, _13792_, _09061_);
  and (_13794_, _13793_, _13789_);
  nor (_13795_, _08573_, _13705_);
  or (_13796_, _13795_, _13706_);
  and (_13797_, _13796_, _06528_);
  or (_13798_, _13797_, _06568_);
  or (_13799_, _13798_, _13794_);
  or (_13800_, _13720_, _06926_);
  and (_13801_, _13800_, _05928_);
  and (_13802_, _13801_, _13799_);
  and (_13803_, _13717_, _05927_);
  or (_13804_, _13803_, _06278_);
  or (_13805_, _13804_, _13802_);
  and (_13806_, _08550_, _07973_);
  or (_13807_, _13706_, _06279_);
  or (_13808_, _13807_, _13806_);
  and (_13809_, _13808_, _01347_);
  and (_13810_, _13809_, _13805_);
  or (_13811_, _13810_, _13704_);
  and (_40594_, _13811_, _42618_);
  not (_13812_, \oc8051_golden_model_1.SP [7]);
  nor (_13813_, _01347_, _13812_);
  and (_13814_, _07602_, \oc8051_golden_model_1.SP [4]);
  and (_13815_, _13814_, \oc8051_golden_model_1.SP [5]);
  and (_13816_, _13815_, \oc8051_golden_model_1.SP [6]);
  or (_13817_, _13816_, \oc8051_golden_model_1.SP [7]);
  nand (_13818_, _13816_, \oc8051_golden_model_1.SP [7]);
  and (_13819_, _13818_, _13817_);
  or (_13820_, _13819_, _07271_);
  nor (_13821_, _07956_, _13812_);
  and (_13822_, _08575_, _08173_);
  or (_13823_, _13822_, _13821_);
  and (_13824_, _13823_, _06536_);
  or (_13825_, _13819_, _07494_);
  and (_13826_, _08768_, _08173_);
  or (_13827_, _13826_, _13821_);
  or (_13828_, _13827_, _07151_);
  and (_13829_, _07956_, \oc8051_golden_model_1.ACC [7]);
  or (_13830_, _13829_, _13821_);
  or (_13831_, _13830_, _07142_);
  or (_13832_, _07141_, \oc8051_golden_model_1.SP [7]);
  and (_13833_, _13832_, _07504_);
  and (_13834_, _13833_, _13831_);
  and (_13835_, _13819_, _06758_);
  or (_13836_, _13835_, _06341_);
  or (_13837_, _13836_, _13834_);
  and (_13838_, _13837_, _06010_);
  and (_13839_, _13838_, _13828_);
  and (_13840_, _13819_, _07611_);
  or (_13841_, _13840_, _06461_);
  or (_13842_, _13841_, _13839_);
  not (_13843_, \oc8051_golden_model_1.SP [6]);
  not (_13844_, \oc8051_golden_model_1.SP [5]);
  not (_13845_, \oc8051_golden_model_1.SP [4]);
  and (_13846_, _08672_, _13845_);
  and (_13847_, _13846_, _13844_);
  and (_13848_, _13847_, _13843_);
  and (_13849_, _13848_, _06800_);
  nor (_13850_, _13849_, _13812_);
  and (_13851_, _13849_, _13812_);
  nor (_13852_, _13851_, _13850_);
  nand (_13853_, _13852_, _06461_);
  and (_13854_, _13853_, _13842_);
  or (_13855_, _13854_, _06464_);
  or (_13856_, _13830_, _06465_);
  and (_13857_, _13856_, _07303_);
  and (_13858_, _13857_, _13855_);
  and (_13859_, _13815_, \oc8051_golden_model_1.SP [0]);
  and (_13860_, _13859_, \oc8051_golden_model_1.SP [6]);
  nor (_13861_, _13860_, _13812_);
  and (_13862_, _13860_, _13812_);
  or (_13863_, _13862_, _13861_);
  nand (_13864_, _13863_, _06267_);
  nand (_13865_, _13864_, _07494_);
  or (_13866_, _13865_, _13858_);
  nand (_13867_, _13866_, _13825_);
  and (_13868_, _06350_, _05944_);
  nor (_13869_, _13868_, _07214_);
  nand (_13870_, _13869_, _13867_);
  and (_13871_, _06337_, _05944_);
  not (_13872_, _08173_);
  nor (_13873_, _08040_, _13872_);
  or (_13874_, _13873_, _13821_);
  nor (_13875_, _13874_, _13869_);
  nor (_13876_, _13875_, _13871_);
  and (_13877_, _13876_, _13870_);
  and (_13878_, _13874_, _13871_);
  or (_13879_, _13878_, _07460_);
  or (_13880_, _13879_, _13877_);
  or (_13881_, _13821_, _07208_);
  and (_13882_, _08755_, _07956_);
  or (_13883_, _13882_, _13881_);
  and (_13884_, _13883_, _05982_);
  and (_13885_, _13884_, _13880_);
  and (_13886_, _09021_, _08173_);
  or (_13887_, _13886_, _13821_);
  and (_13888_, _13887_, _10094_);
  or (_13889_, _13888_, _06218_);
  or (_13890_, _13889_, _13885_);
  and (_13891_, _08825_, _07956_);
  or (_13892_, _13891_, _13821_);
  or (_13893_, _13892_, _06219_);
  and (_13894_, _13893_, _13890_);
  or (_13895_, _13894_, _06217_);
  or (_13896_, _13819_, _05952_);
  and (_13897_, _13896_, _13895_);
  or (_13898_, _13897_, _06369_);
  and (_13899_, _09044_, _07956_);
  or (_13900_, _13899_, _13821_);
  or (_13901_, _13900_, _07237_);
  and (_13902_, _13901_, _07240_);
  and (_13903_, _13902_, _13898_);
  or (_13904_, _13903_, _13824_);
  and (_13905_, _13904_, _07242_);
  or (_13906_, _13821_, _08043_);
  and (_13907_, _13892_, _06375_);
  and (_13908_, _13907_, _13906_);
  or (_13909_, _13908_, _13905_);
  and (_13910_, _13909_, _12772_);
  and (_13911_, _13830_, _06545_);
  and (_13912_, _13911_, _13906_);
  and (_13913_, _13819_, _07233_);
  or (_13914_, _13913_, _06366_);
  or (_13915_, _13914_, _13912_);
  or (_13916_, _13915_, _13910_);
  and (_13917_, _09063_, _07956_);
  or (_13918_, _13917_, _13821_);
  or (_13919_, _13918_, _09056_);
  and (_13920_, _13919_, _13916_);
  or (_13921_, _13920_, _06528_);
  nor (_13922_, _08573_, _13872_);
  or (_13923_, _13821_, _09061_);
  or (_13924_, _13923_, _13922_);
  and (_13925_, _13924_, _06716_);
  and (_13926_, _13925_, _13921_);
  or (_13927_, _13848_, \oc8051_golden_model_1.SP [7]);
  nand (_13928_, _13848_, \oc8051_golden_model_1.SP [7]);
  and (_13929_, _13928_, _13927_);
  and (_13930_, _13929_, _06551_);
  or (_13931_, _13930_, _07253_);
  or (_13932_, _13931_, _13926_);
  or (_13933_, _13819_, _05959_);
  and (_13934_, _13933_, _13932_);
  or (_13935_, _13934_, _06281_);
  or (_13936_, _13929_, _06282_);
  and (_13937_, _13936_, _06926_);
  and (_13938_, _13937_, _13935_);
  and (_13939_, _13827_, _06568_);
  or (_13940_, _13939_, _07695_);
  or (_13941_, _13940_, _13938_);
  and (_13942_, _13941_, _13820_);
  or (_13943_, _13942_, _06278_);
  and (_13944_, _08550_, _08173_);
  or (_13945_, _13821_, _06279_);
  or (_13946_, _13945_, _13944_);
  and (_13947_, _13946_, _01347_);
  and (_13948_, _13947_, _13943_);
  or (_13949_, _13948_, _13813_);
  and (_40595_, _13949_, _42618_);
  and (_13950_, _01351_, \oc8051_golden_model_1.SBUF [7]);
  not (_13951_, _07886_);
  and (_13952_, _13951_, \oc8051_golden_model_1.SBUF [7]);
  nor (_13953_, _08573_, _13951_);
  or (_13954_, _13953_, _13952_);
  and (_13955_, _13954_, _06528_);
  and (_13956_, _08575_, _07886_);
  or (_13957_, _13956_, _13952_);
  and (_13958_, _13957_, _06536_);
  nor (_13959_, _08040_, _13951_);
  or (_13960_, _13959_, _13952_);
  or (_13961_, _13960_, _07215_);
  and (_13962_, _08768_, _07886_);
  or (_13963_, _13962_, _13952_);
  or (_13964_, _13963_, _07151_);
  and (_13965_, _07886_, \oc8051_golden_model_1.ACC [7]);
  or (_13966_, _13965_, _13952_);
  and (_13967_, _13966_, _07141_);
  and (_13968_, _07142_, \oc8051_golden_model_1.SBUF [7]);
  or (_13969_, _13968_, _06341_);
  or (_13970_, _13969_, _13967_);
  and (_13971_, _13970_, _07166_);
  and (_13972_, _13971_, _13964_);
  and (_13973_, _13960_, _06461_);
  or (_13974_, _13973_, _13972_);
  and (_13975_, _13974_, _06465_);
  and (_13976_, _13966_, _06464_);
  or (_13977_, _13976_, _10080_);
  or (_13978_, _13977_, _13975_);
  and (_13979_, _13978_, _13961_);
  or (_13980_, _13979_, _07460_);
  and (_13981_, _08755_, _07886_);
  or (_13982_, _13952_, _07208_);
  or (_13983_, _13982_, _13981_);
  and (_13984_, _13983_, _05982_);
  and (_13985_, _13984_, _13980_);
  and (_13986_, _09021_, _07886_);
  or (_13987_, _13986_, _13952_);
  and (_13988_, _13987_, _10094_);
  or (_13989_, _13988_, _06218_);
  or (_13990_, _13989_, _13985_);
  and (_13991_, _08825_, _07886_);
  or (_13992_, _13991_, _13952_);
  or (_13993_, _13992_, _06219_);
  and (_13994_, _13993_, _13990_);
  or (_13995_, _13994_, _06369_);
  and (_13996_, _09044_, _07886_);
  or (_13997_, _13996_, _13952_);
  or (_13998_, _13997_, _07237_);
  and (_13999_, _13998_, _07240_);
  and (_14000_, _13999_, _13995_);
  or (_14001_, _14000_, _13958_);
  and (_14002_, _14001_, _07242_);
  or (_14003_, _13952_, _08043_);
  and (_14004_, _13992_, _06375_);
  and (_14005_, _14004_, _14003_);
  or (_14006_, _14005_, _14002_);
  and (_14007_, _14006_, _07234_);
  and (_14008_, _13966_, _06545_);
  and (_14009_, _14008_, _14003_);
  or (_14010_, _14009_, _06366_);
  or (_14011_, _14010_, _14007_);
  nor (_14012_, _09043_, _13951_);
  or (_14013_, _13952_, _09056_);
  or (_14014_, _14013_, _14012_);
  and (_14015_, _14014_, _09061_);
  and (_14016_, _14015_, _14011_);
  or (_14017_, _14016_, _13955_);
  and (_14018_, _14017_, _06926_);
  and (_14019_, _13963_, _06568_);
  or (_14020_, _14019_, _06278_);
  or (_14021_, _14020_, _14018_);
  and (_14022_, _08550_, _07886_);
  or (_14023_, _13952_, _06279_);
  or (_14024_, _14023_, _14022_);
  and (_14025_, _14024_, _01347_);
  and (_14026_, _14025_, _14021_);
  or (_14027_, _14026_, _13950_);
  and (_40597_, _14027_, _42618_);
  nor (_14028_, _01347_, _10558_);
  nor (_14029_, _08630_, _10558_);
  and (_14030_, _08649_, _08630_);
  or (_14031_, _14030_, _14029_);
  or (_14032_, _14031_, _05928_);
  and (_14033_, _10664_, _08552_);
  and (_14034_, _10667_, \oc8051_golden_model_1.ACC [7]);
  or (_14035_, _14034_, _11064_);
  or (_14036_, _14035_, _14033_);
  or (_14037_, _14036_, _11037_);
  nor (_14038_, _07935_, _10558_);
  and (_14039_, _08575_, _07935_);
  or (_14040_, _14039_, _14038_);
  and (_14041_, _14040_, _06536_);
  and (_14042_, _09021_, _07935_);
  or (_14043_, _14042_, _14038_);
  and (_14044_, _14043_, _10094_);
  not (_14045_, _07935_);
  nor (_14046_, _08040_, _14045_);
  or (_14047_, _14046_, _14038_);
  or (_14048_, _14047_, _07215_);
  and (_14049_, _10605_, _10601_);
  nor (_14050_, _14049_, _10599_);
  nand (_14051_, _10648_, _10601_);
  or (_14052_, _14051_, _10646_);
  and (_14053_, _14052_, _14050_);
  and (_14054_, _10595_, _08755_);
  or (_14055_, _14054_, _10588_);
  or (_14056_, _14055_, _14053_);
  not (_14057_, _06504_);
  not (_14058_, _06505_);
  nor (_14059_, _13004_, _14058_);
  and (_14060_, _08773_, _08630_);
  or (_14061_, _14060_, _14029_);
  or (_14062_, _14029_, _08789_);
  and (_14063_, _14062_, _06261_);
  and (_14064_, _14063_, _14061_);
  and (_14065_, _12366_, _12362_);
  or (_14066_, _12363_, _14065_);
  and (_14067_, _14066_, _12361_);
  and (_14068_, _12358_, _12356_);
  or (_14069_, _14068_, _12355_);
  or (_14070_, _14069_, _14067_);
  and (_14071_, _14070_, _12354_);
  or (_14072_, _12350_, _12347_);
  and (_14073_, _12345_, _14072_);
  and (_14074_, _14073_, _12346_);
  and (_14075_, _12343_, _08041_);
  or (_14076_, _14075_, _12340_);
  or (_14077_, _14076_, _14074_);
  or (_14078_, _14077_, _14071_);
  nor (_14079_, _12378_, _12371_);
  and (_14080_, _14079_, _14078_);
  and (_14081_, _08768_, _07935_);
  or (_14082_, _14081_, _14038_);
  or (_14083_, _14082_, _07151_);
  and (_14084_, _07935_, \oc8051_golden_model_1.ACC [7]);
  or (_14085_, _14084_, _14038_);
  and (_14086_, _14085_, _07141_);
  nor (_14087_, _07141_, _10558_);
  or (_14088_, _14087_, _06341_);
  or (_14089_, _14088_, _14086_);
  and (_14090_, _14089_, _10776_);
  and (_14091_, _14090_, _14083_);
  nor (_14092_, _10795_, _10776_);
  or (_14093_, _12540_, _06467_);
  or (_14094_, _14093_, _14092_);
  or (_14095_, _14094_, _14091_);
  or (_14096_, _14061_, _06273_);
  or (_14097_, _14047_, _07166_);
  and (_14098_, _14097_, _14096_);
  and (_14099_, _14098_, _14095_);
  or (_14100_, _14099_, _06464_);
  or (_14101_, _14085_, _06465_);
  nor (_14102_, _12559_, _06268_);
  and (_14103_, _14102_, _14101_);
  and (_14104_, _14103_, _14100_);
  and (_14105_, _14031_, _06268_);
  or (_14106_, _14105_, _14104_);
  and (_14107_, _14106_, _12378_);
  or (_14108_, _14107_, _14080_);
  and (_14109_, _14108_, _12177_);
  nand (_14110_, _12329_, _12326_);
  nand (_14111_, _14110_, _12325_);
  and (_14112_, _14111_, _12324_);
  nand (_14113_, _12321_, _12318_);
  and (_14114_, _12319_, _14113_);
  or (_14115_, _14114_, _14112_);
  and (_14116_, _14115_, _12317_);
  nor (_14117_, _12306_, _08802_);
  or (_14118_, _14117_, _12304_);
  nand (_14119_, _12314_, _12311_);
  and (_14120_, _12309_, _14119_);
  and (_14121_, _14120_, _12310_);
  or (_14122_, _14121_, _14118_);
  or (_14123_, _14122_, _14116_);
  and (_14124_, _12335_, _06347_);
  and (_14125_, _14124_, _14123_);
  or (_14126_, _14125_, _14109_);
  and (_14127_, _14126_, _06774_);
  nand (_14128_, _08246_, \oc8051_golden_model_1.ACC [5]);
  nor (_14129_, _08246_, \oc8051_golden_model_1.ACC [5]);
  nor (_14130_, _08543_, \oc8051_golden_model_1.ACC [4]);
  or (_14131_, _14130_, _14129_);
  and (_14132_, _14131_, _14128_);
  and (_14133_, _14132_, _12585_);
  nor (_14134_, _08042_, \oc8051_golden_model_1.ACC [7]);
  or (_14135_, _08144_, \oc8051_golden_model_1.ACC [6]);
  nor (_14136_, _14135_, _08575_);
  or (_14137_, _14136_, _14134_);
  or (_14138_, _14137_, _14133_);
  nand (_14139_, _08291_, \oc8051_golden_model_1.ACC [3]);
  nor (_14140_, _08291_, \oc8051_golden_model_1.ACC [3]);
  nor (_14141_, _08439_, \oc8051_golden_model_1.ACC [2]);
  or (_14142_, _14141_, _14140_);
  and (_14143_, _14142_, _14139_);
  nor (_14144_, _08340_, \oc8051_golden_model_1.ACC [1]);
  nor (_14145_, _08390_, _06097_);
  nor (_14146_, _14145_, _11262_);
  or (_14147_, _14146_, _14144_);
  and (_14148_, _14147_, _12578_);
  or (_14149_, _14148_, _14143_);
  and (_14150_, _14149_, _12586_);
  or (_14151_, _14150_, _14138_);
  nor (_14152_, _12587_, _06774_);
  and (_14153_, _14152_, _14151_);
  or (_14154_, _14153_, _14127_);
  and (_14155_, _14154_, _12176_);
  and (_14156_, _06251_, \oc8051_golden_model_1.ACC [0]);
  nor (_14157_, _14156_, _11303_);
  or (_14158_, _14157_, _11304_);
  and (_14159_, _14158_, _12595_);
  nand (_14160_, _06213_, \oc8051_golden_model_1.ACC [3]);
  nor (_14161_, _06213_, \oc8051_golden_model_1.ACC [3]);
  nor (_14162_, _06656_, \oc8051_golden_model_1.ACC [2]);
  or (_14163_, _14162_, _14161_);
  and (_14164_, _14163_, _14160_);
  or (_14165_, _14164_, _14159_);
  and (_14166_, _14165_, _12603_);
  nand (_14167_, _06611_, \oc8051_golden_model_1.ACC [5]);
  nor (_14168_, _06611_, \oc8051_golden_model_1.ACC [5]);
  nor (_14169_, _06968_, \oc8051_golden_model_1.ACC [4]);
  or (_14170_, _14169_, _14168_);
  and (_14171_, _14170_, _14167_);
  and (_14172_, _14171_, _12602_);
  and (_14173_, _06182_, _08572_);
  or (_14174_, _06317_, \oc8051_golden_model_1.ACC [6]);
  nor (_14175_, _14174_, _10961_);
  or (_14176_, _14175_, _14173_);
  or (_14177_, _14176_, _14172_);
  or (_14178_, _14177_, _14166_);
  nor (_14179_, _12604_, _12176_);
  and (_14180_, _14179_, _14178_);
  or (_14181_, _14180_, _12174_);
  or (_14182_, _14181_, _14155_);
  nand (_14183_, _12174_, \oc8051_golden_model_1.PSW [7]);
  and (_14184_, _14183_, _06262_);
  and (_14185_, _14184_, _14182_);
  nor (_14186_, _14185_, _14064_);
  nor (_14187_, _14186_, _06455_);
  and (_14188_, _06455_, \oc8051_golden_model_1.PSW [7]);
  and (_14189_, _14188_, _13004_);
  or (_14190_, _14189_, _14187_);
  nor (_14191_, _09531_, _06505_);
  and (_14192_, _14191_, _14190_);
  or (_14193_, _14192_, _14059_);
  and (_14194_, _14193_, _14057_);
  and (_14195_, _06886_, _05976_);
  and (_14196_, _06350_, _05976_);
  nor (_14197_, _14196_, _14195_);
  nand (_14198_, _14197_, _10731_);
  or (_14199_, _13004_, \oc8051_golden_model_1.PSW [7]);
  and (_14200_, _14199_, _06504_);
  or (_14201_, _14200_, _14198_);
  or (_14202_, _14201_, _14194_);
  and (_14203_, _06337_, _05976_);
  not (_14204_, _14203_);
  and (_14205_, _10675_, _10670_);
  nor (_14206_, _14205_, _10668_);
  nand (_14207_, _10721_, _10670_);
  or (_14208_, _14207_, _10719_);
  and (_14209_, _14208_, _14206_);
  or (_14210_, _14209_, _14033_);
  and (_14211_, _14210_, _14204_);
  or (_14212_, _14211_, _10735_);
  and (_14213_, _14212_, _14202_);
  and (_14214_, _14210_, _14203_);
  or (_14215_, _14214_, _10656_);
  or (_14216_, _14215_, _14213_);
  and (_14217_, _14216_, _14056_);
  or (_14218_, _14217_, _06512_);
  and (_14219_, _10850_, _10846_);
  nor (_14220_, _14219_, _10844_);
  nand (_14221_, _10892_, _10846_);
  or (_14222_, _14221_, _10890_);
  and (_14223_, _14222_, _14220_);
  and (_14224_, _10840_, _08043_);
  or (_14225_, _14224_, _06517_);
  or (_14226_, _14225_, _14223_);
  and (_14227_, _14226_, _10517_);
  and (_14228_, _14227_, _14218_);
  and (_14229_, _10519_, _07941_);
  and (_14230_, _10531_, _10527_);
  nor (_14231_, _14230_, _10525_);
  nand (_14232_, _10578_, _10527_);
  or (_14233_, _14232_, _10576_);
  and (_14234_, _14233_, _14231_);
  or (_14235_, _14234_, _14229_);
  and (_14236_, _14235_, _10516_);
  or (_14237_, _14236_, _10080_);
  or (_14238_, _14237_, _14228_);
  and (_14239_, _14238_, _14048_);
  or (_14240_, _14239_, _07460_);
  and (_14241_, _08755_, _07935_);
  or (_14242_, _14038_, _07208_);
  or (_14243_, _14242_, _14241_);
  and (_14244_, _14243_, _05982_);
  and (_14245_, _14244_, _14240_);
  or (_14246_, _14245_, _14044_);
  nor (_14247_, _10093_, _06323_);
  and (_14248_, _14247_, _14246_);
  nor (_14249_, _13004_, _10558_);
  and (_14250_, _14249_, _06323_);
  or (_14251_, _14250_, _06218_);
  or (_14252_, _14251_, _14248_);
  and (_14253_, _08825_, _07935_);
  or (_14254_, _14253_, _14038_);
  or (_14255_, _14254_, _06219_);
  and (_14256_, _14255_, _14252_);
  or (_14257_, _14256_, _06322_);
  nand (_14258_, _13004_, _10558_);
  or (_14259_, _14258_, _06881_);
  and (_14260_, _14259_, _14257_);
  or (_14261_, _14260_, _06369_);
  and (_14262_, _09044_, _07935_);
  or (_14263_, _14262_, _14038_);
  or (_14264_, _14263_, _07237_);
  and (_14265_, _14264_, _07240_);
  and (_14266_, _14265_, _14261_);
  or (_14267_, _14266_, _14041_);
  and (_14268_, _14267_, _07242_);
  or (_14269_, _14038_, _08043_);
  and (_14270_, _14254_, _06375_);
  and (_14271_, _14270_, _14269_);
  or (_14272_, _14271_, _14268_);
  and (_14273_, _14272_, _07234_);
  and (_14274_, _14085_, _06545_);
  and (_14275_, _14274_, _14269_);
  or (_14276_, _14275_, _06366_);
  or (_14277_, _14276_, _14273_);
  nor (_14278_, _09043_, _14045_);
  or (_14279_, _14038_, _09056_);
  or (_14280_, _14279_, _14278_);
  and (_14281_, _14280_, _09061_);
  and (_14282_, _14281_, _14277_);
  not (_14283_, _11037_);
  nor (_14284_, _08573_, _14045_);
  or (_14285_, _14284_, _14038_);
  and (_14286_, _14285_, _06528_);
  or (_14287_, _14286_, _14283_);
  or (_14288_, _14287_, _14282_);
  and (_14289_, _14288_, _14037_);
  or (_14290_, _14289_, _11041_);
  or (_14291_, _11069_, _14054_);
  nor (_14292_, _10598_, _08572_);
  or (_14293_, _14292_, _11091_);
  or (_14294_, _14293_, _14291_);
  and (_14295_, _14294_, _06541_);
  and (_14296_, _14295_, _14290_);
  not (_14297_, _12153_);
  nor (_14298_, _10843_, _08572_);
  or (_14299_, _14298_, _11119_);
  or (_14300_, _11097_, _14224_);
  or (_14301_, _14300_, _14299_);
  and (_14302_, _14301_, _14297_);
  or (_14303_, _14302_, _14296_);
  and (_14304_, _10524_, \oc8051_golden_model_1.ACC [7]);
  or (_14305_, _14304_, _11147_);
  or (_14306_, _11127_, _14229_);
  or (_14307_, _14306_, _14305_);
  and (_14308_, _14307_, _11126_);
  and (_14309_, _14308_, _14303_);
  nand (_14310_, _11125_, \oc8051_golden_model_1.ACC [7]);
  nand (_14311_, _14310_, _11157_);
  or (_14312_, _14311_, _14309_);
  and (_14313_, _11192_, _10505_);
  not (_14314_, _10494_);
  or (_14315_, _11160_, _10504_);
  and (_14316_, _14315_, _14314_);
  or (_14317_, _14316_, _11157_);
  or (_14318_, _14317_, _14313_);
  and (_14319_, _14318_, _14312_);
  or (_14320_, _14319_, _11201_);
  and (_14321_, _11235_, _10500_);
  nor (_14322_, _11204_, _10499_);
  nor (_14323_, _14322_, _10498_);
  or (_14324_, _14323_, _11203_);
  or (_14325_, _14324_, _14321_);
  and (_14326_, _14325_, _06285_);
  and (_14327_, _14326_, _14320_);
  not (_14328_, _08573_);
  not (_14329_, _08574_);
  nand (_14330_, _11277_, _14329_);
  and (_14331_, _14330_, _06283_);
  and (_14332_, _14331_, _14328_);
  or (_14333_, _14332_, _11243_);
  or (_14334_, _14333_, _14327_);
  nor (_14335_, _11319_, _10959_);
  or (_14336_, _14335_, _11321_);
  or (_14337_, _14336_, _10960_);
  and (_14338_, _14337_, _14334_);
  or (_14339_, _14338_, _06568_);
  nor (_14340_, _14082_, _06926_);
  nor (_14341_, _14340_, _11335_);
  and (_14342_, _14341_, _14339_);
  and (_14343_, _11335_, \oc8051_golden_model_1.ACC [0]);
  or (_14344_, _14343_, _05927_);
  or (_14345_, _14344_, _14342_);
  and (_14346_, _14345_, _14032_);
  or (_14347_, _14346_, _06278_);
  and (_14348_, _08550_, _07935_);
  or (_14349_, _14038_, _06279_);
  or (_14350_, _14349_, _14348_);
  and (_14351_, _14350_, _01347_);
  and (_14352_, _14351_, _14347_);
  or (_14353_, _14352_, _14028_);
  and (_40598_, _14353_, _42618_);
  and (_14354_, _07535_, _07289_);
  nor (_14355_, _14354_, _07537_);
  nor (_14356_, _07711_, _07536_);
  nor (_14357_, _14356_, _07859_);
  and (_14358_, _14357_, _07535_);
  and (_14359_, _14358_, _14355_);
  not (_14360_, _14359_);
  nand (_14361_, _05940_, _05630_);
  nand (_14362_, _12580_, _09062_);
  or (_14363_, _08390_, _08954_);
  and (_14364_, _08390_, _08954_);
  not (_14365_, _14364_);
  and (_14366_, _14365_, _14363_);
  and (_14367_, _14366_, _07238_);
  nor (_14368_, _05978_, _05630_);
  or (_14369_, _08390_, _06501_);
  nor (_14370_, _12925_, _12901_);
  or (_14371_, _14370_, _08610_);
  nor (_14372_, _08390_, _08652_);
  nand (_14373_, _12387_, _07133_);
  nand (_14374_, _06758_, _05630_);
  or (_14375_, _06758_, \oc8051_golden_model_1.ACC [0]);
  nand (_14376_, _14375_, _14374_);
  and (_14377_, _14376_, _08654_);
  nor (_14378_, _14377_, _07152_);
  and (_14379_, _14378_, _14373_);
  or (_14380_, _14379_, _14372_);
  and (_14381_, _14380_, _08651_);
  nand (_14382_, _12925_, _12902_);
  and (_14383_, _14382_, _06275_);
  or (_14384_, _14383_, _07611_);
  or (_14385_, _14384_, _14381_);
  nor (_14386_, _06010_, \oc8051_golden_model_1.PC [0]);
  nor (_14387_, _14386_, _07167_);
  and (_14388_, _14387_, _14385_);
  and (_14389_, _07167_, _07133_);
  or (_14390_, _14389_, _07179_);
  or (_14391_, _14390_, _14388_);
  and (_14392_, _14391_, _14371_);
  or (_14393_, _14392_, _06267_);
  or (_14394_, _08390_, _07303_);
  and (_14395_, _14394_, _06265_);
  and (_14396_, _14395_, _14393_);
  nand (_14397_, _14382_, _06264_);
  nor (_14398_, _14397_, _12926_);
  or (_14399_, _14398_, _14396_);
  and (_14400_, _14399_, _06007_);
  or (_14401_, _06007_, _05630_);
  nand (_14402_, _06501_, _14401_);
  or (_14403_, _14402_, _14400_);
  and (_14404_, _14403_, _14369_);
  or (_14405_, _14404_, _07197_);
  and (_14406_, _09392_, _06286_);
  nand (_14407_, _08387_, _07197_);
  or (_14408_, _14407_, _14406_);
  and (_14409_, _14408_, _14405_);
  or (_14410_, _14409_, _07196_);
  and (_14411_, _07889_, \oc8051_golden_model_1.PSW [7]);
  and (_14412_, _14411_, _06656_);
  or (_14413_, _14412_, _14370_);
  or (_14414_, _14413_, _08801_);
  and (_14415_, _14414_, _05978_);
  and (_14416_, _14415_, _14410_);
  or (_14417_, _14416_, _14368_);
  and (_14418_, _14417_, _08817_);
  and (_14419_, _08812_, _07133_);
  or (_14420_, _14419_, _08816_);
  or (_14421_, _14420_, _14418_);
  or (_14422_, _09392_, _08821_);
  and (_14423_, _14422_, _07471_);
  and (_14424_, _14423_, _14421_);
  and (_14425_, _08608_, _07133_);
  and (_14426_, _08957_, \oc8051_golden_model_1.TMOD [0]);
  and (_14427_, _08968_, \oc8051_golden_model_1.B [0]);
  or (_14428_, _14427_, _14426_);
  and (_14429_, _08944_, \oc8051_golden_model_1.P0 [0]);
  and (_14430_, _08950_, \oc8051_golden_model_1.ACC [0]);
  or (_14431_, _14430_, _14429_);
  or (_14432_, _14431_, _14428_);
  and (_14433_, _08934_, \oc8051_golden_model_1.TCON [0]);
  and (_14434_, _08965_, \oc8051_golden_model_1.SCON [0]);
  or (_14435_, _14434_, _14433_);
  and (_14436_, _08939_, \oc8051_golden_model_1.TL0 [0]);
  and (_14437_, _09007_, \oc8051_golden_model_1.PSW [0]);
  or (_14438_, _14437_, _14436_);
  or (_14439_, _14438_, _14435_);
  or (_14440_, _14439_, _14432_);
  and (_14441_, _08977_, \oc8051_golden_model_1.PCON [0]);
  and (_14442_, _08979_, \oc8051_golden_model_1.DPH [0]);
  or (_14443_, _14442_, _14441_);
  or (_14444_, _14443_, _14440_);
  and (_14445_, _09013_, \oc8051_golden_model_1.TH0 [0]);
  and (_14446_, _09015_, \oc8051_golden_model_1.TH1 [0]);
  and (_14447_, _08988_, \oc8051_golden_model_1.SP [0]);
  or (_14448_, _14447_, _14446_);
  or (_14449_, _14448_, _14445_);
  and (_14450_, _08999_, \oc8051_golden_model_1.P2 [0]);
  and (_14451_, _08993_, \oc8051_golden_model_1.IE [0]);
  or (_14452_, _14451_, _14450_);
  and (_14453_, _09001_, \oc8051_golden_model_1.P3 [0]);
  and (_14454_, _08996_, \oc8051_golden_model_1.IP [0]);
  or (_14455_, _14454_, _14453_);
  or (_14456_, _14455_, _14452_);
  and (_14457_, _08962_, \oc8051_golden_model_1.P1 [0]);
  and (_14458_, _09005_, \oc8051_golden_model_1.SBUF [0]);
  or (_14459_, _14458_, _14457_);
  or (_14460_, _14459_, _14456_);
  and (_14461_, _08984_, \oc8051_golden_model_1.DPL [0]);
  and (_14462_, _08986_, \oc8051_golden_model_1.TL1 [0]);
  or (_14463_, _14462_, _14461_);
  or (_14464_, _14463_, _14460_);
  or (_14465_, _14464_, _14449_);
  or (_14466_, _14465_, _14444_);
  or (_14467_, _14466_, _14425_);
  and (_14468_, _14467_, _07470_);
  or (_14469_, _14468_, _09031_);
  or (_14470_, _14469_, _14424_);
  and (_14471_, _09031_, _06251_);
  nor (_14472_, _14471_, _06220_);
  and (_14473_, _14472_, _14470_);
  and (_14474_, _08954_, _06220_);
  or (_14475_, _14474_, _06217_);
  or (_14476_, _14475_, _14473_);
  nor (_14477_, _05952_, \oc8051_golden_model_1.PC [0]);
  nor (_14478_, _14477_, _07238_);
  and (_14479_, _14478_, _14476_);
  or (_14480_, _14479_, _14367_);
  and (_14481_, _14480_, _08577_);
  nor (_14482_, _12581_, _08577_);
  or (_14483_, _14482_, _14481_);
  and (_14484_, _14483_, _08571_);
  and (_14485_, _14364_, _07243_);
  or (_14486_, _14485_, _14484_);
  and (_14487_, _14486_, _07236_);
  and (_14488_, _11263_, _07235_);
  or (_14489_, _14488_, _07233_);
  or (_14490_, _14489_, _14487_);
  nor (_14491_, _05961_, \oc8051_golden_model_1.PC [0]);
  nor (_14492_, _14491_, _09057_);
  and (_14493_, _14492_, _14490_);
  and (_14494_, _14363_, _09057_);
  or (_14495_, _14494_, _09062_);
  or (_14496_, _14495_, _14493_);
  and (_14497_, _14496_, _14362_);
  or (_14498_, _14497_, _07253_);
  or (_14499_, _05959_, \oc8051_golden_model_1.PC [0]);
  and (_14500_, _14499_, _08569_);
  and (_14501_, _14500_, _14498_);
  or (_14502_, _08569_, _07133_);
  nand (_14503_, _14502_, _07264_);
  or (_14504_, _14503_, _14501_);
  nand (_14505_, _09392_, _07435_);
  and (_14506_, _14505_, _14504_);
  or (_14507_, _14506_, _07261_);
  not (_14508_, _06361_);
  nand (_14509_, _08390_, _07261_);
  and (_14510_, _14509_, _14508_);
  and (_14511_, _14510_, _14507_);
  and (_14512_, _06361_, _05630_);
  or (_14513_, _14512_, _05940_);
  or (_14514_, _14513_, _14511_);
  and (_14515_, _14514_, _14361_);
  or (_14516_, _14515_, _07270_);
  or (_14517_, _14370_, _07539_);
  and (_14518_, _14517_, _09427_);
  and (_14519_, _14518_, _14516_);
  nor (_14520_, _09427_, _07133_);
  or (_14521_, _14520_, _14519_);
  and (_14522_, _14521_, _07282_);
  nor (_14523_, _09392_, _07282_);
  or (_14524_, _14523_, _07286_);
  or (_14525_, _14524_, _14522_);
  nand (_14526_, _08390_, _07286_);
  and (_14527_, _14526_, _07535_);
  and (_14528_, _14527_, _14525_);
  or (_14529_, _14528_, _14360_);
  or (_14530_, _14359_, \oc8051_golden_model_1.IRAM[0] [0]);
  not (_14531_, _07872_);
  and (_14532_, _07872_, _07866_);
  nor (_14533_, _07873_, _14532_);
  nand (_14534_, _14533_, _07296_);
  or (_14535_, _14534_, _14531_);
  and (_14536_, _14535_, _14530_);
  and (_14537_, _14536_, _14529_);
  and (_14538_, _07872_, _07296_);
  and (_14539_, _14538_, _14533_);
  nand (_14540_, _12276_, _06361_);
  or (_14541_, _12431_, _06361_);
  and (_14542_, _14541_, _14540_);
  and (_14543_, _14542_, _07872_);
  and (_14544_, _14543_, _14539_);
  or (_40612_, _14544_, _14537_);
  nor (_14545_, _09452_, _09394_);
  or (_14546_, _14545_, _07282_);
  not (_14547_, _08565_);
  or (_14548_, _09433_, _08556_);
  and (_14549_, _14548_, _07061_);
  or (_14550_, _14549_, _14547_);
  nor (_14551_, _05959_, \oc8051_golden_model_1.PC [1]);
  or (_14552_, _05952_, _05597_);
  or (_14553_, _09347_, _06182_);
  nand (_14554_, _14553_, _08338_);
  and (_14555_, _14554_, _07197_);
  not (_14556_, _12872_);
  nand (_14557_, _12871_, _12849_);
  and (_14558_, _14557_, _06264_);
  and (_14559_, _14558_, _14556_);
  nor (_14560_, _12871_, _08172_);
  or (_14561_, _14560_, _08610_);
  nor (_14562_, _08761_, _08391_);
  nand (_14563_, _14562_, _07152_);
  and (_14564_, _14548_, _12387_);
  nor (_14565_, _06758_, _06042_);
  and (_14566_, _06758_, _05597_);
  or (_14567_, _14566_, _14565_);
  and (_14568_, _14567_, _08654_);
  or (_14569_, _14568_, _07152_);
  or (_14570_, _14569_, _14564_);
  and (_14571_, _14570_, _14563_);
  or (_14572_, _14571_, _06275_);
  or (_14573_, _14557_, _08651_);
  and (_14574_, _14573_, _14572_);
  or (_14575_, _14574_, _07611_);
  nor (_14576_, _06010_, _05597_);
  nor (_14577_, _14576_, _07167_);
  and (_14578_, _14577_, _14575_);
  and (_14579_, _09432_, _07167_);
  or (_14580_, _14579_, _07179_);
  or (_14581_, _14580_, _14578_);
  and (_14582_, _14581_, _14561_);
  or (_14583_, _14582_, _06267_);
  nand (_14584_, _08340_, _06267_);
  and (_14585_, _14584_, _06265_);
  and (_14586_, _14585_, _14583_);
  or (_14587_, _14586_, _14559_);
  and (_14588_, _14587_, _06007_);
  or (_14589_, _06007_, \oc8051_golden_model_1.PC [1]);
  nand (_14590_, _06501_, _14589_);
  or (_14591_, _14590_, _14588_);
  nand (_14592_, _08340_, _06502_);
  and (_14593_, _14592_, _07198_);
  and (_14594_, _14593_, _14591_);
  or (_14595_, _14594_, _14555_);
  and (_14596_, _14595_, _08801_);
  nand (_14597_, _08172_, _10558_);
  and (_14598_, _14597_, _07196_);
  and (_14599_, _14598_, _14557_);
  or (_14600_, _14599_, _06254_);
  or (_14601_, _14600_, _14596_);
  nor (_14602_, _05978_, _05597_);
  nor (_14603_, _14602_, _08812_);
  and (_14604_, _14603_, _14601_);
  nor (_14605_, _07357_, _08817_);
  or (_14606_, _14605_, _08816_);
  or (_14607_, _14606_, _14604_);
  or (_14608_, _09451_, _08821_);
  and (_14609_, _14608_, _07471_);
  and (_14610_, _14609_, _14607_);
  nor (_14611_, _08825_, _07357_);
  and (_14612_, _08977_, \oc8051_golden_model_1.PCON [1]);
  and (_14613_, _08979_, \oc8051_golden_model_1.DPH [1]);
  or (_14614_, _14613_, _14612_);
  and (_14615_, _08934_, \oc8051_golden_model_1.TCON [1]);
  and (_14616_, _08957_, \oc8051_golden_model_1.TMOD [1]);
  or (_14617_, _14616_, _14615_);
  and (_14618_, _08939_, \oc8051_golden_model_1.TL0 [1]);
  and (_14619_, _08962_, \oc8051_golden_model_1.P1 [1]);
  or (_14620_, _14619_, _14618_);
  or (_14621_, _14620_, _14617_);
  and (_14622_, _08944_, \oc8051_golden_model_1.P0 [1]);
  and (_14623_, _08950_, \oc8051_golden_model_1.ACC [1]);
  or (_14624_, _14623_, _14622_);
  and (_14625_, _08968_, \oc8051_golden_model_1.B [1]);
  and (_14626_, _09007_, \oc8051_golden_model_1.PSW [1]);
  or (_14627_, _14626_, _14625_);
  or (_14628_, _14627_, _14624_);
  or (_14629_, _14628_, _14621_);
  or (_14630_, _14629_, _14614_);
  and (_14631_, _08986_, \oc8051_golden_model_1.TL1 [1]);
  and (_14632_, _09015_, \oc8051_golden_model_1.TH1 [1]);
  and (_14633_, _08988_, \oc8051_golden_model_1.SP [1]);
  or (_14634_, _14633_, _14632_);
  or (_14635_, _14634_, _14631_);
  and (_14636_, _09001_, \oc8051_golden_model_1.P3 [1]);
  and (_14637_, _08996_, \oc8051_golden_model_1.IP [1]);
  or (_14638_, _14637_, _14636_);
  and (_14639_, _08999_, \oc8051_golden_model_1.P2 [1]);
  and (_14640_, _08993_, \oc8051_golden_model_1.IE [1]);
  or (_14641_, _14640_, _14639_);
  or (_14642_, _14641_, _14638_);
  and (_14643_, _08965_, \oc8051_golden_model_1.SCON [1]);
  and (_14644_, _09005_, \oc8051_golden_model_1.SBUF [1]);
  or (_14645_, _14644_, _14643_);
  or (_14646_, _14645_, _14642_);
  and (_14647_, _08984_, \oc8051_golden_model_1.DPL [1]);
  and (_14648_, _09013_, \oc8051_golden_model_1.TH0 [1]);
  or (_14649_, _14648_, _14647_);
  or (_14650_, _14649_, _14646_);
  or (_14651_, _14650_, _14635_);
  or (_14652_, _14651_, _14630_);
  or (_14653_, _14652_, _14611_);
  and (_14654_, _14653_, _07470_);
  or (_14655_, _14654_, _09031_);
  or (_14656_, _14655_, _14610_);
  and (_14657_, _09031_, _07004_);
  nor (_14658_, _14657_, _06220_);
  and (_14659_, _14658_, _14656_);
  and (_14660_, _08936_, _06220_);
  or (_14661_, _14660_, _06217_);
  or (_14662_, _14661_, _14659_);
  and (_14663_, _14662_, _14552_);
  or (_14664_, _14663_, _07238_);
  nand (_14665_, _08340_, _07038_);
  nor (_14666_, _08340_, _07038_);
  not (_14667_, _14666_);
  and (_14668_, _14667_, _14665_);
  or (_14669_, _14668_, _07239_);
  and (_14670_, _14669_, _08577_);
  and (_14671_, _14670_, _14664_);
  and (_14672_, _11262_, _07241_);
  or (_14673_, _14672_, _07243_);
  or (_14674_, _14673_, _14671_);
  or (_14675_, _14666_, _08571_);
  and (_14676_, _14675_, _07236_);
  and (_14677_, _14676_, _14674_);
  and (_14678_, _11260_, _07235_);
  or (_14679_, _14678_, _07233_);
  or (_14680_, _14679_, _14677_);
  nor (_14681_, _05961_, _05597_);
  nor (_14682_, _14681_, _09057_);
  and (_14683_, _14682_, _14680_);
  and (_14684_, _14665_, _09057_);
  or (_14685_, _14684_, _09062_);
  or (_14686_, _14685_, _14683_);
  nand (_14687_, _11261_, _09062_);
  and (_14688_, _14687_, _05959_);
  and (_14689_, _14688_, _14686_);
  nor (_14690_, _14689_, _14551_);
  nor (_14691_, _14690_, _06701_);
  and (_14692_, _14548_, _06701_);
  or (_14693_, _14692_, _06754_);
  or (_14694_, _14693_, _14691_);
  not (_14695_, _06754_);
  or (_14696_, _14548_, _14695_);
  and (_14697_, _14696_, _07062_);
  and (_14698_, _14697_, _14694_);
  or (_14699_, _14698_, _14550_);
  not (_14700_, _07292_);
  or (_14701_, _14548_, _14700_);
  and (_14702_, _14701_, _07264_);
  and (_14703_, _14702_, _14699_);
  nor (_14704_, _14545_, _07264_);
  or (_14705_, _14704_, _14703_);
  and (_14706_, _14705_, _09075_);
  nor (_14707_, _14562_, _09075_);
  or (_14708_, _14707_, _06361_);
  or (_14709_, _14708_, _14706_);
  not (_14710_, _05940_);
  nand (_14711_, _06361_, _06111_);
  and (_14712_, _14711_, _14710_);
  and (_14713_, _14712_, _14709_);
  and (_14714_, _05940_, _05597_);
  or (_14715_, _07270_, _14714_);
  or (_14716_, _14715_, _14713_);
  or (_14717_, _14560_, _07539_);
  and (_14718_, _14717_, _09427_);
  and (_14719_, _14718_, _14716_);
  nor (_14720_, _14548_, _09427_);
  or (_14721_, _14720_, _07281_);
  or (_14722_, _14721_, _14719_);
  and (_14723_, _14722_, _14546_);
  or (_14724_, _14723_, _07286_);
  or (_14725_, _14562_, _09445_);
  and (_14726_, _14725_, _07535_);
  and (_14727_, _14726_, _14724_);
  or (_14728_, _14727_, _14360_);
  or (_14729_, _14359_, \oc8051_golden_model_1.IRAM[0] [1]);
  and (_14730_, _14729_, _14535_);
  and (_14731_, _14730_, _14728_);
  nand (_14732_, _12217_, _06361_);
  or (_14733_, _12426_, _06361_);
  and (_14734_, _14733_, _14732_);
  and (_14735_, _14734_, _07872_);
  and (_14736_, _14735_, _14539_);
  or (_40613_, _14736_, _14731_);
  not (_14737_, _07279_);
  nor (_14738_, _09452_, _09450_);
  nor (_14739_, _14738_, _09453_);
  and (_14740_, _14739_, _07280_);
  not (_14741_, _07280_);
  nor (_14742_, _09433_, _09431_);
  nor (_14743_, _14742_, _09434_);
  and (_14744_, _14743_, _09424_);
  not (_14745_, _07262_);
  not (_14746_, _07263_);
  nor (_14747_, _06085_, _05959_);
  nand (_14748_, _08439_, _06697_);
  nor (_14749_, _08439_, _06697_);
  not (_14750_, _14749_);
  and (_14751_, _14750_, _14748_);
  and (_14752_, _14751_, _07238_);
  or (_14753_, _09302_, _06182_);
  nand (_14754_, _14753_, _08437_);
  and (_14755_, _14754_, _07197_);
  nor (_14756_, _12847_, _07959_);
  or (_14757_, _14756_, _08610_);
  and (_14758_, _08556_, _07776_);
  nor (_14759_, _08556_, _07776_);
  or (_14760_, _14759_, _14758_);
  or (_14761_, _14760_, _08654_);
  nor (_14762_, _06758_, _10213_);
  and (_14763_, _06758_, _06079_);
  nor (_14764_, _14763_, _14762_);
  nand (_14765_, _14764_, _08654_);
  and (_14766_, _14765_, _14761_);
  and (_14767_, _14766_, _08652_);
  and (_14768_, _08761_, _08439_);
  nor (_14769_, _08761_, _08439_);
  or (_14770_, _14769_, _14768_);
  and (_14771_, _14770_, _07152_);
  or (_14772_, _14771_, _14767_);
  and (_14773_, _14772_, _08651_);
  nand (_14774_, _12847_, _12825_);
  and (_14775_, _14774_, _06275_);
  or (_14776_, _14775_, _07611_);
  or (_14777_, _14776_, _14773_);
  nor (_14778_, _06079_, _06010_);
  nor (_14779_, _14778_, _07167_);
  and (_14780_, _14779_, _14777_);
  and (_14781_, _09431_, _07167_);
  or (_14782_, _14781_, _07179_);
  or (_14783_, _14782_, _14780_);
  and (_14784_, _14783_, _14757_);
  or (_14785_, _14784_, _06267_);
  nand (_14786_, _08439_, _06267_);
  and (_14787_, _14786_, _06265_);
  and (_14788_, _14787_, _14785_);
  not (_14789_, _12848_);
  and (_14790_, _14774_, _14789_);
  and (_14791_, _14790_, _06264_);
  or (_14792_, _14791_, _14788_);
  and (_14793_, _14792_, _06007_);
  or (_14794_, _06085_, _06007_);
  nand (_14795_, _06501_, _14794_);
  or (_14796_, _14795_, _14793_);
  nand (_14797_, _08439_, _06502_);
  and (_14798_, _14797_, _07198_);
  and (_14799_, _14798_, _14796_);
  or (_14800_, _14799_, _14755_);
  and (_14801_, _14800_, _08801_);
  and (_14802_, _07917_, \oc8051_golden_model_1.PSW [7]);
  and (_14803_, _14802_, _06656_);
  or (_14804_, _14803_, _14756_);
  and (_14805_, _14804_, _07196_);
  or (_14806_, _14805_, _06254_);
  or (_14807_, _14806_, _14801_);
  nor (_14808_, _06079_, _05978_);
  nor (_14809_, _14808_, _08812_);
  and (_14810_, _14809_, _14807_);
  nor (_14811_, _07776_, _08817_);
  or (_14812_, _14811_, _08816_);
  or (_14813_, _14812_, _14810_);
  or (_14814_, _09450_, _08821_);
  and (_14815_, _14814_, _07471_);
  and (_14816_, _14815_, _14813_);
  nor (_14817_, _08825_, _07776_);
  and (_14818_, _08962_, \oc8051_golden_model_1.P1 [2]);
  and (_14819_, _08965_, \oc8051_golden_model_1.SCON [2]);
  or (_14820_, _14819_, _14818_);
  and (_14821_, _08957_, \oc8051_golden_model_1.TMOD [2]);
  and (_14822_, _08939_, \oc8051_golden_model_1.TL0 [2]);
  or (_14823_, _14822_, _14821_);
  or (_14824_, _14823_, _14820_);
  and (_14825_, _08934_, \oc8051_golden_model_1.TCON [2]);
  and (_14826_, _09007_, \oc8051_golden_model_1.PSW [2]);
  or (_14827_, _14826_, _14825_);
  and (_14828_, _09005_, \oc8051_golden_model_1.SBUF [2]);
  and (_14829_, _08968_, \oc8051_golden_model_1.B [2]);
  or (_14830_, _14829_, _14828_);
  or (_14831_, _14830_, _14827_);
  or (_14832_, _14831_, _14824_);
  and (_14833_, _08977_, \oc8051_golden_model_1.PCON [2]);
  and (_14834_, _08979_, \oc8051_golden_model_1.DPH [2]);
  or (_14835_, _14834_, _14833_);
  or (_14836_, _14835_, _14832_);
  and (_14837_, _08986_, \oc8051_golden_model_1.TL1 [2]);
  and (_14838_, _09015_, \oc8051_golden_model_1.TH1 [2]);
  or (_14839_, _14838_, _14837_);
  and (_14840_, _08988_, \oc8051_golden_model_1.SP [2]);
  or (_14841_, _14840_, _14839_);
  and (_14842_, _08993_, \oc8051_golden_model_1.IE [2]);
  and (_14843_, _08996_, \oc8051_golden_model_1.IP [2]);
  or (_14844_, _14843_, _14842_);
  and (_14845_, _08999_, \oc8051_golden_model_1.P2 [2]);
  and (_14846_, _09001_, \oc8051_golden_model_1.P3 [2]);
  or (_14847_, _14846_, _14845_);
  or (_14848_, _14847_, _14844_);
  and (_14849_, _08944_, \oc8051_golden_model_1.P0 [2]);
  and (_14850_, _08950_, \oc8051_golden_model_1.ACC [2]);
  or (_14851_, _14850_, _14849_);
  or (_14852_, _14851_, _14848_);
  and (_14853_, _08984_, \oc8051_golden_model_1.DPL [2]);
  and (_14854_, _09013_, \oc8051_golden_model_1.TH0 [2]);
  or (_14855_, _14854_, _14853_);
  or (_14856_, _14855_, _14852_);
  or (_14857_, _14856_, _14841_);
  or (_14858_, _14857_, _14836_);
  or (_14859_, _14858_, _14817_);
  and (_14860_, _14859_, _07470_);
  or (_14861_, _14860_, _09031_);
  or (_14862_, _14861_, _14816_);
  and (_14863_, _09031_, _06656_);
  nor (_14864_, _14863_, _06220_);
  and (_14865_, _14864_, _14862_);
  and (_14866_, _08973_, _06220_);
  or (_14867_, _14866_, _06217_);
  or (_14868_, _14867_, _14865_);
  nor (_14869_, _06079_, _05952_);
  nor (_14870_, _14869_, _07238_);
  and (_14871_, _14870_, _14868_);
  or (_14872_, _14871_, _14752_);
  and (_14873_, _14872_, _08577_);
  and (_14874_, _11259_, _07241_);
  or (_14875_, _14874_, _14873_);
  and (_14876_, _14875_, _08571_);
  and (_14877_, _14749_, _07243_);
  or (_14878_, _14877_, _14876_);
  and (_14879_, _14878_, _07236_);
  and (_14880_, _11257_, _07235_);
  or (_14881_, _14880_, _07233_);
  or (_14882_, _14881_, _14879_);
  nor (_14883_, _06079_, _05961_);
  nor (_14884_, _14883_, _09057_);
  and (_14885_, _14884_, _14882_);
  and (_14886_, _14748_, _09057_);
  or (_14887_, _14886_, _09062_);
  or (_14888_, _14887_, _14885_);
  nand (_14889_, _11258_, _09062_);
  and (_14890_, _14889_, _05959_);
  and (_14891_, _14890_, _14888_);
  or (_14892_, _14891_, _14747_);
  and (_14893_, _14892_, _08569_);
  not (_14894_, _08569_);
  and (_14895_, _14760_, _14894_);
  or (_14896_, _14895_, _14893_);
  and (_14897_, _14896_, _14746_);
  nor (_14898_, _09394_, _09302_);
  or (_14899_, _14898_, _09395_);
  and (_14900_, _14899_, _07263_);
  or (_14901_, _14900_, _14897_);
  and (_14902_, _14901_, _14745_);
  and (_14903_, _14899_, _07262_);
  or (_14904_, _14903_, _14902_);
  and (_14905_, _14904_, _09075_);
  and (_14906_, _14770_, _07261_);
  or (_14907_, _14906_, _06361_);
  or (_14908_, _14907_, _14905_);
  nand (_14909_, _12248_, _06361_);
  and (_14910_, _14909_, _14710_);
  and (_14911_, _14910_, _14908_);
  and (_14912_, _06079_, _05940_);
  or (_14913_, _07270_, _14912_);
  or (_14914_, _14913_, _14911_);
  or (_14915_, _14756_, _07539_);
  and (_14916_, _14915_, _09427_);
  and (_14917_, _14916_, _14914_);
  or (_14918_, _14917_, _14744_);
  and (_14919_, _14918_, _14741_);
  or (_14920_, _14919_, _14740_);
  and (_14921_, _14920_, _14737_);
  and (_14922_, _14739_, _07279_);
  or (_14923_, _14922_, _07286_);
  or (_14924_, _14923_, _14921_);
  nor (_14925_, _08440_, _08391_);
  nor (_14926_, _14925_, _08441_);
  or (_14927_, _14926_, _09445_);
  and (_14928_, _14927_, _07535_);
  and (_14929_, _14928_, _14924_);
  or (_14930_, _14929_, _14360_);
  or (_14931_, _14359_, \oc8051_golden_model_1.IRAM[0] [2]);
  and (_14932_, _14931_, _14535_);
  and (_14933_, _14932_, _14930_);
  nand (_14934_, _12203_, _06361_);
  or (_14935_, _12421_, _06361_);
  and (_14936_, _14935_, _14934_);
  and (_14937_, _14936_, _07872_);
  and (_14938_, _14937_, _14539_);
  or (_40614_, _14938_, _14933_);
  nor (_14939_, _05959_, _06033_);
  nand (_14940_, _08291_, _06452_);
  nor (_14941_, _08291_, _06452_);
  not (_14942_, _14941_);
  and (_14943_, _14942_, _14940_);
  and (_14944_, _14943_, _07238_);
  or (_14945_, _09257_, _06182_);
  nand (_14946_, _14945_, _08289_);
  and (_14947_, _14946_, _07197_);
  nor (_14948_, _12975_, _08185_);
  or (_14949_, _14948_, _08610_);
  nand (_14950_, _12975_, _12953_);
  or (_14951_, _14950_, _08651_);
  nor (_14952_, _14768_, _08291_);
  or (_14953_, _14952_, _08763_);
  and (_14954_, _14953_, _07152_);
  nor (_14955_, _14758_, _07594_);
  nor (_14956_, _14955_, _08557_);
  nand (_14957_, _14956_, _12387_);
  and (_14958_, _06758_, _05932_);
  nor (_14959_, _06758_, _06055_);
  nor (_14960_, _14959_, _14958_);
  and (_14961_, _14960_, _08654_);
  nor (_14962_, _14961_, _07152_);
  and (_14963_, _14962_, _14957_);
  or (_14964_, _14963_, _06275_);
  or (_14965_, _14964_, _14954_);
  and (_14966_, _14965_, _14951_);
  or (_14967_, _14966_, _07611_);
  nor (_14968_, _06010_, _05932_);
  nor (_14969_, _14968_, _07167_);
  and (_14970_, _14969_, _14967_);
  and (_14971_, _07595_, _07167_);
  or (_14972_, _14971_, _07179_);
  or (_14973_, _14972_, _14970_);
  and (_14974_, _14973_, _14949_);
  or (_14975_, _14974_, _06267_);
  nand (_14976_, _08291_, _06267_);
  and (_14977_, _14976_, _06265_);
  and (_14978_, _14977_, _14975_);
  not (_14979_, _12976_);
  and (_14980_, _14950_, _14979_);
  and (_14981_, _14980_, _06264_);
  or (_14982_, _14981_, _14978_);
  and (_14983_, _14982_, _06007_);
  or (_14984_, _06007_, _06033_);
  nand (_14985_, _06501_, _14984_);
  or (_14986_, _14985_, _14983_);
  nand (_14987_, _08291_, _06502_);
  and (_14988_, _14987_, _07198_);
  and (_14989_, _14988_, _14986_);
  or (_14990_, _14989_, _14947_);
  and (_14991_, _14990_, _08801_);
  nand (_14992_, _08185_, _10558_);
  and (_14993_, _14992_, _07196_);
  and (_14994_, _14993_, _14950_);
  or (_14995_, _14994_, _06254_);
  or (_14996_, _14995_, _14991_);
  nor (_14997_, _05978_, _05932_);
  nor (_14998_, _14997_, _08812_);
  and (_14999_, _14998_, _14996_);
  nor (_15000_, _07594_, _08817_);
  or (_15001_, _15000_, _08816_);
  or (_15002_, _15001_, _14999_);
  or (_15003_, _09449_, _08821_);
  and (_15004_, _15003_, _07471_);
  and (_15005_, _15004_, _15002_);
  nor (_15006_, _08825_, _07594_);
  and (_15007_, _08944_, \oc8051_golden_model_1.P0 [3]);
  and (_15008_, _08962_, \oc8051_golden_model_1.P1 [3]);
  or (_15009_, _15008_, _15007_);
  and (_15010_, _08939_, \oc8051_golden_model_1.TL0 [3]);
  and (_15011_, _08950_, \oc8051_golden_model_1.ACC [3]);
  or (_15012_, _15011_, _15010_);
  or (_15013_, _15012_, _15009_);
  and (_15014_, _08934_, \oc8051_golden_model_1.TCON [3]);
  and (_15015_, _08957_, \oc8051_golden_model_1.TMOD [3]);
  or (_15016_, _15015_, _15014_);
  and (_15017_, _08965_, \oc8051_golden_model_1.SCON [3]);
  and (_15018_, _09005_, \oc8051_golden_model_1.SBUF [3]);
  or (_15019_, _15018_, _15017_);
  or (_15020_, _15019_, _15016_);
  or (_15021_, _15020_, _15013_);
  and (_15022_, _08977_, \oc8051_golden_model_1.PCON [3]);
  and (_15023_, _08979_, \oc8051_golden_model_1.DPH [3]);
  or (_15024_, _15023_, _15022_);
  or (_15025_, _15024_, _15021_);
  and (_15026_, _09015_, \oc8051_golden_model_1.TH1 [3]);
  and (_15027_, _08984_, \oc8051_golden_model_1.DPL [3]);
  and (_15028_, _08986_, \oc8051_golden_model_1.TL1 [3]);
  or (_15029_, _15028_, _15027_);
  or (_15030_, _15029_, _15026_);
  and (_15031_, _08999_, \oc8051_golden_model_1.P2 [3]);
  and (_15032_, _08996_, \oc8051_golden_model_1.IP [3]);
  or (_15033_, _15032_, _15031_);
  and (_15034_, _08993_, \oc8051_golden_model_1.IE [3]);
  and (_15035_, _09001_, \oc8051_golden_model_1.P3 [3]);
  or (_15036_, _15035_, _15034_);
  or (_15037_, _15036_, _15033_);
  and (_15038_, _08968_, \oc8051_golden_model_1.B [3]);
  and (_15039_, _09007_, \oc8051_golden_model_1.PSW [3]);
  or (_15040_, _15039_, _15038_);
  or (_15041_, _15040_, _15037_);
  and (_15042_, _09013_, \oc8051_golden_model_1.TH0 [3]);
  and (_15043_, _08988_, \oc8051_golden_model_1.SP [3]);
  or (_15044_, _15043_, _15042_);
  or (_15045_, _15044_, _15041_);
  or (_15046_, _15045_, _15030_);
  or (_15047_, _15046_, _15025_);
  or (_15048_, _15047_, _15006_);
  and (_15049_, _15048_, _07470_);
  or (_15050_, _15049_, _09031_);
  or (_15051_, _15050_, _15005_);
  and (_15052_, _09031_, _06213_);
  nor (_15053_, _15052_, _06220_);
  and (_15054_, _15053_, _15051_);
  and (_15055_, _08930_, _06220_);
  or (_15056_, _15055_, _06217_);
  or (_15057_, _15056_, _15054_);
  nor (_15058_, _05952_, _05932_);
  nor (_15059_, _15058_, _07238_);
  and (_15060_, _15059_, _15057_);
  or (_15061_, _15060_, _14944_);
  and (_15062_, _15061_, _08577_);
  and (_15063_, _12577_, _07241_);
  or (_15064_, _15063_, _15062_);
  and (_15065_, _15064_, _08571_);
  and (_15066_, _14941_, _07243_);
  or (_15067_, _15066_, _15065_);
  and (_15068_, _15067_, _07236_);
  and (_15069_, _11255_, _07235_);
  or (_15070_, _15069_, _07233_);
  or (_15071_, _15070_, _15068_);
  nor (_15072_, _05961_, _05932_);
  nor (_15073_, _15072_, _09057_);
  and (_15074_, _15073_, _15071_);
  and (_15075_, _14940_, _09057_);
  or (_15076_, _15075_, _09062_);
  or (_15077_, _15076_, _15074_);
  nand (_15078_, _11256_, _09062_);
  and (_15079_, _15078_, _05959_);
  and (_15080_, _15079_, _15077_);
  or (_15081_, _15080_, _14939_);
  and (_15082_, _15081_, _08568_);
  nor (_15083_, _14956_, _08568_);
  or (_15084_, _15083_, _07292_);
  or (_15085_, _15084_, _15082_);
  nand (_15086_, _14956_, _14547_);
  and (_15087_, _15086_, _14746_);
  and (_15088_, _15087_, _15085_);
  nor (_15089_, _09395_, _09257_);
  or (_15090_, _15089_, _09396_);
  or (_15091_, _15090_, _07262_);
  and (_15092_, _15091_, _07435_);
  or (_15093_, _15092_, _15088_);
  or (_15094_, _15090_, _14745_);
  and (_15095_, _15094_, _09075_);
  and (_15096_, _15095_, _15093_);
  and (_15097_, _14953_, _07261_);
  or (_15098_, _15097_, _06361_);
  or (_15099_, _15098_, _15096_);
  nand (_15100_, _12243_, _06361_);
  and (_15101_, _15100_, _14710_);
  and (_15102_, _15101_, _15099_);
  and (_15103_, _05940_, _05932_);
  or (_15104_, _07270_, _15103_);
  or (_15105_, _15104_, _15102_);
  and (_15106_, _07041_, _05938_);
  nor (_15107_, _15106_, _07510_);
  or (_15108_, _14948_, _07539_);
  and (_15109_, _15108_, _15107_);
  and (_15110_, _15109_, _15105_);
  not (_15111_, _15107_);
  nor (_15112_, _09434_, _07595_);
  nor (_15113_, _15112_, _09435_);
  and (_15114_, _15113_, _15111_);
  and (_15115_, _10732_, _05938_);
  or (_15116_, _15115_, _15114_);
  or (_15117_, _15116_, _15110_);
  not (_15118_, _15115_);
  or (_15119_, _15118_, _15113_);
  and (_15120_, _15119_, _07282_);
  and (_15121_, _15120_, _15117_);
  or (_15122_, _09453_, _09449_);
  nor (_15123_, _09454_, _07282_);
  and (_15124_, _15123_, _15122_);
  or (_15125_, _15124_, _07286_);
  or (_15126_, _15125_, _15121_);
  nor (_15127_, _08441_, _08292_);
  nor (_15128_, _15127_, _08442_);
  or (_15129_, _15128_, _09445_);
  and (_15130_, _15129_, _07535_);
  and (_15131_, _15130_, _15126_);
  or (_15132_, _15131_, _14360_);
  or (_15133_, _14359_, \oc8051_golden_model_1.IRAM[0] [3]);
  and (_15134_, _15133_, _14535_);
  and (_15135_, _15134_, _15132_);
  nand (_15136_, _12208_, _06361_);
  or (_15137_, _12417_, _06361_);
  and (_15138_, _15137_, _15136_);
  and (_15139_, _15138_, _07872_);
  and (_15140_, _15139_, _14539_);
  or (_40615_, _15140_, _15135_);
  nor (_15141_, _09396_, _09212_);
  or (_15142_, _15141_, _09397_);
  and (_15143_, _15142_, _07263_);
  or (_15144_, _12451_, _05952_);
  nor (_15145_, _12452_, _05978_);
  and (_15146_, _12451_, _06758_);
  nor (_15147_, _06758_, _10135_);
  or (_15148_, _15147_, _15146_);
  and (_15149_, _15148_, _08654_);
  and (_15150_, _08557_, _08541_);
  nor (_15151_, _08557_, _08541_);
  or (_15152_, _15151_, _15150_);
  and (_15153_, _15152_, _12387_);
  or (_15154_, _15153_, _15149_);
  and (_15155_, _15154_, _07155_);
  and (_15156_, _09448_, _07154_);
  or (_15157_, _15156_, _15155_);
  and (_15159_, _15157_, _08652_);
  and (_15160_, _08763_, _08543_);
  nor (_15161_, _08763_, _08543_);
  or (_15162_, _15161_, _15160_);
  and (_15163_, _15162_, _07152_);
  or (_15164_, _15163_, _15159_);
  and (_15165_, _15164_, _08651_);
  nand (_15166_, _12897_, _12895_);
  and (_15167_, _15166_, _06275_);
  or (_15168_, _15167_, _07611_);
  or (_15169_, _15168_, _15165_);
  nor (_15170_, _12451_, _06010_);
  nor (_15171_, _15170_, _07167_);
  and (_15172_, _15171_, _15169_);
  and (_15173_, _09430_, _07167_);
  or (_15174_, _15173_, _07179_);
  or (_15175_, _15174_, _15172_);
  nor (_15176_, _12896_, _12895_);
  or (_15177_, _15176_, _08610_);
  and (_15178_, _15177_, _15175_);
  or (_15179_, _15178_, _06267_);
  nand (_15180_, _08543_, _06267_);
  and (_15181_, _15180_, _06265_);
  and (_15182_, _15181_, _15179_);
  not (_15183_, _12898_);
  and (_15184_, _15166_, _15183_);
  and (_15185_, _15184_, _06264_);
  or (_15186_, _15185_, _15182_);
  and (_15187_, _15186_, _06007_);
  or (_15188_, _12452_, _06007_);
  nand (_15189_, _15188_, _06501_);
  or (_15190_, _15189_, _15187_);
  nand (_15191_, _08543_, _06502_);
  and (_15192_, _15191_, _15190_);
  or (_15193_, _15192_, _07197_);
  and (_15194_, _09448_, _06286_);
  nand (_15195_, _08488_, _07197_);
  or (_15196_, _15195_, _15194_);
  and (_15197_, _15196_, _15193_);
  or (_15198_, _15197_, _07196_);
  and (_15199_, _14411_, _06657_);
  or (_15200_, _15199_, _15176_);
  or (_15201_, _15200_, _08801_);
  and (_15202_, _15201_, _05978_);
  and (_15203_, _15202_, _15198_);
  or (_15204_, _15203_, _15145_);
  and (_15205_, _15204_, _08817_);
  nor (_15206_, _08541_, _08817_);
  or (_15207_, _15206_, _08816_);
  or (_15208_, _15207_, _15205_);
  or (_15209_, _09448_, _08821_);
  and (_15210_, _15209_, _07471_);
  and (_15211_, _15210_, _15208_);
  nor (_15212_, _08825_, _08541_);
  and (_15213_, _08962_, \oc8051_golden_model_1.P1 [4]);
  and (_15214_, _08965_, \oc8051_golden_model_1.SCON [4]);
  or (_15215_, _15214_, _15213_);
  and (_15216_, _08944_, \oc8051_golden_model_1.P0 [4]);
  and (_15217_, _08939_, \oc8051_golden_model_1.TL0 [4]);
  or (_15218_, _15217_, _15216_);
  or (_15219_, _15218_, _15215_);
  and (_15220_, _08934_, \oc8051_golden_model_1.TCON [4]);
  and (_15221_, _08957_, \oc8051_golden_model_1.TMOD [4]);
  or (_15222_, _15221_, _15220_);
  and (_15223_, _09005_, \oc8051_golden_model_1.SBUF [4]);
  and (_15224_, _09007_, \oc8051_golden_model_1.PSW [4]);
  or (_15225_, _15224_, _15223_);
  or (_15226_, _15225_, _15222_);
  or (_15227_, _15226_, _15219_);
  and (_15228_, _08977_, \oc8051_golden_model_1.PCON [4]);
  and (_15229_, _08979_, \oc8051_golden_model_1.DPH [4]);
  or (_15230_, _15229_, _15228_);
  or (_15231_, _15230_, _15227_);
  and (_15232_, _09015_, \oc8051_golden_model_1.TH1 [4]);
  and (_15233_, _08986_, \oc8051_golden_model_1.TL1 [4]);
  and (_15234_, _08988_, \oc8051_golden_model_1.SP [4]);
  or (_15235_, _15234_, _15233_);
  or (_15236_, _15235_, _15232_);
  and (_15237_, _08950_, \oc8051_golden_model_1.ACC [4]);
  and (_15238_, _08968_, \oc8051_golden_model_1.B [4]);
  or (_15239_, _15238_, _15237_);
  and (_15240_, _08993_, \oc8051_golden_model_1.IE [4]);
  and (_15241_, _08996_, \oc8051_golden_model_1.IP [4]);
  or (_15242_, _15241_, _15240_);
  and (_15243_, _08999_, \oc8051_golden_model_1.P2 [4]);
  and (_15244_, _09001_, \oc8051_golden_model_1.P3 [4]);
  or (_15245_, _15244_, _15243_);
  or (_15246_, _15245_, _15242_);
  or (_15247_, _15246_, _15239_);
  and (_15248_, _08984_, \oc8051_golden_model_1.DPL [4]);
  and (_15249_, _09013_, \oc8051_golden_model_1.TH0 [4]);
  or (_15250_, _15249_, _15248_);
  or (_15251_, _15250_, _15247_);
  or (_15252_, _15251_, _15236_);
  or (_15253_, _15252_, _15231_);
  or (_15254_, _15253_, _15212_);
  and (_15255_, _15254_, _07470_);
  or (_15256_, _15255_, _09031_);
  or (_15257_, _15256_, _15211_);
  and (_15258_, _09031_, _06968_);
  nor (_15259_, _15258_, _06220_);
  and (_15260_, _15259_, _15257_);
  and (_15261_, _08959_, _06220_);
  or (_15262_, _15261_, _06217_);
  or (_15263_, _15262_, _15260_);
  and (_15264_, _15263_, _15144_);
  or (_15265_, _15264_, _07238_);
  nand (_15266_, _08892_, _08543_);
  nor (_15267_, _08892_, _08543_);
  not (_15268_, _15267_);
  and (_15269_, _15268_, _15266_);
  or (_15270_, _15269_, _07239_);
  and (_15271_, _15270_, _08577_);
  and (_15272_, _15271_, _15265_);
  and (_15273_, _11254_, _07241_);
  or (_15274_, _15273_, _07243_);
  or (_15275_, _15274_, _15272_);
  or (_15276_, _15267_, _08571_);
  and (_15277_, _15276_, _07236_);
  and (_15278_, _15277_, _15275_);
  and (_15279_, _11251_, _07235_);
  or (_15280_, _15279_, _07233_);
  or (_15281_, _15280_, _15278_);
  nor (_15282_, _12451_, _05961_);
  nor (_15283_, _15282_, _09057_);
  and (_15284_, _15283_, _15281_);
  and (_15285_, _15266_, _09057_);
  or (_15286_, _15285_, _09062_);
  or (_15287_, _15286_, _15284_);
  nand (_15288_, _11253_, _09062_);
  and (_15289_, _15288_, _05959_);
  and (_15290_, _15289_, _15287_);
  nor (_15291_, _12452_, _05959_);
  nor (_15292_, _15291_, _07292_);
  nand (_15293_, _15292_, _08568_);
  or (_15294_, _15293_, _15290_);
  or (_15295_, _15152_, _08569_);
  and (_15296_, _15295_, _14746_);
  and (_15297_, _15296_, _15294_);
  or (_15298_, _15297_, _15143_);
  and (_15299_, _15298_, _14745_);
  and (_15300_, _15142_, _07262_);
  or (_15301_, _15300_, _15299_);
  and (_15302_, _15301_, _09075_);
  and (_15303_, _15162_, _07261_);
  or (_15304_, _15303_, _06361_);
  or (_15305_, _15304_, _15302_);
  nand (_15306_, _12239_, _06361_);
  and (_15307_, _15306_, _14710_);
  and (_15308_, _15307_, _15305_);
  and (_15309_, _12451_, _05940_);
  or (_15310_, _15309_, _07270_);
  or (_15311_, _15310_, _15308_);
  or (_15312_, _15176_, _07539_);
  and (_15313_, _15312_, _09427_);
  and (_15314_, _15313_, _15311_);
  or (_15315_, _09435_, _09430_);
  nor (_15316_, _09436_, _09427_);
  and (_15317_, _15316_, _15315_);
  or (_15318_, _15317_, _07280_);
  or (_15319_, _15318_, _15314_);
  nor (_15320_, _09454_, _09448_);
  nor (_15321_, _15320_, _09455_);
  or (_15322_, _15321_, _14741_);
  and (_15323_, _15322_, _14737_);
  and (_15324_, _15323_, _15319_);
  and (_15325_, _15321_, _07279_);
  or (_15326_, _15325_, _07286_);
  or (_15327_, _15326_, _15324_);
  nor (_15328_, _08544_, _08442_);
  nor (_15329_, _15328_, _08545_);
  or (_15330_, _15329_, _09445_);
  and (_15331_, _15330_, _07535_);
  and (_15332_, _15331_, _15327_);
  or (_15333_, _15332_, _14360_);
  or (_15334_, _14359_, \oc8051_golden_model_1.IRAM[0] [4]);
  and (_15335_, _15334_, _14535_);
  and (_15336_, _15335_, _15333_);
  nand (_15337_, _12199_, _06361_);
  or (_15338_, _12414_, _06361_);
  and (_15339_, _15338_, _15337_);
  and (_15340_, _15339_, _07872_);
  and (_15341_, _15340_, _14539_);
  or (_40616_, _15341_, _15336_);
  nor (_15342_, _09397_, _09167_);
  or (_15343_, _15342_, _09398_);
  and (_15344_, _15343_, _07262_);
  not (_15345_, _08563_);
  nor (_15346_, _15150_, _08244_);
  or (_15347_, _15346_, _08558_);
  and (_15348_, _15347_, _15345_);
  or (_15349_, _15348_, _08569_);
  nand (_15350_, _08926_, _08246_);
  nor (_15351_, _08926_, _08246_);
  not (_15352_, _15351_);
  and (_15353_, _15352_, _15350_);
  and (_15354_, _15353_, _07238_);
  nor (_15355_, _12999_, _12998_);
  or (_15356_, _15355_, _08610_);
  nor (_15357_, _15160_, _08246_);
  or (_15358_, _15357_, _08764_);
  and (_15359_, _15358_, _07152_);
  or (_15360_, _09447_, _07155_);
  and (_15361_, _15347_, _12387_);
  nand (_15362_, _12447_, _06758_);
  or (_15363_, _06758_, \oc8051_golden_model_1.ACC [5]);
  and (_15364_, _15363_, _15362_);
  and (_15365_, _15364_, _08654_);
  or (_15366_, _15365_, _07154_);
  or (_15367_, _15366_, _15361_);
  and (_15368_, _15367_, _08652_);
  and (_15369_, _15368_, _15360_);
  or (_15370_, _15369_, _15359_);
  and (_15371_, _15370_, _08651_);
  nand (_15372_, _13000_, _12998_);
  and (_15373_, _15372_, _06275_);
  or (_15374_, _15373_, _07611_);
  or (_15375_, _15374_, _15371_);
  nor (_15376_, _12446_, _06010_);
  nor (_15377_, _15376_, _07167_);
  and (_15378_, _15377_, _15375_);
  and (_15379_, _09429_, _07167_);
  or (_15380_, _15379_, _07179_);
  or (_15381_, _15380_, _15378_);
  and (_15382_, _15381_, _15356_);
  or (_15383_, _15382_, _06267_);
  nand (_15384_, _08246_, _06267_);
  and (_15385_, _15384_, _06265_);
  and (_15386_, _15385_, _15383_);
  not (_15387_, _13001_);
  and (_15388_, _15372_, _06264_);
  and (_15389_, _15388_, _15387_);
  or (_15390_, _15389_, _15386_);
  and (_15391_, _15390_, _06007_);
  or (_15392_, _12447_, _06007_);
  nand (_15393_, _15392_, _06501_);
  or (_15394_, _15393_, _15391_);
  nand (_15395_, _08246_, _06502_);
  and (_15396_, _15395_, _15394_);
  or (_15397_, _15396_, _07197_);
  and (_15398_, _09447_, _06286_);
  nand (_15399_, _08191_, _07197_);
  or (_15400_, _15399_, _15398_);
  and (_15401_, _15400_, _08801_);
  and (_15402_, _15401_, _15397_);
  nand (_15403_, _12999_, _10558_);
  and (_15404_, _15403_, _07196_);
  and (_15405_, _15404_, _15372_);
  or (_15406_, _15405_, _06254_);
  or (_15407_, _15406_, _15402_);
  nor (_15408_, _12446_, _05978_);
  nor (_15409_, _15408_, _08812_);
  and (_15410_, _15409_, _15407_);
  nor (_15411_, _08244_, _08817_);
  or (_15412_, _15411_, _08816_);
  or (_15413_, _15412_, _15410_);
  or (_15414_, _09447_, _08821_);
  and (_15415_, _15414_, _07471_);
  and (_15416_, _15415_, _15413_);
  nor (_15417_, _08825_, _08244_);
  and (_15418_, _09005_, \oc8051_golden_model_1.SBUF [5]);
  and (_15419_, _08968_, \oc8051_golden_model_1.B [5]);
  or (_15420_, _15419_, _15418_);
  and (_15421_, _08934_, \oc8051_golden_model_1.TCON [5]);
  and (_15422_, _09007_, \oc8051_golden_model_1.PSW [5]);
  or (_15423_, _15422_, _15421_);
  or (_15424_, _15423_, _15420_);
  and (_15425_, _08944_, \oc8051_golden_model_1.P0 [5]);
  and (_15426_, _08965_, \oc8051_golden_model_1.SCON [5]);
  or (_15427_, _15426_, _15425_);
  and (_15428_, _08957_, \oc8051_golden_model_1.TMOD [5]);
  and (_15429_, _08962_, \oc8051_golden_model_1.P1 [5]);
  or (_15430_, _15429_, _15428_);
  or (_15431_, _15430_, _15427_);
  or (_15432_, _15431_, _15424_);
  and (_15433_, _08977_, \oc8051_golden_model_1.PCON [5]);
  and (_15434_, _08979_, \oc8051_golden_model_1.DPH [5]);
  or (_15435_, _15434_, _15433_);
  or (_15436_, _15435_, _15432_);
  and (_15437_, _09013_, \oc8051_golden_model_1.TH0 [5]);
  and (_15438_, _08986_, \oc8051_golden_model_1.TL1 [5]);
  and (_15439_, _08988_, \oc8051_golden_model_1.SP [5]);
  or (_15440_, _15439_, _15438_);
  or (_15441_, _15440_, _15437_);
  and (_15442_, _08999_, \oc8051_golden_model_1.P2 [5]);
  and (_15443_, _09001_, \oc8051_golden_model_1.P3 [5]);
  or (_15444_, _15443_, _15442_);
  and (_15445_, _08993_, \oc8051_golden_model_1.IE [5]);
  and (_15446_, _08996_, \oc8051_golden_model_1.IP [5]);
  or (_15447_, _15446_, _15445_);
  or (_15448_, _15447_, _15444_);
  and (_15449_, _08939_, \oc8051_golden_model_1.TL0 [5]);
  and (_15450_, _08950_, \oc8051_golden_model_1.ACC [5]);
  or (_15451_, _15450_, _15449_);
  or (_15452_, _15451_, _15448_);
  and (_15453_, _08984_, \oc8051_golden_model_1.DPL [5]);
  and (_15454_, _09015_, \oc8051_golden_model_1.TH1 [5]);
  or (_15455_, _15454_, _15453_);
  or (_15456_, _15455_, _15452_);
  or (_15457_, _15456_, _15441_);
  or (_15458_, _15457_, _15436_);
  or (_15459_, _15458_, _15417_);
  and (_15460_, _15459_, _07470_);
  or (_15461_, _15460_, _09031_);
  or (_15462_, _15461_, _15416_);
  and (_15463_, _09031_, _06611_);
  nor (_15464_, _15463_, _06220_);
  and (_15465_, _15464_, _15462_);
  and (_15466_, _08946_, _06220_);
  or (_15467_, _15466_, _06217_);
  or (_15468_, _15467_, _15465_);
  nor (_15469_, _12446_, _05952_);
  nor (_15470_, _15469_, _07238_);
  and (_15471_, _15470_, _15468_);
  or (_15472_, _15471_, _15354_);
  and (_15473_, _15472_, _08577_);
  and (_15474_, _11250_, _07241_);
  or (_15475_, _15474_, _15473_);
  and (_15476_, _15475_, _08571_);
  and (_15477_, _15351_, _07243_);
  or (_15478_, _15477_, _15476_);
  and (_15479_, _15478_, _07236_);
  and (_15480_, _11248_, _07235_);
  or (_15481_, _15480_, _07233_);
  or (_15482_, _15481_, _15479_);
  nor (_15483_, _12446_, _05961_);
  nor (_15484_, _15483_, _09057_);
  and (_15485_, _15484_, _15482_);
  and (_15486_, _15350_, _09057_);
  or (_15487_, _15486_, _09062_);
  or (_15488_, _15487_, _15485_);
  nand (_15489_, _11249_, _09062_);
  and (_15490_, _15489_, _05959_);
  and (_15491_, _15490_, _15488_);
  or (_15492_, _08567_, _08564_);
  nor (_15493_, _12447_, _05959_);
  or (_15494_, _15493_, _08566_);
  or (_15495_, _15494_, _15492_);
  or (_15496_, _15495_, _15491_);
  and (_15497_, _15496_, _15349_);
  and (_15498_, _15347_, _08563_);
  or (_15499_, _15498_, _07263_);
  or (_15500_, _15499_, _15497_);
  or (_15501_, _15343_, _14746_);
  and (_15502_, _15501_, _14745_);
  and (_15503_, _15502_, _15500_);
  or (_15504_, _15503_, _15344_);
  and (_15505_, _15504_, _09075_);
  and (_15506_, _15358_, _07261_);
  or (_15507_, _15506_, _06361_);
  or (_15508_, _15507_, _15505_);
  nand (_15509_, _12234_, _06361_);
  and (_15510_, _15509_, _14710_);
  and (_15511_, _15510_, _15508_);
  and (_15512_, _12446_, _05940_);
  or (_15513_, _15512_, _07270_);
  or (_15514_, _15513_, _15511_);
  or (_15515_, _15355_, _07539_);
  and (_15516_, _15515_, _15107_);
  and (_15517_, _15516_, _15514_);
  nor (_15518_, _09436_, _09429_);
  nor (_15519_, _15518_, _09437_);
  and (_15520_, _15519_, _15111_);
  or (_15521_, _15520_, _15115_);
  or (_15522_, _15521_, _15517_);
  or (_15523_, _15519_, _15118_);
  and (_15524_, _15523_, _07282_);
  and (_15525_, _15524_, _15522_);
  or (_15526_, _09455_, _09447_);
  nor (_15527_, _09456_, _07282_);
  and (_15528_, _15527_, _15526_);
  or (_15529_, _15528_, _07286_);
  or (_15530_, _15529_, _15525_);
  nor (_15531_, _08545_, _08247_);
  nor (_15532_, _15531_, _08546_);
  or (_15533_, _15532_, _09445_);
  and (_15534_, _15533_, _07535_);
  and (_15535_, _15534_, _15530_);
  or (_15536_, _15535_, _14360_);
  or (_15537_, _14359_, \oc8051_golden_model_1.IRAM[0] [5]);
  and (_15538_, _15537_, _14535_);
  and (_15539_, _15538_, _15536_);
  nand (_15540_, _12194_, _06361_);
  or (_15541_, _12409_, _06361_);
  and (_15542_, _15541_, _15540_);
  and (_15543_, _15542_, _07872_);
  and (_15544_, _15543_, _14539_);
  or (_40618_, _15544_, _15539_);
  nor (_15545_, _12440_, _05959_);
  nand (_15546_, _08857_, _08144_);
  nor (_15547_, _08857_, _08144_);
  not (_15548_, _15547_);
  and (_15549_, _15548_, _15546_);
  and (_15550_, _15549_, _07238_);
  nor (_15551_, _12949_, _12948_);
  or (_15552_, _15551_, _08610_);
  nor (_15553_, _08764_, _08144_);
  or (_15554_, _15553_, _08765_);
  and (_15555_, _15554_, _07152_);
  or (_15556_, _09446_, _07155_);
  nor (_15557_, _08558_, _08142_);
  or (_15558_, _15557_, _08559_);
  and (_15559_, _15558_, _12387_);
  nand (_15560_, _12440_, _06758_);
  or (_15561_, _06758_, \oc8051_golden_model_1.ACC [6]);
  and (_15562_, _15561_, _15560_);
  and (_15563_, _15562_, _08654_);
  or (_15564_, _15563_, _07154_);
  or (_15565_, _15564_, _15559_);
  and (_15566_, _15565_, _08652_);
  and (_15567_, _15566_, _15556_);
  or (_15568_, _15567_, _15555_);
  and (_15569_, _15568_, _08651_);
  nand (_15570_, _12950_, _12948_);
  and (_15571_, _15570_, _06275_);
  or (_15572_, _15571_, _07611_);
  or (_15573_, _15572_, _15569_);
  nor (_15574_, _12439_, _06010_);
  nor (_15575_, _15574_, _07167_);
  and (_15576_, _15575_, _15573_);
  and (_15577_, _09428_, _07167_);
  or (_15578_, _15577_, _07179_);
  or (_15579_, _15578_, _15576_);
  and (_15580_, _15579_, _15552_);
  or (_15581_, _15580_, _06267_);
  nand (_15582_, _08144_, _06267_);
  and (_15583_, _15582_, _06265_);
  and (_15584_, _15583_, _15581_);
  not (_15585_, _12951_);
  and (_15586_, _15570_, _15585_);
  and (_15587_, _15586_, _06264_);
  or (_15588_, _15587_, _15584_);
  and (_15589_, _15588_, _06007_);
  or (_15590_, _12440_, _06007_);
  nand (_15591_, _15590_, _06501_);
  or (_15592_, _15591_, _15589_);
  nand (_15593_, _08144_, _06502_);
  and (_15594_, _15593_, _15592_);
  or (_15595_, _15594_, _07197_);
  and (_15596_, _09446_, _06286_);
  nand (_15597_, _08089_, _07197_);
  or (_15598_, _15597_, _15596_);
  and (_15599_, _15598_, _08801_);
  and (_15600_, _15599_, _15595_);
  and (_15601_, _14802_, _06657_);
  or (_15602_, _15601_, _15551_);
  and (_15603_, _15602_, _07196_);
  or (_15604_, _15603_, _06254_);
  or (_15605_, _15604_, _15600_);
  nor (_15606_, _12439_, _05978_);
  nor (_15607_, _15606_, _08812_);
  and (_15608_, _15607_, _15605_);
  nor (_15609_, _08142_, _08817_);
  or (_15610_, _15609_, _08816_);
  or (_15611_, _15610_, _15608_);
  or (_15612_, _09446_, _08821_);
  and (_15613_, _15612_, _07471_);
  and (_15614_, _15613_, _15611_);
  nor (_15615_, _08825_, _08142_);
  and (_15616_, _08962_, \oc8051_golden_model_1.P1 [6]);
  and (_15617_, _08965_, \oc8051_golden_model_1.SCON [6]);
  or (_15618_, _15617_, _15616_);
  and (_15619_, _08944_, \oc8051_golden_model_1.P0 [6]);
  and (_15620_, _09005_, \oc8051_golden_model_1.SBUF [6]);
  or (_15621_, _15620_, _15619_);
  or (_15622_, _15621_, _15618_);
  and (_15623_, _08957_, \oc8051_golden_model_1.TMOD [6]);
  and (_15624_, _09007_, \oc8051_golden_model_1.PSW [6]);
  or (_15625_, _15624_, _15623_);
  and (_15626_, _08934_, \oc8051_golden_model_1.TCON [6]);
  and (_15627_, _08950_, \oc8051_golden_model_1.ACC [6]);
  or (_15628_, _15627_, _15626_);
  or (_15629_, _15628_, _15625_);
  or (_15630_, _15629_, _15622_);
  and (_15631_, _08977_, \oc8051_golden_model_1.PCON [6]);
  and (_15632_, _08979_, \oc8051_golden_model_1.DPH [6]);
  or (_15633_, _15632_, _15631_);
  or (_15634_, _15633_, _15630_);
  and (_15635_, _08986_, \oc8051_golden_model_1.TL1 [6]);
  and (_15636_, _08984_, \oc8051_golden_model_1.DPL [6]);
  and (_15637_, _09015_, \oc8051_golden_model_1.TH1 [6]);
  or (_15638_, _15637_, _15636_);
  or (_15639_, _15638_, _15635_);
  and (_15640_, _08999_, \oc8051_golden_model_1.P2 [6]);
  and (_15641_, _09001_, \oc8051_golden_model_1.P3 [6]);
  or (_15642_, _15641_, _15640_);
  and (_15643_, _08993_, \oc8051_golden_model_1.IE [6]);
  and (_15644_, _08996_, \oc8051_golden_model_1.IP [6]);
  or (_15645_, _15644_, _15643_);
  or (_15646_, _15645_, _15642_);
  and (_15647_, _08939_, \oc8051_golden_model_1.TL0 [6]);
  and (_15648_, _08968_, \oc8051_golden_model_1.B [6]);
  or (_15649_, _15648_, _15647_);
  or (_15650_, _15649_, _15646_);
  and (_15651_, _09013_, \oc8051_golden_model_1.TH0 [6]);
  and (_15652_, _08988_, \oc8051_golden_model_1.SP [6]);
  or (_15653_, _15652_, _15651_);
  or (_15654_, _15653_, _15650_);
  or (_15655_, _15654_, _15639_);
  or (_15656_, _15655_, _15634_);
  or (_15657_, _15656_, _15615_);
  and (_15658_, _15657_, _07470_);
  or (_15659_, _15658_, _09031_);
  or (_15660_, _15659_, _15614_);
  and (_15661_, _09031_, _06317_);
  nor (_15662_, _15661_, _06220_);
  and (_15663_, _15662_, _15660_);
  not (_15664_, _08857_);
  and (_15665_, _15664_, _06220_);
  or (_15666_, _15665_, _06217_);
  or (_15667_, _15666_, _15663_);
  nor (_15668_, _12439_, _05952_);
  nor (_15669_, _15668_, _07238_);
  and (_15670_, _15669_, _15667_);
  or (_15671_, _15670_, _15550_);
  and (_15672_, _15671_, _08577_);
  and (_15673_, _11247_, _07241_);
  or (_15674_, _15673_, _15672_);
  and (_15675_, _15674_, _08571_);
  and (_15676_, _15547_, _07243_);
  or (_15677_, _15676_, _15675_);
  and (_15678_, _15677_, _07236_);
  and (_15679_, _11244_, _07235_);
  or (_15680_, _15679_, _07233_);
  or (_15681_, _15680_, _15678_);
  nor (_15682_, _12439_, _05961_);
  nor (_15683_, _15682_, _09057_);
  and (_15684_, _15683_, _15681_);
  and (_15685_, _15546_, _09057_);
  or (_15686_, _15685_, _09062_);
  or (_15687_, _15686_, _15684_);
  nand (_15688_, _11246_, _09062_);
  and (_15689_, _15688_, _05959_);
  and (_15690_, _15689_, _15687_);
  or (_15691_, _15690_, _15545_);
  and (_15692_, _15691_, _08568_);
  not (_15693_, _08568_);
  and (_15694_, _15558_, _15693_);
  or (_15695_, _15694_, _07292_);
  or (_15696_, _15695_, _15692_);
  or (_15697_, _15558_, _08565_);
  and (_15698_, _15697_, _14746_);
  and (_15699_, _15698_, _15696_);
  nor (_15700_, _09398_, _09122_);
  or (_15701_, _15700_, _09399_);
  or (_15702_, _15701_, _07262_);
  and (_15703_, _15702_, _07435_);
  or (_15704_, _15703_, _15699_);
  or (_15705_, _15701_, _14745_);
  and (_15706_, _15705_, _09075_);
  and (_15707_, _15706_, _15704_);
  and (_15708_, _15554_, _07261_);
  or (_15709_, _15708_, _06361_);
  or (_15710_, _15709_, _15707_);
  nand (_15711_, _12226_, _06361_);
  and (_15712_, _15711_, _14710_);
  and (_15713_, _15712_, _15710_);
  and (_15714_, _12439_, _05940_);
  or (_15715_, _15714_, _07270_);
  or (_15716_, _15715_, _15713_);
  or (_15717_, _15551_, _07539_);
  and (_15718_, _15717_, _09427_);
  and (_15719_, _15718_, _15716_);
  nor (_15720_, _09437_, _09428_);
  nor (_15721_, _15720_, _09438_);
  and (_15722_, _15721_, _09424_);
  or (_15723_, _15722_, _07280_);
  or (_15724_, _15723_, _15719_);
  nor (_15725_, _09456_, _09446_);
  nor (_15726_, _15725_, _09457_);
  or (_15727_, _15726_, _14741_);
  and (_15728_, _15727_, _14737_);
  and (_15729_, _15728_, _15724_);
  and (_15730_, _15726_, _07279_);
  or (_15731_, _15730_, _07286_);
  or (_15732_, _15731_, _15729_);
  nor (_15733_, _08546_, _08145_);
  nor (_15734_, _15733_, _08547_);
  or (_15735_, _15734_, _09445_);
  and (_15736_, _15735_, _07535_);
  and (_15737_, _15736_, _15732_);
  or (_15738_, _15737_, _14360_);
  or (_15739_, _14359_, \oc8051_golden_model_1.IRAM[0] [6]);
  and (_15740_, _15739_, _14535_);
  and (_15741_, _15740_, _15738_);
  or (_15742_, _12186_, _14508_);
  or (_15743_, _12403_, _06361_);
  and (_15744_, _15743_, _15742_);
  and (_15745_, _15744_, _07872_);
  and (_15746_, _15745_, _14539_);
  or (_40619_, _15746_, _15741_);
  nand (_15747_, _14359_, _09464_);
  or (_15748_, _14359_, _07980_);
  and (_15749_, _15748_, _14535_);
  nand (_15750_, _15749_, _15747_);
  or (_15751_, _14535_, _09489_);
  and (_40620_, _15751_, _15750_);
  and (_15752_, _14354_, _07453_);
  and (_15753_, _15752_, _14357_);
  not (_15754_, _15753_);
  or (_15755_, _15754_, _14528_);
  or (_15756_, _15753_, \oc8051_golden_model_1.IRAM[1] [0]);
  nand (_15757_, _14533_, _07598_);
  or (_15758_, _15757_, _14531_);
  and (_15759_, _15758_, _15756_);
  and (_15760_, _15759_, _15755_);
  and (_15761_, _07872_, _07598_);
  and (_15762_, _15761_, _14533_);
  and (_15763_, _15762_, _14543_);
  or (_40623_, _15763_, _15760_);
  or (_15764_, _15754_, _14727_);
  or (_15765_, _15753_, \oc8051_golden_model_1.IRAM[1] [1]);
  and (_15766_, _15765_, _15758_);
  and (_15767_, _15766_, _15764_);
  and (_15768_, _15762_, _14735_);
  or (_40626_, _15768_, _15767_);
  or (_15769_, _15754_, _14929_);
  or (_15770_, _15753_, \oc8051_golden_model_1.IRAM[1] [2]);
  and (_15771_, _15770_, _15758_);
  and (_15772_, _15771_, _15769_);
  and (_15773_, _15762_, _14937_);
  or (_40627_, _15773_, _15772_);
  or (_15774_, _15754_, _15131_);
  or (_15775_, _15753_, \oc8051_golden_model_1.IRAM[1] [3]);
  and (_15776_, _15775_, _15758_);
  and (_15777_, _15776_, _15774_);
  and (_15778_, _15762_, _15139_);
  or (_40628_, _15778_, _15777_);
  or (_15779_, _15754_, _15332_);
  or (_15780_, _15753_, \oc8051_golden_model_1.IRAM[1] [4]);
  and (_15781_, _15780_, _15758_);
  and (_15782_, _15781_, _15779_);
  and (_15783_, _15762_, _15340_);
  or (_40629_, _15783_, _15782_);
  or (_15784_, _15754_, _15535_);
  or (_15785_, _15753_, \oc8051_golden_model_1.IRAM[1] [5]);
  and (_15786_, _15785_, _15758_);
  and (_15787_, _15786_, _15784_);
  and (_15788_, _15762_, _15543_);
  or (_40630_, _15788_, _15787_);
  or (_15789_, _15754_, _15737_);
  or (_15790_, _15753_, \oc8051_golden_model_1.IRAM[1] [6]);
  and (_15791_, _15790_, _15758_);
  and (_15792_, _15791_, _15789_);
  and (_15793_, _15762_, _15745_);
  or (_40632_, _15793_, _15792_);
  or (_15794_, _15754_, _09465_);
  or (_15795_, _15753_, \oc8051_golden_model_1.IRAM[1] [7]);
  and (_15796_, _15795_, _15758_);
  and (_15797_, _15796_, _15794_);
  and (_15798_, _15762_, _09490_);
  or (_40633_, _15798_, _15797_);
  not (_15799_, _07537_);
  nor (_15800_, _15799_, _07289_);
  and (_15801_, _15800_, _14357_);
  not (_15802_, _15801_);
  or (_15803_, _15802_, _14528_);
  or (_15804_, _15801_, \oc8051_golden_model_1.IRAM[2] [0]);
  nand (_15805_, _14533_, _08668_);
  or (_15806_, _15805_, _14531_);
  and (_15807_, _15806_, _15804_);
  and (_15808_, _15807_, _15803_);
  and (_15809_, _08668_, _07872_);
  and (_15810_, _15809_, _14533_);
  and (_15811_, _15810_, _14543_);
  or (_40637_, _15811_, _15808_);
  or (_15812_, _15802_, _14727_);
  or (_15813_, _15801_, \oc8051_golden_model_1.IRAM[2] [1]);
  and (_15814_, _15813_, _15806_);
  and (_15815_, _15814_, _15812_);
  and (_15816_, _15810_, _14735_);
  or (_40638_, _15816_, _15815_);
  or (_15817_, _15802_, _14929_);
  or (_15818_, _15801_, \oc8051_golden_model_1.IRAM[2] [2]);
  and (_15819_, _15818_, _15806_);
  and (_15820_, _15819_, _15817_);
  and (_15821_, _15810_, _14937_);
  or (_40640_, _15821_, _15820_);
  or (_15822_, _15802_, _15131_);
  or (_15823_, _15801_, \oc8051_golden_model_1.IRAM[2] [3]);
  and (_15824_, _15823_, _15806_);
  and (_15825_, _15824_, _15822_);
  and (_15826_, _15810_, _15139_);
  or (_40641_, _15826_, _15825_);
  or (_15827_, _15802_, _15332_);
  or (_15828_, _15801_, \oc8051_golden_model_1.IRAM[2] [4]);
  and (_15829_, _15828_, _15806_);
  and (_15830_, _15829_, _15827_);
  and (_15831_, _15810_, _15340_);
  or (_40642_, _15831_, _15830_);
  or (_15832_, _15802_, _15535_);
  or (_15833_, _15801_, \oc8051_golden_model_1.IRAM[2] [5]);
  and (_15834_, _15833_, _15806_);
  and (_15835_, _15834_, _15832_);
  and (_15836_, _15810_, _15543_);
  or (_40643_, _15836_, _15835_);
  or (_15837_, _15802_, _15737_);
  or (_15838_, _15801_, \oc8051_golden_model_1.IRAM[2] [6]);
  and (_15839_, _15838_, _15806_);
  and (_15840_, _15839_, _15837_);
  and (_15841_, _15810_, _15745_);
  or (_40644_, _15841_, _15840_);
  or (_15842_, _15802_, _09465_);
  or (_15843_, _15801_, \oc8051_golden_model_1.IRAM[2] [7]);
  and (_15844_, _15843_, _15806_);
  and (_15845_, _15844_, _15842_);
  and (_15846_, _15810_, _09490_);
  or (_40646_, _15846_, _15845_);
  and (_15847_, _14357_, _07538_);
  or (_15848_, _15847_, \oc8051_golden_model_1.IRAM[3] [0]);
  nand (_15849_, _14533_, _07295_);
  or (_15850_, _15849_, _14531_);
  and (_15851_, _15850_, _15848_);
  not (_15852_, _15847_);
  or (_15853_, _15852_, _14528_);
  and (_15854_, _15853_, _15851_);
  and (_15855_, _07872_, _07295_);
  and (_15856_, _15855_, _14533_);
  and (_15857_, _15856_, _14543_);
  or (_40649_, _15857_, _15854_);
  or (_15858_, _15847_, \oc8051_golden_model_1.IRAM[3] [1]);
  and (_15859_, _15858_, _15850_);
  or (_15860_, _15852_, _14727_);
  and (_15861_, _15860_, _15859_);
  and (_15862_, _15856_, _14735_);
  or (_40651_, _15862_, _15861_);
  nor (_15863_, _15847_, _07728_);
  and (_15864_, _15847_, _14929_);
  or (_15865_, _15864_, _15863_);
  and (_15866_, _15865_, _15850_);
  and (_15867_, _15856_, _14937_);
  or (_40652_, _15867_, _15866_);
  or (_15868_, _15847_, \oc8051_golden_model_1.IRAM[3] [3]);
  and (_15869_, _15868_, _15850_);
  or (_15870_, _15852_, _15131_);
  and (_15871_, _15870_, _15869_);
  and (_15872_, _15856_, _15139_);
  or (_40653_, _15872_, _15871_);
  or (_15873_, _15847_, \oc8051_golden_model_1.IRAM[3] [4]);
  and (_15874_, _15873_, _15850_);
  or (_15875_, _15852_, _15332_);
  and (_15876_, _15875_, _15874_);
  and (_15877_, _15856_, _15340_);
  or (_40654_, _15877_, _15876_);
  or (_15878_, _15847_, \oc8051_golden_model_1.IRAM[3] [5]);
  and (_15879_, _15878_, _15850_);
  or (_15880_, _15852_, _15535_);
  and (_15881_, _15880_, _15879_);
  and (_15882_, _15856_, _15543_);
  or (_40655_, _15882_, _15881_);
  or (_15883_, _15847_, \oc8051_golden_model_1.IRAM[3] [6]);
  and (_15884_, _15883_, _15850_);
  or (_15885_, _15852_, _15737_);
  and (_15886_, _15885_, _15884_);
  and (_15887_, _15856_, _15745_);
  or (_40657_, _15887_, _15886_);
  or (_15888_, _15847_, \oc8051_golden_model_1.IRAM[3] [7]);
  and (_15889_, _15888_, _15850_);
  or (_15890_, _15852_, _09465_);
  and (_15891_, _15890_, _15889_);
  and (_15892_, _15856_, _09490_);
  or (_40658_, _15892_, _15891_);
  and (_15893_, _07859_, _07711_);
  and (_15894_, _15893_, _14355_);
  not (_15895_, _15894_);
  or (_15896_, _15895_, _14528_);
  not (_15897_, _07869_);
  and (_15898_, _14532_, _15897_);
  and (_15899_, _15898_, _07296_);
  not (_15900_, _15899_);
  or (_15901_, _15894_, \oc8051_golden_model_1.IRAM[4] [0]);
  and (_15902_, _15901_, _15900_);
  and (_15903_, _15902_, _15896_);
  and (_15904_, _15899_, _14543_);
  or (_40662_, _15904_, _15903_);
  or (_15905_, _15895_, _14727_);
  or (_15906_, _15894_, \oc8051_golden_model_1.IRAM[4] [1]);
  and (_15907_, _15906_, _15900_);
  and (_15908_, _15907_, _15905_);
  and (_15909_, _15899_, _14735_);
  or (_40663_, _15909_, _15908_);
  or (_15910_, _15895_, _14929_);
  or (_15911_, _15894_, \oc8051_golden_model_1.IRAM[4] [2]);
  and (_15912_, _15911_, _15900_);
  and (_15913_, _15912_, _15910_);
  and (_15914_, _15899_, _14937_);
  or (_40665_, _15914_, _15913_);
  or (_15915_, _15895_, _15131_);
  or (_15916_, _15894_, \oc8051_golden_model_1.IRAM[4] [3]);
  and (_15917_, _15916_, _15900_);
  and (_15918_, _15917_, _15915_);
  and (_15919_, _15899_, _15139_);
  or (_40666_, _15919_, _15918_);
  or (_15920_, _15895_, _15332_);
  or (_15921_, _15894_, \oc8051_golden_model_1.IRAM[4] [4]);
  and (_15922_, _15921_, _15900_);
  and (_15923_, _15922_, _15920_);
  and (_15924_, _15899_, _15340_);
  or (_40667_, _15924_, _15923_);
  or (_15925_, _15895_, _15535_);
  or (_15926_, _15894_, \oc8051_golden_model_1.IRAM[4] [5]);
  and (_15927_, _15926_, _15900_);
  and (_15928_, _15927_, _15925_);
  and (_15929_, _15899_, _15543_);
  or (_40668_, _15929_, _15928_);
  or (_15930_, _15895_, _15737_);
  or (_15931_, _15894_, \oc8051_golden_model_1.IRAM[4] [6]);
  and (_15932_, _15931_, _15900_);
  and (_15933_, _15932_, _15930_);
  and (_15934_, _15899_, _15745_);
  or (_40669_, _15934_, _15933_);
  or (_15935_, _15895_, _09465_);
  or (_15936_, _15894_, \oc8051_golden_model_1.IRAM[4] [7]);
  and (_15937_, _15936_, _15900_);
  and (_15938_, _15937_, _15935_);
  and (_15939_, _15899_, _09490_);
  or (_40671_, _15939_, _15938_);
  and (_15940_, _15893_, _15752_);
  not (_15941_, _15940_);
  or (_15942_, _15941_, _14528_);
  and (_15943_, _15898_, _07598_);
  not (_15944_, _15943_);
  or (_15945_, _15940_, \oc8051_golden_model_1.IRAM[5] [0]);
  and (_15946_, _15945_, _15944_);
  and (_15947_, _15946_, _15942_);
  and (_15948_, _15943_, _14543_);
  or (_40673_, _15948_, _15947_);
  or (_15949_, _15941_, _14727_);
  or (_15950_, _15940_, \oc8051_golden_model_1.IRAM[5] [1]);
  and (_15951_, _15950_, _15944_);
  and (_15952_, _15951_, _15949_);
  and (_15953_, _15943_, _14735_);
  or (_40674_, _15953_, _15952_);
  or (_15954_, _15941_, _14929_);
  or (_15955_, _15940_, \oc8051_golden_model_1.IRAM[5] [2]);
  and (_15956_, _15955_, _15944_);
  and (_15957_, _15956_, _15954_);
  and (_15958_, _15943_, _14937_);
  or (_40677_, _15958_, _15957_);
  or (_15959_, _15941_, _15131_);
  or (_15960_, _15940_, \oc8051_golden_model_1.IRAM[5] [3]);
  and (_15961_, _15960_, _15944_);
  and (_15962_, _15961_, _15959_);
  and (_15963_, _15943_, _15139_);
  or (_40678_, _15963_, _15962_);
  or (_15964_, _15941_, _15332_);
  or (_15965_, _15940_, \oc8051_golden_model_1.IRAM[5] [4]);
  and (_15966_, _15965_, _15944_);
  and (_15967_, _15966_, _15964_);
  and (_15968_, _15943_, _15340_);
  or (_40679_, _15968_, _15967_);
  or (_15969_, _15941_, _15535_);
  or (_15970_, _15940_, \oc8051_golden_model_1.IRAM[5] [5]);
  and (_15971_, _15970_, _15944_);
  and (_15972_, _15971_, _15969_);
  and (_15973_, _15943_, _15543_);
  or (_40680_, _15973_, _15972_);
  or (_15974_, _15941_, _15737_);
  or (_15975_, _15940_, \oc8051_golden_model_1.IRAM[5] [6]);
  and (_15976_, _15975_, _15944_);
  and (_15977_, _15976_, _15974_);
  and (_15978_, _15943_, _15745_);
  or (_40681_, _15978_, _15977_);
  or (_15979_, _15941_, _09465_);
  or (_15980_, _15940_, \oc8051_golden_model_1.IRAM[5] [7]);
  and (_15981_, _15980_, _15944_);
  and (_15982_, _15981_, _15979_);
  and (_15983_, _15943_, _09490_);
  or (_40683_, _15983_, _15982_);
  and (_15984_, _15893_, _15800_);
  not (_15985_, _15984_);
  or (_15986_, _15985_, _14528_);
  and (_15987_, _15898_, _08668_);
  not (_15988_, _15987_);
  or (_15989_, _15984_, \oc8051_golden_model_1.IRAM[6] [0]);
  and (_15990_, _15989_, _15988_);
  and (_15991_, _15990_, _15986_);
  and (_15992_, _15987_, _14543_);
  or (_40685_, _15992_, _15991_);
  or (_15993_, _15985_, _14727_);
  or (_15994_, _15984_, \oc8051_golden_model_1.IRAM[6] [1]);
  and (_15995_, _15994_, _15988_);
  and (_15996_, _15995_, _15993_);
  and (_15997_, _15987_, _14735_);
  or (_40688_, _15997_, _15996_);
  or (_15998_, _15985_, _14929_);
  or (_15999_, _15984_, \oc8051_golden_model_1.IRAM[6] [2]);
  and (_16000_, _15999_, _15988_);
  and (_16001_, _16000_, _15998_);
  and (_16002_, _15987_, _14937_);
  or (_40689_, _16002_, _16001_);
  or (_16003_, _15985_, _15131_);
  or (_16004_, _15984_, \oc8051_golden_model_1.IRAM[6] [3]);
  and (_16005_, _16004_, _15988_);
  and (_16006_, _16005_, _16003_);
  and (_16007_, _15987_, _15139_);
  or (_40690_, _16007_, _16006_);
  or (_16008_, _15985_, _15332_);
  or (_16009_, _15984_, \oc8051_golden_model_1.IRAM[6] [4]);
  and (_16010_, _16009_, _15988_);
  and (_16011_, _16010_, _16008_);
  and (_16012_, _15987_, _15340_);
  or (_40691_, _16012_, _16011_);
  or (_16013_, _15985_, _15535_);
  or (_16014_, _15984_, \oc8051_golden_model_1.IRAM[6] [5]);
  and (_16015_, _16014_, _15988_);
  and (_16016_, _16015_, _16013_);
  and (_16017_, _15987_, _15543_);
  or (_40692_, _16017_, _16016_);
  or (_16018_, _15985_, _15737_);
  or (_16019_, _15984_, \oc8051_golden_model_1.IRAM[6] [6]);
  and (_16020_, _16019_, _15988_);
  and (_16021_, _16020_, _16018_);
  and (_16022_, _15987_, _15745_);
  or (_40694_, _16022_, _16021_);
  or (_16023_, _15985_, _09465_);
  or (_16024_, _15984_, \oc8051_golden_model_1.IRAM[6] [7]);
  and (_16025_, _16024_, _15988_);
  and (_16026_, _16025_, _16023_);
  and (_16027_, _15987_, _09490_);
  or (_40695_, _16027_, _16026_);
  and (_16028_, _15898_, _07295_);
  not (_16029_, _16028_);
  or (_16030_, _16029_, _14543_);
  and (_16031_, _15893_, _07538_);
  and (_16032_, _16031_, _14528_);
  nor (_16033_, _16031_, _07092_);
  or (_16034_, _16033_, _16028_);
  or (_16035_, _16034_, _16032_);
  and (_40698_, _16035_, _16030_);
  or (_16036_, _16031_, \oc8051_golden_model_1.IRAM[7] [1]);
  and (_16037_, _16036_, _16029_);
  not (_16038_, _16031_);
  or (_16039_, _16038_, _14727_);
  and (_16040_, _16039_, _16037_);
  and (_16041_, _16028_, _14735_);
  or (_40700_, _16041_, _16040_);
  nor (_16042_, _16031_, _07736_);
  and (_16043_, _16031_, _14929_);
  or (_16044_, _16043_, _16042_);
  and (_16045_, _16044_, _16029_);
  and (_16046_, _16028_, _14937_);
  or (_40701_, _16046_, _16045_);
  or (_16047_, _16038_, _15131_);
  or (_16048_, _16031_, \oc8051_golden_model_1.IRAM[7] [3]);
  and (_16049_, _16048_, _16029_);
  and (_16050_, _16049_, _16047_);
  and (_16051_, _16028_, _15139_);
  or (_40702_, _16051_, _16050_);
  or (_16052_, _16031_, \oc8051_golden_model_1.IRAM[7] [4]);
  and (_16053_, _16052_, _16029_);
  or (_16054_, _16038_, _15332_);
  and (_16055_, _16054_, _16053_);
  and (_16056_, _16028_, _15340_);
  or (_40703_, _16056_, _16055_);
  or (_16057_, _16038_, _15535_);
  or (_16058_, _16031_, \oc8051_golden_model_1.IRAM[7] [5]);
  and (_16059_, _16058_, _16029_);
  and (_16060_, _16059_, _16057_);
  and (_16061_, _16028_, _15543_);
  or (_40704_, _16061_, _16060_);
  or (_16062_, _16031_, \oc8051_golden_model_1.IRAM[7] [6]);
  and (_16063_, _16062_, _16029_);
  or (_16064_, _16038_, _15737_);
  and (_16065_, _16064_, _16063_);
  and (_16066_, _16028_, _15745_);
  or (_40706_, _16066_, _16065_);
  or (_16067_, _16031_, \oc8051_golden_model_1.IRAM[7] [7]);
  and (_16068_, _16067_, _16029_);
  or (_16069_, _16038_, _09465_);
  and (_16070_, _16069_, _16068_);
  and (_16071_, _16028_, _09490_);
  or (_40707_, _16071_, _16070_);
  and (_16072_, _14356_, _07858_);
  and (_16073_, _16072_, _14355_);
  not (_16074_, _16073_);
  or (_16075_, _16074_, _14528_);
  or (_16076_, _16073_, \oc8051_golden_model_1.IRAM[8] [0]);
  not (_16077_, _07873_);
  or (_16078_, _16077_, _07864_);
  and (_16079_, _16078_, _16076_);
  and (_16080_, _16079_, _16075_);
  not (_16081_, _07866_);
  and (_16082_, _07873_, _16081_);
  and (_16083_, _16082_, _07296_);
  and (_16084_, _16083_, _14543_);
  or (_40711_, _16084_, _16080_);
  or (_16085_, _16074_, _14727_);
  or (_16086_, _16073_, \oc8051_golden_model_1.IRAM[8] [1]);
  and (_16087_, _16086_, _16078_);
  and (_16088_, _16087_, _16085_);
  and (_16089_, _16083_, _14735_);
  or (_40712_, _16089_, _16088_);
  or (_16090_, _16074_, _14929_);
  or (_16091_, _16073_, \oc8051_golden_model_1.IRAM[8] [2]);
  and (_16092_, _16091_, _16078_);
  and (_16093_, _16092_, _16090_);
  and (_16094_, _16083_, _14937_);
  or (_40714_, _16094_, _16093_);
  or (_16095_, _16074_, _15131_);
  or (_16096_, _16073_, \oc8051_golden_model_1.IRAM[8] [3]);
  and (_16097_, _16096_, _16078_);
  and (_16098_, _16097_, _16095_);
  and (_16099_, _16083_, _15139_);
  or (_40715_, _16099_, _16098_);
  or (_16100_, _16074_, _15332_);
  or (_16101_, _16073_, \oc8051_golden_model_1.IRAM[8] [4]);
  and (_16102_, _16101_, _16078_);
  and (_16103_, _16102_, _16100_);
  and (_16104_, _16083_, _15340_);
  or (_40716_, _16104_, _16103_);
  or (_16105_, _16074_, _15535_);
  or (_16106_, _16073_, \oc8051_golden_model_1.IRAM[8] [5]);
  and (_16107_, _16106_, _16078_);
  and (_16108_, _16107_, _16105_);
  and (_16109_, _16083_, _15543_);
  or (_40717_, _16109_, _16108_);
  or (_16110_, _16074_, _15737_);
  or (_16111_, _16073_, \oc8051_golden_model_1.IRAM[8] [6]);
  and (_16112_, _16111_, _16078_);
  and (_16113_, _16112_, _16110_);
  and (_16114_, _16083_, _15745_);
  or (_40718_, _16114_, _16113_);
  or (_16115_, _16074_, _09465_);
  or (_16116_, _16073_, \oc8051_golden_model_1.IRAM[8] [7]);
  and (_16117_, _16116_, _16078_);
  and (_16118_, _16117_, _16115_);
  and (_16119_, _16083_, _09490_);
  or (_40720_, _16119_, _16118_);
  and (_16120_, _16072_, _15752_);
  not (_16121_, _16120_);
  or (_16122_, _16121_, _14528_);
  or (_16123_, _16120_, \oc8051_golden_model_1.IRAM[9] [0]);
  nand (_16124_, _07873_, _07599_);
  and (_16125_, _16124_, _16123_);
  and (_16126_, _16125_, _16122_);
  and (_16127_, _16082_, _07598_);
  and (_16128_, _16127_, _14543_);
  or (_40723_, _16128_, _16126_);
  or (_16129_, _16121_, _14727_);
  or (_16130_, _16120_, \oc8051_golden_model_1.IRAM[9] [1]);
  and (_16131_, _16130_, _16124_);
  and (_16132_, _16131_, _16129_);
  and (_16133_, _16127_, _14735_);
  or (_40724_, _16133_, _16132_);
  or (_16134_, _16121_, _14929_);
  or (_16135_, _16120_, \oc8051_golden_model_1.IRAM[9] [2]);
  and (_16136_, _16135_, _16124_);
  and (_16137_, _16136_, _16134_);
  and (_16138_, _16127_, _14937_);
  or (_40726_, _16138_, _16137_);
  or (_16139_, _16121_, _15131_);
  or (_16140_, _16120_, \oc8051_golden_model_1.IRAM[9] [3]);
  and (_16141_, _16140_, _16124_);
  and (_16142_, _16141_, _16139_);
  and (_16143_, _16127_, _15139_);
  or (_40727_, _16143_, _16142_);
  or (_16144_, _16121_, _15332_);
  or (_16145_, _16120_, \oc8051_golden_model_1.IRAM[9] [4]);
  and (_16146_, _16145_, _16124_);
  and (_16147_, _16146_, _16144_);
  and (_16148_, _16127_, _15340_);
  or (_40728_, _16148_, _16147_);
  or (_16149_, _16121_, _15535_);
  or (_16150_, _16120_, \oc8051_golden_model_1.IRAM[9] [5]);
  and (_16151_, _16150_, _16124_);
  and (_16152_, _16151_, _16149_);
  and (_16153_, _16127_, _15543_);
  or (_40729_, _16153_, _16152_);
  or (_16154_, _16121_, _15737_);
  or (_16155_, _16120_, \oc8051_golden_model_1.IRAM[9] [6]);
  and (_16156_, _16155_, _16124_);
  and (_16157_, _16156_, _16154_);
  and (_16158_, _16127_, _15745_);
  or (_40730_, _16158_, _16157_);
  or (_16159_, _16121_, _09465_);
  or (_16160_, _16120_, \oc8051_golden_model_1.IRAM[9] [7]);
  and (_16161_, _16160_, _16124_);
  and (_16162_, _16161_, _16159_);
  and (_16163_, _16127_, _09490_);
  or (_40732_, _16163_, _16162_);
  and (_16164_, _16072_, _15800_);
  not (_16165_, _16164_);
  or (_16166_, _16165_, _14528_);
  or (_16167_, _16164_, \oc8051_golden_model_1.IRAM[10] [0]);
  and (_16168_, _16082_, _08668_);
  not (_16169_, _16168_);
  and (_16170_, _16169_, _16167_);
  and (_16171_, _16170_, _16166_);
  and (_16172_, _16168_, _14543_);
  or (_40734_, _16172_, _16171_);
  or (_16173_, _16165_, _14727_);
  or (_16174_, _16164_, \oc8051_golden_model_1.IRAM[10] [1]);
  and (_16175_, _16174_, _16169_);
  and (_16176_, _16175_, _16173_);
  and (_16177_, _16168_, _14735_);
  or (_40736_, _16177_, _16176_);
  or (_16178_, _16165_, _14929_);
  or (_16179_, _16164_, \oc8051_golden_model_1.IRAM[10] [2]);
  and (_16180_, _16179_, _16169_);
  and (_16181_, _16180_, _16178_);
  and (_16182_, _16168_, _14937_);
  or (_40737_, _16182_, _16181_);
  or (_16183_, _16165_, _15131_);
  or (_16184_, _16164_, \oc8051_golden_model_1.IRAM[10] [3]);
  and (_16185_, _16184_, _16169_);
  and (_16186_, _16185_, _16183_);
  and (_16187_, _16168_, _15139_);
  or (_40738_, _16187_, _16186_);
  or (_16188_, _16165_, _15332_);
  or (_16189_, _16164_, \oc8051_golden_model_1.IRAM[10] [4]);
  and (_16190_, _16189_, _16169_);
  and (_16191_, _16190_, _16188_);
  and (_16192_, _16168_, _15340_);
  or (_40739_, _16192_, _16191_);
  or (_16193_, _16165_, _15535_);
  or (_16194_, _16164_, \oc8051_golden_model_1.IRAM[10] [5]);
  and (_16195_, _16194_, _16169_);
  and (_16196_, _16195_, _16193_);
  and (_16197_, _16168_, _15543_);
  or (_40740_, _16197_, _16196_);
  or (_16198_, _16165_, _15737_);
  or (_16199_, _16164_, \oc8051_golden_model_1.IRAM[10] [6]);
  and (_16200_, _16199_, _16169_);
  and (_16201_, _16200_, _16198_);
  and (_16202_, _16168_, _15745_);
  or (_40742_, _16202_, _16201_);
  or (_16203_, _16165_, _09465_);
  or (_16204_, _16164_, \oc8051_golden_model_1.IRAM[10] [7]);
  and (_16205_, _16204_, _16169_);
  and (_16206_, _16205_, _16203_);
  and (_16207_, _16168_, _09490_);
  or (_40743_, _16207_, _16206_);
  not (_16208_, _07453_);
  and (_16209_, _14354_, _16208_);
  and (_16210_, _16072_, _16209_);
  not (_16211_, _16210_);
  or (_16212_, _16211_, _14528_);
  and (_16213_, _16082_, _07295_);
  not (_16214_, _16213_);
  or (_16215_, _16210_, \oc8051_golden_model_1.IRAM[11] [0]);
  and (_16216_, _16215_, _16214_);
  and (_16217_, _16216_, _16212_);
  and (_16218_, _16213_, _14543_);
  or (_40746_, _16218_, _16217_);
  and (_16219_, _16072_, _07538_);
  or (_16220_, _16219_, \oc8051_golden_model_1.IRAM[11] [1]);
  and (_16221_, _16220_, _16214_);
  not (_16222_, _16219_);
  or (_16223_, _16222_, _14727_);
  and (_16224_, _16223_, _16221_);
  and (_16225_, _16213_, _14735_);
  or (_40748_, _16225_, _16224_);
  or (_16226_, _16211_, _14929_);
  or (_16227_, _16210_, \oc8051_golden_model_1.IRAM[11] [2]);
  and (_16228_, _16227_, _16214_);
  and (_16229_, _16228_, _16226_);
  and (_16230_, _16213_, _14937_);
  or (_40749_, _16230_, _16229_);
  or (_16231_, _16219_, \oc8051_golden_model_1.IRAM[11] [3]);
  and (_16232_, _16231_, _16214_);
  or (_16233_, _16222_, _15131_);
  and (_16234_, _16233_, _16232_);
  and (_16235_, _16213_, _15139_);
  or (_40750_, _16235_, _16234_);
  or (_16236_, _16219_, \oc8051_golden_model_1.IRAM[11] [4]);
  and (_16237_, _16236_, _16214_);
  or (_16238_, _16222_, _15332_);
  and (_16239_, _16238_, _16237_);
  and (_16240_, _16213_, _15340_);
  or (_40751_, _16240_, _16239_);
  or (_16241_, _16219_, \oc8051_golden_model_1.IRAM[11] [5]);
  and (_16242_, _16241_, _16214_);
  or (_16243_, _16222_, _15535_);
  and (_16244_, _16243_, _16242_);
  and (_16245_, _16213_, _15543_);
  or (_40752_, _16245_, _16244_);
  or (_16246_, _16219_, \oc8051_golden_model_1.IRAM[11] [6]);
  and (_16247_, _16246_, _16214_);
  or (_16248_, _16222_, _15737_);
  and (_16249_, _16248_, _16247_);
  and (_16250_, _16213_, _15745_);
  or (_40754_, _16250_, _16249_);
  or (_16251_, _16219_, \oc8051_golden_model_1.IRAM[11] [7]);
  and (_16252_, _16251_, _16214_);
  or (_16253_, _16222_, _09465_);
  and (_16254_, _16253_, _16252_);
  and (_16255_, _16213_, _09490_);
  or (_40755_, _16255_, _16254_);
  not (_16256_, _07296_);
  nand (_16257_, _14532_, _07869_);
  or (_16258_, _16257_, _16256_);
  nor (_16259_, _16258_, _14543_);
  and (_16260_, _14355_, _07861_);
  nand (_16261_, _16260_, _14528_);
  or (_16262_, _16260_, _07124_);
  and (_16263_, _16262_, _16258_);
  and (_16264_, _16263_, _16261_);
  nor (_40759_, _16264_, _16259_);
  and (_16265_, _07874_, _07296_);
  not (_16266_, _16265_);
  or (_16267_, _16260_, \oc8051_golden_model_1.IRAM[12] [1]);
  and (_16268_, _16267_, _16266_);
  not (_16269_, _16260_);
  or (_16270_, _16269_, _14727_);
  and (_16271_, _16270_, _16268_);
  and (_16272_, _16265_, _14735_);
  or (_40760_, _16272_, _16271_);
  or (_16273_, _16260_, \oc8051_golden_model_1.IRAM[12] [2]);
  and (_16274_, _16273_, _16266_);
  or (_16275_, _16269_, _14929_);
  and (_16276_, _16275_, _16274_);
  and (_16277_, _16265_, _14937_);
  or (_40761_, _16277_, _16276_);
  or (_16278_, _16260_, \oc8051_golden_model_1.IRAM[12] [3]);
  and (_16279_, _16278_, _16266_);
  or (_16280_, _16269_, _15131_);
  and (_16281_, _16280_, _16279_);
  and (_16282_, _16265_, _15139_);
  or (_40762_, _16282_, _16281_);
  or (_16283_, _16260_, \oc8051_golden_model_1.IRAM[12] [4]);
  and (_16284_, _16283_, _16266_);
  or (_16285_, _16269_, _15332_);
  and (_16286_, _16285_, _16284_);
  and (_16287_, _16265_, _15340_);
  or (_40764_, _16287_, _16286_);
  or (_16288_, _16260_, \oc8051_golden_model_1.IRAM[12] [5]);
  and (_16289_, _16288_, _16266_);
  or (_16290_, _16269_, _15535_);
  and (_16291_, _16290_, _16289_);
  and (_16292_, _16265_, _15543_);
  or (_40765_, _16292_, _16291_);
  or (_16293_, _16260_, \oc8051_golden_model_1.IRAM[12] [6]);
  and (_16294_, _16293_, _16266_);
  or (_16295_, _16269_, _15737_);
  and (_16296_, _16295_, _16294_);
  and (_16297_, _16265_, _15745_);
  or (_40766_, _16297_, _16296_);
  or (_16298_, _16260_, \oc8051_golden_model_1.IRAM[12] [7]);
  and (_16299_, _16298_, _16266_);
  or (_16300_, _16269_, _09465_);
  and (_16301_, _16300_, _16299_);
  and (_16302_, _16265_, _09490_);
  or (_40767_, _16302_, _16301_);
  and (_16303_, _15752_, _07861_);
  or (_16304_, _16303_, \oc8051_golden_model_1.IRAM[13] [0]);
  and (_16305_, _07874_, _07598_);
  not (_16306_, _16305_);
  and (_16307_, _16306_, _16304_);
  not (_16308_, _16303_);
  or (_16309_, _16308_, _14528_);
  and (_16310_, _16309_, _16307_);
  and (_16311_, _16305_, _14543_);
  or (_40771_, _16311_, _16310_);
  or (_16312_, _16303_, \oc8051_golden_model_1.IRAM[13] [1]);
  and (_16313_, _16312_, _16306_);
  or (_16314_, _16308_, _14727_);
  and (_16315_, _16314_, _16313_);
  and (_16316_, _16305_, _14735_);
  or (_40772_, _16316_, _16315_);
  or (_16317_, _16303_, \oc8051_golden_model_1.IRAM[13] [2]);
  and (_16318_, _16317_, _16306_);
  or (_16319_, _16308_, _14929_);
  and (_16320_, _16319_, _16318_);
  and (_16321_, _16305_, _14937_);
  or (_40773_, _16321_, _16320_);
  or (_16322_, _16303_, \oc8051_golden_model_1.IRAM[13] [3]);
  and (_16323_, _16322_, _16306_);
  or (_16324_, _16308_, _15131_);
  and (_16325_, _16324_, _16323_);
  and (_16326_, _16305_, _15139_);
  or (_40774_, _16326_, _16325_);
  or (_16327_, _16303_, \oc8051_golden_model_1.IRAM[13] [4]);
  and (_16328_, _16327_, _16306_);
  or (_16329_, _16308_, _15332_);
  and (_16330_, _16329_, _16328_);
  and (_16331_, _16305_, _15340_);
  or (_40776_, _16331_, _16330_);
  or (_16332_, _16303_, \oc8051_golden_model_1.IRAM[13] [5]);
  and (_16333_, _16332_, _16306_);
  or (_16334_, _16308_, _15535_);
  and (_16335_, _16334_, _16333_);
  and (_16336_, _16305_, _15543_);
  or (_40777_, _16336_, _16335_);
  or (_16337_, _16303_, \oc8051_golden_model_1.IRAM[13] [6]);
  and (_16338_, _16337_, _16306_);
  or (_16339_, _16308_, _15737_);
  and (_16340_, _16339_, _16338_);
  and (_16341_, _16305_, _15745_);
  or (_40778_, _16341_, _16340_);
  or (_16342_, _16303_, \oc8051_golden_model_1.IRAM[13] [7]);
  and (_16343_, _16342_, _16306_);
  or (_16344_, _16308_, _09465_);
  and (_16345_, _16344_, _16343_);
  and (_16346_, _16305_, _09490_);
  or (_40779_, _16346_, _16345_);
  and (_16347_, _15800_, _07861_);
  or (_16348_, _16347_, \oc8051_golden_model_1.IRAM[14] [0]);
  and (_16349_, _08668_, _07874_);
  not (_16350_, _16349_);
  and (_16351_, _16350_, _16348_);
  not (_16352_, _16347_);
  or (_16353_, _16352_, _14528_);
  and (_16354_, _16353_, _16351_);
  and (_16355_, _16349_, _14543_);
  or (_40783_, _16355_, _16354_);
  or (_16356_, _16347_, \oc8051_golden_model_1.IRAM[14] [1]);
  and (_16357_, _16356_, _16350_);
  or (_16358_, _16352_, _14727_);
  and (_16359_, _16358_, _16357_);
  and (_16360_, _16349_, _14735_);
  or (_40784_, _16360_, _16359_);
  not (_16361_, _08668_);
  or (_16362_, _16361_, _16257_);
  nor (_16363_, _16347_, _07764_);
  and (_16364_, _16347_, _14929_);
  or (_16365_, _16364_, _16363_);
  and (_16366_, _16365_, _16362_);
  and (_16367_, _16349_, _14937_);
  or (_40785_, _16367_, _16366_);
  or (_16368_, _16347_, \oc8051_golden_model_1.IRAM[14] [3]);
  and (_16369_, _16368_, _16350_);
  or (_16370_, _16352_, _15131_);
  and (_16371_, _16370_, _16369_);
  and (_16372_, _16349_, _15139_);
  or (_40787_, _16372_, _16371_);
  or (_16373_, _16347_, \oc8051_golden_model_1.IRAM[14] [4]);
  and (_16374_, _16373_, _16350_);
  or (_16375_, _16352_, _15332_);
  and (_16376_, _16375_, _16374_);
  and (_16377_, _16349_, _15340_);
  or (_40788_, _16377_, _16376_);
  or (_16378_, _16347_, \oc8051_golden_model_1.IRAM[14] [5]);
  and (_16379_, _16378_, _16350_);
  or (_16380_, _16352_, _15535_);
  and (_16381_, _16380_, _16379_);
  and (_16382_, _16349_, _15543_);
  or (_40789_, _16382_, _16381_);
  or (_16383_, _16347_, \oc8051_golden_model_1.IRAM[14] [6]);
  and (_16384_, _16383_, _16350_);
  or (_16385_, _16352_, _15737_);
  and (_16386_, _16385_, _16384_);
  and (_16387_, _16349_, _15745_);
  or (_40790_, _16387_, _16386_);
  or (_16388_, _16347_, \oc8051_golden_model_1.IRAM[14] [7]);
  and (_16389_, _16388_, _16350_);
  or (_16390_, _16352_, _09465_);
  and (_16391_, _16390_, _16389_);
  and (_16392_, _16349_, _09490_);
  or (_40791_, _16392_, _16391_);
  not (_16393_, _07295_);
  or (_16394_, _16257_, _16393_);
  or (_16395_, _14543_, _16394_);
  and (_16396_, _14528_, _07862_);
  or (_16397_, _07862_, _07119_);
  nand (_16398_, _16397_, _16394_);
  or (_16399_, _16398_, _16396_);
  and (_40795_, _16399_, _16395_);
  or (_16400_, _07862_, \oc8051_golden_model_1.IRAM[15] [1]);
  and (_16401_, _16400_, _07876_);
  or (_16402_, _14727_, _07878_);
  and (_16403_, _16402_, _16401_);
  and (_16404_, _14735_, _07875_);
  or (_40796_, _16404_, _16403_);
  nor (_16405_, _07862_, _07762_);
  and (_16406_, _14929_, _07862_);
  or (_16407_, _16406_, _16405_);
  and (_16408_, _16407_, _16394_);
  and (_16409_, _14937_, _07875_);
  or (_40797_, _16409_, _16408_);
  or (_16410_, _07862_, \oc8051_golden_model_1.IRAM[15] [3]);
  and (_16411_, _16410_, _07876_);
  or (_16412_, _15131_, _07878_);
  and (_16413_, _16412_, _16411_);
  and (_16414_, _15139_, _07875_);
  or (_40799_, _16414_, _16413_);
  or (_16415_, _15332_, _07878_);
  or (_16416_, _07862_, \oc8051_golden_model_1.IRAM[15] [4]);
  and (_16417_, _16416_, _07876_);
  and (_16418_, _16417_, _16415_);
  and (_16419_, _15340_, _07875_);
  or (_40800_, _16419_, _16418_);
  or (_16420_, _07862_, \oc8051_golden_model_1.IRAM[15] [5]);
  and (_16421_, _16420_, _07876_);
  or (_16422_, _15535_, _07878_);
  and (_16423_, _16422_, _16421_);
  and (_16424_, _15543_, _07875_);
  or (_40801_, _16424_, _16423_);
  or (_16425_, _15737_, _07878_);
  or (_16426_, _07862_, \oc8051_golden_model_1.IRAM[15] [6]);
  and (_16427_, _16426_, _07876_);
  and (_16428_, _16427_, _16425_);
  and (_16429_, _15745_, _07875_);
  or (_40802_, _16429_, _16428_);
  nor (_16430_, _01347_, _10106_);
  nand (_16431_, _11263_, _07942_);
  nor (_16432_, _07942_, _10106_);
  nor (_16433_, _16432_, _07234_);
  nand (_16434_, _16433_, _16431_);
  and (_16435_, _07942_, _08954_);
  or (_16436_, _16435_, _16432_);
  or (_16437_, _16436_, _06219_);
  and (_16438_, _07942_, _07133_);
  or (_16439_, _16438_, _16432_);
  or (_16440_, _16439_, _07215_);
  nor (_16441_, _08390_, _09498_);
  or (_16442_, _16441_, _16432_);
  or (_16443_, _16442_, _07151_);
  and (_16444_, _07942_, \oc8051_golden_model_1.ACC [0]);
  or (_16445_, _16444_, _16432_);
  and (_16446_, _16445_, _07141_);
  nor (_16447_, _07141_, _10106_);
  or (_16448_, _16447_, _06341_);
  or (_16449_, _16448_, _16446_);
  and (_16450_, _16449_, _06273_);
  and (_16451_, _16450_, _16443_);
  and (_16452_, _14382_, _08634_);
  nor (_16453_, _08634_, _10106_);
  or (_16454_, _16453_, _16452_);
  and (_16455_, _16454_, _06272_);
  or (_16456_, _16455_, _16451_);
  and (_16457_, _16456_, _07166_);
  and (_16458_, _16439_, _06461_);
  or (_16459_, _16458_, _06464_);
  or (_16460_, _16459_, _16457_);
  or (_16461_, _16445_, _06465_);
  and (_16462_, _16461_, _06269_);
  and (_16463_, _16462_, _16460_);
  and (_16464_, _16432_, _06268_);
  or (_16465_, _16464_, _06261_);
  or (_16466_, _16465_, _16463_);
  or (_16467_, _16442_, _06262_);
  and (_16468_, _16467_, _16466_);
  or (_16469_, _16468_, _09531_);
  nor (_16470_, _10052_, _10050_);
  nor (_16471_, _16470_, _10053_);
  or (_16472_, _16471_, _09537_);
  and (_16473_, _16472_, _06258_);
  and (_16474_, _16473_, _16469_);
  and (_16475_, _14413_, _08634_);
  or (_16476_, _16475_, _16453_);
  and (_16477_, _16476_, _06257_);
  or (_16478_, _16477_, _10080_);
  or (_16479_, _16478_, _16474_);
  and (_16480_, _16479_, _16440_);
  or (_16481_, _16480_, _07460_);
  and (_16482_, _09392_, _07942_);
  or (_16483_, _16432_, _07208_);
  or (_16484_, _16483_, _16482_);
  and (_16485_, _16484_, _16481_);
  or (_16486_, _16485_, _10094_);
  and (_16487_, _14467_, _07942_);
  or (_16488_, _16432_, _05982_);
  or (_16489_, _16488_, _16487_);
  and (_16490_, _16489_, _10100_);
  and (_16491_, _16490_, _16486_);
  nand (_16492_, _10439_, _06097_);
  or (_16493_, _10433_, _10408_);
  or (_16494_, _10439_, _16493_);
  and (_16495_, _16494_, _10093_);
  and (_16496_, _16495_, _16492_);
  or (_16497_, _16496_, _06218_);
  or (_16498_, _16497_, _16491_);
  and (_16499_, _16498_, _16437_);
  or (_16500_, _16499_, _06369_);
  and (_16501_, _14366_, _07942_);
  or (_16502_, _16501_, _16432_);
  or (_16503_, _16502_, _07237_);
  and (_16504_, _16503_, _07240_);
  and (_16505_, _16504_, _16500_);
  nor (_16506_, _12580_, _09498_);
  or (_16507_, _16506_, _16432_);
  and (_16508_, _16431_, _06536_);
  and (_16509_, _16508_, _16507_);
  or (_16510_, _16509_, _16505_);
  and (_16511_, _16510_, _07242_);
  nand (_16512_, _16436_, _06375_);
  nor (_16513_, _16512_, _16441_);
  or (_16514_, _16513_, _06545_);
  or (_16515_, _16514_, _16511_);
  and (_16516_, _16515_, _16434_);
  or (_16517_, _16516_, _06366_);
  and (_16518_, _14363_, _07942_);
  or (_16519_, _16432_, _09056_);
  or (_16520_, _16519_, _16518_);
  and (_16521_, _16520_, _09061_);
  and (_16522_, _16521_, _16517_);
  and (_16523_, _16507_, _06528_);
  or (_16524_, _16523_, _06568_);
  or (_16525_, _16524_, _16522_);
  or (_16526_, _16442_, _06926_);
  and (_16527_, _16526_, _16525_);
  or (_16528_, _16527_, _05927_);
  or (_16529_, _16432_, _05928_);
  and (_16530_, _16529_, _16528_);
  or (_16531_, _16530_, _06278_);
  or (_16532_, _16442_, _06279_);
  and (_16533_, _16532_, _01347_);
  and (_16534_, _16533_, _16531_);
  or (_16535_, _16534_, _16430_);
  and (_43153_, _16535_, _42618_);
  nor (_16536_, _01347_, _10101_);
  nor (_16537_, _07942_, _10101_);
  nor (_16538_, _11261_, _09498_);
  or (_16539_, _16538_, _16537_);
  or (_16540_, _16539_, _09061_);
  or (_16541_, _07942_, \oc8051_golden_model_1.B [1]);
  nand (_16542_, _07942_, _07038_);
  and (_16543_, _16542_, _06218_);
  and (_16544_, _16543_, _16541_);
  nor (_16545_, _08634_, _10101_);
  and (_16546_, _14560_, _08634_);
  or (_16547_, _16546_, _16545_);
  and (_16548_, _16547_, _06268_);
  nor (_16549_, _09498_, _07357_);
  or (_16550_, _16549_, _16537_);
  or (_16551_, _16550_, _07166_);
  and (_16552_, _14562_, _07942_);
  not (_16553_, _16552_);
  and (_16554_, _16553_, _16541_);
  or (_16555_, _16554_, _07151_);
  and (_16556_, _07942_, \oc8051_golden_model_1.ACC [1]);
  or (_16557_, _16556_, _16537_);
  and (_16558_, _16557_, _07141_);
  nor (_16559_, _07141_, _10101_);
  or (_16560_, _16559_, _06341_);
  or (_16561_, _16560_, _16558_);
  and (_16562_, _16561_, _06273_);
  and (_16563_, _16562_, _16555_);
  and (_16564_, _14557_, _08634_);
  or (_16565_, _16564_, _16545_);
  and (_16566_, _16565_, _06272_);
  or (_16567_, _16566_, _06461_);
  or (_16568_, _16567_, _16563_);
  and (_16569_, _16568_, _16551_);
  or (_16570_, _16569_, _06464_);
  or (_16571_, _16557_, _06465_);
  and (_16572_, _16571_, _06269_);
  and (_16573_, _16572_, _16570_);
  or (_16574_, _16573_, _16548_);
  and (_16575_, _16574_, _06262_);
  and (_16576_, _16564_, _14556_);
  or (_16577_, _16576_, _16545_);
  and (_16578_, _16577_, _06261_);
  or (_16579_, _16578_, _09531_);
  or (_16580_, _16579_, _16575_);
  nor (_16581_, _10055_, _09997_);
  nor (_16582_, _16581_, _10056_);
  or (_16583_, _16582_, _09537_);
  and (_16584_, _16583_, _06258_);
  and (_16585_, _16584_, _16580_);
  or (_16586_, _16545_, _14597_);
  and (_16587_, _16586_, _06257_);
  and (_16588_, _16587_, _16565_);
  or (_16589_, _16588_, _10080_);
  or (_16590_, _16589_, _16585_);
  or (_16591_, _16550_, _07215_);
  and (_16592_, _16591_, _16590_);
  or (_16593_, _16592_, _07460_);
  and (_16594_, _09451_, _07942_);
  or (_16595_, _16537_, _07208_);
  or (_16596_, _16595_, _16594_);
  and (_16597_, _16596_, _05982_);
  and (_16598_, _16597_, _16593_);
  or (_16599_, _14653_, _09498_);
  and (_16600_, _16541_, _10094_);
  and (_16601_, _16600_, _16599_);
  or (_16602_, _16601_, _10093_);
  or (_16603_, _16602_, _16598_);
  nor (_16604_, _10434_, _10432_);
  or (_16605_, _16604_, _10435_);
  nor (_16606_, _16605_, _10439_);
  and (_16607_, _10439_, _10405_);
  or (_16608_, _16607_, _16606_);
  or (_16609_, _16608_, _10100_);
  and (_16610_, _16609_, _06219_);
  and (_16611_, _16610_, _16603_);
  or (_16612_, _16611_, _16544_);
  and (_16613_, _16612_, _07237_);
  or (_16614_, _14668_, _09498_);
  and (_16615_, _16541_, _06369_);
  and (_16616_, _16615_, _16614_);
  or (_16617_, _16616_, _06536_);
  or (_16618_, _16617_, _16613_);
  and (_16619_, _11262_, _07942_);
  or (_16620_, _16619_, _16537_);
  or (_16621_, _16620_, _07240_);
  and (_16622_, _16621_, _07242_);
  and (_16623_, _16622_, _16618_);
  or (_16624_, _14666_, _09498_);
  and (_16625_, _16541_, _06375_);
  and (_16626_, _16625_, _16624_);
  or (_16627_, _16626_, _06545_);
  or (_16628_, _16627_, _16623_);
  and (_16629_, _16556_, _08341_);
  or (_16630_, _16537_, _07234_);
  or (_16631_, _16630_, _16629_);
  and (_16632_, _16631_, _09056_);
  and (_16633_, _16632_, _16628_);
  or (_16634_, _16542_, _08341_);
  and (_16635_, _16541_, _06366_);
  and (_16636_, _16635_, _16634_);
  or (_16637_, _16636_, _06528_);
  or (_16638_, _16637_, _16633_);
  and (_16639_, _16638_, _16540_);
  or (_16640_, _16639_, _06568_);
  or (_16641_, _16554_, _06926_);
  and (_16642_, _16641_, _05928_);
  and (_16643_, _16642_, _16640_);
  and (_16644_, _16547_, _05927_);
  or (_16645_, _16644_, _06278_);
  or (_16646_, _16645_, _16643_);
  or (_16647_, _16537_, _06279_);
  or (_16648_, _16647_, _16552_);
  and (_16649_, _16648_, _01347_);
  and (_16650_, _16649_, _16646_);
  or (_16651_, _16650_, _16536_);
  and (_43154_, _16651_, _42618_);
  nor (_16652_, _01347_, _10159_);
  nor (_16653_, _07942_, _10159_);
  and (_16654_, _07942_, _08973_);
  or (_16655_, _16654_, _16653_);
  or (_16656_, _16655_, _06219_);
  nor (_16657_, _09498_, _07776_);
  or (_16658_, _16657_, _16653_);
  or (_16659_, _16658_, _07215_);
  and (_16660_, _14774_, _08634_);
  and (_16661_, _16660_, _14789_);
  nor (_16662_, _08634_, _10159_);
  or (_16663_, _16662_, _06262_);
  or (_16664_, _16663_, _16661_);
  or (_16665_, _16658_, _07166_);
  and (_16666_, _14770_, _07942_);
  or (_16667_, _16666_, _16653_);
  or (_16668_, _16667_, _07151_);
  and (_16669_, _07942_, \oc8051_golden_model_1.ACC [2]);
  or (_16670_, _16669_, _16653_);
  and (_16671_, _16670_, _07141_);
  nor (_16672_, _07141_, _10159_);
  or (_16673_, _16672_, _06341_);
  or (_16674_, _16673_, _16671_);
  and (_16675_, _16674_, _06273_);
  and (_16676_, _16675_, _16668_);
  or (_16677_, _16662_, _16660_);
  and (_16678_, _16677_, _06272_);
  or (_16679_, _16678_, _06461_);
  or (_16680_, _16679_, _16676_);
  and (_16681_, _16680_, _16665_);
  or (_16682_, _16681_, _06464_);
  or (_16683_, _16670_, _06465_);
  and (_16684_, _16683_, _06269_);
  and (_16685_, _16684_, _16682_);
  and (_16686_, _14756_, _08634_);
  or (_16687_, _16686_, _16662_);
  and (_16688_, _16687_, _06268_);
  or (_16689_, _16688_, _06261_);
  or (_16690_, _16689_, _16685_);
  and (_16691_, _16690_, _16664_);
  or (_16692_, _16691_, _09531_);
  or (_16693_, _10057_, _09952_);
  and (_16694_, _16693_, _10058_);
  or (_16695_, _16694_, _09537_);
  and (_16696_, _16695_, _06258_);
  and (_16697_, _16696_, _16692_);
  and (_16698_, _14804_, _08634_);
  or (_16699_, _16698_, _16662_);
  and (_16700_, _16699_, _06257_);
  or (_16701_, _16700_, _10080_);
  or (_16702_, _16701_, _16697_);
  and (_16703_, _16702_, _16659_);
  or (_16704_, _16703_, _07460_);
  and (_16705_, _09450_, _07942_);
  or (_16706_, _16653_, _07208_);
  or (_16707_, _16706_, _16705_);
  and (_16708_, _16707_, _16704_);
  or (_16709_, _16708_, _10094_);
  and (_16710_, _14859_, _07942_);
  or (_16711_, _16653_, _05982_);
  or (_16712_, _16711_, _16710_);
  and (_16713_, _16712_, _10100_);
  and (_16714_, _16713_, _16709_);
  not (_16715_, _10439_);
  or (_16716_, _16715_, _10396_);
  nor (_16717_, _10435_, _10406_);
  not (_16718_, _16717_);
  and (_16719_, _16718_, _10399_);
  nor (_16720_, _16718_, _10399_);
  nor (_16721_, _16720_, _16719_);
  or (_16722_, _16721_, _10439_);
  and (_16723_, _16722_, _10093_);
  and (_16724_, _16723_, _16716_);
  or (_16725_, _16724_, _06218_);
  or (_16726_, _16725_, _16714_);
  and (_16727_, _16726_, _16656_);
  or (_16728_, _16727_, _06369_);
  and (_16729_, _14751_, _07942_);
  or (_16730_, _16729_, _16653_);
  or (_16731_, _16730_, _07237_);
  and (_16732_, _16731_, _07240_);
  and (_16733_, _16732_, _16728_);
  and (_16734_, _11259_, _07942_);
  or (_16735_, _16734_, _16653_);
  and (_16736_, _16735_, _06536_);
  or (_16737_, _16736_, _16733_);
  and (_16738_, _16737_, _07242_);
  or (_16739_, _16653_, _08440_);
  and (_16740_, _16655_, _06375_);
  and (_16741_, _16740_, _16739_);
  or (_16742_, _16741_, _16738_);
  and (_16743_, _16742_, _07234_);
  and (_16744_, _16670_, _06545_);
  and (_16745_, _16744_, _16739_);
  or (_16746_, _16745_, _06366_);
  or (_16747_, _16746_, _16743_);
  and (_16748_, _14748_, _07942_);
  or (_16749_, _16653_, _09056_);
  or (_16750_, _16749_, _16748_);
  and (_16751_, _16750_, _09061_);
  and (_16752_, _16751_, _16747_);
  nor (_16753_, _11258_, _09498_);
  or (_16754_, _16753_, _16653_);
  and (_16755_, _16754_, _06528_);
  or (_16756_, _16755_, _06568_);
  or (_16757_, _16756_, _16752_);
  or (_16758_, _16667_, _06926_);
  and (_16759_, _16758_, _05928_);
  and (_16760_, _16759_, _16757_);
  and (_16761_, _16687_, _05927_);
  or (_16762_, _16761_, _06278_);
  or (_16763_, _16762_, _16760_);
  and (_16764_, _14926_, _07942_);
  or (_16765_, _16653_, _06279_);
  or (_16766_, _16765_, _16764_);
  and (_16767_, _16766_, _01347_);
  and (_16768_, _16767_, _16763_);
  or (_16769_, _16768_, _16652_);
  and (_43155_, _16769_, _42618_);
  nor (_16770_, _01347_, _10145_);
  nor (_16771_, _07942_, _10145_);
  and (_16772_, _07942_, _08930_);
  or (_16773_, _16772_, _16771_);
  or (_16774_, _16773_, _06219_);
  and (_16775_, _15048_, _07942_);
  or (_16776_, _16775_, _16771_);
  and (_16777_, _16776_, _10094_);
  nor (_16778_, _08634_, _10145_);
  and (_16779_, _14950_, _08634_);
  or (_16780_, _16779_, _16778_);
  or (_16781_, _16778_, _14979_);
  and (_16782_, _16781_, _16780_);
  or (_16783_, _16782_, _06262_);
  and (_16784_, _14953_, _07942_);
  or (_16785_, _16784_, _16771_);
  or (_16786_, _16785_, _07151_);
  and (_16787_, _07942_, \oc8051_golden_model_1.ACC [3]);
  or (_16788_, _16787_, _16771_);
  and (_16789_, _16788_, _07141_);
  nor (_16790_, _07141_, _10145_);
  or (_16791_, _16790_, _06341_);
  or (_16792_, _16791_, _16789_);
  and (_16793_, _16792_, _06273_);
  and (_16794_, _16793_, _16786_);
  and (_16795_, _16780_, _06272_);
  or (_16796_, _16795_, _06461_);
  or (_16797_, _16796_, _16794_);
  nor (_16798_, _09498_, _07594_);
  or (_16799_, _16798_, _16771_);
  or (_16800_, _16799_, _07166_);
  and (_16801_, _16800_, _16797_);
  or (_16802_, _16801_, _06464_);
  or (_16803_, _16788_, _06465_);
  and (_16804_, _16803_, _06269_);
  and (_16805_, _16804_, _16802_);
  and (_16806_, _14948_, _08634_);
  or (_16807_, _16806_, _16778_);
  and (_16808_, _16807_, _06268_);
  or (_16809_, _16808_, _06261_);
  or (_16810_, _16809_, _16805_);
  and (_16811_, _16810_, _16783_);
  or (_16812_, _16811_, _09531_);
  nor (_16813_, _10060_, _09894_);
  nor (_16814_, _16813_, _10061_);
  or (_16815_, _16814_, _09537_);
  and (_16816_, _16815_, _06258_);
  and (_16817_, _16816_, _16812_);
  or (_16818_, _16778_, _14992_);
  and (_16819_, _16818_, _06257_);
  and (_16820_, _16819_, _16780_);
  or (_16821_, _16820_, _10080_);
  or (_16822_, _16821_, _16817_);
  or (_16823_, _16799_, _07215_);
  and (_16824_, _16823_, _16822_);
  or (_16825_, _16824_, _07460_);
  and (_16826_, _09449_, _07942_);
  or (_16827_, _16771_, _07208_);
  or (_16828_, _16827_, _16826_);
  and (_16829_, _16828_, _05982_);
  and (_16830_, _16829_, _16825_);
  or (_16831_, _16830_, _16777_);
  and (_16832_, _16831_, _10100_);
  nor (_16833_, _16719_, _10398_);
  nor (_16834_, _16833_, _10391_);
  and (_16835_, _16833_, _10391_);
  or (_16836_, _16835_, _16834_);
  or (_16837_, _16836_, _10439_);
  or (_16838_, _16715_, _10388_);
  and (_16839_, _16838_, _10093_);
  and (_16840_, _16839_, _16837_);
  or (_16841_, _16840_, _06218_);
  or (_16842_, _16841_, _16832_);
  and (_16843_, _16842_, _16774_);
  or (_16844_, _16843_, _06369_);
  and (_16845_, _14943_, _07942_);
  or (_16846_, _16845_, _16771_);
  or (_16847_, _16846_, _07237_);
  and (_16848_, _16847_, _07240_);
  and (_16849_, _16848_, _16844_);
  and (_16850_, _12577_, _07942_);
  or (_16851_, _16850_, _16771_);
  and (_16852_, _16851_, _06536_);
  or (_16853_, _16852_, _16849_);
  and (_16854_, _16853_, _07242_);
  or (_16855_, _16771_, _08292_);
  and (_16856_, _16773_, _06375_);
  and (_16857_, _16856_, _16855_);
  or (_16858_, _16857_, _16854_);
  and (_16859_, _16858_, _07234_);
  and (_16860_, _16788_, _06545_);
  and (_16861_, _16860_, _16855_);
  or (_16862_, _16861_, _06366_);
  or (_16863_, _16862_, _16859_);
  and (_16864_, _14940_, _07942_);
  or (_16865_, _16771_, _09056_);
  or (_16866_, _16865_, _16864_);
  and (_16867_, _16866_, _09061_);
  and (_16868_, _16867_, _16863_);
  nor (_16869_, _11256_, _09498_);
  or (_16870_, _16869_, _16771_);
  and (_16871_, _16870_, _06528_);
  or (_16872_, _16871_, _06568_);
  or (_16873_, _16872_, _16868_);
  or (_16874_, _16785_, _06926_);
  and (_16875_, _16874_, _05928_);
  and (_16876_, _16875_, _16873_);
  and (_16877_, _16807_, _05927_);
  or (_16878_, _16877_, _06278_);
  or (_16879_, _16878_, _16876_);
  and (_16880_, _15128_, _07942_);
  or (_16881_, _16771_, _06279_);
  or (_16882_, _16881_, _16880_);
  and (_16883_, _16882_, _01347_);
  and (_16884_, _16883_, _16879_);
  or (_16885_, _16884_, _16770_);
  and (_43156_, _16885_, _42618_);
  nor (_16886_, _01347_, _10241_);
  nor (_16887_, _07942_, _10241_);
  and (_16888_, _08959_, _07942_);
  or (_16889_, _16888_, _16887_);
  or (_16890_, _16889_, _06219_);
  and (_16891_, _15254_, _07942_);
  or (_16892_, _16891_, _16887_);
  and (_16893_, _16892_, _10094_);
  nor (_16894_, _08541_, _09498_);
  or (_16895_, _16894_, _16887_);
  or (_16896_, _16895_, _07215_);
  nor (_16897_, _08634_, _10241_);
  and (_16898_, _15176_, _08634_);
  or (_16899_, _16898_, _16897_);
  and (_16900_, _16899_, _06268_);
  and (_16901_, _15162_, _07942_);
  or (_16902_, _16901_, _16887_);
  or (_16903_, _16902_, _07151_);
  and (_16904_, _07942_, \oc8051_golden_model_1.ACC [4]);
  or (_16905_, _16904_, _16887_);
  and (_16906_, _16905_, _07141_);
  nor (_16907_, _07141_, _10241_);
  or (_16908_, _16907_, _06341_);
  or (_16909_, _16908_, _16906_);
  and (_16910_, _16909_, _06273_);
  and (_16911_, _16910_, _16903_);
  and (_16912_, _15166_, _08634_);
  or (_16913_, _16912_, _16897_);
  and (_16914_, _16913_, _06272_);
  or (_16915_, _16914_, _06461_);
  or (_16916_, _16915_, _16911_);
  or (_16917_, _16895_, _07166_);
  and (_16918_, _16917_, _16916_);
  or (_16919_, _16918_, _06464_);
  or (_16920_, _16905_, _06465_);
  and (_16921_, _16920_, _06269_);
  and (_16922_, _16921_, _16919_);
  or (_16923_, _16922_, _16900_);
  and (_16924_, _16923_, _06262_);
  or (_16925_, _16897_, _15183_);
  and (_16926_, _16925_, _06261_);
  and (_16927_, _16926_, _16913_);
  or (_16928_, _16927_, _09531_);
  or (_16929_, _16928_, _16924_);
  or (_16930_, _10064_, _10062_);
  and (_16931_, _16930_, _10065_);
  or (_16932_, _16931_, _09537_);
  and (_16933_, _16932_, _06258_);
  and (_16934_, _16933_, _16929_);
  and (_16935_, _15200_, _08634_);
  or (_16936_, _16935_, _16897_);
  and (_16937_, _16936_, _06257_);
  or (_16938_, _16937_, _10080_);
  or (_16939_, _16938_, _16934_);
  and (_16940_, _16939_, _16896_);
  or (_16941_, _16940_, _07460_);
  and (_16942_, _09448_, _07942_);
  or (_16943_, _16887_, _07208_);
  or (_16944_, _16943_, _16942_);
  and (_16945_, _16944_, _05982_);
  and (_16946_, _16945_, _16941_);
  or (_16947_, _16946_, _16893_);
  and (_16948_, _16947_, _10100_);
  or (_16949_, _16715_, _10380_);
  nor (_16950_, _16833_, _10390_);
  or (_16951_, _16950_, _10389_);
  nand (_16952_, _16951_, _10426_);
  or (_16953_, _16951_, _10426_);
  and (_16954_, _16953_, _16952_);
  or (_16955_, _16954_, _10439_);
  and (_16956_, _16955_, _10093_);
  and (_16957_, _16956_, _16949_);
  or (_16958_, _16957_, _06218_);
  or (_16959_, _16958_, _16948_);
  and (_16960_, _16959_, _16890_);
  or (_16961_, _16960_, _06369_);
  and (_16962_, _15269_, _07942_);
  or (_16963_, _16962_, _16887_);
  or (_16964_, _16963_, _07237_);
  and (_16965_, _16964_, _07240_);
  and (_16966_, _16965_, _16961_);
  and (_16967_, _11254_, _07942_);
  or (_16968_, _16967_, _16887_);
  and (_16969_, _16968_, _06536_);
  or (_16970_, _16969_, _16966_);
  and (_16971_, _16970_, _07242_);
  or (_16972_, _16887_, _08544_);
  and (_16973_, _16889_, _06375_);
  and (_16974_, _16973_, _16972_);
  or (_16975_, _16974_, _16971_);
  and (_16976_, _16975_, _07234_);
  and (_16977_, _16905_, _06545_);
  and (_16978_, _16977_, _16972_);
  or (_16979_, _16978_, _06366_);
  or (_16980_, _16979_, _16976_);
  and (_16981_, _15266_, _07942_);
  or (_16982_, _16887_, _09056_);
  or (_16983_, _16982_, _16981_);
  and (_16984_, _16983_, _09061_);
  and (_16985_, _16984_, _16980_);
  nor (_16986_, _11253_, _09498_);
  or (_16987_, _16986_, _16887_);
  and (_16988_, _16987_, _06528_);
  or (_16989_, _16988_, _06568_);
  or (_16990_, _16989_, _16985_);
  or (_16991_, _16902_, _06926_);
  and (_16992_, _16991_, _05928_);
  and (_16993_, _16992_, _16990_);
  and (_16994_, _16899_, _05927_);
  or (_16995_, _16994_, _06278_);
  or (_16996_, _16995_, _16993_);
  and (_16997_, _15329_, _07942_);
  or (_16998_, _16887_, _06279_);
  or (_16999_, _16998_, _16997_);
  and (_17000_, _16999_, _01347_);
  and (_17001_, _17000_, _16996_);
  or (_17002_, _17001_, _16886_);
  and (_43157_, _17002_, _42618_);
  nor (_17003_, _01347_, _10229_);
  nor (_17004_, _07942_, _10229_);
  and (_17005_, _15459_, _07942_);
  or (_17006_, _17005_, _17004_);
  and (_17007_, _17006_, _10094_);
  nor (_17008_, _08244_, _09498_);
  or (_17009_, _17008_, _17004_);
  or (_17010_, _17009_, _07215_);
  nor (_17011_, _08634_, _10229_);
  and (_17012_, _15355_, _08634_);
  or (_17013_, _17012_, _17011_);
  and (_17014_, _17013_, _06268_);
  and (_17015_, _15358_, _07942_);
  or (_17016_, _17015_, _17004_);
  or (_17017_, _17016_, _07151_);
  and (_17018_, _07942_, \oc8051_golden_model_1.ACC [5]);
  or (_17019_, _17018_, _17004_);
  and (_17020_, _17019_, _07141_);
  nor (_17021_, _07141_, _10229_);
  or (_17022_, _17021_, _06341_);
  or (_17023_, _17022_, _17020_);
  and (_17024_, _17023_, _06273_);
  and (_17025_, _17024_, _17017_);
  and (_17026_, _15372_, _08634_);
  or (_17027_, _17026_, _17011_);
  and (_17028_, _17027_, _06272_);
  or (_17029_, _17028_, _06461_);
  or (_17030_, _17029_, _17025_);
  or (_17031_, _17009_, _07166_);
  and (_17032_, _17031_, _17030_);
  or (_17033_, _17032_, _06464_);
  or (_17034_, _17019_, _06465_);
  and (_17035_, _17034_, _06269_);
  and (_17036_, _17035_, _17033_);
  or (_17037_, _17036_, _17014_);
  and (_17038_, _17037_, _06262_);
  or (_17039_, _17011_, _15387_);
  and (_17040_, _17039_, _06261_);
  and (_17041_, _17040_, _17027_);
  or (_17042_, _17041_, _09531_);
  or (_17043_, _17042_, _17038_);
  nor (_17044_, _10067_, _09757_);
  nor (_17045_, _17044_, _10068_);
  or (_17046_, _17045_, _09537_);
  and (_17047_, _17046_, _06258_);
  and (_17048_, _17047_, _17043_);
  or (_17049_, _17011_, _15403_);
  and (_17050_, _17049_, _06257_);
  and (_17051_, _17050_, _17027_);
  or (_17052_, _17051_, _10080_);
  or (_17053_, _17052_, _17048_);
  and (_17054_, _17053_, _17010_);
  or (_17055_, _17054_, _07460_);
  and (_17056_, _09447_, _07942_);
  or (_17057_, _17004_, _07208_);
  or (_17058_, _17057_, _17056_);
  and (_17059_, _17058_, _05982_);
  and (_17060_, _17059_, _17055_);
  or (_17061_, _17060_, _17007_);
  and (_17062_, _17061_, _10100_);
  or (_17063_, _16715_, _10372_);
  not (_17064_, _10417_);
  and (_17065_, _16952_, _17064_);
  nor (_17066_, _17065_, _10427_);
  and (_17067_, _17065_, _10427_);
  or (_17068_, _17067_, _17066_);
  or (_17069_, _17068_, _10439_);
  and (_17070_, _17069_, _10093_);
  and (_17071_, _17070_, _17063_);
  or (_17072_, _17071_, _06218_);
  or (_17073_, _17072_, _17062_);
  and (_17074_, _08946_, _07942_);
  or (_17075_, _17074_, _17004_);
  or (_17076_, _17075_, _06219_);
  and (_17077_, _17076_, _17073_);
  or (_17078_, _17077_, _06369_);
  and (_17079_, _15353_, _07942_);
  or (_17080_, _17079_, _17004_);
  or (_17081_, _17080_, _07237_);
  and (_17082_, _17081_, _07240_);
  and (_17083_, _17082_, _17078_);
  and (_17084_, _11250_, _07942_);
  or (_17085_, _17084_, _17004_);
  and (_17086_, _17085_, _06536_);
  or (_17087_, _17086_, _17083_);
  and (_17088_, _17087_, _07242_);
  or (_17089_, _17004_, _08247_);
  and (_17090_, _17075_, _06375_);
  and (_17091_, _17090_, _17089_);
  or (_17092_, _17091_, _17088_);
  and (_17093_, _17092_, _07234_);
  and (_17094_, _17019_, _06545_);
  and (_17095_, _17094_, _17089_);
  or (_17096_, _17095_, _06366_);
  or (_17097_, _17096_, _17093_);
  and (_17098_, _15350_, _07942_);
  or (_17099_, _17004_, _09056_);
  or (_17100_, _17099_, _17098_);
  and (_17101_, _17100_, _09061_);
  and (_17102_, _17101_, _17097_);
  nor (_17103_, _11249_, _09498_);
  or (_17104_, _17103_, _17004_);
  and (_17105_, _17104_, _06528_);
  or (_17106_, _17105_, _06568_);
  or (_17107_, _17106_, _17102_);
  or (_17108_, _17016_, _06926_);
  and (_17109_, _17108_, _05928_);
  and (_17110_, _17109_, _17107_);
  and (_17111_, _17013_, _05927_);
  or (_17112_, _17111_, _06278_);
  or (_17113_, _17112_, _17110_);
  and (_17114_, _15532_, _07942_);
  or (_17115_, _17004_, _06279_);
  or (_17116_, _17115_, _17114_);
  and (_17117_, _17116_, _01347_);
  and (_17118_, _17117_, _17113_);
  or (_17119_, _17118_, _17003_);
  and (_43159_, _17119_, _42618_);
  nor (_17120_, _01347_, _10357_);
  nor (_17121_, _07942_, _10357_);
  and (_17122_, _15664_, _07942_);
  or (_17123_, _17122_, _17121_);
  or (_17124_, _17123_, _06219_);
  and (_17125_, _15657_, _07942_);
  or (_17126_, _17125_, _17121_);
  and (_17127_, _17126_, _10094_);
  nor (_17128_, _08142_, _09498_);
  or (_17129_, _17128_, _17121_);
  or (_17130_, _17129_, _07215_);
  nor (_17131_, _08634_, _10357_);
  and (_17132_, _15551_, _08634_);
  or (_17133_, _17132_, _17131_);
  and (_17134_, _17133_, _06268_);
  and (_17135_, _15554_, _07942_);
  or (_17136_, _17135_, _17121_);
  or (_17137_, _17136_, _07151_);
  and (_17138_, _07942_, \oc8051_golden_model_1.ACC [6]);
  or (_17139_, _17138_, _17121_);
  and (_17140_, _17139_, _07141_);
  nor (_17141_, _07141_, _10357_);
  or (_17142_, _17141_, _06341_);
  or (_17143_, _17142_, _17140_);
  and (_17144_, _17143_, _06273_);
  and (_17145_, _17144_, _17137_);
  and (_17146_, _15570_, _08634_);
  or (_17147_, _17146_, _17131_);
  and (_17148_, _17147_, _06272_);
  or (_17149_, _17148_, _06461_);
  or (_17150_, _17149_, _17145_);
  or (_17151_, _17129_, _07166_);
  and (_17152_, _17151_, _17150_);
  or (_17153_, _17152_, _06464_);
  or (_17154_, _17139_, _06465_);
  and (_17155_, _17154_, _06269_);
  and (_17156_, _17155_, _17153_);
  or (_17157_, _17156_, _17134_);
  and (_17158_, _17157_, _06262_);
  or (_17159_, _17131_, _15585_);
  and (_17160_, _17159_, _06261_);
  and (_17161_, _17160_, _17147_);
  or (_17162_, _17161_, _09531_);
  or (_17163_, _17162_, _17158_);
  nor (_17164_, _10073_, _10069_);
  nor (_17165_, _17164_, _10074_);
  or (_17166_, _17165_, _09537_);
  and (_17167_, _17166_, _06258_);
  and (_17168_, _17167_, _17163_);
  and (_17169_, _15602_, _08634_);
  or (_17170_, _17169_, _17131_);
  and (_17171_, _17170_, _06257_);
  or (_17172_, _17171_, _10080_);
  or (_17173_, _17172_, _17168_);
  and (_17174_, _17173_, _17130_);
  or (_17175_, _17174_, _07460_);
  and (_17176_, _09446_, _07942_);
  or (_17177_, _17121_, _07208_);
  or (_17178_, _17177_, _17176_);
  and (_17179_, _17178_, _05982_);
  and (_17180_, _17179_, _17175_);
  or (_17181_, _17180_, _17127_);
  and (_17182_, _17181_, _10100_);
  nor (_17183_, _17065_, _10373_);
  or (_17184_, _17183_, _10374_);
  or (_17185_, _17184_, _10429_);
  nand (_17186_, _17184_, _10429_);
  and (_17187_, _17186_, _17185_);
  or (_17188_, _17187_, _10439_);
  nor (_17189_, _10439_, _10100_);
  and (_17190_, _10363_, _10093_);
  or (_17191_, _17190_, _17189_);
  and (_17192_, _17191_, _17188_);
  or (_17193_, _17192_, _06218_);
  or (_17194_, _17193_, _17182_);
  and (_17195_, _17194_, _17124_);
  or (_17196_, _17195_, _06369_);
  and (_17197_, _15549_, _07942_);
  or (_17198_, _17197_, _17121_);
  or (_17199_, _17198_, _07237_);
  and (_17200_, _17199_, _07240_);
  and (_17201_, _17200_, _17196_);
  and (_17202_, _11247_, _07942_);
  or (_17203_, _17202_, _17121_);
  and (_17204_, _17203_, _06536_);
  or (_17205_, _17204_, _17201_);
  and (_17206_, _17205_, _07242_);
  or (_17207_, _17121_, _08145_);
  and (_17208_, _17123_, _06375_);
  and (_17209_, _17208_, _17207_);
  or (_17210_, _17209_, _17206_);
  and (_17211_, _17210_, _07234_);
  and (_17212_, _17139_, _06545_);
  and (_17213_, _17212_, _17207_);
  or (_17214_, _17213_, _06366_);
  or (_17215_, _17214_, _17211_);
  and (_17216_, _15546_, _07942_);
  or (_17217_, _17121_, _09056_);
  or (_17218_, _17217_, _17216_);
  and (_17219_, _17218_, _09061_);
  and (_17220_, _17219_, _17215_);
  nor (_17221_, _11246_, _09498_);
  or (_17222_, _17221_, _17121_);
  and (_17223_, _17222_, _06528_);
  or (_17224_, _17223_, _06568_);
  or (_17225_, _17224_, _17220_);
  or (_17226_, _17136_, _06926_);
  and (_17227_, _17226_, _05928_);
  and (_17228_, _17227_, _17225_);
  and (_17229_, _17133_, _05927_);
  or (_17230_, _17229_, _06278_);
  or (_17231_, _17230_, _17228_);
  and (_17232_, _15734_, _07942_);
  or (_17233_, _17121_, _06279_);
  or (_17234_, _17233_, _17232_);
  and (_17235_, _17234_, _01347_);
  and (_17236_, _17235_, _17231_);
  or (_17237_, _17236_, _17120_);
  and (_43160_, _17237_, _42618_);
  nor (_17238_, _01347_, _06097_);
  nand (_17239_, _11284_, _08572_);
  nand (_17240_, _12581_, _06283_);
  and (_17241_, _17240_, _11321_);
  nor (_17242_, _07133_, \oc8051_golden_model_1.ACC [0]);
  nor (_17243_, _17242_, _11179_);
  and (_17244_, _11154_, _17243_);
  and (_17245_, _11156_, _17243_);
  nor (_17246_, _10634_, _06097_);
  or (_17247_, _17246_, _10635_);
  or (_17248_, _11069_, _17247_);
  nand (_17249_, _11021_, _12596_);
  nand (_17250_, _12581_, _06533_);
  and (_17251_, _17250_, _10955_);
  nand (_17252_, _06251_, _05974_);
  nor (_17253_, _07939_, _06097_);
  and (_17254_, _14467_, _07939_);
  or (_17255_, _17254_, _17253_);
  and (_17256_, _17255_, _10094_);
  and (_17257_, _07939_, _07133_);
  or (_17258_, _17257_, _17253_);
  or (_17259_, _17258_, _07215_);
  or (_17260_, _17247_, _10588_);
  or (_17261_, _10743_, _07133_);
  or (_17262_, _10755_, _07133_);
  nor (_17263_, _06781_, _06097_);
  and (_17264_, _06781_, _06097_);
  nor (_17265_, _17264_, _17263_);
  nand (_17266_, _17265_, _10755_);
  and (_17267_, _17266_, _10759_);
  and (_17268_, _17267_, _17262_);
  and (_17269_, _17268_, _07155_);
  or (_17270_, _17269_, _09392_);
  or (_17271_, _17268_, _10758_);
  and (_17272_, _17271_, _06015_);
  or (_17273_, _17272_, _07154_);
  and (_17274_, _17273_, _07151_);
  and (_17275_, _17274_, _17270_);
  nor (_17276_, _08390_, _10490_);
  or (_17277_, _17276_, _17253_);
  and (_17278_, _17277_, _06341_);
  or (_17279_, _17278_, _06272_);
  or (_17280_, _17279_, _17275_);
  and (_17281_, _14382_, _08636_);
  nor (_17282_, _08636_, _06097_);
  or (_17283_, _17282_, _06273_);
  or (_17284_, _17283_, _17281_);
  and (_17285_, _17284_, _07166_);
  and (_17286_, _17285_, _17280_);
  and (_17287_, _17258_, _06461_);
  or (_17288_, _17287_, _10744_);
  or (_17289_, _17288_, _17286_);
  and (_17290_, _17289_, _17261_);
  or (_17291_, _17290_, _07174_);
  or (_17292_, _09392_, _07175_);
  and (_17293_, _17292_, _06465_);
  and (_17294_, _17293_, _17291_);
  and (_17295_, _08390_, _06464_);
  or (_17296_, _17295_, _10811_);
  or (_17297_, _17296_, _17294_);
  nand (_17298_, _10811_, _10135_);
  and (_17299_, _17298_, _17297_);
  or (_17300_, _17299_, _06268_);
  or (_17301_, _17253_, _06269_);
  and (_17302_, _17301_, _06262_);
  and (_17303_, _17302_, _17300_);
  and (_17304_, _17277_, _06261_);
  or (_17305_, _17304_, _09531_);
  or (_17306_, _17305_, _17303_);
  nor (_17307_, _07211_, _05977_);
  nor (_17308_, _17307_, _14203_);
  not (_17309_, _14197_);
  or (_17310_, _17309_, _10729_);
  nor (_17311_, _17310_, _06705_);
  nand (_17312_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [0]);
  nand (_17313_, _17312_, _09531_);
  and (_17314_, _17313_, _17311_);
  and (_17315_, _17314_, _17308_);
  and (_17316_, _17315_, _17306_);
  nor (_17317_, _10709_, _06097_);
  or (_17318_, _17317_, _10710_);
  and (_17319_, _10737_, _17318_);
  or (_17320_, _17319_, _10656_);
  or (_17321_, _17320_, _17316_);
  and (_17322_, _17321_, _17260_);
  or (_17323_, _17322_, _06512_);
  nor (_17324_, _10881_, _06097_);
  or (_17325_, _17324_, _10882_);
  or (_17326_, _17325_, _06517_);
  and (_17327_, _17326_, _10517_);
  and (_17328_, _17327_, _17323_);
  nor (_17329_, _10564_, _06097_);
  or (_17330_, _17329_, _10565_);
  and (_17331_, _17330_, _10516_);
  or (_17332_, _17331_, _10515_);
  or (_17333_, _17332_, _17328_);
  nand (_17334_, _06251_, _10515_);
  and (_17335_, _17334_, _06258_);
  and (_17336_, _17335_, _17333_);
  and (_17337_, _14413_, _08636_);
  or (_17338_, _17337_, _17282_);
  and (_17340_, _17338_, _06257_);
  or (_17341_, _17340_, _10080_);
  or (_17342_, _17341_, _17336_);
  and (_17343_, _17342_, _17259_);
  or (_17344_, _17343_, _07460_);
  and (_17345_, _09392_, _07939_);
  or (_17346_, _17253_, _07208_);
  or (_17347_, _17346_, _17345_);
  and (_17348_, _17347_, _05982_);
  and (_17349_, _17348_, _17344_);
  or (_17351_, _17349_, _17256_);
  and (_17352_, _17351_, _10100_);
  or (_17353_, _17189_, _05974_);
  or (_17354_, _17353_, _17352_);
  and (_17355_, _17354_, _17252_);
  or (_17356_, _17355_, _06218_);
  and (_17357_, _07939_, _08954_);
  or (_17358_, _17357_, _17253_);
  or (_17359_, _17358_, _06219_);
  and (_17360_, _17359_, _10930_);
  and (_17362_, _17360_, _17356_);
  nor (_17363_, _10930_, _06251_);
  or (_17364_, _17363_, _10937_);
  or (_17365_, _17364_, _17362_);
  or (_17366_, _10940_, _17243_);
  and (_17367_, _10946_, _10508_);
  and (_17368_, _17367_, _17366_);
  and (_17369_, _17368_, _17365_);
  not (_17370_, _17367_);
  and (_17371_, _17370_, _17243_);
  or (_17373_, _17371_, _10501_);
  or (_17374_, _17373_, _17369_);
  not (_17375_, _10501_);
  nor (_17376_, _09392_, \oc8051_golden_model_1.ACC [0]);
  nor (_17377_, _11223_, _17376_);
  or (_17378_, _17377_, _17375_);
  and (_17379_, _17378_, _06885_);
  and (_17380_, _17379_, _17374_);
  and (_17381_, _17377_, _06884_);
  or (_17382_, _17381_, _06533_);
  or (_17384_, _17382_, _17380_);
  and (_17385_, _17384_, _17251_);
  and (_17386_, _10954_, _12597_);
  or (_17387_, _17386_, _06369_);
  or (_17388_, _17387_, _17385_);
  and (_17389_, _14366_, _07939_);
  or (_17390_, _17389_, _17253_);
  or (_17391_, _17390_, _07237_);
  and (_17392_, _17391_, _17388_);
  or (_17393_, _17392_, _06536_);
  or (_17395_, _17253_, _07240_);
  and (_17396_, _17395_, _10977_);
  and (_17397_, _17396_, _17393_);
  or (_17398_, _10985_, _11179_);
  and (_17399_, _17398_, _10987_);
  or (_17400_, _17399_, _17397_);
  not (_17401_, _10983_);
  not (_17402_, _10985_);
  or (_17403_, _17402_, _11179_);
  and (_17404_, _17403_, _17401_);
  and (_17405_, _17404_, _17400_);
  and (_17406_, _10983_, _11223_);
  or (_17407_, _17406_, _06542_);
  or (_17408_, _17407_, _17405_);
  or (_17409_, _11263_, _06543_);
  and (_17410_, _17409_, _10497_);
  and (_17411_, _17410_, _17408_);
  and (_17412_, _11302_, _10496_);
  or (_17413_, _17412_, _17411_);
  and (_17414_, _17413_, _07242_);
  nand (_17415_, _17358_, _06375_);
  nor (_17416_, _17415_, _17276_);
  or (_17417_, _17416_, _06711_);
  or (_17418_, _17417_, _17414_);
  nor (_17419_, _17242_, _06755_);
  or (_17420_, _17419_, _10998_);
  and (_17421_, _17420_, _17418_);
  and (_17422_, _06350_, _06527_);
  nor (_17423_, _17422_, _07040_);
  and (_17424_, _17423_, _12156_);
  not (_17425_, _17242_);
  nand (_17426_, _17425_, _06755_);
  nand (_17427_, _17426_, _17424_);
  or (_17428_, _17427_, _17421_);
  and (_17429_, _06337_, _06527_);
  not (_17430_, _17429_);
  or (_17431_, _17424_, _17425_);
  and (_17432_, _17431_, _17430_);
  and (_17433_, _17432_, _17428_);
  nor (_17434_, _17242_, _17430_);
  or (_17435_, _17434_, _11014_);
  or (_17436_, _17435_, _17433_);
  nand (_17437_, _11014_, _17376_);
  and (_17438_, _17437_, _06531_);
  and (_17439_, _17438_, _17436_);
  nand (_17440_, _11024_, _12580_);
  and (_17441_, _17440_, _11023_);
  or (_17442_, _17441_, _17439_);
  and (_17443_, _17442_, _17249_);
  or (_17444_, _17443_, _06366_);
  and (_17445_, _14363_, _07939_);
  or (_17446_, _17253_, _09056_);
  or (_17447_, _17446_, _17445_);
  and (_17448_, _17447_, _11037_);
  and (_17449_, _17448_, _17444_);
  and (_17450_, _14283_, _17318_);
  or (_17451_, _17450_, _11041_);
  or (_17452_, _17451_, _17449_);
  and (_17453_, _17452_, _17248_);
  or (_17454_, _17453_, _06540_);
  or (_17455_, _17325_, _06541_);
  and (_17456_, _17455_, _11127_);
  and (_17457_, _17456_, _17454_);
  and (_17458_, _11097_, _17330_);
  or (_17459_, _17458_, _11125_);
  or (_17460_, _17459_, _17457_);
  and (_17461_, _11125_, _10558_);
  or (_17462_, _17461_, _07045_);
  nor (_17463_, _17462_, _11155_);
  and (_17464_, _17463_, _17460_);
  nor (_17465_, _17464_, _17245_);
  nor (_17466_, _17465_, _11154_);
  or (_17467_, _17466_, _17244_);
  and (_17468_, _17467_, _11203_);
  and (_17469_, _11201_, _17377_);
  or (_17470_, _17469_, _06283_);
  or (_17471_, _17470_, _17468_);
  and (_17472_, _17471_, _17241_);
  and (_17473_, _11243_, _12597_);
  or (_17474_, _17473_, _11284_);
  or (_17475_, _17474_, _17472_);
  and (_17476_, _17475_, _17239_);
  or (_17477_, _17476_, _06568_);
  or (_17478_, _17277_, _06926_);
  and (_17479_, _17478_, _11331_);
  and (_17480_, _17479_, _17477_);
  nor (_17481_, _11335_, _06097_);
  nor (_17482_, _17481_, _13037_);
  or (_17483_, _17482_, _17480_);
  nand (_17484_, _11335_, _06042_);
  and (_17485_, _17484_, _05928_);
  and (_17486_, _17485_, _17483_);
  and (_17487_, _17253_, _05927_);
  or (_17488_, _17487_, _06278_);
  or (_17489_, _17488_, _17486_);
  or (_17490_, _17277_, _06279_);
  and (_17491_, _17490_, _11354_);
  and (_17492_, _17491_, _17489_);
  nor (_17493_, _11360_, _06097_);
  nor (_17494_, _17493_, _12141_);
  or (_17495_, _17494_, _17492_);
  nand (_17496_, _11360_, _06042_);
  and (_17497_, _17496_, _01347_);
  and (_17498_, _17497_, _17495_);
  or (_17499_, _17498_, _17238_);
  and (_43161_, _17499_, _42618_);
  nor (_17500_, _01347_, _06042_);
  or (_17501_, _11106_, _11105_);
  nor (_17502_, _11107_, _06541_);
  and (_17503_, _17502_, _17501_);
  and (_17504_, _06886_, _06364_);
  nor (_17505_, _11035_, _17504_);
  not (_17506_, _17423_);
  not (_17507_, _12157_);
  nand (_17508_, _17507_, _11177_);
  or (_17509_, _17401_, _11220_);
  not (_17510_, _06888_);
  and (_17511_, _06350_, _06535_);
  not (_17512_, _17511_);
  and (_17513_, _17512_, _10508_);
  nor (_17514_, _07939_, _06042_);
  nor (_17515_, _10490_, _07357_);
  or (_17516_, _17515_, _17514_);
  or (_17517_, _17516_, _07215_);
  nor (_17518_, _08636_, _06042_);
  and (_17519_, _14557_, _08636_);
  or (_17520_, _17519_, _17518_);
  or (_17521_, _17518_, _14556_);
  and (_17522_, _17521_, _06261_);
  and (_17523_, _17522_, _17520_);
  nand (_17524_, _10744_, _07357_);
  nand (_17525_, _10756_, _07357_);
  nor (_17526_, _06781_, _06042_);
  and (_17527_, _06781_, _06042_);
  nor (_17528_, _17527_, _17526_);
  nand (_17529_, _17528_, _10755_);
  and (_17530_, _17529_, _10759_);
  and (_17531_, _17530_, _17525_);
  or (_17532_, _17531_, _10758_);
  and (_17533_, _17532_, _06015_);
  or (_17534_, _17533_, _07154_);
  and (_17535_, _17531_, _07155_);
  or (_17536_, _17535_, _09451_);
  and (_17537_, _17536_, _17534_);
  or (_17538_, _17537_, _06341_);
  or (_17539_, _07939_, \oc8051_golden_model_1.ACC [1]);
  and (_17540_, _14562_, _07939_);
  not (_17541_, _17540_);
  and (_17542_, _17541_, _17539_);
  or (_17543_, _17542_, _07151_);
  and (_17544_, _17543_, _17538_);
  or (_17545_, _17544_, _10775_);
  nor (_17546_, _10779_, \oc8051_golden_model_1.PSW [6]);
  nor (_17547_, _17546_, \oc8051_golden_model_1.ACC [1]);
  and (_17548_, _17546_, \oc8051_golden_model_1.ACC [1]);
  nor (_17549_, _17548_, _17547_);
  nand (_17550_, _17549_, _10775_);
  and (_17551_, _17550_, _06466_);
  and (_17552_, _17551_, _17545_);
  and (_17553_, _17520_, _06272_);
  and (_17554_, _17516_, _06461_);
  or (_17555_, _17554_, _10744_);
  or (_17556_, _17555_, _17553_);
  or (_17557_, _17556_, _17552_);
  and (_17558_, _17557_, _17524_);
  or (_17559_, _17558_, _07174_);
  or (_17560_, _09451_, _07175_);
  and (_17561_, _17560_, _06465_);
  and (_17562_, _17561_, _17559_);
  nor (_17563_, _08340_, _06465_);
  or (_17564_, _17563_, _10811_);
  or (_17565_, _17564_, _17562_);
  nand (_17566_, _10811_, _10170_);
  and (_17567_, _17566_, _17565_);
  or (_17568_, _17567_, _06268_);
  and (_17569_, _14560_, _08636_);
  or (_17570_, _17569_, _17518_);
  or (_17571_, _17570_, _06269_);
  and (_17572_, _17571_, _06262_);
  and (_17573_, _17572_, _17568_);
  or (_17574_, _17573_, _17523_);
  and (_17575_, _17574_, _09537_);
  nor (_17576_, _10031_, _10030_);
  nor (_17577_, _17576_, _10032_);
  nand (_17578_, _17577_, _09531_);
  nand (_17579_, _17578_, _10735_);
  or (_17580_, _17579_, _17575_);
  nor (_17581_, _10657_, _06097_);
  or (_17582_, _17581_, _10708_);
  nor (_17583_, _17582_, _11178_);
  and (_17584_, _17582_, _11178_);
  or (_17585_, _17584_, _10735_);
  or (_17586_, _17585_, _17583_);
  and (_17587_, _17586_, _10588_);
  and (_17588_, _17587_, _17580_);
  not (_17589_, _11222_);
  nor (_17590_, _10589_, _06097_);
  or (_17591_, _17590_, _10633_);
  nand (_17592_, _17591_, _17589_);
  or (_17593_, _17591_, _17589_);
  and (_17594_, _17593_, _10656_);
  and (_17595_, _17594_, _17592_);
  or (_17596_, _17595_, _06512_);
  or (_17597_, _17596_, _17588_);
  nor (_17598_, _10834_, _06097_);
  or (_17599_, _17598_, _10880_);
  nor (_17600_, _17599_, _11262_);
  and (_17601_, _17599_, _11262_);
  or (_17602_, _17601_, _06517_);
  or (_17603_, _17602_, _17600_);
  and (_17604_, _17603_, _10517_);
  and (_17605_, _17604_, _17597_);
  nor (_17606_, _06251_, \oc8051_golden_model_1.ACC [0]);
  not (_17607_, _17606_);
  and (_17608_, _11305_, _17607_);
  nor (_17609_, _11305_, _17607_);
  nor (_17610_, _17609_, _17608_);
  or (_17611_, _12597_, _10558_);
  and (_17612_, _17611_, _17610_);
  and (_17613_, _12598_, \oc8051_golden_model_1.PSW [7]);
  or (_17614_, _17613_, _17612_);
  and (_17615_, _17614_, _10516_);
  or (_17616_, _17615_, _10515_);
  or (_17617_, _17616_, _17605_);
  nand (_17618_, _07004_, _10515_);
  and (_17619_, _17618_, _06258_);
  and (_17620_, _17619_, _17617_);
  or (_17621_, _17518_, _14597_);
  and (_17622_, _17621_, _06257_);
  and (_17623_, _17622_, _17520_);
  or (_17624_, _17623_, _10080_);
  or (_17625_, _17624_, _17620_);
  and (_17626_, _17625_, _17517_);
  or (_17627_, _17626_, _07460_);
  and (_17628_, _09451_, _07939_);
  or (_17629_, _17514_, _07208_);
  or (_17630_, _17629_, _17628_);
  and (_17631_, _17630_, _05982_);
  and (_17632_, _17631_, _17627_);
  or (_17633_, _14653_, _10490_);
  and (_17634_, _17539_, _10094_);
  and (_17635_, _17634_, _17633_);
  or (_17636_, _17635_, _10093_);
  or (_17637_, _17636_, _17632_);
  nand (_17638_, _10350_, _10093_);
  and (_17639_, _17638_, _17637_);
  or (_17640_, _17639_, _05974_);
  nand (_17641_, _07004_, _05974_);
  and (_17642_, _17641_, _06219_);
  and (_17643_, _17642_, _17640_);
  nand (_17644_, _07939_, _07038_);
  and (_17645_, _17539_, _06218_);
  and (_17646_, _17645_, _17644_);
  or (_17647_, _17646_, _10929_);
  or (_17648_, _17647_, _17643_);
  nand (_17649_, _10929_, _07004_);
  and (_17650_, _17649_, _10940_);
  and (_17651_, _17650_, _17648_);
  and (_17652_, _10937_, _11178_);
  or (_17653_, _17652_, _17651_);
  and (_17654_, _17653_, _17513_);
  not (_17655_, _17513_);
  and (_17656_, _17655_, _11178_);
  or (_17657_, _17656_, _17654_);
  and (_17658_, _17657_, _17510_);
  and (_17659_, _11178_, _06888_);
  or (_17660_, _17659_, _10948_);
  or (_17661_, _17660_, _17658_);
  or (_17662_, _11222_, _10502_);
  and (_17663_, _17662_, _17661_);
  or (_17664_, _17663_, _06533_);
  or (_17665_, _11262_, _06534_);
  and (_17666_, _17665_, _10955_);
  and (_17667_, _17666_, _17664_);
  nor (_17668_, _10955_, _11305_);
  or (_17669_, _17668_, _17667_);
  and (_17670_, _17669_, _07237_);
  or (_17671_, _14668_, _10490_);
  and (_17672_, _17539_, _06369_);
  and (_17673_, _17672_, _17671_);
  or (_17674_, _17673_, _06536_);
  or (_17675_, _17674_, _17670_);
  or (_17676_, _17514_, _07240_);
  and (_17677_, _17676_, _10986_);
  and (_17678_, _17677_, _17675_);
  and (_17679_, _10987_, _11176_);
  or (_17680_, _17679_, _10983_);
  or (_17681_, _17680_, _17678_);
  and (_17682_, _17681_, _17509_);
  or (_17683_, _17682_, _06542_);
  or (_17684_, _11260_, _06543_);
  and (_17685_, _17684_, _10497_);
  and (_17686_, _17685_, _17683_);
  and (_17687_, _11301_, _10496_);
  or (_17688_, _17687_, _17686_);
  and (_17689_, _17688_, _07242_);
  or (_17690_, _14666_, _10490_);
  and (_17691_, _17539_, _06375_);
  and (_17692_, _17691_, _17690_);
  or (_17693_, _17692_, _17507_);
  or (_17694_, _17693_, _17689_);
  and (_17695_, _17694_, _17508_);
  or (_17696_, _17695_, _17506_);
  nand (_17697_, _17506_, _11177_);
  and (_17698_, _17697_, _17430_);
  and (_17699_, _17698_, _17696_);
  nor (_17700_, _11177_, _17430_);
  or (_17701_, _17700_, _11014_);
  or (_17702_, _17701_, _17699_);
  nand (_17703_, _11014_, _11221_);
  and (_17704_, _17703_, _06531_);
  and (_17705_, _17704_, _17702_);
  nand (_17706_, _11024_, _11261_);
  and (_17707_, _17706_, _11023_);
  or (_17708_, _17707_, _17705_);
  and (_17709_, _11021_, _06042_);
  nand (_17710_, _17709_, _07004_);
  and (_17711_, _17710_, _09056_);
  and (_17712_, _17711_, _17708_);
  or (_17713_, _17644_, _08341_);
  and (_17714_, _17539_, _06366_);
  and (_17715_, _17714_, _17713_);
  or (_17716_, _17715_, _17712_);
  and (_17717_, _17716_, _17505_);
  nor (_17718_, _11050_, _11049_);
  nor (_17719_, _17718_, _11051_);
  and (_17720_, _17719_, _14283_);
  or (_17721_, _17720_, _17717_);
  not (_17722_, _11040_);
  and (_17723_, _07209_, _06364_);
  not (_17724_, _17723_);
  or (_17725_, _17719_, _17724_);
  and (_17726_, _17725_, _17722_);
  and (_17727_, _17726_, _17721_);
  nor (_17728_, _11078_, _11077_);
  nor (_17729_, _17728_, _11079_);
  and (_17730_, _17729_, _11040_);
  or (_17731_, _17730_, _11039_);
  or (_17732_, _17731_, _17727_);
  not (_17733_, _11039_);
  or (_17734_, _17729_, _17733_);
  and (_17735_, _17734_, _06541_);
  and (_17736_, _17735_, _17732_);
  or (_17737_, _17736_, _17503_);
  and (_17738_, _17737_, _11127_);
  or (_17739_, _11134_, _10568_);
  nor (_17740_, _11135_, _11127_);
  and (_17741_, _17740_, _17739_);
  or (_17742_, _17741_, _11125_);
  or (_17743_, _17742_, _17738_);
  nand (_17744_, _11125_, _06097_);
  and (_17745_, _17744_, _11157_);
  and (_17746_, _17745_, _17743_);
  or (_17747_, _11179_, _11178_);
  nor (_17748_, _11180_, _11157_);
  and (_17749_, _17748_, _17747_);
  or (_17750_, _17749_, _11201_);
  or (_17751_, _17750_, _17746_);
  nor (_17752_, _11223_, _11222_);
  nor (_17753_, _17752_, _11224_);
  or (_17754_, _17753_, _11203_);
  and (_17755_, _17754_, _06285_);
  and (_17756_, _17755_, _17751_);
  nor (_17757_, _11263_, _11262_);
  nor (_17758_, _17757_, _11264_);
  and (_17759_, _17758_, _06283_);
  or (_17760_, _17759_, _11243_);
  or (_17761_, _17760_, _17756_);
  nor (_17762_, _11306_, _11302_);
  nor (_17763_, _17762_, _11307_);
  or (_17764_, _17763_, _11321_);
  and (_17765_, _17764_, _11285_);
  and (_17766_, _17765_, _17761_);
  and (_17767_, _11284_, \oc8051_golden_model_1.ACC [0]);
  or (_17768_, _17767_, _06568_);
  or (_17769_, _17768_, _17766_);
  or (_17770_, _17542_, _06926_);
  and (_17771_, _17770_, _11331_);
  and (_17772_, _17771_, _17769_);
  nor (_17773_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.ACC [0]);
  nor (_17774_, _11361_, _17773_);
  nor (_17775_, _17774_, _11331_);
  or (_17776_, _17775_, _11335_);
  or (_17777_, _17776_, _17772_);
  nand (_17778_, _11335_, _10213_);
  and (_17779_, _17778_, _05928_);
  and (_17780_, _17779_, _17777_);
  and (_17781_, _17570_, _05927_);
  or (_17782_, _17781_, _06278_);
  or (_17783_, _17782_, _17780_);
  or (_17784_, _17540_, _17514_);
  or (_17785_, _17784_, _06279_);
  and (_17786_, _17785_, _11354_);
  and (_17787_, _17786_, _17783_);
  and (_17788_, _17774_, _11353_);
  or (_17789_, _17788_, _11360_);
  or (_17790_, _17789_, _17787_);
  nand (_17791_, _11360_, _10213_);
  and (_17792_, _17791_, _01347_);
  and (_17793_, _17792_, _17790_);
  or (_17794_, _17793_, _17500_);
  and (_43163_, _17794_, _42618_);
  nor (_17795_, _01347_, _10213_);
  nand (_17796_, _11284_, _06042_);
  or (_17797_, _11266_, _11259_);
  nor (_17798_, _11267_, _06285_);
  and (_17799_, _17798_, _17797_);
  not (_17800_, _11200_);
  nor (_17801_, _11226_, _11219_);
  nor (_17802_, _17801_, _11227_);
  or (_17803_, _17802_, _17800_);
  and (_17804_, _11136_, _10556_);
  nor (_17805_, _17804_, _11137_);
  or (_17806_, _17805_, _11127_);
  nand (_17807_, _11014_, _11218_);
  or (_17808_, _11219_, _10502_);
  nand (_17809_, _06656_, _05974_);
  nor (_17810_, _07939_, _10213_);
  nor (_17811_, _10490_, _07776_);
  or (_17812_, _17811_, _17810_);
  or (_17813_, _17812_, _07215_);
  nand (_17814_, _10744_, _07776_);
  nor (_17815_, _10758_, _07154_);
  or (_17816_, _17815_, _09450_);
  nor (_17817_, _10755_, _07776_);
  or (_17818_, _06781_, \oc8051_golden_model_1.ACC [2]);
  nand (_17819_, _06781_, \oc8051_golden_model_1.ACC [2]);
  and (_17820_, _17819_, _17818_);
  and (_17821_, _17820_, _10755_);
  or (_17822_, _17821_, _10758_);
  or (_17823_, _17822_, _17817_);
  and (_17824_, _17823_, _06015_);
  or (_17825_, _17824_, _07154_);
  and (_17826_, _17825_, _17816_);
  or (_17827_, _17826_, _06341_);
  and (_17828_, _14770_, _07939_);
  or (_17829_, _17828_, _17810_);
  or (_17830_, _17829_, _07151_);
  and (_17831_, _17830_, _17827_);
  or (_17832_, _17831_, _10775_);
  nor (_17833_, _17547_, _10213_);
  and (_17834_, _10778_, \oc8051_golden_model_1.PSW [6]);
  nor (_17835_, _17834_, _17833_);
  nand (_17836_, _17835_, _10775_);
  and (_17837_, _17836_, _06466_);
  and (_17838_, _17837_, _17832_);
  nor (_17839_, _08636_, _10213_);
  and (_17840_, _14774_, _08636_);
  or (_17841_, _17840_, _17839_);
  and (_17842_, _17841_, _06272_);
  and (_17843_, _17812_, _06461_);
  or (_17844_, _17843_, _10744_);
  or (_17845_, _17844_, _17842_);
  or (_17846_, _17845_, _17838_);
  and (_17847_, _17846_, _17814_);
  or (_17848_, _17847_, _07174_);
  or (_17849_, _09450_, _07175_);
  and (_17850_, _17849_, _06465_);
  and (_17851_, _17850_, _17848_);
  nor (_17852_, _08439_, _06465_);
  or (_17853_, _17852_, _10811_);
  or (_17854_, _17853_, _17851_);
  nand (_17855_, _10811_, _10116_);
  and (_17856_, _17855_, _17854_);
  or (_17857_, _17856_, _06268_);
  and (_17858_, _14756_, _08636_);
  or (_17859_, _17858_, _17839_);
  or (_17860_, _17859_, _06269_);
  and (_17861_, _17860_, _06262_);
  and (_17862_, _17861_, _17857_);
  or (_17863_, _17839_, _14789_);
  and (_17864_, _17841_, _06261_);
  and (_17865_, _17864_, _17863_);
  or (_17866_, _17865_, _09531_);
  or (_17867_, _17866_, _17862_);
  nor (_17868_, _10034_, _10032_);
  or (_17869_, _17868_, _10035_);
  nand (_17870_, _17869_, _09531_);
  and (_17871_, _17870_, _10735_);
  and (_17872_, _17871_, _17867_);
  and (_17873_, _07357_, \oc8051_golden_model_1.ACC [1]);
  and (_17874_, _07133_, _06097_);
  nor (_17875_, _17874_, _11178_);
  nor (_17876_, _17875_, _17873_);
  nor (_17877_, _11175_, _17876_);
  and (_17878_, _11175_, _17876_);
  nor (_17879_, _17878_, _17877_);
  nor (_17880_, _17243_, _11178_);
  and (_17881_, _17880_, \oc8051_golden_model_1.PSW [7]);
  or (_17882_, _17881_, _17879_);
  nand (_17883_, _17881_, _17879_);
  and (_17884_, _17883_, _10737_);
  and (_17885_, _17884_, _17882_);
  or (_17886_, _17885_, _17872_);
  and (_17887_, _17886_, _10588_);
  and (_17888_, _09347_, \oc8051_golden_model_1.ACC [1]);
  and (_17889_, _09392_, _06097_);
  nor (_17890_, _17889_, _11222_);
  nor (_17891_, _17890_, _17888_);
  nor (_17892_, _11219_, _17891_);
  and (_17893_, _11219_, _17891_);
  nor (_17894_, _17893_, _17892_);
  nor (_17895_, _17377_, _11222_);
  not (_17896_, _17895_);
  or (_17897_, _17896_, _17894_);
  and (_17898_, _17897_, \oc8051_golden_model_1.PSW [7]);
  nor (_17899_, _17894_, \oc8051_golden_model_1.PSW [7]);
  nor (_17900_, _17899_, _17898_);
  and (_17901_, _17896_, _17894_);
  or (_17902_, _17901_, _17900_);
  and (_17903_, _17902_, _10656_);
  or (_17904_, _17903_, _12644_);
  or (_17905_, _17904_, _17887_);
  and (_17906_, _08340_, \oc8051_golden_model_1.ACC [1]);
  and (_17907_, _08390_, _06097_);
  nor (_17908_, _14144_, _17907_);
  nor (_17909_, _17908_, _17906_);
  nor (_17910_, _11259_, _17909_);
  and (_17911_, _11259_, _17909_);
  nor (_17912_, _17911_, _17910_);
  and (_17913_, _12582_, \oc8051_golden_model_1.PSW [7]);
  nand (_17914_, _17913_, _17912_);
  or (_17915_, _17913_, _17912_);
  and (_17916_, _17915_, _17914_);
  or (_17917_, _17916_, _06517_);
  nor (_17918_, _17608_, _11303_);
  nor (_17919_, _11300_, _17918_);
  and (_17920_, _11300_, _17918_);
  nor (_17921_, _17920_, _17919_);
  not (_17922_, _17613_);
  nor (_17923_, _17922_, _17921_);
  and (_17924_, _17922_, _17921_);
  or (_17925_, _17924_, _10517_);
  or (_17926_, _17925_, _17923_);
  and (_17927_, _17926_, _17917_);
  and (_17928_, _17927_, _17905_);
  or (_17929_, _17928_, _10515_);
  nand (_17930_, _06656_, _10515_);
  and (_17931_, _17930_, _06258_);
  and (_17932_, _17931_, _17929_);
  and (_17933_, _14804_, _08636_);
  or (_17934_, _17933_, _17839_);
  and (_17935_, _17934_, _06257_);
  or (_17936_, _17935_, _10080_);
  or (_17937_, _17936_, _17932_);
  and (_17938_, _17937_, _17813_);
  or (_17939_, _17938_, _07460_);
  and (_17940_, _09450_, _07939_);
  or (_17941_, _17810_, _07208_);
  or (_17942_, _17941_, _17940_);
  and (_17943_, _17942_, _05982_);
  and (_17944_, _17943_, _17939_);
  and (_17945_, _14859_, _07939_);
  or (_17946_, _17945_, _17810_);
  and (_17947_, _17946_, _10094_);
  or (_17948_, _17947_, _10093_);
  or (_17949_, _17948_, _17944_);
  or (_17950_, _10286_, _10100_);
  and (_17951_, _17950_, _17949_);
  or (_17952_, _17951_, _05974_);
  and (_17953_, _17952_, _17809_);
  or (_17954_, _17953_, _06218_);
  and (_17955_, _07939_, _08973_);
  or (_17956_, _17955_, _17810_);
  or (_17957_, _17956_, _06219_);
  and (_17958_, _17957_, _10930_);
  and (_17959_, _17958_, _17954_);
  nor (_17960_, _10930_, _06656_);
  or (_17961_, _17960_, _17959_);
  nor (_17962_, _10937_, _06703_);
  and (_17964_, _17962_, _17961_);
  not (_17965_, _17962_);
  and (_17966_, _17965_, _11175_);
  or (_17967_, _17966_, _10506_);
  or (_17968_, _17967_, _17964_);
  not (_17969_, _10506_);
  or (_17970_, _11175_, _17969_);
  and (_17971_, _10732_, _06535_);
  not (_17972_, _17971_);
  and (_17973_, _17972_, _17970_);
  and (_17974_, _17973_, _17968_);
  and (_17975_, _17971_, _11175_);
  or (_17976_, _17975_, _10948_);
  or (_17977_, _17976_, _17974_);
  and (_17978_, _17977_, _17808_);
  or (_17979_, _17978_, _06533_);
  or (_17980_, _11259_, _06534_);
  and (_17981_, _17980_, _10955_);
  and (_17982_, _17981_, _17979_);
  and (_17983_, _10954_, _11300_);
  or (_17984_, _17983_, _06369_);
  or (_17985_, _17984_, _17982_);
  and (_17986_, _14751_, _07939_);
  or (_17987_, _17986_, _17810_);
  or (_17988_, _17987_, _07237_);
  and (_17989_, _17988_, _17985_);
  or (_17990_, _17989_, _06536_);
  or (_17991_, _17810_, _07240_);
  and (_17992_, _17991_, _10977_);
  and (_17993_, _17992_, _17990_);
  or (_17994_, _10985_, _11173_);
  and (_17995_, _17994_, _10987_);
  or (_17996_, _17995_, _17993_);
  or (_17997_, _17402_, _11173_);
  and (_17998_, _17997_, _17401_);
  and (_17999_, _17998_, _17996_);
  and (_18000_, _10983_, _11217_);
  or (_18001_, _18000_, _06542_);
  or (_18002_, _18001_, _17999_);
  or (_18003_, _11257_, _06543_);
  and (_18004_, _18003_, _10497_);
  and (_18005_, _18004_, _18002_);
  and (_18006_, _11298_, _10496_);
  or (_18007_, _18006_, _18005_);
  and (_18008_, _18007_, _07242_);
  nand (_18009_, _17956_, _06375_);
  nor (_18010_, _18009_, _11258_);
  or (_18011_, _18010_, _06711_);
  or (_18012_, _18011_, _18008_);
  nor (_18013_, _07042_, _06755_);
  nand (_18014_, _11174_, _06711_);
  and (_18015_, _18014_, _18013_);
  and (_18016_, _18015_, _18012_);
  nor (_18017_, _18013_, _11174_);
  or (_18018_, _18017_, _17506_);
  or (_18019_, _18018_, _18016_);
  nand (_18020_, _17506_, _11174_);
  and (_18021_, _18020_, _17430_);
  and (_18022_, _18021_, _18019_);
  nor (_18023_, _11174_, _17430_);
  or (_18024_, _18023_, _11014_);
  or (_18025_, _18024_, _18022_);
  and (_18026_, _18025_, _17807_);
  or (_18027_, _18026_, _06530_);
  nand (_18028_, _11258_, _06530_);
  and (_18029_, _18028_, _11024_);
  and (_18030_, _18029_, _18027_);
  nor (_18031_, _11024_, _11299_);
  or (_18032_, _18031_, _06366_);
  or (_18033_, _18032_, _18030_);
  and (_18034_, _14748_, _07939_);
  or (_18035_, _17810_, _09056_);
  or (_18036_, _18035_, _18034_);
  and (_18037_, _18036_, _11037_);
  and (_18038_, _18037_, _18033_);
  and (_18039_, _11052_, _10701_);
  nor (_18040_, _18039_, _11053_);
  and (_18041_, _18040_, _14283_);
  or (_18042_, _18041_, _11041_);
  or (_18043_, _18042_, _18038_);
  and (_18044_, _11080_, _10627_);
  nor (_18045_, _18044_, _11081_);
  or (_18046_, _18045_, _11069_);
  and (_18047_, _18046_, _06541_);
  and (_18048_, _18047_, _18043_);
  nand (_18049_, _11108_, _10874_);
  nor (_18050_, _11109_, _06541_);
  and (_18051_, _18050_, _18049_);
  or (_18052_, _18051_, _11097_);
  or (_18053_, _18052_, _18048_);
  and (_18054_, _18053_, _17806_);
  or (_18055_, _18054_, _11125_);
  nand (_18056_, _11125_, _06042_);
  and (_18057_, _18056_, _11157_);
  and (_18058_, _18057_, _18055_);
  not (_18059_, _11157_);
  nor (_18060_, _11182_, _11175_);
  nor (_18061_, _18060_, _11183_);
  and (_18062_, _18061_, _18059_);
  or (_18063_, _18062_, _11200_);
  or (_18064_, _18063_, _18058_);
  and (_18065_, _18064_, _17803_);
  or (_18066_, _18065_, _11199_);
  not (_18067_, _11199_);
  or (_18068_, _17802_, _18067_);
  and (_18069_, _18068_, _06285_);
  and (_18070_, _18069_, _18066_);
  or (_18071_, _18070_, _17799_);
  and (_18072_, _18071_, _11321_);
  or (_18073_, _11309_, _11300_);
  nor (_18074_, _11310_, _11321_);
  and (_18075_, _18074_, _18073_);
  or (_18076_, _18075_, _11284_);
  or (_18077_, _18076_, _18072_);
  and (_18078_, _18077_, _17796_);
  or (_18079_, _18078_, _06568_);
  or (_18080_, _17829_, _06926_);
  and (_18081_, _18080_, _11331_);
  and (_18082_, _18081_, _18079_);
  nor (_18083_, _17773_, _10213_);
  or (_18084_, _18083_, _11336_);
  and (_18085_, _18084_, _11330_);
  or (_18086_, _18085_, _11335_);
  or (_18087_, _18086_, _18082_);
  nand (_18088_, _11335_, _06055_);
  and (_18089_, _18088_, _05928_);
  and (_18090_, _18089_, _18087_);
  and (_18091_, _17859_, _05927_);
  or (_18092_, _18091_, _06278_);
  or (_18093_, _18092_, _18090_);
  and (_18094_, _14926_, _07939_);
  or (_18095_, _18094_, _17810_);
  or (_18096_, _18095_, _06279_);
  and (_18097_, _18096_, _11354_);
  and (_18098_, _18097_, _18093_);
  nor (_18099_, _11361_, \oc8051_golden_model_1.ACC [2]);
  nor (_18100_, _18099_, _11362_);
  and (_18101_, _18100_, _11353_);
  or (_18102_, _18101_, _11360_);
  or (_18103_, _18102_, _18098_);
  nand (_18104_, _11360_, _06055_);
  and (_18105_, _18104_, _01347_);
  and (_18106_, _18105_, _18103_);
  or (_18107_, _18106_, _17795_);
  and (_43164_, _18107_, _42618_);
  nor (_18108_, _01347_, _06055_);
  and (_18109_, _11054_, _10696_);
  nor (_18110_, _18109_, _11055_);
  and (_18111_, _18110_, _17724_);
  or (_18112_, _18111_, _11037_);
  nor (_18113_, _11215_, _11216_);
  or (_18114_, _18113_, _06885_);
  nand (_18115_, _06213_, _05974_);
  nor (_18116_, _07939_, _06055_);
  nor (_18117_, _10490_, _07594_);
  or (_18118_, _18117_, _18116_);
  or (_18119_, _18118_, _07215_);
  and (_18120_, _06656_, \oc8051_golden_model_1.ACC [2]);
  nor (_18121_, _17919_, _18120_);
  nor (_18122_, _12594_, _18121_);
  and (_18123_, _12594_, _18121_);
  nor (_18124_, _18123_, _18122_);
  or (_18125_, _17923_, _18124_);
  nand (_18126_, _17923_, _18124_);
  and (_18127_, _18126_, _18125_);
  or (_18128_, _18127_, _10517_);
  nor (_18129_, _08636_, _06055_);
  and (_18130_, _14950_, _08636_);
  or (_18131_, _18130_, _18129_);
  or (_18132_, _18129_, _14979_);
  and (_18133_, _18132_, _06261_);
  and (_18134_, _18133_, _18131_);
  nand (_18135_, _10744_, _07594_);
  or (_18136_, _18131_, _06273_);
  and (_18137_, _18136_, _07166_);
  and (_18138_, _14953_, _07939_);
  or (_18139_, _18138_, _18116_);
  and (_18140_, _18139_, _06341_);
  nand (_18141_, _10756_, _07594_);
  nor (_18142_, _06781_, _06055_);
  and (_18143_, _06781_, _06055_);
  nor (_18144_, _18143_, _18142_);
  nand (_18145_, _18144_, _10755_);
  and (_18146_, _18145_, _10759_);
  and (_18147_, _18146_, _18141_);
  and (_18148_, _18147_, _07155_);
  or (_18149_, _18148_, _09449_);
  or (_18150_, _18147_, _10758_);
  and (_18151_, _18150_, _06015_);
  or (_18152_, _18151_, _07154_);
  and (_18153_, _18152_, _07151_);
  and (_18154_, _18153_, _18149_);
  or (_18155_, _18154_, _18140_);
  and (_18156_, _18155_, _10776_);
  not (_18157_, \oc8051_golden_model_1.PSW [6]);
  nor (_18158_, _10778_, _18157_);
  nor (_18159_, _18158_, \oc8051_golden_model_1.ACC [3]);
  nor (_18160_, _18159_, _10779_);
  and (_18161_, _18160_, _10775_);
  or (_18162_, _18161_, _06272_);
  or (_18163_, _18162_, _18156_);
  and (_18164_, _18163_, _18137_);
  and (_18165_, _18118_, _06461_);
  or (_18166_, _18165_, _10744_);
  or (_18167_, _18166_, _18164_);
  and (_18168_, _18167_, _18135_);
  or (_18169_, _18168_, _07174_);
  or (_18170_, _09449_, _07175_);
  and (_18171_, _18170_, _06465_);
  and (_18172_, _18171_, _18169_);
  nor (_18173_, _08291_, _06465_);
  or (_18174_, _18173_, _10811_);
  or (_18175_, _18174_, _18172_);
  nand (_18176_, _10811_, _08572_);
  and (_18177_, _18176_, _18175_);
  or (_18178_, _18177_, _06268_);
  and (_18179_, _14948_, _08636_);
  or (_18180_, _18179_, _18129_);
  or (_18181_, _18180_, _06269_);
  and (_18182_, _18181_, _06262_);
  and (_18183_, _18182_, _18178_);
  or (_18184_, _18183_, _18134_);
  and (_18185_, _18184_, _09537_);
  or (_18186_, _10037_, _10035_);
  nor (_18187_, _10038_, _09537_);
  nand (_18188_, _18187_, _18186_);
  nand (_18189_, _18188_, _10731_);
  or (_18190_, _18189_, _18185_);
  and (_18191_, _07776_, \oc8051_golden_model_1.ACC [2]);
  nor (_18192_, _17877_, _18191_);
  nor (_18193_, _11171_, _11172_);
  not (_18194_, _18193_);
  and (_18195_, _18194_, _18192_);
  nor (_18196_, _18194_, _18192_);
  nor (_18197_, _18196_, _18195_);
  nor (_18198_, _18197_, _10558_);
  and (_18199_, _18197_, _10558_);
  nor (_18200_, _18199_, _18198_);
  and (_18201_, _17879_, \oc8051_golden_model_1.PSW [7]);
  nor (_18202_, _17880_, _10558_);
  nor (_18203_, _18202_, _18201_);
  not (_18204_, _18203_);
  and (_18205_, _18204_, _18200_);
  nor (_18206_, _18204_, _18200_);
  nor (_18207_, _18206_, _18205_);
  and (_18208_, _18207_, _10734_);
  or (_18209_, _18208_, _10735_);
  and (_18210_, _18209_, _18190_);
  and (_18211_, _18207_, _10733_);
  or (_18212_, _18211_, _10656_);
  or (_18213_, _18212_, _18210_);
  and (_18214_, _09302_, \oc8051_golden_model_1.ACC [2]);
  nor (_18215_, _17892_, _18214_);
  nor (_18216_, _18113_, _18215_);
  and (_18217_, _18113_, _18215_);
  nor (_18218_, _18217_, _18216_);
  and (_18219_, _18218_, \oc8051_golden_model_1.PSW [7]);
  nor (_18220_, _18218_, \oc8051_golden_model_1.PSW [7]);
  nor (_18221_, _18220_, _18219_);
  and (_18222_, _18221_, _17898_);
  nor (_18223_, _18221_, _17898_);
  nor (_18224_, _18223_, _18222_);
  or (_18225_, _18224_, _10588_);
  and (_18226_, _18225_, _06517_);
  and (_18227_, _18226_, _18213_);
  and (_18228_, _12583_, \oc8051_golden_model_1.PSW [7]);
  and (_18229_, _08439_, \oc8051_golden_model_1.ACC [2]);
  nor (_18230_, _17910_, _18229_);
  nor (_18231_, _12577_, _18230_);
  and (_18232_, _12577_, _18230_);
  nor (_18233_, _18232_, _18231_);
  not (_18234_, _12582_);
  or (_18235_, _18234_, _17912_);
  or (_18236_, _18235_, _10558_);
  and (_18237_, _18236_, _18233_);
  or (_18238_, _18237_, _10516_);
  or (_18239_, _18238_, _18228_);
  and (_18240_, _18239_, _12644_);
  or (_18241_, _18240_, _18227_);
  and (_18242_, _18241_, _18128_);
  or (_18243_, _18242_, _10515_);
  nand (_18244_, _06213_, _10515_);
  and (_18245_, _18244_, _06258_);
  and (_18246_, _18245_, _18243_);
  or (_18247_, _18129_, _14992_);
  and (_18248_, _18247_, _06257_);
  and (_18249_, _18248_, _18131_);
  or (_18250_, _18249_, _10080_);
  or (_18251_, _18250_, _18246_);
  and (_18252_, _18251_, _18119_);
  or (_18253_, _18252_, _07460_);
  and (_18254_, _09449_, _07939_);
  or (_18255_, _18116_, _07208_);
  or (_18256_, _18255_, _18254_);
  and (_18257_, _18256_, _05982_);
  and (_18258_, _18257_, _18253_);
  and (_18259_, _15048_, _07939_);
  or (_18260_, _18259_, _18116_);
  and (_18261_, _18260_, _10094_);
  or (_18262_, _18261_, _10093_);
  or (_18263_, _18262_, _18258_);
  or (_18264_, _10235_, _10100_);
  and (_18265_, _18264_, _18263_);
  or (_18266_, _18265_, _05974_);
  and (_18267_, _18266_, _18115_);
  or (_18268_, _18267_, _06218_);
  and (_18269_, _07939_, _08930_);
  or (_18270_, _18269_, _18116_);
  or (_18271_, _18270_, _06219_);
  and (_18272_, _18271_, _10930_);
  and (_18273_, _18272_, _18268_);
  or (_18274_, _10930_, _06213_);
  or (_18275_, _06734_, _06328_);
  and (_18276_, _18275_, _06535_);
  and (_18277_, _06335_, _06535_);
  or (_18278_, _10506_, _18277_);
  nor (_18279_, _18278_, _18276_);
  nand (_18280_, _18279_, _18274_);
  or (_18281_, _18280_, _18273_);
  nor (_18282_, _17511_, _06887_);
  or (_18283_, _18279_, _18193_);
  and (_18284_, _18283_, _18282_);
  and (_18285_, _18284_, _18281_);
  not (_18286_, _18282_);
  and (_18287_, _18286_, _18193_);
  or (_18288_, _18287_, _06888_);
  or (_18289_, _18288_, _18285_);
  or (_18290_, _18193_, _17510_);
  and (_18291_, _18290_, _17375_);
  and (_18292_, _18291_, _18289_);
  or (_18293_, _18113_, _06884_);
  and (_18294_, _18293_, _10948_);
  or (_18295_, _18294_, _18292_);
  and (_18296_, _18295_, _18114_);
  or (_18297_, _18296_, _06533_);
  or (_18298_, _12577_, _06534_);
  and (_18299_, _18298_, _10955_);
  and (_18300_, _18299_, _18297_);
  and (_18301_, _10954_, _12594_);
  or (_18302_, _18301_, _06369_);
  or (_18303_, _18302_, _18300_);
  and (_18304_, _14943_, _07939_);
  or (_18305_, _18304_, _18116_);
  or (_18306_, _18305_, _07237_);
  and (_18307_, _18306_, _18303_);
  or (_18308_, _18307_, _06536_);
  or (_18309_, _18116_, _07240_);
  and (_18310_, _18309_, _10977_);
  and (_18311_, _18310_, _18308_);
  or (_18312_, _10985_, _11171_);
  and (_18313_, _18312_, _10987_);
  or (_18314_, _18313_, _18311_);
  or (_18315_, _17402_, _11171_);
  and (_18316_, _18315_, _17401_);
  and (_18317_, _18316_, _18314_);
  and (_18318_, _10983_, _11215_);
  or (_18319_, _18318_, _06542_);
  or (_18320_, _18319_, _18317_);
  or (_18321_, _11255_, _06543_);
  and (_18322_, _18321_, _10497_);
  and (_18323_, _18322_, _18320_);
  and (_18324_, _11296_, _10496_);
  or (_18325_, _18324_, _18323_);
  and (_18326_, _18325_, _07242_);
  nand (_18327_, _18270_, _06375_);
  nor (_18328_, _18327_, _11256_);
  or (_18329_, _18328_, _10999_);
  or (_18330_, _18329_, _18326_);
  nand (_18331_, _10999_, _11172_);
  and (_18332_, _18331_, _07043_);
  and (_18333_, _18332_, _11009_);
  and (_18334_, _18333_, _18330_);
  and (_18335_, _11009_, _07043_);
  nor (_18336_, _18335_, _11172_);
  or (_18337_, _18336_, _11014_);
  or (_18338_, _18337_, _18334_);
  nand (_18339_, _11014_, _11216_);
  and (_18340_, _18339_, _06531_);
  and (_18341_, _18340_, _18338_);
  nand (_18342_, _11024_, _11256_);
  and (_18343_, _18342_, _11023_);
  or (_18344_, _18343_, _18341_);
  nand (_18345_, _11021_, _11297_);
  and (_18346_, _18345_, _09056_);
  and (_18347_, _18346_, _18344_);
  and (_18348_, _14940_, _07939_);
  or (_18349_, _18348_, _18116_);
  nand (_18350_, _18349_, _06366_);
  nand (_18351_, _18350_, _17505_);
  or (_18352_, _18351_, _18347_);
  and (_18353_, _18352_, _18112_);
  and (_18354_, _18110_, _17723_);
  or (_18355_, _18354_, _11041_);
  or (_18356_, _18355_, _18353_);
  and (_18357_, _11082_, _10622_);
  nor (_18358_, _18357_, _11083_);
  or (_18359_, _18358_, _11069_);
  and (_18360_, _18359_, _06541_);
  and (_18361_, _18360_, _18356_);
  and (_18362_, _11110_, _10869_);
  nor (_18363_, _18362_, _11111_);
  or (_18364_, _18363_, _11097_);
  and (_18365_, _18364_, _14297_);
  or (_18366_, _18365_, _18361_);
  and (_18367_, _11138_, _10551_);
  nor (_18368_, _18367_, _11139_);
  or (_18369_, _18368_, _11127_);
  and (_18370_, _18369_, _11126_);
  and (_18371_, _18370_, _18366_);
  and (_18372_, _11125_, \oc8051_golden_model_1.ACC [2]);
  nor (_18373_, _18372_, _11201_);
  nand (_18374_, _18373_, _11157_);
  or (_18375_, _18374_, _18371_);
  nor (_18376_, _11228_, _18113_);
  and (_18377_, _11228_, _18113_);
  or (_18378_, _18377_, _18376_);
  or (_18379_, _18378_, _11203_);
  or (_18380_, _11184_, _18194_);
  nand (_18381_, _11184_, _18194_);
  and (_18382_, _18381_, _18380_);
  or (_18383_, _18382_, _11157_);
  and (_18384_, _18383_, _06285_);
  and (_18385_, _18384_, _18379_);
  and (_18386_, _18385_, _18375_);
  and (_18387_, _11268_, _12577_);
  nor (_18388_, _11268_, _12577_);
  or (_18389_, _18388_, _18387_);
  and (_18390_, _18389_, _06283_);
  or (_18391_, _18390_, _11243_);
  or (_18392_, _18391_, _18386_);
  and (_18393_, _11311_, _12594_);
  nor (_18394_, _11311_, _12594_);
  or (_18395_, _18394_, _11321_);
  or (_18396_, _18395_, _18393_);
  and (_18397_, _18396_, _11285_);
  and (_18398_, _18397_, _18392_);
  and (_18399_, _11284_, \oc8051_golden_model_1.ACC [2]);
  or (_18400_, _18399_, _06568_);
  or (_18401_, _18400_, _18398_);
  or (_18402_, _18139_, _06926_);
  and (_18403_, _18402_, _11331_);
  and (_18404_, _18403_, _18401_);
  nor (_18405_, _11336_, _06055_);
  or (_18406_, _18405_, _11337_);
  and (_18407_, _18406_, _11330_);
  or (_18408_, _18407_, _11335_);
  or (_18409_, _18408_, _18404_);
  nand (_18410_, _11335_, _10135_);
  and (_18411_, _18410_, _05928_);
  and (_18412_, _18411_, _18409_);
  and (_18413_, _18180_, _05927_);
  or (_18414_, _18413_, _06278_);
  or (_18415_, _18414_, _18412_);
  and (_18416_, _15128_, _07939_);
  or (_18417_, _18416_, _18116_);
  or (_18418_, _18417_, _06279_);
  and (_18419_, _18418_, _11354_);
  and (_18420_, _18419_, _18415_);
  nor (_18421_, _11362_, \oc8051_golden_model_1.ACC [3]);
  nor (_18422_, _18421_, _11363_);
  and (_18423_, _18422_, _11353_);
  or (_18424_, _18423_, _11360_);
  or (_18425_, _18424_, _18420_);
  nand (_18426_, _11360_, _10135_);
  and (_18427_, _18426_, _01347_);
  and (_18428_, _18427_, _18425_);
  or (_18429_, _18428_, _18108_);
  and (_43165_, _18429_, _42618_);
  nor (_18430_, _01347_, _10135_);
  or (_18431_, _11230_, _11214_);
  and (_18432_, _18431_, _11231_);
  or (_18433_, _18432_, _17800_);
  or (_18434_, _11056_, _10689_);
  and (_18435_, _18434_, _11057_);
  and (_18436_, _18435_, _14283_);
  nand (_18437_, _11021_, _11294_);
  or (_18438_, _12157_, _11169_);
  or (_18439_, _17401_, _11211_);
  or (_18440_, _11214_, _10502_);
  nand (_18441_, _06968_, _05974_);
  nor (_18442_, _07939_, _10135_);
  nor (_18443_, _08541_, _10490_);
  or (_18444_, _18443_, _18442_);
  or (_18445_, _18444_, _07215_);
  nor (_18446_, _12583_, _10558_);
  or (_18447_, _18230_, _14140_);
  and (_18448_, _18447_, _14139_);
  nor (_18449_, _11254_, _18448_);
  and (_18450_, _11254_, _18448_);
  nor (_18451_, _18450_, _18449_);
  and (_18452_, _18451_, \oc8051_golden_model_1.PSW [7]);
  nor (_18453_, _18451_, \oc8051_golden_model_1.PSW [7]);
  nor (_18454_, _18453_, _18452_);
  or (_18455_, _18454_, _18446_);
  and (_18456_, _18454_, _18446_);
  nor (_18457_, _18456_, _06517_);
  and (_18458_, _18457_, _18455_);
  or (_18459_, _18205_, _18198_);
  nor (_18460_, _07594_, \oc8051_golden_model_1.ACC [3]);
  nand (_18461_, _07594_, \oc8051_golden_model_1.ACC [3]);
  and (_18462_, _18461_, _18192_);
  or (_18463_, _18462_, _18460_);
  nor (_18464_, _11170_, _18463_);
  and (_18465_, _11170_, _18463_);
  nor (_18466_, _18465_, _18464_);
  and (_18467_, _18466_, \oc8051_golden_model_1.PSW [7]);
  nor (_18468_, _18466_, \oc8051_golden_model_1.PSW [7]);
  nor (_18469_, _18468_, _18467_);
  or (_18470_, _18469_, _18459_);
  and (_18471_, _18469_, _18459_);
  nor (_18472_, _10735_, _18471_);
  and (_18473_, _18472_, _18470_);
  nand (_18474_, _10744_, _08541_);
  nor (_18475_, _08636_, _10135_);
  and (_18476_, _15166_, _08636_);
  or (_18477_, _18476_, _18475_);
  or (_18478_, _18477_, _06273_);
  and (_18479_, _18478_, _07166_);
  nand (_18480_, _10756_, _08541_);
  nor (_18481_, _06781_, _10135_);
  and (_18482_, _06781_, _10135_);
  nor (_18483_, _18482_, _18481_);
  nand (_18484_, _18483_, _10755_);
  and (_18485_, _18484_, _10759_);
  and (_18486_, _18485_, _18480_);
  and (_18487_, _10758_, _09448_);
  or (_18488_, _18487_, _18486_);
  and (_18489_, _18488_, _10769_);
  and (_18490_, _15162_, _07939_);
  or (_18491_, _18490_, _18442_);
  and (_18492_, _18491_, _06341_);
  or (_18493_, _18492_, _18489_);
  and (_18494_, _18493_, _10776_);
  nor (_18495_, _10779_, \oc8051_golden_model_1.ACC [4]);
  nor (_18496_, _18495_, _10780_);
  and (_18497_, _18496_, _10775_);
  or (_18498_, _18497_, _06272_);
  or (_18499_, _18498_, _18494_);
  and (_18500_, _18499_, _18479_);
  and (_18501_, _18444_, _06461_);
  or (_18502_, _18501_, _10744_);
  or (_18503_, _18502_, _18500_);
  and (_18504_, _18503_, _18474_);
  or (_18505_, _18504_, _07174_);
  or (_18506_, _09448_, _07175_);
  and (_18507_, _18506_, _06465_);
  and (_18508_, _18507_, _18505_);
  nor (_18509_, _08543_, _06465_);
  or (_18510_, _18509_, _10811_);
  or (_18511_, _18510_, _18508_);
  nand (_18512_, _10811_, _06097_);
  and (_18513_, _18512_, _18511_);
  or (_18514_, _18513_, _06268_);
  and (_18515_, _15176_, _08636_);
  or (_18516_, _18515_, _18475_);
  or (_18517_, _18516_, _06269_);
  and (_18518_, _18517_, _06262_);
  and (_18519_, _18518_, _18514_);
  or (_18520_, _18475_, _15183_);
  and (_18521_, _18520_, _06261_);
  and (_18522_, _18521_, _18477_);
  or (_18523_, _18522_, _09531_);
  or (_18524_, _18523_, _18519_);
  nor (_18525_, _10040_, _10038_);
  nor (_18526_, _18525_, _10041_);
  or (_18527_, _18526_, _09537_);
  and (_18528_, _18527_, _10735_);
  and (_18529_, _18528_, _18524_);
  nor (_18530_, _18529_, _18473_);
  nor (_18531_, _18530_, _10587_);
  or (_18532_, _18222_, _18219_);
  and (_18533_, _09449_, _06055_);
  or (_18534_, _09449_, _06055_);
  and (_18535_, _18534_, _18215_);
  or (_18536_, _18535_, _18533_);
  nor (_18537_, _11214_, _18536_);
  and (_18538_, _11214_, _18536_);
  nor (_18539_, _18538_, _18537_);
  and (_18540_, _18539_, \oc8051_golden_model_1.PSW [7]);
  nor (_18541_, _18539_, \oc8051_golden_model_1.PSW [7]);
  nor (_18542_, _18541_, _18540_);
  and (_18543_, _18542_, _18532_);
  nor (_18544_, _18542_, _18532_);
  nor (_18545_, _18544_, _18543_);
  and (_18546_, _18545_, _10587_);
  or (_18547_, _18546_, _18531_);
  or (_18548_, _18547_, _10586_);
  not (_18549_, _10586_);
  or (_18550_, _18545_, _18549_);
  and (_18551_, _18550_, _06517_);
  and (_18552_, _18551_, _18548_);
  or (_18553_, _18552_, _18458_);
  and (_18554_, _18553_, _10517_);
  nor (_18555_, _12599_, _10558_);
  or (_18556_, _18121_, _14161_);
  and (_18557_, _18556_, _14160_);
  nor (_18558_, _11295_, _18557_);
  and (_18559_, _11295_, _18557_);
  nor (_18560_, _18559_, _18558_);
  and (_18561_, _18560_, \oc8051_golden_model_1.PSW [7]);
  nor (_18562_, _18560_, \oc8051_golden_model_1.PSW [7]);
  nor (_18563_, _18562_, _18561_);
  or (_18564_, _18563_, _18555_);
  and (_18565_, _18563_, _18555_);
  nor (_18566_, _18565_, _10517_);
  and (_18567_, _18566_, _18564_);
  or (_18568_, _18567_, _10515_);
  or (_18569_, _18568_, _18554_);
  nand (_18570_, _06968_, _10515_);
  and (_18571_, _18570_, _06258_);
  and (_18572_, _18571_, _18569_);
  and (_18573_, _15200_, _08636_);
  or (_18574_, _18573_, _18475_);
  and (_18575_, _18574_, _06257_);
  or (_18576_, _18575_, _10080_);
  or (_18577_, _18576_, _18572_);
  and (_18578_, _18577_, _18445_);
  or (_18579_, _18578_, _07460_);
  and (_18580_, _09448_, _07939_);
  or (_18581_, _18442_, _07208_);
  or (_18582_, _18581_, _18580_);
  and (_18583_, _18582_, _05982_);
  and (_18584_, _18583_, _18579_);
  and (_18585_, _15254_, _07939_);
  or (_18586_, _18585_, _18442_);
  and (_18587_, _18586_, _10094_);
  or (_18588_, _18587_, _10093_);
  or (_18589_, _18588_, _18584_);
  or (_18590_, _10181_, _10100_);
  and (_18591_, _18590_, _18589_);
  or (_18592_, _18591_, _05974_);
  and (_18593_, _18592_, _18441_);
  or (_18594_, _18593_, _06218_);
  and (_18595_, _08959_, _07939_);
  or (_18596_, _18595_, _18442_);
  or (_18597_, _18596_, _06219_);
  and (_18598_, _18597_, _10930_);
  and (_18599_, _18598_, _18594_);
  nor (_18600_, _10930_, _06968_);
  or (_18601_, _18600_, _18277_);
  or (_18602_, _18601_, _18599_);
  not (_18603_, _18277_);
  or (_18604_, _11170_, _18603_);
  and (_18605_, _18604_, _18602_);
  or (_18606_, _18605_, _06891_);
  not (_18607_, _06891_);
  or (_18608_, _11170_, _18607_);
  and (_18609_, _18608_, _06745_);
  and (_18610_, _18609_, _18606_);
  and (_18611_, _11170_, _06744_);
  or (_18612_, _18611_, _10507_);
  or (_18613_, _18612_, _18610_);
  not (_18614_, _10507_);
  or (_18615_, _11170_, _18614_);
  and (_18616_, _18615_, _17972_);
  and (_18617_, _18616_, _18613_);
  and (_18618_, _17971_, _11170_);
  or (_18619_, _18618_, _10948_);
  or (_18620_, _18619_, _18617_);
  and (_18621_, _18620_, _18440_);
  or (_18622_, _18621_, _06533_);
  or (_18623_, _11254_, _06534_);
  and (_18624_, _18623_, _10955_);
  and (_18625_, _18624_, _18622_);
  and (_18626_, _10954_, _11295_);
  or (_18627_, _18626_, _06369_);
  or (_18628_, _18627_, _18625_);
  and (_18629_, _15269_, _07939_);
  or (_18630_, _18629_, _18442_);
  or (_18631_, _18630_, _07237_);
  and (_18632_, _18631_, _18628_);
  or (_18633_, _18632_, _06536_);
  or (_18634_, _18442_, _07240_);
  and (_18635_, _18634_, _10986_);
  and (_18636_, _18635_, _18633_);
  and (_18637_, _10987_, _11167_);
  or (_18638_, _18637_, _10983_);
  or (_18639_, _18638_, _18636_);
  and (_18640_, _18639_, _18439_);
  or (_18641_, _18640_, _06542_);
  or (_18642_, _11251_, _06543_);
  and (_18643_, _18642_, _10497_);
  and (_18644_, _18643_, _18641_);
  and (_18645_, _11292_, _10496_);
  or (_18646_, _18645_, _18644_);
  and (_18647_, _18646_, _07242_);
  nand (_18648_, _18596_, _06375_);
  nor (_18649_, _18648_, _11253_);
  or (_18650_, _18649_, _17507_);
  or (_18651_, _18650_, _18647_);
  and (_18652_, _18651_, _18438_);
  or (_18653_, _18652_, _17506_);
  or (_18654_, _17423_, _11169_);
  and (_18655_, _18654_, _17430_);
  and (_18656_, _18655_, _18653_);
  and (_18657_, _11169_, _17429_);
  or (_18658_, _18657_, _11014_);
  or (_18659_, _18658_, _18656_);
  or (_18660_, _11013_, _11213_);
  and (_18661_, _18660_, _06531_);
  and (_18662_, _18661_, _18659_);
  nand (_18663_, _11024_, _11253_);
  and (_18664_, _18663_, _11023_);
  or (_18665_, _18664_, _18662_);
  and (_18666_, _18665_, _18437_);
  or (_18667_, _18666_, _06366_);
  and (_18668_, _15266_, _07939_);
  or (_18669_, _18442_, _09056_);
  or (_18670_, _18669_, _18668_);
  and (_18671_, _18670_, _11037_);
  and (_18672_, _18671_, _18667_);
  or (_18673_, _18672_, _18436_);
  and (_18674_, _18673_, _17722_);
  or (_18675_, _11084_, _10616_);
  and (_18676_, _18675_, _11085_);
  and (_18677_, _18676_, _11040_);
  or (_18678_, _18677_, _11039_);
  or (_18679_, _18678_, _18674_);
  or (_18680_, _18676_, _17733_);
  and (_18681_, _18680_, _06541_);
  and (_18682_, _18681_, _18679_);
  or (_18683_, _11112_, _10863_);
  and (_18684_, _18683_, _11113_);
  or (_18685_, _18684_, _11097_);
  and (_18686_, _18685_, _14297_);
  or (_18687_, _18686_, _18682_);
  or (_18688_, _11140_, _10545_);
  and (_18689_, _18688_, _11141_);
  or (_18690_, _18689_, _11127_);
  and (_18691_, _18690_, _18687_);
  or (_18692_, _18691_, _11125_);
  nand (_18693_, _11125_, _06055_);
  and (_18694_, _18693_, _11157_);
  and (_18695_, _18694_, _18692_);
  nor (_18696_, _11186_, _11170_);
  nor (_18697_, _18696_, _11187_);
  and (_18698_, _18697_, _18059_);
  or (_18699_, _18698_, _11200_);
  or (_18700_, _18699_, _18695_);
  and (_18701_, _18700_, _18433_);
  or (_18702_, _18701_, _11199_);
  or (_18703_, _18432_, _18067_);
  and (_18704_, _18703_, _13012_);
  and (_18705_, _18704_, _18702_);
  or (_18706_, _11313_, _11295_);
  and (_18707_, _18706_, _11314_);
  and (_18708_, _18707_, _11243_);
  or (_18709_, _18708_, _11284_);
  or (_18710_, _11270_, _11254_);
  and (_18711_, _11271_, _06283_);
  and (_18712_, _18711_, _18710_);
  or (_18713_, _18712_, _18709_);
  or (_18714_, _18713_, _18705_);
  nand (_18715_, _11284_, _06055_);
  and (_18716_, _18715_, _18714_);
  or (_18717_, _18716_, _06568_);
  or (_18718_, _18491_, _06926_);
  and (_18719_, _18718_, _11331_);
  and (_18720_, _18719_, _18717_);
  nor (_18721_, _11337_, _10135_);
  or (_18722_, _18721_, _11338_);
  and (_18723_, _18722_, _11330_);
  or (_18724_, _18723_, _11335_);
  or (_18725_, _18724_, _18720_);
  nand (_18726_, _11335_, _10170_);
  and (_18727_, _18726_, _05928_);
  and (_18728_, _18727_, _18725_);
  and (_18729_, _18516_, _05927_);
  or (_18730_, _18729_, _06278_);
  or (_18731_, _18730_, _18728_);
  and (_18732_, _15329_, _07939_);
  or (_18733_, _18732_, _18442_);
  or (_18734_, _18733_, _06279_);
  and (_18735_, _18734_, _11354_);
  and (_18736_, _18735_, _18731_);
  nor (_18737_, _11363_, \oc8051_golden_model_1.ACC [4]);
  nor (_18738_, _18737_, _11364_);
  and (_18739_, _18738_, _11353_);
  or (_18740_, _18739_, _11360_);
  or (_18741_, _18740_, _18736_);
  nand (_18742_, _11360_, _10170_);
  and (_18743_, _18742_, _01347_);
  and (_18744_, _18743_, _18741_);
  or (_18745_, _18744_, _18430_);
  and (_43166_, _18745_, _42618_);
  nor (_18746_, _01347_, _10170_);
  and (_18747_, _11058_, _10686_);
  nor (_18748_, _18747_, _11059_);
  or (_18749_, _18748_, _11037_);
  or (_18750_, _11248_, _06543_);
  and (_18752_, _18750_, _10497_);
  nand (_18753_, _11210_, _10948_);
  or (_18754_, _11166_, _06704_);
  and (_18755_, _18754_, _17969_);
  and (_18756_, _11166_, _06891_);
  nand (_18757_, _06611_, _05974_);
  nor (_18758_, _07939_, _10170_);
  nor (_18759_, _08244_, _10490_);
  or (_18760_, _18759_, _18758_);
  or (_18761_, _18760_, _07215_);
  and (_18762_, _06968_, \oc8051_golden_model_1.ACC [4]);
  nor (_18763_, _18558_, _18762_);
  nor (_18764_, _12600_, _18763_);
  and (_18765_, _12600_, _18763_);
  nor (_18766_, _18765_, _18764_);
  and (_18767_, _18766_, \oc8051_golden_model_1.PSW [7]);
  nor (_18768_, _18766_, \oc8051_golden_model_1.PSW [7]);
  nor (_18769_, _18768_, _18767_);
  nor (_18770_, _18565_, _18561_);
  not (_18771_, _18770_);
  and (_18774_, _18771_, _18769_);
  nor (_18775_, _18771_, _18769_);
  nor (_18776_, _18775_, _18774_);
  or (_18777_, _18776_, _10517_);
  not (_18778_, _10730_);
  and (_18779_, _08541_, \oc8051_golden_model_1.ACC [4]);
  nor (_18780_, _18464_, _18779_);
  nor (_18781_, _11166_, _18780_);
  and (_18782_, _11166_, _18780_);
  nor (_18783_, _18782_, _18781_);
  and (_18785_, _18783_, \oc8051_golden_model_1.PSW [7]);
  nor (_18786_, _18783_, \oc8051_golden_model_1.PSW [7]);
  nor (_18787_, _18786_, _18785_);
  nor (_18788_, _18471_, _18467_);
  not (_18789_, _18788_);
  and (_18790_, _18789_, _18787_);
  nor (_18791_, _18789_, _18787_);
  nor (_18792_, _18791_, _18790_);
  or (_18793_, _18792_, _18778_);
  nor (_18794_, _08636_, _10170_);
  and (_18796_, _15372_, _08636_);
  or (_18797_, _18796_, _18794_);
  or (_18798_, _18794_, _15387_);
  and (_18799_, _18798_, _06261_);
  and (_18800_, _18799_, _18797_);
  nand (_18801_, _10744_, _08244_);
  nand (_18802_, _10756_, _08244_);
  nor (_18803_, _06781_, _10170_);
  and (_18804_, _06781_, _10170_);
  nor (_18805_, _18804_, _18803_);
  nand (_18807_, _18805_, _10755_);
  and (_18808_, _18807_, _10759_);
  and (_18809_, _18808_, _18802_);
  and (_18810_, _10758_, _09447_);
  or (_18811_, _18810_, _18809_);
  and (_18812_, _18811_, _10769_);
  and (_18813_, _15358_, _07939_);
  or (_18814_, _18813_, _18758_);
  and (_18815_, _18814_, _06341_);
  or (_18816_, _18815_, _10775_);
  or (_18818_, _18816_, _18812_);
  nor (_18819_, _10795_, _10787_);
  nand (_18820_, _10795_, _10787_);
  nand (_18821_, _18820_, _10775_);
  or (_18822_, _18821_, _18819_);
  and (_18823_, _18822_, _06466_);
  and (_18824_, _18823_, _18818_);
  and (_18825_, _18797_, _06272_);
  and (_18826_, _18760_, _06461_);
  or (_18827_, _18826_, _10744_);
  or (_18829_, _18827_, _18825_);
  or (_18830_, _18829_, _18824_);
  and (_18831_, _18830_, _18801_);
  or (_18832_, _18831_, _07174_);
  or (_18833_, _09447_, _07175_);
  and (_18834_, _18833_, _06465_);
  and (_18835_, _18834_, _18832_);
  nor (_18836_, _08246_, _06465_);
  or (_18837_, _18836_, _10811_);
  or (_18838_, _18837_, _18835_);
  nand (_18840_, _10811_, _06042_);
  and (_18841_, _18840_, _18838_);
  or (_18842_, _18841_, _06268_);
  and (_18843_, _15355_, _08636_);
  or (_18844_, _18843_, _18794_);
  or (_18845_, _18844_, _06269_);
  and (_18846_, _18845_, _06262_);
  and (_18847_, _18846_, _18842_);
  or (_18848_, _18847_, _18800_);
  and (_18849_, _18848_, _09537_);
  or (_18851_, _10043_, _10041_);
  nor (_18852_, _10044_, _09537_);
  and (_18853_, _18852_, _18851_);
  or (_18854_, _18853_, _10730_);
  or (_18855_, _18854_, _18849_);
  and (_18856_, _18855_, _18793_);
  or (_18857_, _18856_, _17310_);
  not (_18858_, _17310_);
  or (_18859_, _18792_, _18858_);
  and (_18860_, _18859_, _14204_);
  and (_18862_, _18860_, _18857_);
  and (_18863_, _18792_, _14203_);
  or (_18864_, _18863_, _10656_);
  or (_18865_, _18864_, _18862_);
  and (_18866_, _09212_, \oc8051_golden_model_1.ACC [4]);
  nor (_18867_, _18537_, _18866_);
  nor (_18868_, _11210_, _18867_);
  and (_18869_, _11210_, _18867_);
  nor (_18870_, _18869_, _18868_);
  nor (_18871_, _18870_, _10558_);
  and (_18873_, _18870_, _10558_);
  nor (_18874_, _18873_, _18871_);
  nor (_18875_, _18543_, _18540_);
  not (_18876_, _18875_);
  and (_18877_, _18876_, _18874_);
  nor (_18878_, _18876_, _18874_);
  nor (_18879_, _18878_, _18877_);
  or (_18880_, _18879_, _10588_);
  and (_18881_, _18880_, _06517_);
  and (_18882_, _18881_, _18865_);
  and (_18884_, _08543_, \oc8051_golden_model_1.ACC [4]);
  nor (_18885_, _18449_, _18884_);
  nor (_18886_, _11250_, _18885_);
  and (_18887_, _11250_, _18885_);
  nor (_18888_, _18887_, _18886_);
  and (_18889_, _18888_, \oc8051_golden_model_1.PSW [7]);
  nor (_18890_, _18888_, \oc8051_golden_model_1.PSW [7]);
  nor (_18891_, _18890_, _18889_);
  nor (_18892_, _18456_, _18452_);
  not (_18893_, _18892_);
  and (_18895_, _18893_, _18891_);
  nor (_18896_, _18893_, _18891_);
  nor (_18897_, _18896_, _18895_);
  or (_18898_, _18897_, _10516_);
  and (_18899_, _18898_, _12644_);
  or (_18900_, _18899_, _18882_);
  and (_18901_, _18900_, _18777_);
  or (_18902_, _18901_, _10515_);
  nand (_18903_, _06611_, _10515_);
  and (_18904_, _18903_, _06258_);
  and (_18906_, _18904_, _18902_);
  or (_18907_, _18794_, _15403_);
  and (_18908_, _18907_, _06257_);
  and (_18909_, _18908_, _18797_);
  or (_18910_, _18909_, _10080_);
  or (_18911_, _18910_, _18906_);
  and (_18912_, _18911_, _18761_);
  or (_18913_, _18912_, _07460_);
  and (_18914_, _09447_, _07939_);
  or (_18915_, _18758_, _07208_);
  or (_18917_, _18915_, _18914_);
  and (_18918_, _18917_, _05982_);
  and (_18919_, _18918_, _18913_);
  and (_18920_, _15459_, _07939_);
  or (_18921_, _18920_, _18758_);
  and (_18922_, _18921_, _10094_);
  or (_18923_, _18922_, _10093_);
  or (_18924_, _18923_, _18919_);
  or (_18925_, _10153_, _10100_);
  and (_18926_, _18925_, _18924_);
  or (_18927_, _18926_, _05974_);
  and (_18928_, _18927_, _18757_);
  or (_18929_, _18928_, _06218_);
  and (_18930_, _08946_, _07939_);
  or (_18931_, _18930_, _18758_);
  or (_18932_, _18931_, _06219_);
  and (_18933_, _18932_, _10930_);
  and (_18934_, _18933_, _18929_);
  nor (_18935_, _10930_, _06611_);
  or (_18936_, _18935_, _18277_);
  or (_18938_, _18936_, _18934_);
  or (_18939_, _11166_, _18603_);
  and (_18940_, _18939_, _18607_);
  and (_18941_, _18940_, _18938_);
  or (_18942_, _18941_, _18756_);
  and (_18943_, _18942_, _06745_);
  and (_18944_, _11166_, _06744_);
  or (_18945_, _18944_, _06703_);
  or (_18946_, _18945_, _18943_);
  and (_18947_, _18946_, _18755_);
  and (_18949_, _11166_, _10506_);
  or (_18950_, _18949_, _06887_);
  or (_18951_, _18950_, _18947_);
  not (_18952_, _06887_);
  or (_18953_, _11166_, _18952_);
  and (_18954_, _18953_, _10946_);
  and (_18955_, _18954_, _18951_);
  and (_18956_, _10945_, _11166_);
  or (_18957_, _18956_, _10948_);
  or (_18958_, _18957_, _18955_);
  and (_18960_, _18958_, _18753_);
  or (_18961_, _18960_, _06533_);
  or (_18962_, _11250_, _06534_);
  and (_18963_, _18962_, _10955_);
  and (_18964_, _18963_, _18961_);
  and (_18965_, _10954_, _12600_);
  or (_18966_, _18965_, _06369_);
  or (_18967_, _18966_, _18964_);
  and (_18968_, _15353_, _07939_);
  or (_18969_, _18968_, _18758_);
  or (_18971_, _18969_, _07237_);
  and (_18972_, _18971_, _18967_);
  or (_18973_, _18972_, _06536_);
  and (_18974_, _11032_, _07211_);
  or (_18975_, _18974_, _05960_);
  or (_18976_, _18758_, _07240_);
  and (_18977_, _18976_, _18975_);
  and (_18978_, _18977_, _18973_);
  and (_18979_, _10987_, _11164_);
  or (_18980_, _18979_, _18978_);
  nand (_18982_, _10732_, _06544_);
  or (_18983_, _18982_, _11164_);
  and (_18984_, _18983_, _17401_);
  and (_18985_, _18984_, _18980_);
  and (_18986_, _10983_, _11208_);
  or (_18987_, _18986_, _06542_);
  or (_18988_, _18987_, _18985_);
  and (_18989_, _18988_, _18752_);
  and (_18990_, _11290_, _10496_);
  or (_18991_, _18990_, _18989_);
  and (_18993_, _18991_, _07242_);
  nand (_18994_, _18931_, _06375_);
  nor (_18995_, _18994_, _11249_);
  or (_18996_, _18995_, _17507_);
  or (_18997_, _18996_, _18993_);
  nand (_18998_, _17507_, _11165_);
  and (_18999_, _18998_, _18997_);
  or (_19000_, _18999_, _17506_);
  nand (_19001_, _17506_, _11165_);
  and (_19002_, _19001_, _17430_);
  and (_19004_, _19002_, _19000_);
  nor (_19005_, _11165_, _17430_);
  or (_19006_, _19005_, _11014_);
  or (_19007_, _19006_, _19004_);
  or (_19008_, _11013_, \oc8051_golden_model_1.ACC [5]);
  or (_19009_, _19008_, _09447_);
  and (_19010_, _19009_, _06531_);
  and (_19011_, _19010_, _19007_);
  nand (_19012_, _11024_, _11249_);
  and (_19013_, _19012_, _11023_);
  or (_19015_, _19013_, _19011_);
  nand (_19016_, _11021_, _11291_);
  and (_19017_, _19016_, _09056_);
  and (_19018_, _19017_, _19015_);
  and (_19019_, _15350_, _07939_);
  or (_19020_, _19019_, _18758_);
  and (_19021_, _19020_, _06366_);
  or (_19022_, _19021_, _14283_);
  or (_19023_, _19022_, _19018_);
  and (_19024_, _19023_, _18749_);
  or (_19026_, _19024_, _11041_);
  and (_19027_, _11086_, _10610_);
  nor (_19028_, _19027_, _11087_);
  or (_19029_, _19028_, _11069_);
  and (_19030_, _19029_, _06541_);
  and (_19031_, _19030_, _19026_);
  nand (_19032_, _11114_, _10860_);
  nor (_19033_, _11115_, _06541_);
  and (_19034_, _19033_, _19032_);
  or (_19035_, _19034_, _11097_);
  or (_19037_, _19035_, _19031_);
  and (_19038_, _11142_, _10542_);
  nor (_19039_, _19038_, _11143_);
  or (_19040_, _19039_, _11127_);
  and (_19041_, _19040_, _11126_);
  and (_19042_, _19041_, _19037_);
  nand (_19043_, _11125_, \oc8051_golden_model_1.ACC [4]);
  nand (_19044_, _19043_, _12151_);
  or (_19045_, _19044_, _19042_);
  and (_19046_, _11232_, _11210_);
  nor (_19048_, _19046_, _11233_);
  or (_19049_, _19048_, _11203_);
  nor (_19050_, _11189_, _11166_);
  nor (_19051_, _19050_, _11190_);
  or (_19052_, _19051_, _11157_);
  and (_19053_, _19052_, _06285_);
  and (_19054_, _19053_, _19049_);
  and (_19055_, _19054_, _19045_);
  not (_19056_, _13012_);
  nor (_19057_, _11273_, _11250_);
  nor (_19059_, _19057_, _11274_);
  or (_19060_, _19059_, _11243_);
  and (_19061_, _19060_, _19056_);
  or (_19062_, _19061_, _19055_);
  and (_19063_, _11315_, _12600_);
  nor (_19064_, _11315_, _12600_);
  or (_19065_, _19064_, _11321_);
  or (_19066_, _19065_, _19063_);
  and (_19067_, _19066_, _11285_);
  and (_19068_, _19067_, _19062_);
  and (_19070_, _11284_, \oc8051_golden_model_1.ACC [4]);
  or (_19071_, _19070_, _06568_);
  or (_19072_, _19071_, _19068_);
  or (_19073_, _18814_, _06926_);
  and (_19074_, _19073_, _11331_);
  and (_19075_, _19074_, _19072_);
  nor (_19076_, _11338_, _10170_);
  or (_19077_, _19076_, _11339_);
  and (_19078_, _19077_, _11330_);
  or (_19079_, _19078_, _11335_);
  or (_19081_, _19079_, _19075_);
  nand (_19082_, _11335_, _10116_);
  and (_19083_, _19082_, _05928_);
  and (_19084_, _19083_, _19081_);
  and (_19085_, _18844_, _05927_);
  or (_19086_, _19085_, _06278_);
  or (_19087_, _19086_, _19084_);
  and (_19088_, _15532_, _07939_);
  or (_19089_, _19088_, _18758_);
  or (_19090_, _19089_, _06279_);
  and (_19092_, _19090_, _11354_);
  and (_19093_, _19092_, _19087_);
  nor (_19094_, _11364_, \oc8051_golden_model_1.ACC [5]);
  nor (_19095_, _19094_, _11365_);
  and (_19096_, _19095_, _11353_);
  or (_19097_, _19096_, _11360_);
  or (_19098_, _19097_, _19093_);
  nand (_19099_, _11360_, _10116_);
  and (_19100_, _19099_, _01347_);
  and (_19101_, _19100_, _19098_);
  or (_19103_, _19101_, _18746_);
  and (_43167_, _19103_, _42618_);
  nor (_19104_, _01347_, _10116_);
  or (_19105_, _11116_, _10893_);
  and (_19106_, _11117_, _06540_);
  and (_19107_, _19106_, _19105_);
  nand (_19108_, _11021_, _11288_);
  or (_19109_, _17401_, _11204_);
  or (_19110_, _11207_, _10502_);
  nor (_19111_, _07939_, _10116_);
  and (_19113_, _15657_, _07939_);
  or (_19114_, _19113_, _19111_);
  and (_19115_, _19114_, _10094_);
  nor (_19116_, _08142_, _10490_);
  or (_19117_, _19116_, _19111_);
  or (_19118_, _19117_, _07215_);
  or (_19119_, _09447_, _10170_);
  and (_19120_, _09447_, _10170_);
  or (_19121_, _18867_, _19120_);
  and (_19122_, _19121_, _19119_);
  nor (_19124_, _19122_, _11207_);
  and (_19125_, _19122_, _11207_);
  nor (_19126_, _19125_, _19124_);
  nor (_19127_, _18877_, _18871_);
  and (_19128_, _19127_, \oc8051_golden_model_1.PSW [7]);
  or (_19129_, _19128_, _19126_);
  nand (_19130_, _19128_, _19126_);
  and (_19131_, _19130_, _19129_);
  or (_19132_, _19131_, _10588_);
  nand (_19133_, _10744_, _08142_);
  nand (_19135_, _10756_, _08142_);
  nor (_19136_, _06781_, _10116_);
  and (_19137_, _06781_, _10116_);
  nor (_19138_, _19137_, _19136_);
  nand (_19139_, _19138_, _10755_);
  and (_19140_, _19139_, _10759_);
  and (_19141_, _19140_, _19135_);
  and (_19142_, _10758_, _09446_);
  or (_19143_, _19142_, _19141_);
  and (_19144_, _19143_, _10769_);
  and (_19146_, _15554_, _07939_);
  or (_19147_, _19146_, _19111_);
  and (_19148_, _19147_, _06341_);
  or (_19149_, _19148_, _10775_);
  or (_19150_, _19149_, _19144_);
  not (_19151_, _18819_);
  nor (_19152_, _19151_, _10789_);
  and (_19153_, _19151_, _10789_);
  or (_19154_, _19153_, _19152_);
  or (_19155_, _19154_, _10776_);
  and (_19157_, _19155_, _06466_);
  and (_19158_, _19157_, _19150_);
  nor (_19159_, _08636_, _10116_);
  and (_19160_, _15570_, _08636_);
  or (_19161_, _19160_, _19159_);
  and (_19162_, _19161_, _06272_);
  and (_19163_, _19117_, _06461_);
  or (_19164_, _19163_, _10744_);
  or (_19165_, _19164_, _19162_);
  or (_19166_, _19165_, _19158_);
  and (_19168_, _19166_, _19133_);
  or (_19169_, _19168_, _07174_);
  or (_19170_, _09446_, _07175_);
  and (_19171_, _19170_, _06465_);
  and (_19172_, _19171_, _19169_);
  nor (_19173_, _08144_, _06465_);
  or (_19174_, _19173_, _10811_);
  or (_19175_, _19174_, _19172_);
  nand (_19176_, _10811_, _10213_);
  and (_19177_, _19176_, _19175_);
  or (_19179_, _19177_, _06268_);
  and (_19180_, _15551_, _08636_);
  or (_19181_, _19180_, _19159_);
  or (_19182_, _19181_, _06269_);
  and (_19183_, _19182_, _06262_);
  and (_19184_, _19183_, _19179_);
  or (_19185_, _19159_, _15585_);
  and (_19186_, _19185_, _06261_);
  and (_19187_, _19186_, _19161_);
  or (_19188_, _19187_, _09531_);
  or (_19190_, _19188_, _19184_);
  nor (_19191_, _10046_, _10044_);
  nor (_19192_, _19191_, _10047_);
  or (_19193_, _19192_, _09537_);
  and (_19194_, _19193_, _10735_);
  and (_19195_, _19194_, _19190_);
  nand (_19196_, _08244_, \oc8051_golden_model_1.ACC [5]);
  nor (_19197_, _08244_, \oc8051_golden_model_1.ACC [5]);
  or (_19198_, _18780_, _19197_);
  and (_19199_, _19198_, _19196_);
  nor (_19201_, _19199_, _11163_);
  and (_19202_, _19199_, _11163_);
  nor (_19203_, _19202_, _19201_);
  nor (_19204_, _18790_, _18785_);
  and (_19205_, _19204_, \oc8051_golden_model_1.PSW [7]);
  or (_19206_, _19205_, _19203_);
  nand (_19207_, _19205_, _19203_);
  and (_19208_, _19207_, _10737_);
  and (_19209_, _19208_, _19206_);
  or (_19210_, _19209_, _10656_);
  or (_19212_, _19210_, _19195_);
  and (_19213_, _19212_, _06517_);
  and (_19214_, _19213_, _19132_);
  or (_19215_, _18885_, _14129_);
  and (_19216_, _19215_, _14128_);
  nor (_19217_, _19216_, _11247_);
  and (_19218_, _19216_, _11247_);
  nor (_19219_, _19218_, _19217_);
  nor (_19220_, _18895_, _18889_);
  and (_19221_, _19220_, \oc8051_golden_model_1.PSW [7]);
  nand (_19223_, _19221_, _19219_);
  or (_19224_, _19221_, _19219_);
  and (_19225_, _19224_, _06512_);
  and (_19226_, _19225_, _19223_);
  or (_19227_, _19226_, _19214_);
  and (_19228_, _19227_, _10517_);
  or (_19229_, _18763_, _14168_);
  and (_19230_, _19229_, _14167_);
  nor (_19231_, _19230_, _11289_);
  and (_19232_, _19230_, _11289_);
  nor (_19234_, _19232_, _19231_);
  nor (_19235_, _18774_, _18767_);
  and (_19236_, _19235_, \oc8051_golden_model_1.PSW [7]);
  or (_19237_, _19236_, _19234_);
  nand (_19238_, _19236_, _19234_);
  and (_19239_, _19238_, _10516_);
  and (_19240_, _19239_, _19237_);
  or (_19241_, _19240_, _10515_);
  or (_19242_, _19241_, _19228_);
  nand (_19243_, _06317_, _10515_);
  and (_19245_, _19243_, _06258_);
  and (_19246_, _19245_, _19242_);
  and (_19247_, _15602_, _08636_);
  or (_19248_, _19247_, _19159_);
  and (_19249_, _19248_, _06257_);
  or (_19250_, _19249_, _10080_);
  or (_19251_, _19250_, _19246_);
  and (_19252_, _19251_, _19118_);
  or (_19253_, _19252_, _07460_);
  and (_19254_, _09446_, _07939_);
  or (_19256_, _19111_, _07208_);
  or (_19257_, _19256_, _19254_);
  and (_19258_, _19257_, _05982_);
  and (_19259_, _19258_, _19253_);
  or (_19260_, _19259_, _19115_);
  and (_19261_, _19260_, _12172_);
  nor (_19262_, _06317_, _05975_);
  not (_19263_, _10122_);
  nor (_19264_, _19263_, _10117_);
  and (_19265_, _19264_, _05973_);
  and (_19267_, _19265_, _10093_);
  or (_19268_, _19267_, _19262_);
  or (_19269_, _19268_, _19261_);
  and (_19270_, _19269_, _06219_);
  and (_19271_, _15664_, _07939_);
  or (_19272_, _19271_, _19111_);
  and (_19273_, _19272_, _06218_);
  or (_19274_, _19273_, _10929_);
  or (_19275_, _19274_, _19270_);
  nand (_19276_, _10929_, _06317_);
  and (_19278_, _19276_, _17962_);
  and (_19279_, _19278_, _19275_);
  and (_19280_, _17965_, _11163_);
  or (_19281_, _19280_, _10506_);
  or (_19282_, _19281_, _19279_);
  or (_19283_, _11163_, _17969_);
  and (_19284_, _19283_, _18952_);
  and (_19285_, _19284_, _19282_);
  or (_19286_, _17511_, _11163_);
  and (_19287_, _19286_, _18286_);
  or (_19289_, _19287_, _19285_);
  or (_19290_, _17512_, _11163_);
  and (_19291_, _19290_, _17510_);
  and (_19292_, _19291_, _19289_);
  and (_19293_, _11163_, _06888_);
  or (_19294_, _19293_, _10948_);
  or (_19295_, _19294_, _19292_);
  and (_19296_, _19295_, _19110_);
  or (_19297_, _19296_, _06533_);
  or (_19298_, _11247_, _06534_);
  and (_19300_, _19298_, _10955_);
  and (_19301_, _19300_, _19297_);
  and (_19302_, _10954_, _11289_);
  or (_19303_, _19302_, _06369_);
  or (_19304_, _19303_, _19301_);
  and (_19305_, _15549_, _07939_);
  or (_19306_, _19305_, _19111_);
  or (_19307_, _19306_, _07237_);
  and (_19308_, _19307_, _19304_);
  or (_19309_, _19308_, _06536_);
  or (_19311_, _19111_, _07240_);
  and (_19312_, _19311_, _10986_);
  and (_19313_, _19312_, _19309_);
  and (_19314_, _10987_, _11160_);
  or (_19315_, _19314_, _10983_);
  or (_19316_, _19315_, _19313_);
  and (_19317_, _19316_, _19109_);
  or (_19318_, _19317_, _06542_);
  or (_19319_, _11244_, _06543_);
  and (_19320_, _19319_, _10497_);
  and (_19322_, _19320_, _19318_);
  and (_19323_, _11286_, _10496_);
  or (_19324_, _19323_, _19322_);
  and (_19325_, _19324_, _07242_);
  and (_19326_, _10998_, _07043_);
  nand (_19327_, _19272_, _06375_);
  or (_19328_, _19327_, _11246_);
  nand (_19329_, _19328_, _19326_);
  or (_19330_, _19329_, _19325_);
  or (_19331_, _19326_, _11162_);
  and (_19333_, _19331_, _11009_);
  and (_19334_, _19333_, _19330_);
  and (_19335_, _11008_, _11162_);
  or (_19336_, _19335_, _11014_);
  or (_19337_, _19336_, _19334_);
  or (_19338_, _11013_, _11205_);
  and (_19339_, _19338_, _06531_);
  and (_19340_, _19339_, _19337_);
  nand (_19341_, _11024_, _11246_);
  and (_19342_, _19341_, _11023_);
  or (_19344_, _19342_, _19340_);
  and (_19345_, _19344_, _19108_);
  or (_19346_, _19345_, _06366_);
  and (_19347_, _15546_, _07939_);
  or (_19348_, _19111_, _09056_);
  or (_19349_, _19348_, _19347_);
  and (_19350_, _19349_, _11037_);
  and (_19351_, _19350_, _19346_);
  nor (_19352_, _11060_, _10722_);
  nor (_19353_, _19352_, _11061_);
  and (_19355_, _19353_, _14283_);
  or (_19356_, _19355_, _11041_);
  or (_19357_, _19356_, _19351_);
  or (_19358_, _11088_, _10649_);
  and (_19359_, _19358_, _11089_);
  or (_19360_, _19359_, _11069_);
  and (_19361_, _19360_, _06541_);
  and (_19362_, _19361_, _19357_);
  or (_19363_, _19362_, _19107_);
  and (_19364_, _19363_, _11127_);
  or (_19366_, _11144_, _10579_);
  nor (_19367_, _11145_, _11127_);
  and (_19368_, _19367_, _19366_);
  or (_19369_, _19368_, _11125_);
  or (_19370_, _19369_, _19364_);
  nand (_19371_, _11125_, _10170_);
  and (_19372_, _19371_, _11157_);
  and (_19373_, _19372_, _19370_);
  nor (_19374_, _11191_, _11163_);
  nor (_19375_, _19374_, _11192_);
  and (_19377_, _19375_, _18059_);
  or (_19378_, _19377_, _11201_);
  or (_19379_, _19378_, _19373_);
  nor (_19380_, _11234_, _11207_);
  nor (_19381_, _19380_, _11235_);
  or (_19382_, _19381_, _11203_);
  and (_19383_, _19382_, _06285_);
  and (_19384_, _19383_, _19379_);
  or (_19385_, _11275_, _11247_);
  and (_19386_, _19385_, _11276_);
  or (_19388_, _19386_, _11243_);
  and (_19389_, _19388_, _19056_);
  or (_19390_, _19389_, _19384_);
  or (_19391_, _11317_, _11289_);
  and (_19392_, _19391_, _11318_);
  or (_19393_, _19392_, _11321_);
  and (_19394_, _19393_, _11285_);
  and (_19395_, _19394_, _19390_);
  and (_19396_, _11284_, \oc8051_golden_model_1.ACC [5]);
  or (_19397_, _19396_, _06568_);
  or (_19399_, _19397_, _19395_);
  or (_19400_, _19147_, _06926_);
  and (_19401_, _19400_, _11331_);
  and (_19402_, _19401_, _19399_);
  nor (_19403_, _11339_, _10116_);
  or (_19404_, _19403_, _11340_);
  and (_19405_, _19404_, _11330_);
  or (_19406_, _19405_, _11335_);
  or (_19407_, _19406_, _19402_);
  nand (_19408_, _11335_, _08572_);
  and (_19410_, _19408_, _05928_);
  and (_19411_, _19410_, _19407_);
  and (_19412_, _19181_, _05927_);
  or (_19413_, _19412_, _06278_);
  or (_19414_, _19413_, _19411_);
  and (_19415_, _15734_, _07939_);
  or (_19416_, _19415_, _19111_);
  or (_19417_, _19416_, _06279_);
  and (_19418_, _19417_, _11354_);
  and (_19419_, _19418_, _19414_);
  nor (_19421_, _11365_, \oc8051_golden_model_1.ACC [6]);
  nor (_19422_, _19421_, _11366_);
  and (_19423_, _19422_, _11353_);
  or (_19424_, _19423_, _11360_);
  or (_19425_, _19424_, _19419_);
  nand (_19426_, _11360_, _08572_);
  and (_19427_, _19426_, _01347_);
  and (_19428_, _19427_, _19425_);
  or (_19429_, _19428_, _19104_);
  and (_43168_, _19429_, _42618_);
  not (_19431_, \oc8051_golden_model_1.PCON [0]);
  nor (_19432_, _01347_, _19431_);
  nand (_19433_, _11263_, _07951_);
  nor (_19434_, _07951_, _19431_);
  nor (_19435_, _19434_, _07234_);
  nand (_19436_, _19435_, _19433_);
  and (_19437_, _07951_, _07133_);
  or (_19438_, _19437_, _19434_);
  or (_19439_, _19438_, _07215_);
  nor (_19440_, _08390_, _11380_);
  or (_19442_, _19440_, _19434_);
  or (_19443_, _19442_, _07151_);
  and (_19444_, _07951_, \oc8051_golden_model_1.ACC [0]);
  or (_19445_, _19444_, _19434_);
  and (_19446_, _19445_, _07141_);
  nor (_19447_, _07141_, _19431_);
  or (_19448_, _19447_, _06341_);
  or (_19449_, _19448_, _19446_);
  and (_19450_, _19449_, _07166_);
  and (_19451_, _19450_, _19443_);
  and (_19453_, _19438_, _06461_);
  or (_19454_, _19453_, _19451_);
  and (_19455_, _19454_, _06465_);
  and (_19456_, _19445_, _06464_);
  or (_19457_, _19456_, _10080_);
  or (_19458_, _19457_, _19455_);
  and (_19459_, _19458_, _19439_);
  or (_19460_, _19459_, _07460_);
  and (_19461_, _09392_, _07951_);
  or (_19462_, _19434_, _07208_);
  or (_19464_, _19462_, _19461_);
  and (_19465_, _19464_, _19460_);
  or (_19466_, _19465_, _10094_);
  and (_19467_, _14467_, _07951_);
  or (_19468_, _19434_, _05982_);
  or (_19469_, _19468_, _19467_);
  and (_19470_, _19469_, _06219_);
  and (_19471_, _19470_, _19466_);
  and (_19472_, _07951_, _08954_);
  or (_19473_, _19472_, _19434_);
  and (_19475_, _19473_, _06218_);
  or (_19476_, _19475_, _06369_);
  or (_19477_, _19476_, _19471_);
  and (_19478_, _14366_, _07951_);
  or (_19479_, _19478_, _19434_);
  or (_19480_, _19479_, _07237_);
  and (_19481_, _19480_, _07240_);
  and (_19482_, _19481_, _19477_);
  nor (_19483_, _12580_, _11380_);
  or (_19484_, _19483_, _19434_);
  and (_19486_, _19433_, _06536_);
  and (_19487_, _19486_, _19484_);
  or (_19488_, _19487_, _19482_);
  and (_19489_, _19488_, _07242_);
  nand (_19490_, _19473_, _06375_);
  nor (_19491_, _19490_, _19440_);
  or (_19492_, _19491_, _06545_);
  or (_19493_, _19492_, _19489_);
  and (_19494_, _19493_, _19436_);
  or (_19495_, _19494_, _06366_);
  and (_19497_, _14363_, _07951_);
  or (_19498_, _19497_, _19434_);
  or (_19499_, _19498_, _09056_);
  and (_19500_, _19499_, _09061_);
  and (_19501_, _19500_, _19495_);
  not (_19502_, _06661_);
  and (_19503_, _19484_, _06528_);
  or (_19504_, _19503_, _19502_);
  or (_19505_, _19504_, _19501_);
  or (_19506_, _19442_, _06661_);
  and (_19508_, _19506_, _01347_);
  and (_19509_, _19508_, _19505_);
  or (_19510_, _19509_, _19432_);
  and (_43170_, _19510_, _42618_);
  not (_19511_, \oc8051_golden_model_1.PCON [1]);
  nor (_19512_, _01347_, _19511_);
  nand (_19513_, _07951_, _07038_);
  or (_19514_, _07951_, \oc8051_golden_model_1.PCON [1]);
  and (_19515_, _19514_, _06218_);
  and (_19516_, _19515_, _19513_);
  nor (_19518_, _07951_, _19511_);
  nor (_19519_, _11380_, _07357_);
  or (_19520_, _19519_, _19518_);
  or (_19521_, _19520_, _07215_);
  and (_19522_, _14562_, _07951_);
  not (_19523_, _19522_);
  and (_19524_, _19523_, _19514_);
  or (_19525_, _19524_, _07151_);
  and (_19526_, _07951_, \oc8051_golden_model_1.ACC [1]);
  or (_19527_, _19526_, _19518_);
  and (_19529_, _19527_, _07141_);
  nor (_19530_, _07141_, _19511_);
  or (_19531_, _19530_, _06341_);
  or (_19532_, _19531_, _19529_);
  and (_19533_, _19532_, _07166_);
  and (_19534_, _19533_, _19525_);
  and (_19535_, _19520_, _06461_);
  or (_19536_, _19535_, _19534_);
  and (_19537_, _19536_, _06465_);
  and (_19538_, _19527_, _06464_);
  or (_19540_, _19538_, _10080_);
  or (_19541_, _19540_, _19537_);
  and (_19542_, _19541_, _19521_);
  or (_19543_, _19542_, _07460_);
  and (_19544_, _09451_, _07951_);
  or (_19545_, _19518_, _07208_);
  or (_19546_, _19545_, _19544_);
  and (_19547_, _19546_, _05982_);
  and (_19548_, _19547_, _19543_);
  or (_19549_, _14653_, _11380_);
  and (_19551_, _19514_, _10094_);
  and (_19552_, _19551_, _19549_);
  or (_19553_, _19552_, _19548_);
  and (_19554_, _19553_, _06219_);
  or (_19555_, _19554_, _19516_);
  and (_19556_, _19555_, _07237_);
  or (_19557_, _14668_, _11380_);
  and (_19558_, _19514_, _06369_);
  and (_19559_, _19558_, _19557_);
  or (_19560_, _19559_, _06536_);
  or (_19562_, _19560_, _19556_);
  nor (_19563_, _11261_, _11380_);
  or (_19564_, _19563_, _19518_);
  nand (_19565_, _11260_, _07951_);
  and (_19566_, _19565_, _19564_);
  or (_19567_, _19566_, _07240_);
  and (_19568_, _19567_, _07242_);
  and (_19569_, _19568_, _19562_);
  or (_19570_, _14666_, _11380_);
  and (_19571_, _19514_, _06375_);
  and (_19573_, _19571_, _19570_);
  or (_19574_, _19573_, _06545_);
  or (_19575_, _19574_, _19569_);
  nor (_19576_, _19518_, _07234_);
  nand (_19577_, _19576_, _19565_);
  and (_19578_, _19577_, _09056_);
  and (_19579_, _19578_, _19575_);
  or (_19580_, _19513_, _08341_);
  and (_19581_, _19514_, _06366_);
  and (_19582_, _19581_, _19580_);
  or (_19584_, _19582_, _06528_);
  or (_19585_, _19584_, _19579_);
  or (_19586_, _19564_, _09061_);
  and (_19587_, _19586_, _06926_);
  and (_19588_, _19587_, _19585_);
  and (_19589_, _19524_, _06568_);
  or (_19590_, _19589_, _06278_);
  or (_19591_, _19590_, _19588_);
  or (_19592_, _19518_, _06279_);
  or (_19593_, _19592_, _19522_);
  and (_19595_, _19593_, _01347_);
  and (_19596_, _19595_, _19591_);
  or (_19597_, _19596_, _19512_);
  and (_43171_, _19597_, _42618_);
  not (_19598_, \oc8051_golden_model_1.PCON [2]);
  nor (_19599_, _01347_, _19598_);
  nor (_19600_, _07951_, _19598_);
  nor (_19601_, _11380_, _07776_);
  or (_19602_, _19601_, _19600_);
  or (_19603_, _19602_, _07215_);
  and (_19605_, _14770_, _07951_);
  or (_19606_, _19605_, _19600_);
  and (_19607_, _19606_, _06341_);
  nor (_19608_, _07141_, _19598_);
  and (_19609_, _07951_, \oc8051_golden_model_1.ACC [2]);
  or (_19610_, _19609_, _19600_);
  and (_19611_, _19610_, _07141_);
  or (_19612_, _19611_, _19608_);
  and (_19613_, _19612_, _07151_);
  or (_19614_, _19613_, _06461_);
  or (_19616_, _19614_, _19607_);
  or (_19617_, _19602_, _07166_);
  and (_19618_, _19617_, _06465_);
  and (_19619_, _19618_, _19616_);
  and (_19620_, _19610_, _06464_);
  or (_19621_, _19620_, _10080_);
  or (_19622_, _19621_, _19619_);
  and (_19623_, _19622_, _19603_);
  or (_19624_, _19623_, _07460_);
  and (_19625_, _09450_, _07951_);
  or (_19627_, _19600_, _07208_);
  or (_19628_, _19627_, _19625_);
  and (_19629_, _19628_, _19624_);
  or (_19630_, _19629_, _10094_);
  and (_19631_, _14859_, _07951_);
  or (_19632_, _19600_, _05982_);
  or (_19633_, _19632_, _19631_);
  and (_19634_, _19633_, _06219_);
  and (_19635_, _19634_, _19630_);
  and (_19636_, _07951_, _08973_);
  or (_19638_, _19636_, _19600_);
  and (_19639_, _19638_, _06218_);
  or (_19640_, _19639_, _06369_);
  or (_19641_, _19640_, _19635_);
  and (_19642_, _14751_, _07951_);
  or (_19643_, _19642_, _19600_);
  or (_19644_, _19643_, _07237_);
  and (_19645_, _19644_, _07240_);
  and (_19646_, _19645_, _19641_);
  and (_19647_, _11259_, _07951_);
  or (_19649_, _19647_, _19600_);
  and (_19650_, _19649_, _06536_);
  or (_19651_, _19650_, _19646_);
  and (_19652_, _19651_, _07242_);
  or (_19653_, _19600_, _08440_);
  and (_19654_, _19638_, _06375_);
  and (_19655_, _19654_, _19653_);
  or (_19656_, _19655_, _19652_);
  and (_19657_, _19656_, _07234_);
  and (_19658_, _19610_, _06545_);
  and (_19660_, _19658_, _19653_);
  or (_19661_, _19660_, _06366_);
  or (_19662_, _19661_, _19657_);
  and (_19663_, _14748_, _07951_);
  or (_19664_, _19600_, _09056_);
  or (_19665_, _19664_, _19663_);
  and (_19666_, _19665_, _09061_);
  and (_19667_, _19666_, _19662_);
  nor (_19668_, _11258_, _11380_);
  or (_19669_, _19668_, _19600_);
  and (_19671_, _19669_, _06528_);
  or (_19672_, _19671_, _19667_);
  and (_19673_, _19672_, _06926_);
  and (_19674_, _19606_, _06568_);
  or (_19675_, _19674_, _06278_);
  or (_19676_, _19675_, _19673_);
  and (_19677_, _14926_, _07951_);
  or (_19678_, _19600_, _06279_);
  or (_19679_, _19678_, _19677_);
  and (_19680_, _19679_, _01347_);
  and (_19682_, _19680_, _19676_);
  or (_19683_, _19682_, _19599_);
  and (_43172_, _19683_, _42618_);
  not (_19684_, \oc8051_golden_model_1.PCON [3]);
  nor (_19685_, _01347_, _19684_);
  nor (_19686_, _07951_, _19684_);
  and (_19687_, _14953_, _07951_);
  or (_19688_, _19687_, _19686_);
  or (_19689_, _19688_, _07151_);
  and (_19690_, _07951_, \oc8051_golden_model_1.ACC [3]);
  or (_19692_, _19690_, _19686_);
  and (_19693_, _19692_, _07141_);
  nor (_19694_, _07141_, _19684_);
  or (_19695_, _19694_, _06341_);
  or (_19696_, _19695_, _19693_);
  and (_19697_, _19696_, _07166_);
  and (_19698_, _19697_, _19689_);
  nor (_19699_, _11380_, _07594_);
  or (_19700_, _19699_, _19686_);
  and (_19701_, _19700_, _06461_);
  or (_19703_, _19701_, _19698_);
  and (_19704_, _19703_, _06465_);
  and (_19705_, _19692_, _06464_);
  or (_19706_, _19705_, _10080_);
  or (_19707_, _19706_, _19704_);
  or (_19708_, _19700_, _07215_);
  and (_19709_, _19708_, _07208_);
  and (_19710_, _19709_, _19707_);
  and (_19711_, _09449_, _07951_);
  or (_19712_, _19711_, _19686_);
  and (_19714_, _19712_, _07460_);
  or (_19715_, _19714_, _10094_);
  or (_19716_, _19715_, _19710_);
  and (_19717_, _15048_, _07951_);
  or (_19718_, _19686_, _05982_);
  or (_19719_, _19718_, _19717_);
  and (_19720_, _19719_, _06219_);
  and (_19721_, _19720_, _19716_);
  and (_19722_, _07951_, _08930_);
  or (_19723_, _19722_, _19686_);
  and (_19725_, _19723_, _06218_);
  or (_19726_, _19725_, _06369_);
  or (_19727_, _19726_, _19721_);
  and (_19728_, _14943_, _07951_);
  or (_19729_, _19728_, _19686_);
  or (_19730_, _19729_, _07237_);
  and (_19731_, _19730_, _07240_);
  and (_19732_, _19731_, _19727_);
  and (_19733_, _12577_, _07951_);
  or (_19734_, _19733_, _19686_);
  and (_19736_, _19734_, _06536_);
  or (_19737_, _19736_, _19732_);
  and (_19738_, _19737_, _07242_);
  or (_19739_, _19686_, _08292_);
  and (_19740_, _19723_, _06375_);
  and (_19741_, _19740_, _19739_);
  or (_19742_, _19741_, _19738_);
  and (_19743_, _19742_, _07234_);
  and (_19744_, _19692_, _06545_);
  and (_19745_, _19744_, _19739_);
  or (_19747_, _19745_, _06366_);
  or (_19748_, _19747_, _19743_);
  and (_19749_, _14940_, _07951_);
  or (_19750_, _19686_, _09056_);
  or (_19751_, _19750_, _19749_);
  and (_19752_, _19751_, _09061_);
  and (_19753_, _19752_, _19748_);
  nor (_19754_, _11256_, _11380_);
  or (_19755_, _19754_, _19686_);
  and (_19756_, _19755_, _06528_);
  or (_19758_, _19756_, _19753_);
  and (_19759_, _19758_, _06926_);
  and (_19760_, _19688_, _06568_);
  or (_19761_, _19760_, _06278_);
  or (_19762_, _19761_, _19759_);
  and (_19763_, _15128_, _07951_);
  or (_19764_, _19686_, _06279_);
  or (_19765_, _19764_, _19763_);
  and (_19766_, _19765_, _01347_);
  and (_19767_, _19766_, _19762_);
  or (_19770_, _19767_, _19685_);
  and (_43173_, _19770_, _42618_);
  not (_19771_, \oc8051_golden_model_1.PCON [4]);
  nor (_19772_, _01347_, _19771_);
  nor (_19773_, _07951_, _19771_);
  nor (_19774_, _08541_, _11380_);
  or (_19775_, _19774_, _19773_);
  or (_19776_, _19775_, _07215_);
  and (_19777_, _15162_, _07951_);
  or (_19778_, _19777_, _19773_);
  or (_19781_, _19778_, _07151_);
  and (_19782_, _07951_, \oc8051_golden_model_1.ACC [4]);
  or (_19783_, _19782_, _19773_);
  and (_19784_, _19783_, _07141_);
  nor (_19785_, _07141_, _19771_);
  or (_19786_, _19785_, _06341_);
  or (_19787_, _19786_, _19784_);
  and (_19788_, _19787_, _07166_);
  and (_19789_, _19788_, _19781_);
  and (_19790_, _19775_, _06461_);
  or (_19793_, _19790_, _19789_);
  and (_19794_, _19793_, _06465_);
  and (_19795_, _19783_, _06464_);
  or (_19796_, _19795_, _10080_);
  or (_19797_, _19796_, _19794_);
  and (_19798_, _19797_, _19776_);
  or (_19799_, _19798_, _07460_);
  and (_19800_, _09448_, _07951_);
  or (_19801_, _19773_, _07208_);
  or (_19802_, _19801_, _19800_);
  and (_19805_, _19802_, _19799_);
  or (_19806_, _19805_, _10094_);
  and (_19807_, _15254_, _07951_);
  or (_19808_, _19773_, _05982_);
  or (_19809_, _19808_, _19807_);
  and (_19810_, _19809_, _06219_);
  and (_19811_, _19810_, _19806_);
  and (_19812_, _08959_, _07951_);
  or (_19813_, _19812_, _19773_);
  and (_19814_, _19813_, _06218_);
  or (_19817_, _19814_, _06369_);
  or (_19818_, _19817_, _19811_);
  and (_19819_, _15269_, _07951_);
  or (_19820_, _19819_, _19773_);
  or (_19821_, _19820_, _07237_);
  and (_19822_, _19821_, _07240_);
  and (_19823_, _19822_, _19818_);
  and (_19824_, _11254_, _07951_);
  or (_19825_, _19824_, _19773_);
  and (_19826_, _19825_, _06536_);
  or (_19829_, _19826_, _19823_);
  and (_19830_, _19829_, _07242_);
  or (_19831_, _19773_, _08544_);
  and (_19832_, _19813_, _06375_);
  and (_19833_, _19832_, _19831_);
  or (_19834_, _19833_, _19830_);
  and (_19835_, _19834_, _07234_);
  and (_19836_, _19783_, _06545_);
  and (_19837_, _19836_, _19831_);
  or (_19838_, _19837_, _06366_);
  or (_19841_, _19838_, _19835_);
  and (_19842_, _15266_, _07951_);
  or (_19843_, _19773_, _09056_);
  or (_19844_, _19843_, _19842_);
  and (_19845_, _19844_, _09061_);
  and (_19846_, _19845_, _19841_);
  nor (_19847_, _11253_, _11380_);
  or (_19848_, _19847_, _19773_);
  and (_19849_, _19848_, _06528_);
  or (_19850_, _19849_, _19846_);
  and (_19852_, _19850_, _06926_);
  and (_19853_, _19778_, _06568_);
  or (_19854_, _19853_, _06278_);
  or (_19855_, _19854_, _19852_);
  and (_19856_, _15329_, _07951_);
  or (_19857_, _19773_, _06279_);
  or (_19858_, _19857_, _19856_);
  and (_19859_, _19858_, _01347_);
  and (_19860_, _19859_, _19855_);
  or (_19861_, _19860_, _19772_);
  and (_43174_, _19861_, _42618_);
  not (_19863_, \oc8051_golden_model_1.PCON [5]);
  nor (_19864_, _01347_, _19863_);
  nor (_19865_, _07951_, _19863_);
  nor (_19866_, _08244_, _11380_);
  or (_19867_, _19866_, _19865_);
  or (_19868_, _19867_, _07215_);
  and (_19869_, _15358_, _07951_);
  or (_19870_, _19869_, _19865_);
  or (_19871_, _19870_, _07151_);
  and (_19873_, _07951_, \oc8051_golden_model_1.ACC [5]);
  or (_19874_, _19873_, _19865_);
  and (_19875_, _19874_, _07141_);
  nor (_19876_, _07141_, _19863_);
  or (_19877_, _19876_, _06341_);
  or (_19878_, _19877_, _19875_);
  and (_19879_, _19878_, _07166_);
  and (_19880_, _19879_, _19871_);
  and (_19881_, _19867_, _06461_);
  or (_19882_, _19881_, _19880_);
  and (_19884_, _19882_, _06465_);
  and (_19885_, _19874_, _06464_);
  or (_19886_, _19885_, _10080_);
  or (_19887_, _19886_, _19884_);
  and (_19888_, _19887_, _19868_);
  or (_19889_, _19888_, _07460_);
  and (_19890_, _09447_, _07951_);
  or (_19891_, _19865_, _07208_);
  or (_19892_, _19891_, _19890_);
  and (_19893_, _19892_, _05982_);
  and (_19895_, _19893_, _19889_);
  and (_19896_, _15459_, _07951_);
  or (_19897_, _19896_, _19865_);
  and (_19898_, _19897_, _10094_);
  or (_19899_, _19898_, _06218_);
  or (_19900_, _19899_, _19895_);
  and (_19901_, _08946_, _07951_);
  or (_19902_, _19901_, _19865_);
  or (_19903_, _19902_, _06219_);
  and (_19904_, _19903_, _19900_);
  or (_19906_, _19904_, _06369_);
  and (_19907_, _15353_, _07951_);
  or (_19908_, _19907_, _19865_);
  or (_19909_, _19908_, _07237_);
  and (_19910_, _19909_, _07240_);
  and (_19911_, _19910_, _19906_);
  and (_19912_, _11250_, _07951_);
  or (_19913_, _19912_, _19865_);
  and (_19914_, _19913_, _06536_);
  or (_19915_, _19914_, _19911_);
  and (_19917_, _19915_, _07242_);
  or (_19918_, _19865_, _08247_);
  and (_19919_, _19902_, _06375_);
  and (_19920_, _19919_, _19918_);
  or (_19921_, _19920_, _19917_);
  and (_19922_, _19921_, _07234_);
  and (_19923_, _19874_, _06545_);
  and (_19924_, _19923_, _19918_);
  or (_19925_, _19924_, _06366_);
  or (_19926_, _19925_, _19922_);
  and (_19928_, _15350_, _07951_);
  or (_19929_, _19865_, _09056_);
  or (_19930_, _19929_, _19928_);
  and (_19931_, _19930_, _09061_);
  and (_19932_, _19931_, _19926_);
  nor (_19933_, _11249_, _11380_);
  or (_19934_, _19933_, _19865_);
  and (_19935_, _19934_, _06528_);
  or (_19936_, _19935_, _19932_);
  and (_19937_, _19936_, _06926_);
  and (_19939_, _19870_, _06568_);
  or (_19940_, _19939_, _06278_);
  or (_19941_, _19940_, _19937_);
  and (_19942_, _15532_, _07951_);
  or (_19943_, _19865_, _06279_);
  or (_19944_, _19943_, _19942_);
  and (_19945_, _19944_, _01347_);
  and (_19946_, _19945_, _19941_);
  or (_19947_, _19946_, _19864_);
  and (_43175_, _19947_, _42618_);
  not (_19949_, \oc8051_golden_model_1.PCON [6]);
  nor (_19950_, _01347_, _19949_);
  nor (_19951_, _07951_, _19949_);
  nor (_19952_, _08142_, _11380_);
  or (_19953_, _19952_, _19951_);
  or (_19954_, _19953_, _07215_);
  and (_19955_, _15554_, _07951_);
  or (_19956_, _19955_, _19951_);
  or (_19957_, _19956_, _07151_);
  and (_19958_, _07951_, \oc8051_golden_model_1.ACC [6]);
  or (_19960_, _19958_, _19951_);
  and (_19961_, _19960_, _07141_);
  nor (_19962_, _07141_, _19949_);
  or (_19963_, _19962_, _06341_);
  or (_19964_, _19963_, _19961_);
  and (_19965_, _19964_, _07166_);
  and (_19966_, _19965_, _19957_);
  and (_19967_, _19953_, _06461_);
  or (_19968_, _19967_, _19966_);
  and (_19969_, _19968_, _06465_);
  and (_19971_, _19960_, _06464_);
  or (_19972_, _19971_, _10080_);
  or (_19973_, _19972_, _19969_);
  and (_19974_, _19973_, _19954_);
  or (_19975_, _19974_, _07460_);
  and (_19976_, _09446_, _07951_);
  or (_19977_, _19951_, _07208_);
  or (_19978_, _19977_, _19976_);
  and (_19979_, _19978_, _05982_);
  and (_19980_, _19979_, _19975_);
  and (_19982_, _15657_, _07951_);
  or (_19983_, _19982_, _19951_);
  and (_19984_, _19983_, _10094_);
  or (_19985_, _19984_, _06218_);
  or (_19986_, _19985_, _19980_);
  and (_19987_, _15664_, _07951_);
  or (_19988_, _19987_, _19951_);
  or (_19989_, _19988_, _06219_);
  and (_19990_, _19989_, _19986_);
  or (_19991_, _19990_, _06369_);
  and (_19993_, _15549_, _07951_);
  or (_19994_, _19993_, _19951_);
  or (_19995_, _19994_, _07237_);
  and (_19996_, _19995_, _07240_);
  and (_19997_, _19996_, _19991_);
  and (_19998_, _11247_, _07951_);
  or (_19999_, _19998_, _19951_);
  and (_20000_, _19999_, _06536_);
  or (_20001_, _20000_, _19997_);
  and (_20002_, _20001_, _07242_);
  or (_20004_, _19951_, _08145_);
  and (_20005_, _19988_, _06375_);
  and (_20006_, _20005_, _20004_);
  or (_20007_, _20006_, _20002_);
  and (_20008_, _20007_, _07234_);
  and (_20009_, _19960_, _06545_);
  and (_20010_, _20009_, _20004_);
  or (_20011_, _20010_, _06366_);
  or (_20012_, _20011_, _20008_);
  and (_20013_, _15546_, _07951_);
  or (_20015_, _19951_, _09056_);
  or (_20016_, _20015_, _20013_);
  and (_20017_, _20016_, _09061_);
  and (_20018_, _20017_, _20012_);
  nor (_20019_, _11246_, _11380_);
  or (_20020_, _20019_, _19951_);
  and (_20021_, _20020_, _06528_);
  or (_20022_, _20021_, _20018_);
  and (_20023_, _20022_, _06926_);
  and (_20024_, _19956_, _06568_);
  or (_20026_, _20024_, _06278_);
  or (_20027_, _20026_, _20023_);
  and (_20028_, _15734_, _07951_);
  or (_20029_, _19951_, _06279_);
  or (_20030_, _20029_, _20028_);
  and (_20031_, _20030_, _01347_);
  and (_20032_, _20031_, _20027_);
  or (_20033_, _20032_, _19950_);
  and (_43176_, _20033_, _42618_);
  not (_20034_, \oc8051_golden_model_1.TMOD [0]);
  nor (_20036_, _01347_, _20034_);
  nand (_20037_, _11263_, _07914_);
  nor (_20038_, _07914_, _20034_);
  nor (_20039_, _20038_, _07234_);
  nand (_20040_, _20039_, _20037_);
  and (_20041_, _07914_, _07133_);
  or (_20042_, _20041_, _20038_);
  or (_20043_, _20042_, _07215_);
  nor (_20044_, _08390_, _11457_);
  or (_20045_, _20044_, _20038_);
  or (_20047_, _20045_, _07151_);
  and (_20048_, _07914_, \oc8051_golden_model_1.ACC [0]);
  or (_20049_, _20048_, _20038_);
  and (_20050_, _20049_, _07141_);
  nor (_20051_, _07141_, _20034_);
  or (_20052_, _20051_, _06341_);
  or (_20053_, _20052_, _20050_);
  and (_20054_, _20053_, _07166_);
  and (_20055_, _20054_, _20047_);
  and (_20056_, _20042_, _06461_);
  or (_20058_, _20056_, _20055_);
  and (_20059_, _20058_, _06465_);
  and (_20060_, _20049_, _06464_);
  or (_20061_, _20060_, _10080_);
  or (_20062_, _20061_, _20059_);
  and (_20063_, _20062_, _20043_);
  or (_20064_, _20063_, _07460_);
  and (_20065_, _09392_, _07914_);
  or (_20066_, _20038_, _07208_);
  or (_20067_, _20066_, _20065_);
  and (_20069_, _20067_, _20064_);
  or (_20070_, _20069_, _10094_);
  and (_20071_, _14467_, _07914_);
  or (_20072_, _20038_, _05982_);
  or (_20073_, _20072_, _20071_);
  and (_20074_, _20073_, _06219_);
  and (_20075_, _20074_, _20070_);
  and (_20076_, _07914_, _08954_);
  or (_20077_, _20076_, _20038_);
  and (_20078_, _20077_, _06218_);
  or (_20080_, _20078_, _06369_);
  or (_20081_, _20080_, _20075_);
  and (_20082_, _14366_, _07914_);
  or (_20083_, _20082_, _20038_);
  or (_20084_, _20083_, _07237_);
  and (_20085_, _20084_, _07240_);
  and (_20086_, _20085_, _20081_);
  nor (_20087_, _12580_, _11457_);
  or (_20088_, _20087_, _20038_);
  and (_20089_, _20037_, _06536_);
  and (_20091_, _20089_, _20088_);
  or (_20092_, _20091_, _20086_);
  and (_20093_, _20092_, _07242_);
  nand (_20094_, _20077_, _06375_);
  nor (_20095_, _20094_, _20044_);
  or (_20096_, _20095_, _06545_);
  or (_20097_, _20096_, _20093_);
  and (_20098_, _20097_, _20040_);
  or (_20099_, _20098_, _06366_);
  and (_20100_, _14363_, _07914_);
  or (_20102_, _20038_, _09056_);
  or (_20103_, _20102_, _20100_);
  and (_20104_, _20103_, _09061_);
  and (_20105_, _20104_, _20099_);
  and (_20106_, _20088_, _06528_);
  or (_20107_, _20106_, _19502_);
  or (_20108_, _20107_, _20105_);
  or (_20109_, _20045_, _06661_);
  and (_20110_, _20109_, _01347_);
  and (_20111_, _20110_, _20108_);
  or (_20113_, _20111_, _20036_);
  and (_43178_, _20113_, _42618_);
  and (_20114_, _01351_, \oc8051_golden_model_1.TMOD [1]);
  nand (_20115_, _07914_, _07038_);
  or (_20116_, _07914_, \oc8051_golden_model_1.TMOD [1]);
  and (_20117_, _20116_, _06218_);
  and (_20118_, _20117_, _20115_);
  and (_20119_, _11457_, \oc8051_golden_model_1.TMOD [1]);
  nor (_20120_, _11457_, _07357_);
  or (_20121_, _20120_, _20119_);
  or (_20123_, _20121_, _07215_);
  and (_20124_, _14562_, _07914_);
  not (_20125_, _20124_);
  and (_20126_, _20125_, _20116_);
  or (_20127_, _20126_, _07151_);
  and (_20128_, _07914_, \oc8051_golden_model_1.ACC [1]);
  or (_20129_, _20128_, _20119_);
  and (_20130_, _20129_, _07141_);
  and (_20131_, _07142_, \oc8051_golden_model_1.TMOD [1]);
  or (_20132_, _20131_, _06341_);
  or (_20134_, _20132_, _20130_);
  and (_20135_, _20134_, _07166_);
  and (_20136_, _20135_, _20127_);
  and (_20137_, _20121_, _06461_);
  or (_20138_, _20137_, _20136_);
  and (_20139_, _20138_, _06465_);
  and (_20140_, _20129_, _06464_);
  or (_20141_, _20140_, _10080_);
  or (_20142_, _20141_, _20139_);
  and (_20143_, _20142_, _20123_);
  or (_20145_, _20143_, _07460_);
  and (_20146_, _09451_, _07914_);
  or (_20147_, _20119_, _07208_);
  or (_20148_, _20147_, _20146_);
  and (_20149_, _20148_, _05982_);
  and (_20150_, _20149_, _20145_);
  or (_20151_, _14653_, _11457_);
  and (_20152_, _20116_, _10094_);
  and (_20153_, _20152_, _20151_);
  or (_20154_, _20153_, _20150_);
  and (_20156_, _20154_, _06219_);
  or (_20157_, _20156_, _20118_);
  and (_20158_, _20157_, _07237_);
  or (_20159_, _14668_, _11457_);
  and (_20160_, _20116_, _06369_);
  and (_20161_, _20160_, _20159_);
  or (_20162_, _20161_, _06536_);
  or (_20163_, _20162_, _20158_);
  and (_20164_, _11262_, _07914_);
  or (_20165_, _20164_, _20119_);
  or (_20167_, _20165_, _07240_);
  and (_20168_, _20167_, _07242_);
  and (_20169_, _20168_, _20163_);
  or (_20170_, _14666_, _11457_);
  and (_20171_, _20116_, _06375_);
  and (_20172_, _20171_, _20170_);
  or (_20173_, _20172_, _06545_);
  or (_20174_, _20173_, _20169_);
  and (_20175_, _20128_, _08341_);
  or (_20176_, _20119_, _07234_);
  or (_20178_, _20176_, _20175_);
  and (_20179_, _20178_, _09056_);
  and (_20180_, _20179_, _20174_);
  or (_20181_, _20115_, _08341_);
  and (_20182_, _20116_, _06366_);
  and (_20183_, _20182_, _20181_);
  or (_20184_, _20183_, _06528_);
  or (_20185_, _20184_, _20180_);
  nor (_20186_, _11261_, _11457_);
  or (_20187_, _20186_, _20119_);
  or (_20189_, _20187_, _09061_);
  and (_20190_, _20189_, _06926_);
  and (_20191_, _20190_, _20185_);
  and (_20192_, _20126_, _06568_);
  or (_20193_, _20192_, _06278_);
  or (_20194_, _20193_, _20191_);
  or (_20195_, _20119_, _06279_);
  or (_20196_, _20195_, _20124_);
  and (_20197_, _20196_, _01347_);
  and (_20198_, _20197_, _20194_);
  or (_20200_, _20198_, _20114_);
  and (_43179_, _20200_, _42618_);
  and (_20201_, _01351_, \oc8051_golden_model_1.TMOD [2]);
  and (_20202_, _11457_, \oc8051_golden_model_1.TMOD [2]);
  and (_20203_, _09450_, _07914_);
  or (_20204_, _20203_, _20202_);
  and (_20205_, _20204_, _07460_);
  and (_20206_, _14770_, _07914_);
  or (_20207_, _20206_, _20202_);
  or (_20208_, _20207_, _07151_);
  and (_20210_, _07914_, \oc8051_golden_model_1.ACC [2]);
  or (_20211_, _20210_, _20202_);
  and (_20212_, _20211_, _07141_);
  and (_20213_, _07142_, \oc8051_golden_model_1.TMOD [2]);
  or (_20214_, _20213_, _06341_);
  or (_20215_, _20214_, _20212_);
  and (_20216_, _20215_, _07166_);
  and (_20217_, _20216_, _20208_);
  nor (_20218_, _11457_, _07776_);
  or (_20219_, _20218_, _20202_);
  and (_20221_, _20219_, _06461_);
  or (_20222_, _20221_, _20217_);
  and (_20223_, _20222_, _06465_);
  and (_20224_, _20211_, _06464_);
  or (_20225_, _20224_, _10080_);
  or (_20226_, _20225_, _20223_);
  or (_20227_, _20219_, _07215_);
  and (_20228_, _20227_, _07208_);
  and (_20229_, _20228_, _20226_);
  or (_20230_, _20229_, _10094_);
  or (_20232_, _20230_, _20205_);
  and (_20233_, _14859_, _07914_);
  or (_20234_, _20202_, _05982_);
  or (_20235_, _20234_, _20233_);
  and (_20236_, _20235_, _06219_);
  and (_20237_, _20236_, _20232_);
  and (_20238_, _07914_, _08973_);
  or (_20239_, _20238_, _20202_);
  and (_20240_, _20239_, _06218_);
  or (_20241_, _20240_, _06369_);
  or (_20243_, _20241_, _20237_);
  and (_20244_, _14751_, _07914_);
  or (_20245_, _20244_, _20202_);
  or (_20246_, _20245_, _07237_);
  and (_20247_, _20246_, _07240_);
  and (_20248_, _20247_, _20243_);
  and (_20249_, _11259_, _07914_);
  or (_20250_, _20249_, _20202_);
  and (_20251_, _20250_, _06536_);
  or (_20252_, _20251_, _20248_);
  and (_20254_, _20252_, _07242_);
  or (_20255_, _20202_, _08440_);
  and (_20256_, _20239_, _06375_);
  and (_20257_, _20256_, _20255_);
  or (_20258_, _20257_, _20254_);
  and (_20259_, _20258_, _07234_);
  and (_20260_, _20211_, _06545_);
  and (_20261_, _20260_, _20255_);
  or (_20262_, _20261_, _06366_);
  or (_20263_, _20262_, _20259_);
  and (_20265_, _14748_, _07914_);
  or (_20266_, _20202_, _09056_);
  or (_20267_, _20266_, _20265_);
  and (_20268_, _20267_, _09061_);
  and (_20269_, _20268_, _20263_);
  nor (_20270_, _11258_, _11457_);
  or (_20271_, _20270_, _20202_);
  and (_20272_, _20271_, _06528_);
  or (_20273_, _20272_, _20269_);
  and (_20274_, _20273_, _06926_);
  and (_20276_, _20207_, _06568_);
  or (_20277_, _20276_, _06278_);
  or (_20278_, _20277_, _20274_);
  and (_20279_, _14926_, _07914_);
  or (_20280_, _20202_, _06279_);
  or (_20281_, _20280_, _20279_);
  and (_20282_, _20281_, _01347_);
  and (_20283_, _20282_, _20278_);
  or (_20284_, _20283_, _20201_);
  and (_43180_, _20284_, _42618_);
  and (_20286_, _01351_, \oc8051_golden_model_1.TMOD [3]);
  and (_20287_, _11457_, \oc8051_golden_model_1.TMOD [3]);
  and (_20288_, _14953_, _07914_);
  or (_20289_, _20288_, _20287_);
  or (_20290_, _20289_, _07151_);
  and (_20291_, _07914_, \oc8051_golden_model_1.ACC [3]);
  or (_20292_, _20291_, _20287_);
  and (_20293_, _20292_, _07141_);
  and (_20294_, _07142_, \oc8051_golden_model_1.TMOD [3]);
  or (_20295_, _20294_, _06341_);
  or (_20297_, _20295_, _20293_);
  and (_20298_, _20297_, _07166_);
  and (_20299_, _20298_, _20290_);
  nor (_20300_, _11457_, _07594_);
  or (_20301_, _20300_, _20287_);
  and (_20302_, _20301_, _06461_);
  or (_20303_, _20302_, _20299_);
  and (_20304_, _20303_, _06465_);
  and (_20305_, _20292_, _06464_);
  or (_20306_, _20305_, _10080_);
  or (_20308_, _20306_, _20304_);
  or (_20309_, _20301_, _07215_);
  and (_20310_, _20309_, _07208_);
  and (_20311_, _20310_, _20308_);
  and (_20312_, _09449_, _07914_);
  or (_20313_, _20312_, _20287_);
  and (_20314_, _20313_, _07460_);
  or (_20315_, _20314_, _10094_);
  or (_20316_, _20315_, _20311_);
  and (_20317_, _15048_, _07914_);
  or (_20319_, _20287_, _05982_);
  or (_20320_, _20319_, _20317_);
  and (_20321_, _20320_, _06219_);
  and (_20322_, _20321_, _20316_);
  and (_20323_, _07914_, _08930_);
  or (_20324_, _20323_, _20287_);
  and (_20325_, _20324_, _06218_);
  or (_20326_, _20325_, _06369_);
  or (_20327_, _20326_, _20322_);
  and (_20328_, _14943_, _07914_);
  or (_20330_, _20328_, _20287_);
  or (_20331_, _20330_, _07237_);
  and (_20332_, _20331_, _07240_);
  and (_20333_, _20332_, _20327_);
  and (_20334_, _12577_, _07914_);
  or (_20335_, _20334_, _20287_);
  and (_20336_, _20335_, _06536_);
  or (_20337_, _20336_, _20333_);
  and (_20338_, _20337_, _07242_);
  or (_20339_, _20287_, _08292_);
  and (_20341_, _20324_, _06375_);
  and (_20342_, _20341_, _20339_);
  or (_20343_, _20342_, _20338_);
  and (_20344_, _20343_, _07234_);
  and (_20345_, _20292_, _06545_);
  and (_20346_, _20345_, _20339_);
  or (_20347_, _20346_, _06366_);
  or (_20348_, _20347_, _20344_);
  and (_20349_, _14940_, _07914_);
  or (_20350_, _20287_, _09056_);
  or (_20352_, _20350_, _20349_);
  and (_20353_, _20352_, _09061_);
  and (_20354_, _20353_, _20348_);
  nor (_20355_, _11256_, _11457_);
  or (_20356_, _20355_, _20287_);
  and (_20357_, _20356_, _06528_);
  or (_20358_, _20357_, _20354_);
  and (_20359_, _20358_, _06926_);
  and (_20360_, _20289_, _06568_);
  or (_20361_, _20360_, _06278_);
  or (_20363_, _20361_, _20359_);
  and (_20364_, _15128_, _07914_);
  or (_20365_, _20287_, _06279_);
  or (_20366_, _20365_, _20364_);
  and (_20367_, _20366_, _01347_);
  and (_20368_, _20367_, _20363_);
  or (_20369_, _20368_, _20286_);
  and (_43182_, _20369_, _42618_);
  and (_20370_, _01351_, \oc8051_golden_model_1.TMOD [4]);
  and (_20371_, _11457_, \oc8051_golden_model_1.TMOD [4]);
  nor (_20373_, _08541_, _11457_);
  or (_20374_, _20373_, _20371_);
  or (_20375_, _20374_, _07215_);
  and (_20376_, _15162_, _07914_);
  or (_20377_, _20376_, _20371_);
  or (_20378_, _20377_, _07151_);
  and (_20379_, _07914_, \oc8051_golden_model_1.ACC [4]);
  or (_20380_, _20379_, _20371_);
  and (_20381_, _20380_, _07141_);
  and (_20382_, _07142_, \oc8051_golden_model_1.TMOD [4]);
  or (_20384_, _20382_, _06341_);
  or (_20385_, _20384_, _20381_);
  and (_20386_, _20385_, _07166_);
  and (_20387_, _20386_, _20378_);
  and (_20388_, _20374_, _06461_);
  or (_20389_, _20388_, _20387_);
  and (_20390_, _20389_, _06465_);
  and (_20391_, _20380_, _06464_);
  or (_20392_, _20391_, _10080_);
  or (_20393_, _20392_, _20390_);
  and (_20395_, _20393_, _20375_);
  or (_20396_, _20395_, _07460_);
  and (_20397_, _09448_, _07914_);
  or (_20398_, _20371_, _07208_);
  or (_20399_, _20398_, _20397_);
  and (_20400_, _20399_, _20396_);
  or (_20401_, _20400_, _10094_);
  and (_20402_, _15254_, _07914_);
  or (_20403_, _20371_, _05982_);
  or (_20404_, _20403_, _20402_);
  and (_20406_, _20404_, _06219_);
  and (_20407_, _20406_, _20401_);
  and (_20408_, _08959_, _07914_);
  or (_20409_, _20408_, _20371_);
  and (_20410_, _20409_, _06218_);
  or (_20411_, _20410_, _06369_);
  or (_20412_, _20411_, _20407_);
  and (_20413_, _15269_, _07914_);
  or (_20414_, _20413_, _20371_);
  or (_20415_, _20414_, _07237_);
  and (_20417_, _20415_, _07240_);
  and (_20418_, _20417_, _20412_);
  and (_20419_, _11254_, _07914_);
  or (_20420_, _20419_, _20371_);
  and (_20421_, _20420_, _06536_);
  or (_20422_, _20421_, _20418_);
  and (_20423_, _20422_, _07242_);
  or (_20424_, _20371_, _08544_);
  and (_20425_, _20409_, _06375_);
  and (_20426_, _20425_, _20424_);
  or (_20428_, _20426_, _20423_);
  and (_20429_, _20428_, _07234_);
  and (_20430_, _20380_, _06545_);
  and (_20431_, _20430_, _20424_);
  or (_20432_, _20431_, _06366_);
  or (_20433_, _20432_, _20429_);
  and (_20434_, _15266_, _07914_);
  or (_20435_, _20371_, _09056_);
  or (_20436_, _20435_, _20434_);
  and (_20437_, _20436_, _09061_);
  and (_20439_, _20437_, _20433_);
  nor (_20440_, _11253_, _11457_);
  or (_20441_, _20440_, _20371_);
  and (_20442_, _20441_, _06528_);
  or (_20443_, _20442_, _20439_);
  and (_20444_, _20443_, _06926_);
  and (_20445_, _20377_, _06568_);
  or (_20446_, _20445_, _06278_);
  or (_20447_, _20446_, _20444_);
  and (_20448_, _15329_, _07914_);
  or (_20450_, _20371_, _06279_);
  or (_20451_, _20450_, _20448_);
  and (_20452_, _20451_, _01347_);
  and (_20453_, _20452_, _20447_);
  or (_20454_, _20453_, _20370_);
  and (_43183_, _20454_, _42618_);
  and (_20455_, _01351_, \oc8051_golden_model_1.TMOD [5]);
  and (_20456_, _11457_, \oc8051_golden_model_1.TMOD [5]);
  nor (_20457_, _08244_, _11457_);
  or (_20458_, _20457_, _20456_);
  or (_20460_, _20458_, _07215_);
  and (_20461_, _15358_, _07914_);
  or (_20462_, _20461_, _20456_);
  or (_20463_, _20462_, _07151_);
  and (_20464_, _07914_, \oc8051_golden_model_1.ACC [5]);
  or (_20465_, _20464_, _20456_);
  and (_20466_, _20465_, _07141_);
  and (_20467_, _07142_, \oc8051_golden_model_1.TMOD [5]);
  or (_20468_, _20467_, _06341_);
  or (_20469_, _20468_, _20466_);
  and (_20471_, _20469_, _07166_);
  and (_20472_, _20471_, _20463_);
  and (_20473_, _20458_, _06461_);
  or (_20474_, _20473_, _20472_);
  and (_20475_, _20474_, _06465_);
  and (_20476_, _20465_, _06464_);
  or (_20477_, _20476_, _10080_);
  or (_20478_, _20477_, _20475_);
  and (_20479_, _20478_, _20460_);
  or (_20480_, _20479_, _07460_);
  and (_20482_, _09447_, _07914_);
  or (_20483_, _20456_, _07208_);
  or (_20484_, _20483_, _20482_);
  and (_20485_, _20484_, _05982_);
  and (_20486_, _20485_, _20480_);
  and (_20487_, _15459_, _07914_);
  or (_20488_, _20487_, _20456_);
  and (_20489_, _20488_, _10094_);
  or (_20490_, _20489_, _06218_);
  or (_20491_, _20490_, _20486_);
  and (_20493_, _08946_, _07914_);
  or (_20494_, _20493_, _20456_);
  or (_20495_, _20494_, _06219_);
  and (_20496_, _20495_, _20491_);
  or (_20497_, _20496_, _06369_);
  and (_20498_, _15353_, _07914_);
  or (_20499_, _20498_, _20456_);
  or (_20500_, _20499_, _07237_);
  and (_20501_, _20500_, _07240_);
  and (_20502_, _20501_, _20497_);
  and (_20504_, _11250_, _07914_);
  or (_20505_, _20504_, _20456_);
  and (_20506_, _20505_, _06536_);
  or (_20507_, _20506_, _20502_);
  and (_20508_, _20507_, _07242_);
  or (_20509_, _20456_, _08247_);
  and (_20510_, _20494_, _06375_);
  and (_20511_, _20510_, _20509_);
  or (_20512_, _20511_, _20508_);
  and (_20513_, _20512_, _07234_);
  and (_20515_, _20465_, _06545_);
  and (_20516_, _20515_, _20509_);
  or (_20517_, _20516_, _06366_);
  or (_20518_, _20517_, _20513_);
  and (_20519_, _15350_, _07914_);
  or (_20520_, _20456_, _09056_);
  or (_20521_, _20520_, _20519_);
  and (_20522_, _20521_, _09061_);
  and (_20523_, _20522_, _20518_);
  nor (_20524_, _11249_, _11457_);
  or (_20526_, _20524_, _20456_);
  and (_20527_, _20526_, _06528_);
  or (_20528_, _20527_, _20523_);
  and (_20529_, _20528_, _06926_);
  and (_20530_, _20462_, _06568_);
  or (_20531_, _20530_, _06278_);
  or (_20532_, _20531_, _20529_);
  and (_20533_, _15532_, _07914_);
  or (_20534_, _20456_, _06279_);
  or (_20535_, _20534_, _20533_);
  and (_20537_, _20535_, _01347_);
  and (_20538_, _20537_, _20532_);
  or (_20539_, _20538_, _20455_);
  and (_43184_, _20539_, _42618_);
  and (_20540_, _01351_, \oc8051_golden_model_1.TMOD [6]);
  and (_20541_, _11457_, \oc8051_golden_model_1.TMOD [6]);
  and (_20542_, _15554_, _07914_);
  or (_20543_, _20542_, _20541_);
  or (_20544_, _20543_, _07151_);
  and (_20545_, _07914_, \oc8051_golden_model_1.ACC [6]);
  or (_20547_, _20545_, _20541_);
  and (_20548_, _20547_, _07141_);
  and (_20549_, _07142_, \oc8051_golden_model_1.TMOD [6]);
  or (_20550_, _20549_, _06341_);
  or (_20551_, _20550_, _20548_);
  and (_20552_, _20551_, _07166_);
  and (_20553_, _20552_, _20544_);
  nor (_20554_, _08142_, _11457_);
  or (_20555_, _20554_, _20541_);
  and (_20556_, _20555_, _06461_);
  or (_20558_, _20556_, _20553_);
  and (_20559_, _20558_, _06465_);
  and (_20560_, _20547_, _06464_);
  or (_20561_, _20560_, _10080_);
  or (_20562_, _20561_, _20559_);
  or (_20563_, _20555_, _07215_);
  and (_20564_, _20563_, _20562_);
  or (_20565_, _20564_, _07460_);
  and (_20566_, _09446_, _07914_);
  or (_20567_, _20541_, _07208_);
  or (_20569_, _20567_, _20566_);
  and (_20570_, _20569_, _05982_);
  and (_20571_, _20570_, _20565_);
  and (_20572_, _15657_, _07914_);
  or (_20573_, _20572_, _20541_);
  and (_20574_, _20573_, _10094_);
  or (_20575_, _20574_, _06218_);
  or (_20576_, _20575_, _20571_);
  and (_20577_, _15664_, _07914_);
  or (_20578_, _20577_, _20541_);
  or (_20580_, _20578_, _06219_);
  and (_20581_, _20580_, _20576_);
  or (_20582_, _20581_, _06369_);
  and (_20583_, _15549_, _07914_);
  or (_20584_, _20583_, _20541_);
  or (_20585_, _20584_, _07237_);
  and (_20586_, _20585_, _07240_);
  and (_20587_, _20586_, _20582_);
  and (_20588_, _11247_, _07914_);
  or (_20589_, _20588_, _20541_);
  and (_20591_, _20589_, _06536_);
  or (_20592_, _20591_, _20587_);
  and (_20593_, _20592_, _07242_);
  or (_20594_, _20541_, _08145_);
  and (_20595_, _20578_, _06375_);
  and (_20596_, _20595_, _20594_);
  or (_20597_, _20596_, _20593_);
  and (_20598_, _20597_, _07234_);
  and (_20599_, _20547_, _06545_);
  and (_20600_, _20599_, _20594_);
  or (_20602_, _20600_, _06366_);
  or (_20603_, _20602_, _20598_);
  and (_20604_, _15546_, _07914_);
  or (_20605_, _20541_, _09056_);
  or (_20606_, _20605_, _20604_);
  and (_20607_, _20606_, _09061_);
  and (_20608_, _20607_, _20603_);
  nor (_20609_, _11246_, _11457_);
  or (_20610_, _20609_, _20541_);
  and (_20611_, _20610_, _06528_);
  or (_20613_, _20611_, _20608_);
  and (_20614_, _20613_, _06926_);
  and (_20615_, _20543_, _06568_);
  or (_20616_, _20615_, _06278_);
  or (_20617_, _20616_, _20614_);
  and (_20618_, _15734_, _07914_);
  or (_20619_, _20541_, _06279_);
  or (_20620_, _20619_, _20618_);
  and (_20621_, _20620_, _01347_);
  and (_20622_, _20621_, _20617_);
  or (_20624_, _20622_, _20540_);
  and (_43185_, _20624_, _42618_);
  not (_20625_, \oc8051_golden_model_1.DPL [0]);
  nor (_20626_, _01347_, _20625_);
  and (_20627_, _07960_, \oc8051_golden_model_1.ACC [0]);
  and (_20628_, _20627_, _08390_);
  nor (_20629_, _07960_, _20625_);
  or (_20630_, _20629_, _07234_);
  or (_20631_, _20630_, _20628_);
  and (_20632_, _09392_, _07960_);
  or (_20634_, _20632_, _20629_);
  and (_20635_, _20634_, _07460_);
  and (_20636_, _07960_, _07133_);
  or (_20637_, _20636_, _20629_);
  or (_20638_, _20637_, _07166_);
  nor (_20639_, _08390_, _11537_);
  or (_20640_, _20639_, _20629_);
  and (_20641_, _20640_, _06341_);
  nor (_20642_, _07141_, _20625_);
  or (_20643_, _20629_, _20627_);
  and (_20645_, _20643_, _07141_);
  or (_20646_, _20645_, _20642_);
  and (_20647_, _20646_, _07151_);
  or (_20648_, _20647_, _06461_);
  or (_20649_, _20648_, _20641_);
  and (_20650_, _20649_, _20638_);
  or (_20651_, _20650_, _06464_);
  or (_20652_, _20643_, _06465_);
  and (_20653_, _20652_, _11562_);
  and (_20654_, _20653_, _20651_);
  and (_20656_, _11561_, _20625_);
  or (_20657_, _20656_, _20654_);
  and (_20658_, _20657_, _06374_);
  nor (_20659_, _06872_, _06374_);
  or (_20660_, _20659_, _10080_);
  or (_20661_, _20660_, _20658_);
  or (_20662_, _20637_, _07215_);
  and (_20663_, _20662_, _07208_);
  and (_20664_, _20663_, _20661_);
  or (_20665_, _20664_, _10094_);
  or (_20666_, _20665_, _20635_);
  and (_20667_, _14467_, _07960_);
  or (_20668_, _20629_, _05982_);
  or (_20669_, _20668_, _20667_);
  and (_20670_, _20669_, _06219_);
  and (_20671_, _20670_, _20666_);
  and (_20672_, _07960_, _08954_);
  or (_20673_, _20672_, _20629_);
  and (_20674_, _20673_, _06218_);
  or (_20675_, _20674_, _06369_);
  or (_20677_, _20675_, _20671_);
  and (_20678_, _14366_, _07960_);
  or (_20679_, _20678_, _20629_);
  or (_20680_, _20679_, _07237_);
  and (_20681_, _20680_, _07240_);
  and (_20682_, _20681_, _20677_);
  nor (_20683_, _12580_, _11537_);
  or (_20684_, _20683_, _20629_);
  nor (_20685_, _20628_, _07240_);
  and (_20686_, _20685_, _20684_);
  or (_20689_, _20686_, _20682_);
  and (_20690_, _20689_, _07242_);
  nand (_20691_, _20673_, _06375_);
  nor (_20692_, _20691_, _20639_);
  or (_20693_, _20692_, _06545_);
  or (_20694_, _20693_, _20690_);
  and (_20695_, _20694_, _20631_);
  or (_20696_, _20695_, _06366_);
  and (_20697_, _14363_, _07960_);
  or (_20698_, _20697_, _20629_);
  or (_20700_, _20698_, _09056_);
  and (_20701_, _20700_, _09061_);
  and (_20702_, _20701_, _20696_);
  and (_20703_, _20684_, _06528_);
  or (_20704_, _20703_, _19502_);
  or (_20705_, _20704_, _20702_);
  or (_20706_, _20640_, _06661_);
  and (_20707_, _20706_, _01347_);
  and (_20708_, _20707_, _20705_);
  or (_20709_, _20708_, _20626_);
  and (_43187_, _20709_, _42618_);
  not (_20710_, \oc8051_golden_model_1.DPL [1]);
  nor (_20711_, _01347_, _20710_);
  or (_20712_, _09451_, _11537_);
  or (_20713_, _07960_, \oc8051_golden_model_1.DPL [1]);
  and (_20714_, _20713_, _07460_);
  and (_20715_, _20714_, _20712_);
  nor (_20716_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.DPL [0]);
  nor (_20717_, _20716_, _11566_);
  and (_20718_, _20717_, _11561_);
  and (_20720_, _14562_, _07960_);
  not (_20721_, _20720_);
  and (_20722_, _20721_, _20713_);
  or (_20723_, _20722_, _07151_);
  nor (_20724_, _07960_, _20710_);
  and (_20725_, _07960_, \oc8051_golden_model_1.ACC [1]);
  or (_20726_, _20725_, _20724_);
  and (_20727_, _20726_, _07141_);
  nor (_20728_, _07141_, _20710_);
  or (_20729_, _20728_, _06341_);
  or (_20732_, _20729_, _20727_);
  and (_20733_, _20732_, _07166_);
  and (_20734_, _20733_, _20723_);
  nor (_20735_, _11537_, _07357_);
  or (_20736_, _20735_, _20724_);
  and (_20737_, _20736_, _06461_);
  or (_20738_, _20737_, _06464_);
  or (_20739_, _20738_, _20734_);
  or (_20740_, _20726_, _06465_);
  and (_20741_, _20740_, _11562_);
  and (_20742_, _20741_, _20739_);
  or (_20743_, _20742_, _20718_);
  and (_20744_, _20743_, _06374_);
  nor (_20745_, _07038_, _06374_);
  or (_20746_, _20745_, _10080_);
  or (_20747_, _20746_, _20744_);
  or (_20748_, _20736_, _07215_);
  and (_20749_, _20748_, _07208_);
  and (_20750_, _20749_, _20747_);
  or (_20751_, _20750_, _20715_);
  and (_20753_, _20751_, _05982_);
  or (_20754_, _14653_, _11537_);
  and (_20755_, _20713_, _10094_);
  and (_20756_, _20755_, _20754_);
  or (_20757_, _20756_, _20753_);
  and (_20758_, _20757_, _06219_);
  nand (_20759_, _07960_, _07038_);
  and (_20760_, _20713_, _06218_);
  and (_20761_, _20760_, _20759_);
  or (_20762_, _20761_, _20758_);
  and (_20765_, _20762_, _07237_);
  or (_20766_, _14668_, _11537_);
  and (_20767_, _20713_, _06369_);
  and (_20768_, _20767_, _20766_);
  or (_20769_, _20768_, _06536_);
  or (_20770_, _20769_, _20765_);
  nor (_20771_, _11261_, _11537_);
  or (_20772_, _20771_, _20724_);
  nand (_20773_, _11260_, _07960_);
  and (_20774_, _20773_, _20772_);
  or (_20776_, _20774_, _07240_);
  and (_20777_, _20776_, _07242_);
  and (_20778_, _20777_, _20770_);
  or (_20779_, _14666_, _11537_);
  and (_20780_, _20713_, _06375_);
  and (_20781_, _20780_, _20779_);
  or (_20782_, _20781_, _06545_);
  or (_20783_, _20782_, _20778_);
  nor (_20784_, _20724_, _07234_);
  nand (_20785_, _20784_, _20773_);
  and (_20787_, _20785_, _09056_);
  and (_20788_, _20787_, _20783_);
  or (_20789_, _20759_, _08341_);
  and (_20790_, _20713_, _06366_);
  and (_20791_, _20790_, _20789_);
  or (_20792_, _20791_, _06528_);
  or (_20793_, _20792_, _20788_);
  or (_20794_, _20772_, _09061_);
  and (_20795_, _20794_, _06926_);
  and (_20796_, _20795_, _20793_);
  and (_20798_, _20722_, _06568_);
  or (_20799_, _20798_, _06278_);
  or (_20800_, _20799_, _20796_);
  or (_20801_, _20724_, _06279_);
  or (_20802_, _20801_, _20720_);
  and (_20803_, _20802_, _01347_);
  and (_20804_, _20803_, _20800_);
  or (_20805_, _20804_, _20711_);
  and (_43188_, _20805_, _42618_);
  not (_20806_, \oc8051_golden_model_1.DPL [2]);
  nor (_20807_, _01347_, _20806_);
  nor (_20808_, _07960_, _20806_);
  nor (_20809_, _11537_, _07776_);
  or (_20810_, _20809_, _20808_);
  or (_20811_, _20810_, _07215_);
  or (_20812_, _20810_, _07166_);
  and (_20813_, _14770_, _07960_);
  or (_20814_, _20813_, _20808_);
  and (_20815_, _20814_, _06341_);
  nor (_20816_, _07141_, _20806_);
  and (_20819_, _07960_, \oc8051_golden_model_1.ACC [2]);
  or (_20820_, _20819_, _20808_);
  and (_20821_, _20820_, _07141_);
  or (_20822_, _20821_, _20816_);
  and (_20823_, _20822_, _07151_);
  or (_20824_, _20823_, _06461_);
  or (_20825_, _20824_, _20815_);
  and (_20826_, _20825_, _20812_);
  or (_20827_, _20826_, _06464_);
  or (_20828_, _20820_, _06465_);
  and (_20830_, _20828_, _11562_);
  and (_20831_, _20830_, _20827_);
  nor (_20832_, _11566_, \oc8051_golden_model_1.DPL [2]);
  nor (_20833_, _20832_, _11567_);
  and (_20834_, _20833_, _11561_);
  or (_20835_, _20834_, _20831_);
  and (_20836_, _20835_, _06374_);
  nor (_20837_, _06697_, _06374_);
  or (_20838_, _20837_, _10080_);
  or (_20839_, _20838_, _20836_);
  and (_20841_, _20839_, _20811_);
  or (_20842_, _20841_, _07460_);
  and (_20843_, _09450_, _07960_);
  or (_20844_, _20808_, _07208_);
  or (_20845_, _20844_, _20843_);
  and (_20846_, _20845_, _05982_);
  and (_20847_, _20846_, _20842_);
  and (_20848_, _14859_, _07960_);
  or (_20849_, _20848_, _20808_);
  and (_20850_, _20849_, _10094_);
  or (_20852_, _20850_, _06218_);
  or (_20853_, _20852_, _20847_);
  and (_20854_, _07960_, _08973_);
  or (_20855_, _20854_, _20808_);
  or (_20856_, _20855_, _06219_);
  and (_20857_, _20856_, _20853_);
  or (_20858_, _20857_, _06369_);
  and (_20859_, _14751_, _07960_);
  or (_20860_, _20859_, _20808_);
  or (_20861_, _20860_, _07237_);
  and (_20863_, _20861_, _07240_);
  and (_20864_, _20863_, _20858_);
  and (_20865_, _11259_, _07960_);
  or (_20866_, _20865_, _20808_);
  and (_20867_, _20866_, _06536_);
  or (_20868_, _20867_, _20864_);
  and (_20869_, _20868_, _07242_);
  or (_20870_, _20808_, _08440_);
  and (_20871_, _20855_, _06375_);
  and (_20872_, _20871_, _20870_);
  or (_20874_, _20872_, _20869_);
  and (_20875_, _20874_, _07234_);
  and (_20876_, _20820_, _06545_);
  and (_20877_, _20876_, _20870_);
  or (_20878_, _20877_, _06366_);
  or (_20879_, _20878_, _20875_);
  and (_20880_, _14748_, _07960_);
  or (_20881_, _20808_, _09056_);
  or (_20882_, _20881_, _20880_);
  and (_20883_, _20882_, _09061_);
  and (_20885_, _20883_, _20879_);
  nor (_20886_, _11258_, _11537_);
  or (_20887_, _20886_, _20808_);
  and (_20888_, _20887_, _06528_);
  or (_20889_, _20888_, _20885_);
  and (_20890_, _20889_, _06926_);
  and (_20891_, _20814_, _06568_);
  or (_20892_, _20891_, _06278_);
  or (_20893_, _20892_, _20890_);
  and (_20894_, _14926_, _07960_);
  or (_20896_, _20808_, _06279_);
  or (_20897_, _20896_, _20894_);
  and (_20898_, _20897_, _01347_);
  and (_20899_, _20898_, _20893_);
  or (_20900_, _20899_, _20807_);
  and (_43189_, _20900_, _42618_);
  not (_20901_, \oc8051_golden_model_1.DPL [3]);
  nor (_20902_, _01347_, _20901_);
  nor (_20903_, _07960_, _20901_);
  nor (_20904_, _11537_, _07594_);
  or (_20906_, _20904_, _20903_);
  or (_20907_, _20906_, _07215_);
  and (_20908_, _14953_, _07960_);
  or (_20909_, _20908_, _20903_);
  or (_20910_, _20909_, _07151_);
  and (_20911_, _07960_, \oc8051_golden_model_1.ACC [3]);
  or (_20912_, _20911_, _20903_);
  and (_20913_, _20912_, _07141_);
  nor (_20914_, _07141_, _20901_);
  or (_20915_, _20914_, _06341_);
  or (_20917_, _20915_, _20913_);
  and (_20918_, _20917_, _07166_);
  and (_20919_, _20918_, _20910_);
  and (_20920_, _20906_, _06461_);
  or (_20921_, _20920_, _06464_);
  or (_20922_, _20921_, _20919_);
  or (_20923_, _20912_, _06465_);
  and (_20924_, _20923_, _11562_);
  and (_20925_, _20924_, _20922_);
  nor (_20926_, _11567_, \oc8051_golden_model_1.DPL [3]);
  nor (_20928_, _20926_, _11568_);
  and (_20929_, _20928_, _11561_);
  or (_20930_, _20929_, _20925_);
  and (_20931_, _20930_, _06374_);
  nor (_20932_, _06452_, _06374_);
  or (_20933_, _20932_, _10080_);
  or (_20934_, _20933_, _20931_);
  and (_20935_, _20934_, _20907_);
  or (_20936_, _20935_, _07460_);
  and (_20937_, _09449_, _07960_);
  or (_20938_, _20903_, _07208_);
  or (_20939_, _20938_, _20937_);
  and (_20940_, _20939_, _05982_);
  and (_20941_, _20940_, _20936_);
  and (_20942_, _15048_, _07960_);
  or (_20943_, _20942_, _20903_);
  and (_20944_, _20943_, _10094_);
  or (_20945_, _20944_, _06218_);
  or (_20946_, _20945_, _20941_);
  and (_20947_, _07960_, _08930_);
  or (_20950_, _20947_, _20903_);
  or (_20951_, _20950_, _06219_);
  and (_20952_, _20951_, _20946_);
  or (_20953_, _20952_, _06369_);
  and (_20954_, _14943_, _07960_);
  or (_20955_, _20954_, _20903_);
  or (_20956_, _20955_, _07237_);
  and (_20957_, _20956_, _07240_);
  and (_20958_, _20957_, _20953_);
  and (_20959_, _12577_, _07960_);
  or (_20961_, _20959_, _20903_);
  and (_20962_, _20961_, _06536_);
  or (_20963_, _20962_, _20958_);
  and (_20964_, _20963_, _07242_);
  or (_20965_, _20903_, _08292_);
  and (_20966_, _20950_, _06375_);
  and (_20967_, _20966_, _20965_);
  or (_20968_, _20967_, _20964_);
  and (_20969_, _20968_, _07234_);
  and (_20970_, _20912_, _06545_);
  and (_20972_, _20970_, _20965_);
  or (_20973_, _20972_, _06366_);
  or (_20974_, _20973_, _20969_);
  and (_20975_, _14940_, _07960_);
  or (_20976_, _20903_, _09056_);
  or (_20977_, _20976_, _20975_);
  and (_20978_, _20977_, _09061_);
  and (_20979_, _20978_, _20974_);
  nor (_20980_, _11256_, _11537_);
  or (_20981_, _20980_, _20903_);
  and (_20983_, _20981_, _06528_);
  or (_20984_, _20983_, _20979_);
  and (_20985_, _20984_, _06926_);
  and (_20986_, _20909_, _06568_);
  or (_20987_, _20986_, _06278_);
  or (_20988_, _20987_, _20985_);
  and (_20989_, _15128_, _07960_);
  or (_20990_, _20903_, _06279_);
  or (_20991_, _20990_, _20989_);
  and (_20992_, _20991_, _01347_);
  and (_20994_, _20992_, _20988_);
  or (_20995_, _20994_, _20902_);
  and (_43190_, _20995_, _42618_);
  not (_20996_, \oc8051_golden_model_1.DPL [4]);
  nor (_20997_, _01347_, _20996_);
  nor (_20998_, _07960_, _20996_);
  nor (_20999_, _08541_, _11537_);
  or (_21000_, _20999_, _20998_);
  or (_21001_, _21000_, _07215_);
  and (_21002_, _15162_, _07960_);
  or (_21004_, _21002_, _20998_);
  or (_21005_, _21004_, _07151_);
  and (_21006_, _07960_, \oc8051_golden_model_1.ACC [4]);
  or (_21007_, _21006_, _20998_);
  and (_21008_, _21007_, _07141_);
  nor (_21009_, _07141_, _20996_);
  or (_21010_, _21009_, _06341_);
  or (_21011_, _21010_, _21008_);
  and (_21012_, _21011_, _07166_);
  and (_21013_, _21012_, _21005_);
  and (_21015_, _21000_, _06461_);
  or (_21016_, _21015_, _06464_);
  or (_21017_, _21016_, _21013_);
  or (_21018_, _21007_, _06465_);
  and (_21019_, _21018_, _11562_);
  and (_21020_, _21019_, _21017_);
  nor (_21021_, _11568_, \oc8051_golden_model_1.DPL [4]);
  nor (_21022_, _21021_, _11569_);
  and (_21023_, _21022_, _11561_);
  or (_21024_, _21023_, _21020_);
  and (_21026_, _21024_, _06374_);
  nor (_21027_, _08892_, _06374_);
  or (_21028_, _21027_, _10080_);
  or (_21029_, _21028_, _21026_);
  and (_21030_, _21029_, _21001_);
  or (_21031_, _21030_, _07460_);
  and (_21032_, _09448_, _07960_);
  or (_21033_, _20998_, _07208_);
  or (_21034_, _21033_, _21032_);
  and (_21035_, _21034_, _05982_);
  and (_21037_, _21035_, _21031_);
  and (_21038_, _15254_, _07960_);
  or (_21039_, _21038_, _20998_);
  and (_21040_, _21039_, _10094_);
  or (_21041_, _21040_, _06218_);
  or (_21042_, _21041_, _21037_);
  and (_21043_, _08959_, _07960_);
  or (_21044_, _21043_, _20998_);
  or (_21045_, _21044_, _06219_);
  and (_21046_, _21045_, _21042_);
  or (_21048_, _21046_, _06369_);
  and (_21049_, _15269_, _07960_);
  or (_21050_, _21049_, _20998_);
  or (_21051_, _21050_, _07237_);
  and (_21052_, _21051_, _07240_);
  and (_21053_, _21052_, _21048_);
  and (_21054_, _11254_, _07960_);
  or (_21055_, _21054_, _20998_);
  and (_21056_, _21055_, _06536_);
  or (_21057_, _21056_, _21053_);
  and (_21059_, _21057_, _07242_);
  or (_21060_, _20998_, _08544_);
  and (_21061_, _21044_, _06375_);
  and (_21062_, _21061_, _21060_);
  or (_21063_, _21062_, _21059_);
  and (_21064_, _21063_, _07234_);
  and (_21065_, _21007_, _06545_);
  and (_21066_, _21065_, _21060_);
  or (_21067_, _21066_, _06366_);
  or (_21068_, _21067_, _21064_);
  and (_21070_, _15266_, _07960_);
  or (_21071_, _20998_, _09056_);
  or (_21072_, _21071_, _21070_);
  and (_21073_, _21072_, _09061_);
  and (_21074_, _21073_, _21068_);
  nor (_21075_, _11253_, _11537_);
  or (_21076_, _21075_, _20998_);
  and (_21077_, _21076_, _06528_);
  or (_21078_, _21077_, _21074_);
  and (_21079_, _21078_, _06926_);
  and (_21081_, _21004_, _06568_);
  or (_21082_, _21081_, _06278_);
  or (_21083_, _21082_, _21079_);
  and (_21084_, _15329_, _07960_);
  or (_21085_, _20998_, _06279_);
  or (_21086_, _21085_, _21084_);
  and (_21087_, _21086_, _01347_);
  and (_21088_, _21087_, _21083_);
  or (_21089_, _21088_, _20997_);
  and (_43191_, _21089_, _42618_);
  not (_21091_, \oc8051_golden_model_1.DPL [5]);
  nor (_21092_, _01347_, _21091_);
  nor (_21093_, _07960_, _21091_);
  nor (_21094_, _08244_, _11537_);
  or (_21095_, _21094_, _21093_);
  or (_21096_, _21095_, _07215_);
  and (_21097_, _15358_, _07960_);
  or (_21098_, _21097_, _21093_);
  or (_21099_, _21098_, _07151_);
  and (_21100_, _07960_, \oc8051_golden_model_1.ACC [5]);
  or (_21102_, _21100_, _21093_);
  and (_21103_, _21102_, _07141_);
  nor (_21104_, _07141_, _21091_);
  or (_21105_, _21104_, _06341_);
  or (_21106_, _21105_, _21103_);
  and (_21107_, _21106_, _07166_);
  and (_21108_, _21107_, _21099_);
  and (_21109_, _21095_, _06461_);
  or (_21110_, _21109_, _06464_);
  or (_21111_, _21110_, _21108_);
  or (_21112_, _21102_, _06465_);
  and (_21113_, _21112_, _11562_);
  and (_21114_, _21113_, _21111_);
  nor (_21115_, _11569_, \oc8051_golden_model_1.DPL [5]);
  nor (_21116_, _21115_, _11570_);
  and (_21117_, _21116_, _11561_);
  or (_21118_, _21117_, _21114_);
  and (_21119_, _21118_, _06374_);
  nor (_21120_, _08926_, _06374_);
  or (_21121_, _21120_, _10080_);
  or (_21124_, _21121_, _21119_);
  and (_21125_, _21124_, _21096_);
  or (_21126_, _21125_, _07460_);
  and (_21127_, _09447_, _07960_);
  or (_21128_, _21093_, _07208_);
  or (_21129_, _21128_, _21127_);
  and (_21130_, _21129_, _05982_);
  and (_21131_, _21130_, _21126_);
  and (_21132_, _15459_, _07960_);
  or (_21133_, _21132_, _21093_);
  and (_21135_, _21133_, _10094_);
  or (_21136_, _21135_, _06218_);
  or (_21137_, _21136_, _21131_);
  and (_21138_, _08946_, _07960_);
  or (_21139_, _21138_, _21093_);
  or (_21140_, _21139_, _06219_);
  and (_21141_, _21140_, _21137_);
  or (_21142_, _21141_, _06369_);
  and (_21143_, _15353_, _07960_);
  or (_21144_, _21143_, _21093_);
  or (_21146_, _21144_, _07237_);
  and (_21147_, _21146_, _07240_);
  and (_21148_, _21147_, _21142_);
  and (_21149_, _11250_, _07960_);
  or (_21150_, _21149_, _21093_);
  and (_21151_, _21150_, _06536_);
  or (_21152_, _21151_, _21148_);
  and (_21153_, _21152_, _07242_);
  or (_21154_, _21093_, _08247_);
  and (_21155_, _21139_, _06375_);
  and (_21157_, _21155_, _21154_);
  or (_21158_, _21157_, _21153_);
  and (_21159_, _21158_, _07234_);
  and (_21160_, _21102_, _06545_);
  and (_21161_, _21160_, _21154_);
  or (_21162_, _21161_, _06366_);
  or (_21163_, _21162_, _21159_);
  and (_21164_, _15350_, _07960_);
  or (_21165_, _21093_, _09056_);
  or (_21166_, _21165_, _21164_);
  and (_21168_, _21166_, _09061_);
  and (_21169_, _21168_, _21163_);
  nor (_21170_, _11249_, _11537_);
  or (_21171_, _21170_, _21093_);
  and (_21172_, _21171_, _06528_);
  or (_21173_, _21172_, _21169_);
  and (_21174_, _21173_, _06926_);
  and (_21175_, _21098_, _06568_);
  or (_21176_, _21175_, _06278_);
  or (_21177_, _21176_, _21174_);
  and (_21179_, _15532_, _07960_);
  or (_21180_, _21093_, _06279_);
  or (_21181_, _21180_, _21179_);
  and (_21182_, _21181_, _01347_);
  and (_21183_, _21182_, _21177_);
  or (_21184_, _21183_, _21092_);
  and (_43192_, _21184_, _42618_);
  not (_21185_, \oc8051_golden_model_1.DPL [6]);
  nor (_21186_, _01347_, _21185_);
  nor (_21187_, _07960_, _21185_);
  nor (_21189_, _08142_, _11537_);
  or (_21190_, _21189_, _21187_);
  or (_21191_, _21190_, _07215_);
  and (_21192_, _15554_, _07960_);
  or (_21193_, _21192_, _21187_);
  or (_21194_, _21193_, _07151_);
  and (_21195_, _07960_, \oc8051_golden_model_1.ACC [6]);
  or (_21196_, _21195_, _21187_);
  and (_21197_, _21196_, _07141_);
  nor (_21198_, _07141_, _21185_);
  or (_21200_, _21198_, _06341_);
  or (_21201_, _21200_, _21197_);
  and (_21202_, _21201_, _07166_);
  and (_21203_, _21202_, _21194_);
  and (_21204_, _21190_, _06461_);
  or (_21205_, _21204_, _06464_);
  or (_21206_, _21205_, _21203_);
  or (_21207_, _21196_, _06465_);
  and (_21208_, _21207_, _11562_);
  and (_21209_, _21208_, _21206_);
  nor (_21211_, _11570_, \oc8051_golden_model_1.DPL [6]);
  nor (_21212_, _21211_, _11571_);
  and (_21213_, _21212_, _11561_);
  or (_21214_, _21213_, _21209_);
  and (_21215_, _21214_, _06374_);
  nor (_21216_, _08857_, _06374_);
  or (_21217_, _21216_, _10080_);
  or (_21218_, _21217_, _21215_);
  and (_21219_, _21218_, _21191_);
  or (_21220_, _21219_, _07460_);
  and (_21222_, _09446_, _07960_);
  or (_21223_, _21187_, _07208_);
  or (_21224_, _21223_, _21222_);
  and (_21225_, _21224_, _05982_);
  and (_21226_, _21225_, _21220_);
  and (_21227_, _15657_, _07960_);
  or (_21228_, _21227_, _21187_);
  and (_21229_, _21228_, _10094_);
  or (_21230_, _21229_, _06218_);
  or (_21231_, _21230_, _21226_);
  and (_21233_, _15664_, _07960_);
  or (_21234_, _21233_, _21187_);
  or (_21235_, _21234_, _06219_);
  and (_21236_, _21235_, _21231_);
  or (_21237_, _21236_, _06369_);
  and (_21238_, _15549_, _07960_);
  or (_21239_, _21238_, _21187_);
  or (_21240_, _21239_, _07237_);
  and (_21241_, _21240_, _07240_);
  and (_21242_, _21241_, _21237_);
  and (_21244_, _11247_, _07960_);
  or (_21245_, _21244_, _21187_);
  and (_21246_, _21245_, _06536_);
  or (_21247_, _21246_, _21242_);
  and (_21248_, _21247_, _07242_);
  or (_21249_, _21187_, _08145_);
  and (_21250_, _21234_, _06375_);
  and (_21251_, _21250_, _21249_);
  or (_21252_, _21251_, _21248_);
  and (_21253_, _21252_, _07234_);
  and (_21255_, _21196_, _06545_);
  and (_21256_, _21255_, _21249_);
  or (_21257_, _21256_, _06366_);
  or (_21258_, _21257_, _21253_);
  and (_21259_, _15546_, _07960_);
  or (_21260_, _21187_, _09056_);
  or (_21261_, _21260_, _21259_);
  and (_21262_, _21261_, _09061_);
  and (_21263_, _21262_, _21258_);
  nor (_21264_, _11246_, _11537_);
  or (_21266_, _21264_, _21187_);
  and (_21267_, _21266_, _06528_);
  or (_21268_, _21267_, _21263_);
  and (_21269_, _21268_, _06926_);
  and (_21270_, _21193_, _06568_);
  or (_21271_, _21270_, _06278_);
  or (_21272_, _21271_, _21269_);
  and (_21273_, _15734_, _07960_);
  or (_21274_, _21187_, _06279_);
  or (_21275_, _21274_, _21273_);
  and (_21277_, _21275_, _01347_);
  and (_21278_, _21277_, _21272_);
  or (_21279_, _21278_, _21186_);
  and (_43193_, _21279_, _42618_);
  nor (_21280_, _01347_, _12693_);
  nor (_21281_, _07963_, _12693_);
  and (_21282_, _07963_, \oc8051_golden_model_1.ACC [0]);
  and (_21283_, _21282_, _08390_);
  or (_21284_, _21283_, _21281_);
  or (_21285_, _21284_, _07234_);
  and (_21287_, _09392_, _07963_);
  or (_21288_, _21287_, _21281_);
  and (_21289_, _21288_, _07460_);
  and (_21290_, _08186_, _07133_);
  or (_21291_, _21290_, _21281_);
  or (_21292_, _21291_, _07166_);
  nor (_21293_, _08390_, _11633_);
  or (_21294_, _21293_, _21281_);
  and (_21295_, _21294_, _06341_);
  nor (_21296_, _07141_, _12693_);
  or (_21298_, _21282_, _21281_);
  and (_21299_, _21298_, _07141_);
  or (_21300_, _21299_, _21296_);
  and (_21301_, _21300_, _07151_);
  or (_21302_, _21301_, _06461_);
  or (_21303_, _21302_, _21295_);
  and (_21304_, _21303_, _21292_);
  or (_21305_, _21304_, _06464_);
  or (_21306_, _21298_, _06465_);
  and (_21307_, _21306_, _11562_);
  and (_21308_, _21307_, _21305_);
  or (_21309_, _11573_, \oc8051_golden_model_1.DPH [0]);
  nor (_21310_, _11660_, _11562_);
  and (_21311_, _21310_, _21309_);
  or (_21312_, _21311_, _21308_);
  and (_21313_, _21312_, _06374_);
  nor (_21314_, _06374_, _06251_);
  or (_21315_, _21314_, _10080_);
  or (_21316_, _21315_, _21313_);
  or (_21317_, _21291_, _07215_);
  and (_21320_, _21317_, _07208_);
  and (_21321_, _21320_, _21316_);
  or (_21322_, _21321_, _10094_);
  or (_21323_, _21322_, _21289_);
  and (_21324_, _14467_, _08186_);
  or (_21325_, _21281_, _05982_);
  or (_21326_, _21325_, _21324_);
  and (_21327_, _21326_, _06219_);
  and (_21328_, _21327_, _21323_);
  and (_21329_, _07963_, _08954_);
  or (_21331_, _21329_, _21281_);
  and (_21332_, _21331_, _06218_);
  or (_21333_, _21332_, _06369_);
  or (_21334_, _21333_, _21328_);
  and (_21335_, _14366_, _07963_);
  or (_21336_, _21335_, _21281_);
  or (_21337_, _21336_, _07237_);
  and (_21338_, _21337_, _07240_);
  and (_21339_, _21338_, _21334_);
  nor (_21340_, _12580_, _11633_);
  or (_21342_, _21340_, _21281_);
  nor (_21343_, _21283_, _07240_);
  and (_21344_, _21343_, _21342_);
  or (_21345_, _21344_, _21339_);
  and (_21346_, _21345_, _07242_);
  nand (_21347_, _21331_, _06375_);
  nor (_21348_, _21347_, _21293_);
  or (_21349_, _21348_, _06545_);
  or (_21350_, _21349_, _21346_);
  and (_21351_, _21350_, _21285_);
  or (_21353_, _21351_, _06366_);
  and (_21354_, _14363_, _07963_);
  or (_21355_, _21354_, _21281_);
  or (_21356_, _21355_, _09056_);
  and (_21357_, _21356_, _09061_);
  and (_21358_, _21357_, _21353_);
  and (_21359_, _21342_, _06528_);
  or (_21360_, _21359_, _19502_);
  or (_21361_, _21360_, _21358_);
  or (_21362_, _21294_, _06661_);
  and (_21364_, _21362_, _01347_);
  and (_21365_, _21364_, _21361_);
  or (_21366_, _21365_, _21280_);
  and (_43195_, _21366_, _42618_);
  not (_21367_, \oc8051_golden_model_1.DPH [1]);
  nor (_21368_, _01347_, _21367_);
  or (_21369_, _07963_, \oc8051_golden_model_1.DPH [1]);
  and (_21370_, _21369_, _06218_);
  nand (_21371_, _08186_, _07038_);
  and (_21372_, _21371_, _21370_);
  or (_21374_, _09451_, _11633_);
  and (_21375_, _21369_, _07460_);
  and (_21376_, _21375_, _21374_);
  nor (_21377_, _11660_, \oc8051_golden_model_1.DPH [1]);
  nor (_21378_, _21377_, _11661_);
  and (_21379_, _21378_, _11561_);
  and (_21380_, _14562_, _08186_);
  not (_21381_, _21380_);
  and (_21382_, _21381_, _21369_);
  or (_21383_, _21382_, _07151_);
  nor (_21385_, _07963_, _21367_);
  and (_21386_, _07963_, \oc8051_golden_model_1.ACC [1]);
  or (_21387_, _21386_, _21385_);
  and (_21388_, _21387_, _07141_);
  nor (_21389_, _07141_, _21367_);
  or (_21390_, _21389_, _06341_);
  or (_21391_, _21390_, _21388_);
  and (_21392_, _21391_, _07166_);
  and (_21393_, _21392_, _21383_);
  nor (_21394_, _11633_, _07357_);
  or (_21396_, _21394_, _21385_);
  and (_21397_, _21396_, _06461_);
  or (_21398_, _21397_, _06464_);
  or (_21399_, _21398_, _21393_);
  or (_21400_, _21387_, _06465_);
  and (_21401_, _21400_, _11562_);
  and (_21402_, _21401_, _21399_);
  or (_21403_, _21402_, _21379_);
  and (_21404_, _21403_, _06374_);
  nor (_21405_, _07004_, _06374_);
  or (_21407_, _21405_, _10080_);
  or (_21408_, _21407_, _21404_);
  or (_21409_, _21396_, _07215_);
  and (_21410_, _21409_, _07208_);
  and (_21411_, _21410_, _21408_);
  or (_21412_, _21411_, _21376_);
  and (_21413_, _21412_, _05982_);
  and (_21414_, _14653_, _07963_);
  or (_21415_, _21414_, _21385_);
  and (_21416_, _21415_, _10094_);
  or (_21418_, _21416_, _21413_);
  and (_21419_, _21418_, _06219_);
  or (_21420_, _21419_, _21372_);
  and (_21421_, _21420_, _07237_);
  or (_21422_, _14668_, _11633_);
  and (_21423_, _21369_, _06369_);
  and (_21424_, _21423_, _21422_);
  or (_21425_, _21424_, _06536_);
  or (_21426_, _21425_, _21421_);
  nor (_21427_, _11261_, _11633_);
  or (_21429_, _21427_, _21385_);
  nand (_21430_, _11260_, _08186_);
  and (_21431_, _21430_, _21429_);
  or (_21432_, _21431_, _07240_);
  and (_21433_, _21432_, _07242_);
  and (_21434_, _21433_, _21426_);
  or (_21435_, _14666_, _11633_);
  and (_21436_, _21369_, _06375_);
  and (_21437_, _21436_, _21435_);
  or (_21438_, _21437_, _06545_);
  or (_21440_, _21438_, _21434_);
  nor (_21441_, _21385_, _07234_);
  nand (_21442_, _21441_, _21430_);
  and (_21443_, _21442_, _09056_);
  and (_21444_, _21443_, _21440_);
  or (_21445_, _21371_, _08341_);
  and (_21446_, _21369_, _06366_);
  and (_21447_, _21446_, _21445_);
  or (_21448_, _21447_, _06528_);
  or (_21449_, _21448_, _21444_);
  or (_21451_, _21429_, _09061_);
  and (_21452_, _21451_, _06926_);
  and (_21453_, _21452_, _21449_);
  and (_21454_, _21382_, _06568_);
  or (_21455_, _21454_, _06278_);
  or (_21456_, _21455_, _21453_);
  or (_21457_, _21385_, _06279_);
  or (_21458_, _21457_, _21380_);
  and (_21459_, _21458_, _01347_);
  and (_21460_, _21459_, _21456_);
  or (_21462_, _21460_, _21368_);
  and (_43196_, _21462_, _42618_);
  and (_21463_, _01351_, \oc8051_golden_model_1.DPH [2]);
  and (_21464_, _11633_, \oc8051_golden_model_1.DPH [2]);
  nor (_21465_, _11633_, _07776_);
  or (_21466_, _21465_, _21464_);
  or (_21467_, _21466_, _07215_);
  or (_21468_, _11661_, \oc8051_golden_model_1.DPH [2]);
  nor (_21469_, _11662_, _11562_);
  and (_21470_, _21469_, _21468_);
  and (_21472_, _14770_, _08186_);
  or (_21473_, _21472_, _21464_);
  or (_21474_, _21473_, _07151_);
  and (_21475_, _07963_, \oc8051_golden_model_1.ACC [2]);
  or (_21476_, _21475_, _21464_);
  and (_21477_, _21476_, _07141_);
  and (_21478_, _07142_, \oc8051_golden_model_1.DPH [2]);
  or (_21479_, _21478_, _06341_);
  or (_21480_, _21479_, _21477_);
  and (_21481_, _21480_, _07166_);
  and (_21483_, _21481_, _21474_);
  and (_21484_, _21466_, _06461_);
  or (_21485_, _21484_, _06464_);
  or (_21486_, _21485_, _21483_);
  or (_21487_, _21476_, _06465_);
  and (_21488_, _21487_, _11562_);
  and (_21489_, _21488_, _21486_);
  or (_21490_, _21489_, _21470_);
  and (_21491_, _21490_, _06374_);
  nor (_21492_, _06656_, _06374_);
  or (_21494_, _21492_, _10080_);
  or (_21495_, _21494_, _21491_);
  and (_21496_, _21495_, _21467_);
  or (_21497_, _21496_, _07460_);
  or (_21498_, _21464_, _07208_);
  and (_21499_, _09450_, _07963_);
  or (_21500_, _21499_, _21498_);
  and (_21501_, _21500_, _05982_);
  and (_21502_, _21501_, _21497_);
  and (_21503_, _14859_, _07963_);
  or (_21505_, _21503_, _21464_);
  and (_21506_, _21505_, _10094_);
  or (_21507_, _21506_, _06218_);
  or (_21508_, _21507_, _21502_);
  and (_21509_, _07963_, _08973_);
  or (_21510_, _21509_, _21464_);
  or (_21511_, _21510_, _06219_);
  and (_21512_, _21511_, _21508_);
  or (_21513_, _21512_, _06369_);
  and (_21514_, _14751_, _07963_);
  or (_21516_, _21514_, _21464_);
  or (_21517_, _21516_, _07237_);
  and (_21518_, _21517_, _07240_);
  and (_21519_, _21518_, _21513_);
  and (_21520_, _11259_, _07963_);
  or (_21521_, _21520_, _21464_);
  and (_21522_, _21521_, _06536_);
  or (_21523_, _21522_, _21519_);
  and (_21524_, _21523_, _07242_);
  or (_21525_, _21464_, _08440_);
  and (_21527_, _21510_, _06375_);
  and (_21528_, _21527_, _21525_);
  or (_21529_, _21528_, _21524_);
  and (_21530_, _21529_, _07234_);
  and (_21531_, _21476_, _06545_);
  and (_21532_, _21531_, _21525_);
  or (_21533_, _21532_, _06366_);
  or (_21534_, _21533_, _21530_);
  and (_21535_, _14748_, _08186_);
  or (_21536_, _21464_, _09056_);
  or (_21538_, _21536_, _21535_);
  and (_21539_, _21538_, _09061_);
  and (_21540_, _21539_, _21534_);
  nor (_21541_, _11258_, _11633_);
  or (_21542_, _21541_, _21464_);
  and (_21543_, _21542_, _06528_);
  or (_21544_, _21543_, _21540_);
  and (_21545_, _21544_, _06926_);
  and (_21546_, _21473_, _06568_);
  or (_21547_, _21546_, _06278_);
  or (_21549_, _21547_, _21545_);
  and (_21550_, _14926_, _08186_);
  or (_21551_, _21464_, _06279_);
  or (_21552_, _21551_, _21550_);
  and (_21553_, _21552_, _01347_);
  and (_21554_, _21553_, _21549_);
  or (_21555_, _21554_, _21463_);
  and (_43197_, _21555_, _42618_);
  and (_21556_, _01351_, \oc8051_golden_model_1.DPH [3]);
  and (_21557_, _11633_, \oc8051_golden_model_1.DPH [3]);
  nor (_21559_, _11633_, _07594_);
  or (_21560_, _21559_, _21557_);
  or (_21561_, _21560_, _07215_);
  or (_21562_, _11662_, \oc8051_golden_model_1.DPH [3]);
  nor (_21563_, _11663_, _11562_);
  and (_21564_, _21563_, _21562_);
  and (_21565_, _14953_, _08186_);
  or (_21566_, _21565_, _21557_);
  or (_21567_, _21566_, _07151_);
  and (_21568_, _07963_, \oc8051_golden_model_1.ACC [3]);
  or (_21570_, _21568_, _21557_);
  and (_21571_, _21570_, _07141_);
  and (_21572_, _07142_, \oc8051_golden_model_1.DPH [3]);
  or (_21573_, _21572_, _06341_);
  or (_21574_, _21573_, _21571_);
  and (_21575_, _21574_, _07166_);
  and (_21576_, _21575_, _21567_);
  and (_21577_, _21560_, _06461_);
  or (_21578_, _21577_, _06464_);
  or (_21579_, _21578_, _21576_);
  or (_21581_, _21570_, _06465_);
  and (_21582_, _21581_, _11562_);
  and (_21583_, _21582_, _21579_);
  or (_21584_, _21583_, _21564_);
  and (_21585_, _21584_, _06374_);
  nor (_21586_, _06374_, _06213_);
  or (_21587_, _21586_, _10080_);
  or (_21588_, _21587_, _21585_);
  and (_21589_, _21588_, _21561_);
  or (_21590_, _21589_, _07460_);
  or (_21592_, _21557_, _07208_);
  and (_21593_, _09449_, _07963_);
  or (_21594_, _21593_, _21592_);
  and (_21595_, _21594_, _05982_);
  and (_21596_, _21595_, _21590_);
  and (_21597_, _15048_, _07963_);
  or (_21598_, _21597_, _21557_);
  and (_21599_, _21598_, _10094_);
  or (_21600_, _21599_, _06218_);
  or (_21601_, _21600_, _21596_);
  and (_21603_, _07963_, _08930_);
  or (_21604_, _21603_, _21557_);
  or (_21605_, _21604_, _06219_);
  and (_21606_, _21605_, _21601_);
  or (_21607_, _21606_, _06369_);
  and (_21608_, _14943_, _07963_);
  or (_21609_, _21608_, _21557_);
  or (_21610_, _21609_, _07237_);
  and (_21611_, _21610_, _07240_);
  and (_21612_, _21611_, _21607_);
  and (_21614_, _12577_, _07963_);
  or (_21615_, _21614_, _21557_);
  and (_21616_, _21615_, _06536_);
  or (_21617_, _21616_, _21612_);
  and (_21618_, _21617_, _07242_);
  or (_21619_, _21557_, _08292_);
  and (_21620_, _21604_, _06375_);
  and (_21621_, _21620_, _21619_);
  or (_21622_, _21621_, _21618_);
  and (_21623_, _21622_, _07234_);
  and (_21625_, _21570_, _06545_);
  and (_21626_, _21625_, _21619_);
  or (_21627_, _21626_, _06366_);
  or (_21628_, _21627_, _21623_);
  and (_21629_, _14940_, _08186_);
  or (_21630_, _21557_, _09056_);
  or (_21631_, _21630_, _21629_);
  and (_21632_, _21631_, _09061_);
  and (_21633_, _21632_, _21628_);
  nor (_21634_, _11256_, _11633_);
  or (_21636_, _21634_, _21557_);
  and (_21637_, _21636_, _06528_);
  or (_21638_, _21637_, _21633_);
  and (_21639_, _21638_, _06926_);
  and (_21640_, _21566_, _06568_);
  or (_21641_, _21640_, _06278_);
  or (_21642_, _21641_, _21639_);
  and (_21643_, _15128_, _08186_);
  or (_21644_, _21557_, _06279_);
  or (_21645_, _21644_, _21643_);
  and (_21647_, _21645_, _01347_);
  and (_21648_, _21647_, _21642_);
  or (_21649_, _21648_, _21556_);
  and (_43198_, _21649_, _42618_);
  not (_21650_, \oc8051_golden_model_1.DPH [4]);
  nor (_21651_, _01347_, _21650_);
  nor (_21652_, _07963_, _21650_);
  nor (_21653_, _08541_, _11633_);
  or (_21654_, _21653_, _21652_);
  or (_21655_, _21654_, _07215_);
  and (_21656_, _15162_, _08186_);
  or (_21657_, _21656_, _21652_);
  or (_21658_, _21657_, _07151_);
  and (_21659_, _07963_, \oc8051_golden_model_1.ACC [4]);
  or (_21660_, _21659_, _21652_);
  and (_21661_, _21660_, _07141_);
  nor (_21662_, _07141_, _21650_);
  or (_21663_, _21662_, _06341_);
  or (_21664_, _21663_, _21661_);
  and (_21665_, _21664_, _07166_);
  and (_21668_, _21665_, _21658_);
  and (_21669_, _21654_, _06461_);
  or (_21670_, _21669_, _06464_);
  or (_21671_, _21670_, _21668_);
  or (_21672_, _21660_, _06465_);
  and (_21673_, _21672_, _11562_);
  and (_21674_, _21673_, _21671_);
  or (_21675_, _11663_, \oc8051_golden_model_1.DPH [4]);
  nor (_21676_, _11664_, _11562_);
  and (_21677_, _21676_, _21675_);
  or (_21679_, _21677_, _21674_);
  and (_21680_, _21679_, _06374_);
  nor (_21681_, _06968_, _06374_);
  or (_21682_, _21681_, _10080_);
  or (_21683_, _21682_, _21680_);
  and (_21684_, _21683_, _21655_);
  or (_21685_, _21684_, _07460_);
  or (_21686_, _21652_, _07208_);
  and (_21687_, _09448_, _07963_);
  or (_21688_, _21687_, _21686_);
  and (_21690_, _21688_, _05982_);
  and (_21691_, _21690_, _21685_);
  and (_21692_, _15254_, _07963_);
  or (_21693_, _21692_, _21652_);
  and (_21694_, _21693_, _10094_);
  or (_21695_, _21694_, _06218_);
  or (_21696_, _21695_, _21691_);
  and (_21697_, _08959_, _07963_);
  or (_21698_, _21697_, _21652_);
  or (_21699_, _21698_, _06219_);
  and (_21701_, _21699_, _21696_);
  or (_21702_, _21701_, _06369_);
  and (_21703_, _15269_, _07963_);
  or (_21704_, _21703_, _21652_);
  or (_21705_, _21704_, _07237_);
  and (_21706_, _21705_, _07240_);
  and (_21707_, _21706_, _21702_);
  and (_21708_, _11254_, _07963_);
  or (_21709_, _21708_, _21652_);
  and (_21710_, _21709_, _06536_);
  or (_21712_, _21710_, _21707_);
  and (_21713_, _21712_, _07242_);
  or (_21714_, _21652_, _08544_);
  and (_21715_, _21698_, _06375_);
  and (_21716_, _21715_, _21714_);
  or (_21717_, _21716_, _21713_);
  and (_21718_, _21717_, _07234_);
  and (_21719_, _21660_, _06545_);
  and (_21720_, _21719_, _21714_);
  or (_21721_, _21720_, _06366_);
  or (_21723_, _21721_, _21718_);
  and (_21724_, _15266_, _08186_);
  or (_21725_, _21652_, _09056_);
  or (_21726_, _21725_, _21724_);
  and (_21727_, _21726_, _09061_);
  and (_21728_, _21727_, _21723_);
  nor (_21729_, _11253_, _11633_);
  or (_21730_, _21729_, _21652_);
  and (_21731_, _21730_, _06528_);
  or (_21732_, _21731_, _21728_);
  and (_21734_, _21732_, _06926_);
  and (_21735_, _21657_, _06568_);
  or (_21736_, _21735_, _06278_);
  or (_21737_, _21736_, _21734_);
  and (_21738_, _15329_, _08186_);
  or (_21739_, _21652_, _06279_);
  or (_21740_, _21739_, _21738_);
  and (_21741_, _21740_, _01347_);
  and (_21742_, _21741_, _21737_);
  or (_21743_, _21742_, _21651_);
  and (_43199_, _21743_, _42618_);
  and (_21745_, _01351_, \oc8051_golden_model_1.DPH [5]);
  and (_21746_, _11633_, \oc8051_golden_model_1.DPH [5]);
  nor (_21747_, _08244_, _11633_);
  or (_21748_, _21747_, _21746_);
  or (_21749_, _21748_, _07215_);
  and (_21750_, _15358_, _08186_);
  or (_21751_, _21750_, _21746_);
  or (_21752_, _21751_, _07151_);
  and (_21753_, _07963_, \oc8051_golden_model_1.ACC [5]);
  or (_21755_, _21753_, _21746_);
  and (_21756_, _21755_, _07141_);
  and (_21757_, _07142_, \oc8051_golden_model_1.DPH [5]);
  or (_21758_, _21757_, _06341_);
  or (_21759_, _21758_, _21756_);
  and (_21760_, _21759_, _07166_);
  and (_21761_, _21760_, _21752_);
  and (_21762_, _21748_, _06461_);
  or (_21763_, _21762_, _06464_);
  or (_21764_, _21763_, _21761_);
  or (_21765_, _21755_, _06465_);
  and (_21766_, _21765_, _11562_);
  and (_21767_, _21766_, _21764_);
  or (_21768_, _11664_, \oc8051_golden_model_1.DPH [5]);
  nor (_21769_, _11665_, _11562_);
  and (_21770_, _21769_, _21768_);
  or (_21771_, _21770_, _21767_);
  and (_21772_, _21771_, _06374_);
  nor (_21773_, _06611_, _06374_);
  or (_21774_, _21773_, _10080_);
  or (_21777_, _21774_, _21772_);
  and (_21778_, _21777_, _21749_);
  or (_21779_, _21778_, _07460_);
  or (_21780_, _21746_, _07208_);
  and (_21781_, _09447_, _07963_);
  or (_21782_, _21781_, _21780_);
  and (_21783_, _21782_, _05982_);
  and (_21784_, _21783_, _21779_);
  and (_21785_, _15459_, _07963_);
  or (_21786_, _21785_, _21746_);
  and (_21788_, _21786_, _10094_);
  or (_21789_, _21788_, _06218_);
  or (_21790_, _21789_, _21784_);
  and (_21791_, _08946_, _07963_);
  or (_21792_, _21791_, _21746_);
  or (_21793_, _21792_, _06219_);
  and (_21794_, _21793_, _21790_);
  or (_21795_, _21794_, _06369_);
  and (_21796_, _15353_, _07963_);
  or (_21797_, _21796_, _21746_);
  or (_21799_, _21797_, _07237_);
  and (_21800_, _21799_, _07240_);
  and (_21801_, _21800_, _21795_);
  and (_21802_, _11250_, _07963_);
  or (_21803_, _21802_, _21746_);
  and (_21804_, _21803_, _06536_);
  or (_21805_, _21804_, _21801_);
  and (_21806_, _21805_, _07242_);
  or (_21807_, _21746_, _08247_);
  and (_21808_, _21792_, _06375_);
  and (_21810_, _21808_, _21807_);
  or (_21811_, _21810_, _21806_);
  and (_21812_, _21811_, _07234_);
  and (_21813_, _21755_, _06545_);
  and (_21814_, _21813_, _21807_);
  or (_21815_, _21814_, _06366_);
  or (_21816_, _21815_, _21812_);
  and (_21817_, _15350_, _08186_);
  or (_21818_, _21746_, _09056_);
  or (_21819_, _21818_, _21817_);
  and (_21821_, _21819_, _09061_);
  and (_21822_, _21821_, _21816_);
  nor (_21823_, _11249_, _11633_);
  or (_21824_, _21823_, _21746_);
  and (_21825_, _21824_, _06528_);
  or (_21826_, _21825_, _21822_);
  and (_21827_, _21826_, _06926_);
  and (_21828_, _21751_, _06568_);
  or (_21829_, _21828_, _06278_);
  or (_21830_, _21829_, _21827_);
  and (_21832_, _15532_, _08186_);
  or (_21833_, _21746_, _06279_);
  or (_21834_, _21833_, _21832_);
  and (_21835_, _21834_, _01347_);
  and (_21836_, _21835_, _21830_);
  or (_21837_, _21836_, _21745_);
  and (_43200_, _21837_, _42618_);
  not (_21838_, \oc8051_golden_model_1.DPH [6]);
  nor (_21839_, _01347_, _21838_);
  nor (_21840_, _07963_, _21838_);
  nor (_21842_, _08142_, _11633_);
  or (_21843_, _21842_, _21840_);
  or (_21844_, _21843_, _07215_);
  and (_21845_, _15554_, _08186_);
  or (_21846_, _21845_, _21840_);
  or (_21847_, _21846_, _07151_);
  and (_21848_, _07963_, \oc8051_golden_model_1.ACC [6]);
  or (_21849_, _21848_, _21840_);
  and (_21850_, _21849_, _07141_);
  nor (_21851_, _07141_, _21838_);
  or (_21853_, _21851_, _06341_);
  or (_21854_, _21853_, _21850_);
  and (_21855_, _21854_, _07166_);
  and (_21856_, _21855_, _21847_);
  and (_21857_, _21843_, _06461_);
  or (_21858_, _21857_, _06464_);
  or (_21859_, _21858_, _21856_);
  or (_21860_, _21849_, _06465_);
  and (_21861_, _21860_, _11562_);
  and (_21862_, _21861_, _21859_);
  or (_21864_, _11665_, \oc8051_golden_model_1.DPH [6]);
  nor (_21865_, _11666_, _11562_);
  and (_21866_, _21865_, _21864_);
  or (_21867_, _21866_, _21862_);
  and (_21868_, _21867_, _06374_);
  nor (_21869_, _06374_, _06317_);
  or (_21870_, _21869_, _10080_);
  or (_21871_, _21870_, _21868_);
  and (_21872_, _21871_, _21844_);
  or (_21873_, _21872_, _07460_);
  or (_21875_, _21840_, _07208_);
  and (_21876_, _09446_, _07963_);
  or (_21877_, _21876_, _21875_);
  and (_21878_, _21877_, _05982_);
  and (_21879_, _21878_, _21873_);
  and (_21880_, _15657_, _07963_);
  or (_21881_, _21880_, _21840_);
  and (_21882_, _21881_, _10094_);
  or (_21883_, _21882_, _06218_);
  or (_21884_, _21883_, _21879_);
  and (_21886_, _15664_, _07963_);
  or (_21887_, _21886_, _21840_);
  or (_21888_, _21887_, _06219_);
  and (_21889_, _21888_, _21884_);
  or (_21890_, _21889_, _06369_);
  and (_21891_, _15549_, _07963_);
  or (_21892_, _21891_, _21840_);
  or (_21893_, _21892_, _07237_);
  and (_21894_, _21893_, _07240_);
  and (_21895_, _21894_, _21890_);
  and (_21897_, _11247_, _07963_);
  or (_21898_, _21897_, _21840_);
  and (_21899_, _21898_, _06536_);
  or (_21900_, _21899_, _21895_);
  and (_21901_, _21900_, _07242_);
  or (_21902_, _21840_, _08145_);
  and (_21903_, _21887_, _06375_);
  and (_21904_, _21903_, _21902_);
  or (_21905_, _21904_, _21901_);
  and (_21906_, _21905_, _07234_);
  and (_21908_, _21849_, _06545_);
  and (_21909_, _21908_, _21902_);
  or (_21910_, _21909_, _06366_);
  or (_21911_, _21910_, _21906_);
  and (_21912_, _15546_, _08186_);
  or (_21913_, _21840_, _09056_);
  or (_21914_, _21913_, _21912_);
  and (_21915_, _21914_, _09061_);
  and (_21916_, _21915_, _21911_);
  nor (_21917_, _11246_, _11633_);
  or (_21919_, _21917_, _21840_);
  and (_21920_, _21919_, _06528_);
  or (_21921_, _21920_, _21916_);
  and (_21922_, _21921_, _06926_);
  and (_21923_, _21846_, _06568_);
  or (_21924_, _21923_, _06278_);
  or (_21925_, _21924_, _21922_);
  and (_21926_, _15734_, _08186_);
  or (_21927_, _21840_, _06279_);
  or (_21928_, _21927_, _21926_);
  and (_21930_, _21928_, _01347_);
  and (_21931_, _21930_, _21925_);
  or (_21932_, _21931_, _21839_);
  and (_43201_, _21932_, _42618_);
  not (_21933_, \oc8051_golden_model_1.TL1 [0]);
  nor (_21934_, _01347_, _21933_);
  nand (_21935_, _11263_, _07968_);
  nor (_21936_, _07968_, _21933_);
  nor (_21937_, _21936_, _07234_);
  nand (_21938_, _21937_, _21935_);
  and (_21940_, _07968_, _07133_);
  or (_21941_, _21940_, _21936_);
  or (_21942_, _21941_, _07215_);
  nor (_21943_, _08390_, _11726_);
  or (_21944_, _21943_, _21936_);
  or (_21945_, _21944_, _07151_);
  and (_21946_, _07968_, \oc8051_golden_model_1.ACC [0]);
  or (_21947_, _21946_, _21936_);
  and (_21948_, _21947_, _07141_);
  nor (_21949_, _07141_, _21933_);
  or (_21951_, _21949_, _06341_);
  or (_21952_, _21951_, _21948_);
  and (_21953_, _21952_, _07166_);
  and (_21954_, _21953_, _21945_);
  and (_21955_, _21941_, _06461_);
  or (_21956_, _21955_, _21954_);
  and (_21957_, _21956_, _06465_);
  and (_21958_, _21947_, _06464_);
  or (_21959_, _21958_, _10080_);
  or (_21960_, _21959_, _21957_);
  and (_21962_, _21960_, _21942_);
  or (_21963_, _21962_, _07460_);
  and (_21964_, _09392_, _07968_);
  or (_21965_, _21936_, _07208_);
  or (_21966_, _21965_, _21964_);
  and (_21967_, _21966_, _21963_);
  or (_21968_, _21967_, _10094_);
  and (_21969_, _14467_, _07968_);
  or (_21970_, _21936_, _05982_);
  or (_21971_, _21970_, _21969_);
  and (_21973_, _21971_, _06219_);
  and (_21974_, _21973_, _21968_);
  and (_21975_, _07968_, _08954_);
  or (_21976_, _21975_, _21936_);
  and (_21977_, _21976_, _06218_);
  or (_21978_, _21977_, _06369_);
  or (_21979_, _21978_, _21974_);
  and (_21980_, _14366_, _07968_);
  or (_21981_, _21980_, _21936_);
  or (_21982_, _21981_, _07237_);
  and (_21984_, _21982_, _07240_);
  and (_21985_, _21984_, _21979_);
  nor (_21986_, _12580_, _11726_);
  or (_21987_, _21986_, _21936_);
  and (_21988_, _21935_, _06536_);
  and (_21989_, _21988_, _21987_);
  or (_21990_, _21989_, _21985_);
  and (_21991_, _21990_, _07242_);
  nand (_21992_, _21976_, _06375_);
  nor (_21993_, _21992_, _21943_);
  or (_21995_, _21993_, _06545_);
  or (_21996_, _21995_, _21991_);
  and (_21997_, _21996_, _21938_);
  or (_21998_, _21997_, _06366_);
  and (_21999_, _14363_, _07968_);
  or (_22000_, _21936_, _09056_);
  or (_22001_, _22000_, _21999_);
  and (_22002_, _22001_, _09061_);
  and (_22003_, _22002_, _21998_);
  and (_22004_, _21987_, _06528_);
  or (_22006_, _22004_, _19502_);
  or (_22007_, _22006_, _22003_);
  or (_22008_, _21944_, _06661_);
  and (_22009_, _22008_, _01347_);
  and (_22010_, _22009_, _22007_);
  or (_22011_, _22010_, _21934_);
  and (_43202_, _22011_, _42618_);
  not (_22012_, \oc8051_golden_model_1.TL1 [1]);
  nor (_22013_, _01347_, _22012_);
  or (_22014_, _07968_, \oc8051_golden_model_1.TL1 [1]);
  and (_22016_, _14562_, _07968_);
  not (_22017_, _22016_);
  and (_22018_, _22017_, _22014_);
  or (_22019_, _22018_, _07151_);
  nor (_22020_, _07968_, _22012_);
  and (_22021_, _07968_, \oc8051_golden_model_1.ACC [1]);
  or (_22022_, _22021_, _22020_);
  and (_22023_, _22022_, _07141_);
  nor (_22024_, _07141_, _22012_);
  or (_22025_, _22024_, _06341_);
  or (_22027_, _22025_, _22023_);
  and (_22028_, _22027_, _07166_);
  and (_22029_, _22028_, _22019_);
  nor (_22030_, _11726_, _07357_);
  or (_22031_, _22030_, _22020_);
  and (_22032_, _22031_, _06461_);
  or (_22033_, _22032_, _22029_);
  and (_22034_, _22033_, _06465_);
  and (_22035_, _22022_, _06464_);
  or (_22036_, _22035_, _10080_);
  or (_22038_, _22036_, _22034_);
  or (_22039_, _22031_, _07215_);
  and (_22040_, _22039_, _22038_);
  or (_22041_, _22040_, _07460_);
  and (_22042_, _09451_, _07968_);
  or (_22043_, _22020_, _07208_);
  or (_22044_, _22043_, _22042_);
  and (_22045_, _22044_, _05982_);
  and (_22046_, _22045_, _22041_);
  or (_22047_, _14653_, _11726_);
  and (_22049_, _22014_, _10094_);
  and (_22050_, _22049_, _22047_);
  or (_22051_, _22050_, _22046_);
  and (_22052_, _22051_, _06219_);
  nand (_22053_, _07968_, _07038_);
  and (_22054_, _22014_, _06218_);
  and (_22055_, _22054_, _22053_);
  or (_22056_, _22055_, _22052_);
  and (_22057_, _22056_, _07237_);
  or (_22058_, _14668_, _11726_);
  and (_22060_, _22014_, _06369_);
  and (_22061_, _22060_, _22058_);
  or (_22062_, _22061_, _06536_);
  or (_22063_, _22062_, _22057_);
  nor (_22064_, _11261_, _11726_);
  or (_22065_, _22064_, _22020_);
  nand (_22066_, _11260_, _07968_);
  and (_22067_, _22066_, _22065_);
  or (_22068_, _22067_, _07240_);
  and (_22069_, _22068_, _07242_);
  and (_22071_, _22069_, _22063_);
  or (_22072_, _14666_, _11726_);
  and (_22073_, _22014_, _06375_);
  and (_22074_, _22073_, _22072_);
  or (_22075_, _22074_, _06545_);
  or (_22076_, _22075_, _22071_);
  nor (_22077_, _22020_, _07234_);
  nand (_22078_, _22077_, _22066_);
  and (_22079_, _22078_, _09056_);
  and (_22080_, _22079_, _22076_);
  or (_22082_, _22053_, _08341_);
  and (_22083_, _22014_, _06366_);
  and (_22084_, _22083_, _22082_);
  or (_22085_, _22084_, _06528_);
  or (_22086_, _22085_, _22080_);
  or (_22087_, _22065_, _09061_);
  and (_22088_, _22087_, _06926_);
  and (_22089_, _22088_, _22086_);
  and (_22090_, _22018_, _06568_);
  or (_22091_, _22090_, _06278_);
  or (_22093_, _22091_, _22089_);
  or (_22094_, _22020_, _06279_);
  or (_22095_, _22094_, _22016_);
  and (_22096_, _22095_, _01347_);
  and (_22097_, _22096_, _22093_);
  or (_22098_, _22097_, _22013_);
  and (_43204_, _22098_, _42618_);
  and (_22099_, _01351_, \oc8051_golden_model_1.TL1 [2]);
  and (_22100_, _11726_, \oc8051_golden_model_1.TL1 [2]);
  nor (_22101_, _11726_, _07776_);
  or (_22103_, _22101_, _22100_);
  or (_22104_, _22103_, _07215_);
  and (_22105_, _14770_, _07968_);
  or (_22106_, _22105_, _22100_);
  and (_22107_, _22106_, _06341_);
  and (_22108_, _07142_, \oc8051_golden_model_1.TL1 [2]);
  and (_22109_, _07968_, \oc8051_golden_model_1.ACC [2]);
  or (_22110_, _22109_, _22100_);
  and (_22111_, _22110_, _07141_);
  or (_22112_, _22111_, _22108_);
  and (_22114_, _22112_, _07151_);
  or (_22115_, _22114_, _06461_);
  or (_22116_, _22115_, _22107_);
  or (_22117_, _22103_, _07166_);
  and (_22118_, _22117_, _06465_);
  and (_22119_, _22118_, _22116_);
  and (_22120_, _22110_, _06464_);
  or (_22121_, _22120_, _10080_);
  or (_22122_, _22121_, _22119_);
  and (_22123_, _22122_, _22104_);
  or (_22126_, _22123_, _07460_);
  and (_22127_, _09450_, _07968_);
  or (_22128_, _22100_, _07208_);
  or (_22129_, _22128_, _22127_);
  and (_22130_, _22129_, _22126_);
  or (_22131_, _22130_, _10094_);
  and (_22132_, _14859_, _07968_);
  or (_22133_, _22100_, _05982_);
  or (_22134_, _22133_, _22132_);
  and (_22135_, _22134_, _06219_);
  and (_22137_, _22135_, _22131_);
  and (_22138_, _07968_, _08973_);
  or (_22139_, _22138_, _22100_);
  and (_22140_, _22139_, _06218_);
  or (_22141_, _22140_, _06369_);
  or (_22142_, _22141_, _22137_);
  and (_22143_, _14751_, _07968_);
  or (_22144_, _22143_, _22100_);
  or (_22145_, _22144_, _07237_);
  and (_22146_, _22145_, _07240_);
  and (_22148_, _22146_, _22142_);
  and (_22149_, _11259_, _07968_);
  or (_22150_, _22149_, _22100_);
  and (_22151_, _22150_, _06536_);
  or (_22152_, _22151_, _22148_);
  and (_22153_, _22152_, _07242_);
  or (_22154_, _22100_, _08440_);
  and (_22155_, _22139_, _06375_);
  and (_22156_, _22155_, _22154_);
  or (_22157_, _22156_, _22153_);
  and (_22159_, _22157_, _07234_);
  and (_22160_, _22110_, _06545_);
  and (_22161_, _22160_, _22154_);
  or (_22162_, _22161_, _06366_);
  or (_22163_, _22162_, _22159_);
  and (_22164_, _14748_, _07968_);
  or (_22165_, _22100_, _09056_);
  or (_22166_, _22165_, _22164_);
  and (_22167_, _22166_, _09061_);
  and (_22168_, _22167_, _22163_);
  nor (_22170_, _11258_, _11726_);
  or (_22171_, _22170_, _22100_);
  and (_22172_, _22171_, _06528_);
  or (_22173_, _22172_, _22168_);
  and (_22174_, _22173_, _06926_);
  and (_22175_, _22106_, _06568_);
  or (_22176_, _22175_, _06278_);
  or (_22177_, _22176_, _22174_);
  and (_22178_, _14926_, _07968_);
  or (_22179_, _22100_, _06279_);
  or (_22181_, _22179_, _22178_);
  and (_22182_, _22181_, _01347_);
  and (_22183_, _22182_, _22177_);
  or (_22184_, _22183_, _22099_);
  and (_43205_, _22184_, _42618_);
  and (_22185_, _01351_, \oc8051_golden_model_1.TL1 [3]);
  and (_22186_, _11726_, \oc8051_golden_model_1.TL1 [3]);
  and (_22187_, _14953_, _07968_);
  or (_22188_, _22187_, _22186_);
  or (_22189_, _22188_, _07151_);
  and (_22191_, _07968_, \oc8051_golden_model_1.ACC [3]);
  or (_22192_, _22191_, _22186_);
  and (_22193_, _22192_, _07141_);
  and (_22194_, _07142_, \oc8051_golden_model_1.TL1 [3]);
  or (_22195_, _22194_, _06341_);
  or (_22196_, _22195_, _22193_);
  and (_22197_, _22196_, _07166_);
  and (_22198_, _22197_, _22189_);
  nor (_22199_, _11726_, _07594_);
  or (_22200_, _22199_, _22186_);
  and (_22202_, _22200_, _06461_);
  or (_22203_, _22202_, _22198_);
  and (_22204_, _22203_, _06465_);
  and (_22205_, _22192_, _06464_);
  or (_22206_, _22205_, _10080_);
  or (_22207_, _22206_, _22204_);
  or (_22208_, _22200_, _07215_);
  and (_22209_, _22208_, _22207_);
  or (_22210_, _22209_, _07460_);
  and (_22211_, _09449_, _07968_);
  or (_22212_, _22186_, _07208_);
  or (_22213_, _22212_, _22211_);
  and (_22214_, _22213_, _05982_);
  and (_22215_, _22214_, _22210_);
  and (_22216_, _15048_, _07968_);
  or (_22217_, _22216_, _22186_);
  and (_22218_, _22217_, _10094_);
  or (_22219_, _22218_, _06218_);
  or (_22220_, _22219_, _22215_);
  and (_22221_, _07968_, _08930_);
  or (_22224_, _22221_, _22186_);
  or (_22225_, _22224_, _06219_);
  and (_22226_, _22225_, _22220_);
  or (_22227_, _22226_, _06369_);
  and (_22228_, _14943_, _07968_);
  or (_22229_, _22228_, _22186_);
  or (_22230_, _22229_, _07237_);
  and (_22231_, _22230_, _07240_);
  and (_22232_, _22231_, _22227_);
  and (_22233_, _12577_, _07968_);
  or (_22235_, _22233_, _22186_);
  and (_22236_, _22235_, _06536_);
  or (_22237_, _22236_, _22232_);
  and (_22238_, _22237_, _07242_);
  or (_22239_, _22186_, _08292_);
  and (_22240_, _22224_, _06375_);
  and (_22241_, _22240_, _22239_);
  or (_22242_, _22241_, _22238_);
  and (_22243_, _22242_, _07234_);
  and (_22244_, _22192_, _06545_);
  and (_22246_, _22244_, _22239_);
  or (_22247_, _22246_, _06366_);
  or (_22248_, _22247_, _22243_);
  and (_22249_, _14940_, _07968_);
  or (_22250_, _22186_, _09056_);
  or (_22251_, _22250_, _22249_);
  and (_22252_, _22251_, _09061_);
  and (_22253_, _22252_, _22248_);
  nor (_22254_, _11256_, _11726_);
  or (_22255_, _22254_, _22186_);
  and (_22257_, _22255_, _06528_);
  or (_22258_, _22257_, _22253_);
  and (_22259_, _22258_, _06926_);
  and (_22260_, _22188_, _06568_);
  or (_22261_, _22260_, _06278_);
  or (_22262_, _22261_, _22259_);
  and (_22263_, _15128_, _07968_);
  or (_22264_, _22186_, _06279_);
  or (_22265_, _22264_, _22263_);
  and (_22266_, _22265_, _01347_);
  and (_22268_, _22266_, _22262_);
  or (_22269_, _22268_, _22185_);
  and (_43206_, _22269_, _42618_);
  and (_22270_, _01351_, \oc8051_golden_model_1.TL1 [4]);
  and (_22271_, _11726_, \oc8051_golden_model_1.TL1 [4]);
  and (_22272_, _15162_, _07968_);
  or (_22273_, _22272_, _22271_);
  or (_22274_, _22273_, _07151_);
  and (_22275_, _07968_, \oc8051_golden_model_1.ACC [4]);
  or (_22276_, _22275_, _22271_);
  and (_22278_, _22276_, _07141_);
  and (_22279_, _07142_, \oc8051_golden_model_1.TL1 [4]);
  or (_22280_, _22279_, _06341_);
  or (_22281_, _22280_, _22278_);
  and (_22282_, _22281_, _07166_);
  and (_22283_, _22282_, _22274_);
  nor (_22284_, _08541_, _11726_);
  or (_22285_, _22284_, _22271_);
  and (_22286_, _22285_, _06461_);
  or (_22287_, _22286_, _22283_);
  and (_22289_, _22287_, _06465_);
  and (_22290_, _22276_, _06464_);
  or (_22291_, _22290_, _10080_);
  or (_22292_, _22291_, _22289_);
  or (_22293_, _22285_, _07215_);
  and (_22294_, _22293_, _22292_);
  or (_22295_, _22294_, _07460_);
  and (_22296_, _09448_, _07968_);
  or (_22297_, _22271_, _07208_);
  or (_22298_, _22297_, _22296_);
  and (_22300_, _22298_, _22295_);
  or (_22301_, _22300_, _10094_);
  and (_22302_, _15254_, _07968_);
  or (_22303_, _22271_, _05982_);
  or (_22304_, _22303_, _22302_);
  and (_22305_, _22304_, _06219_);
  and (_22306_, _22305_, _22301_);
  and (_22307_, _08959_, _07968_);
  or (_22308_, _22307_, _22271_);
  and (_22309_, _22308_, _06218_);
  or (_22311_, _22309_, _06369_);
  or (_22312_, _22311_, _22306_);
  and (_22313_, _15269_, _07968_);
  or (_22314_, _22313_, _22271_);
  or (_22315_, _22314_, _07237_);
  and (_22316_, _22315_, _07240_);
  and (_22317_, _22316_, _22312_);
  and (_22318_, _11254_, _07968_);
  or (_22319_, _22318_, _22271_);
  and (_22320_, _22319_, _06536_);
  or (_22322_, _22320_, _22317_);
  and (_22323_, _22322_, _07242_);
  or (_22324_, _22271_, _08544_);
  and (_22325_, _22308_, _06375_);
  and (_22326_, _22325_, _22324_);
  or (_22327_, _22326_, _22323_);
  and (_22328_, _22327_, _07234_);
  and (_22329_, _22276_, _06545_);
  and (_22330_, _22329_, _22324_);
  or (_22331_, _22330_, _06366_);
  or (_22333_, _22331_, _22328_);
  and (_22334_, _15266_, _07968_);
  or (_22335_, _22271_, _09056_);
  or (_22336_, _22335_, _22334_);
  and (_22337_, _22336_, _09061_);
  and (_22338_, _22337_, _22333_);
  nor (_22339_, _11253_, _11726_);
  or (_22340_, _22339_, _22271_);
  and (_22341_, _22340_, _06528_);
  or (_22342_, _22341_, _22338_);
  and (_22344_, _22342_, _06926_);
  and (_22345_, _22273_, _06568_);
  or (_22346_, _22345_, _06278_);
  or (_22347_, _22346_, _22344_);
  and (_22348_, _15329_, _07968_);
  or (_22349_, _22271_, _06279_);
  or (_22350_, _22349_, _22348_);
  and (_22351_, _22350_, _01347_);
  and (_22352_, _22351_, _22347_);
  or (_22353_, _22352_, _22270_);
  and (_43207_, _22353_, _42618_);
  and (_22355_, _01351_, \oc8051_golden_model_1.TL1 [5]);
  and (_22356_, _11726_, \oc8051_golden_model_1.TL1 [5]);
  nor (_22357_, _08244_, _11726_);
  or (_22358_, _22357_, _22356_);
  or (_22359_, _22358_, _07215_);
  and (_22360_, _15358_, _07968_);
  or (_22361_, _22360_, _22356_);
  or (_22362_, _22361_, _07151_);
  and (_22363_, _07968_, \oc8051_golden_model_1.ACC [5]);
  or (_22365_, _22363_, _22356_);
  and (_22366_, _22365_, _07141_);
  and (_22367_, _07142_, \oc8051_golden_model_1.TL1 [5]);
  or (_22368_, _22367_, _06341_);
  or (_22369_, _22368_, _22366_);
  and (_22370_, _22369_, _07166_);
  and (_22371_, _22370_, _22362_);
  and (_22372_, _22358_, _06461_);
  or (_22373_, _22372_, _22371_);
  and (_22374_, _22373_, _06465_);
  and (_22376_, _22365_, _06464_);
  or (_22377_, _22376_, _10080_);
  or (_22378_, _22377_, _22374_);
  and (_22379_, _22378_, _22359_);
  or (_22380_, _22379_, _07460_);
  and (_22381_, _09447_, _07968_);
  or (_22382_, _22356_, _07208_);
  or (_22383_, _22382_, _22381_);
  and (_22384_, _22383_, _05982_);
  and (_22385_, _22384_, _22380_);
  and (_22387_, _15459_, _07968_);
  or (_22388_, _22387_, _22356_);
  and (_22389_, _22388_, _10094_);
  or (_22390_, _22389_, _06218_);
  or (_22391_, _22390_, _22385_);
  and (_22392_, _08946_, _07968_);
  or (_22393_, _22392_, _22356_);
  or (_22394_, _22393_, _06219_);
  and (_22395_, _22394_, _22391_);
  or (_22396_, _22395_, _06369_);
  and (_22398_, _15353_, _07968_);
  or (_22399_, _22398_, _22356_);
  or (_22400_, _22399_, _07237_);
  and (_22401_, _22400_, _07240_);
  and (_22402_, _22401_, _22396_);
  and (_22403_, _11250_, _07968_);
  or (_22404_, _22403_, _22356_);
  and (_22405_, _22404_, _06536_);
  or (_22406_, _22405_, _22402_);
  and (_22407_, _22406_, _07242_);
  or (_22409_, _22356_, _08247_);
  and (_22410_, _22393_, _06375_);
  and (_22411_, _22410_, _22409_);
  or (_22412_, _22411_, _22407_);
  and (_22413_, _22412_, _07234_);
  and (_22414_, _22365_, _06545_);
  and (_22415_, _22414_, _22409_);
  or (_22416_, _22415_, _06366_);
  or (_22417_, _22416_, _22413_);
  and (_22418_, _15350_, _07968_);
  or (_22420_, _22356_, _09056_);
  or (_22421_, _22420_, _22418_);
  and (_22422_, _22421_, _09061_);
  and (_22423_, _22422_, _22417_);
  nor (_22424_, _11249_, _11726_);
  or (_22425_, _22424_, _22356_);
  and (_22426_, _22425_, _06528_);
  or (_22427_, _22426_, _22423_);
  and (_22428_, _22427_, _06926_);
  and (_22429_, _22361_, _06568_);
  or (_22431_, _22429_, _06278_);
  or (_22432_, _22431_, _22428_);
  and (_22433_, _15532_, _07968_);
  or (_22434_, _22356_, _06279_);
  or (_22435_, _22434_, _22433_);
  and (_22436_, _22435_, _01347_);
  and (_22437_, _22436_, _22432_);
  or (_22438_, _22437_, _22355_);
  and (_43208_, _22438_, _42618_);
  and (_22439_, _01351_, \oc8051_golden_model_1.TL1 [6]);
  and (_22441_, _11726_, \oc8051_golden_model_1.TL1 [6]);
  and (_22442_, _15554_, _07968_);
  or (_22443_, _22442_, _22441_);
  or (_22444_, _22443_, _07151_);
  and (_22445_, _07968_, \oc8051_golden_model_1.ACC [6]);
  or (_22446_, _22445_, _22441_);
  and (_22447_, _22446_, _07141_);
  and (_22448_, _07142_, \oc8051_golden_model_1.TL1 [6]);
  or (_22449_, _22448_, _06341_);
  or (_22450_, _22449_, _22447_);
  and (_22452_, _22450_, _07166_);
  and (_22453_, _22452_, _22444_);
  nor (_22454_, _08142_, _11726_);
  or (_22455_, _22454_, _22441_);
  and (_22456_, _22455_, _06461_);
  or (_22457_, _22456_, _22453_);
  and (_22458_, _22457_, _06465_);
  and (_22459_, _22446_, _06464_);
  or (_22460_, _22459_, _10080_);
  or (_22461_, _22460_, _22458_);
  or (_22463_, _22455_, _07215_);
  and (_22464_, _22463_, _22461_);
  or (_22465_, _22464_, _07460_);
  and (_22466_, _09446_, _07968_);
  or (_22467_, _22441_, _07208_);
  or (_22468_, _22467_, _22466_);
  and (_22469_, _22468_, _05982_);
  and (_22470_, _22469_, _22465_);
  and (_22471_, _15657_, _07968_);
  or (_22472_, _22471_, _22441_);
  and (_22474_, _22472_, _10094_);
  or (_22475_, _22474_, _06218_);
  or (_22476_, _22475_, _22470_);
  and (_22477_, _15664_, _07968_);
  or (_22478_, _22477_, _22441_);
  or (_22479_, _22478_, _06219_);
  and (_22480_, _22479_, _22476_);
  or (_22481_, _22480_, _06369_);
  and (_22482_, _15549_, _07968_);
  or (_22483_, _22482_, _22441_);
  or (_22485_, _22483_, _07237_);
  and (_22486_, _22485_, _07240_);
  and (_22487_, _22486_, _22481_);
  and (_22488_, _11247_, _07968_);
  or (_22489_, _22488_, _22441_);
  and (_22490_, _22489_, _06536_);
  or (_22491_, _22490_, _22487_);
  and (_22492_, _22491_, _07242_);
  or (_22493_, _22441_, _08145_);
  and (_22494_, _22478_, _06375_);
  and (_22496_, _22494_, _22493_);
  or (_22497_, _22496_, _22492_);
  and (_22498_, _22497_, _07234_);
  and (_22499_, _22446_, _06545_);
  and (_22500_, _22499_, _22493_);
  or (_22501_, _22500_, _06366_);
  or (_22502_, _22501_, _22498_);
  and (_22503_, _15546_, _07968_);
  or (_22504_, _22441_, _09056_);
  or (_22505_, _22504_, _22503_);
  and (_22506_, _22505_, _09061_);
  and (_22507_, _22506_, _22502_);
  nor (_22508_, _11246_, _11726_);
  or (_22509_, _22508_, _22441_);
  and (_22510_, _22509_, _06528_);
  or (_22511_, _22510_, _22507_);
  and (_22512_, _22511_, _06926_);
  and (_22513_, _22443_, _06568_);
  or (_22514_, _22513_, _06278_);
  or (_22515_, _22514_, _22512_);
  and (_22518_, _15734_, _07968_);
  or (_22519_, _22441_, _06279_);
  or (_22520_, _22519_, _22518_);
  and (_22521_, _22520_, _01347_);
  and (_22522_, _22521_, _22515_);
  or (_22523_, _22522_, _22439_);
  and (_43209_, _22523_, _42618_);
  not (_22524_, \oc8051_golden_model_1.TL0 [0]);
  nor (_22525_, _01347_, _22524_);
  nand (_22526_, _11263_, _07919_);
  nor (_22528_, _07919_, _22524_);
  nor (_22529_, _22528_, _07234_);
  nand (_22530_, _22529_, _22526_);
  nor (_22531_, _08390_, _11804_);
  or (_22532_, _22531_, _22528_);
  or (_22533_, _22532_, _07151_);
  and (_22534_, _07919_, \oc8051_golden_model_1.ACC [0]);
  or (_22535_, _22534_, _22528_);
  and (_22536_, _22535_, _07141_);
  nor (_22537_, _07141_, _22524_);
  or (_22539_, _22537_, _06341_);
  or (_22540_, _22539_, _22536_);
  and (_22541_, _22540_, _07166_);
  and (_22542_, _22541_, _22533_);
  and (_22543_, _07919_, _07133_);
  or (_22544_, _22543_, _22528_);
  and (_22545_, _22544_, _06461_);
  or (_22546_, _22545_, _22542_);
  and (_22547_, _22546_, _06465_);
  and (_22548_, _22535_, _06464_);
  or (_22550_, _22548_, _10080_);
  or (_22551_, _22550_, _22547_);
  or (_22552_, _22544_, _07215_);
  and (_22553_, _22552_, _22551_);
  or (_22554_, _22553_, _07460_);
  and (_22555_, _09392_, _07919_);
  or (_22556_, _22528_, _07208_);
  or (_22557_, _22556_, _22555_);
  and (_22558_, _22557_, _22554_);
  or (_22559_, _22558_, _10094_);
  and (_22561_, _14467_, _07919_);
  or (_22562_, _22528_, _05982_);
  or (_22563_, _22562_, _22561_);
  and (_22564_, _22563_, _06219_);
  and (_22565_, _22564_, _22559_);
  and (_22566_, _07919_, _08954_);
  or (_22567_, _22566_, _22528_);
  and (_22568_, _22567_, _06218_);
  or (_22569_, _22568_, _06369_);
  or (_22570_, _22569_, _22565_);
  and (_22572_, _14366_, _07919_);
  or (_22573_, _22572_, _22528_);
  or (_22574_, _22573_, _07237_);
  and (_22575_, _22574_, _07240_);
  and (_22576_, _22575_, _22570_);
  nor (_22577_, _12580_, _11804_);
  or (_22578_, _22577_, _22528_);
  and (_22579_, _22526_, _06536_);
  and (_22580_, _22579_, _22578_);
  or (_22581_, _22580_, _22576_);
  and (_22583_, _22581_, _07242_);
  nand (_22584_, _22567_, _06375_);
  nor (_22585_, _22584_, _22531_);
  or (_22586_, _22585_, _06545_);
  or (_22587_, _22586_, _22583_);
  and (_22588_, _22587_, _22530_);
  or (_22589_, _22588_, _06366_);
  and (_22590_, _14363_, _07919_);
  or (_22591_, _22528_, _09056_);
  or (_22592_, _22591_, _22590_);
  and (_22594_, _22592_, _09061_);
  and (_22595_, _22594_, _22589_);
  and (_22596_, _22578_, _06528_);
  or (_22597_, _22596_, _19502_);
  or (_22598_, _22597_, _22595_);
  or (_22599_, _22532_, _06661_);
  and (_22600_, _22599_, _01347_);
  and (_22601_, _22600_, _22598_);
  or (_22602_, _22601_, _22525_);
  and (_43211_, _22602_, _42618_);
  not (_22604_, \oc8051_golden_model_1.TL0 [1]);
  nor (_22605_, _01347_, _22604_);
  and (_22606_, _09451_, _07919_);
  nor (_22607_, _07919_, _22604_);
  or (_22608_, _22607_, _07208_);
  or (_22609_, _22608_, _22606_);
  nor (_22610_, _11804_, _07357_);
  and (_22611_, _07215_, _07166_);
  or (_22612_, _22611_, _22607_);
  or (_22613_, _22612_, _22610_);
  and (_22614_, _07919_, \oc8051_golden_model_1.ACC [1]);
  or (_22615_, _22614_, _22607_);
  and (_22616_, _22615_, _06464_);
  or (_22617_, _22616_, _10080_);
  or (_22618_, _07919_, \oc8051_golden_model_1.TL0 [1]);
  and (_22619_, _14562_, _07919_);
  not (_22620_, _22619_);
  and (_22621_, _22620_, _22618_);
  and (_22622_, _22621_, _06341_);
  nor (_22623_, _07141_, _22604_);
  and (_22626_, _22615_, _07141_);
  or (_22627_, _22626_, _22623_);
  and (_22628_, _22627_, _07151_);
  or (_22629_, _22628_, _06461_);
  or (_22630_, _22629_, _22622_);
  and (_22631_, _22630_, _06465_);
  or (_22632_, _22631_, _22617_);
  and (_22633_, _22632_, _22613_);
  or (_22634_, _22633_, _07460_);
  and (_22635_, _22634_, _05982_);
  and (_22637_, _22635_, _22609_);
  or (_22638_, _14653_, _11804_);
  and (_22639_, _22618_, _10094_);
  and (_22640_, _22639_, _22638_);
  or (_22641_, _22640_, _22637_);
  and (_22642_, _22641_, _06219_);
  nand (_22643_, _07919_, _07038_);
  and (_22644_, _22618_, _06218_);
  and (_22645_, _22644_, _22643_);
  or (_22646_, _22645_, _22642_);
  and (_22648_, _22646_, _07237_);
  or (_22649_, _14668_, _11804_);
  and (_22650_, _22618_, _06369_);
  and (_22651_, _22650_, _22649_);
  or (_22652_, _22651_, _06536_);
  or (_22653_, _22652_, _22648_);
  nor (_22654_, _11261_, _11804_);
  or (_22655_, _22654_, _22607_);
  nand (_22656_, _11260_, _07919_);
  and (_22657_, _22656_, _22655_);
  or (_22659_, _22657_, _07240_);
  and (_22660_, _22659_, _07242_);
  and (_22661_, _22660_, _22653_);
  or (_22662_, _14666_, _11804_);
  and (_22663_, _22618_, _06375_);
  and (_22664_, _22663_, _22662_);
  or (_22665_, _22664_, _06545_);
  or (_22666_, _22665_, _22661_);
  nor (_22667_, _22607_, _07234_);
  nand (_22668_, _22667_, _22656_);
  and (_22670_, _22668_, _09056_);
  and (_22671_, _22670_, _22666_);
  or (_22672_, _22643_, _08341_);
  and (_22673_, _22618_, _06366_);
  and (_22674_, _22673_, _22672_);
  or (_22675_, _22674_, _06528_);
  or (_22676_, _22675_, _22671_);
  or (_22677_, _22655_, _09061_);
  and (_22678_, _22677_, _06926_);
  and (_22679_, _22678_, _22676_);
  and (_22681_, _22621_, _06568_);
  or (_22682_, _22681_, _06278_);
  or (_22683_, _22682_, _22679_);
  or (_22684_, _22607_, _06279_);
  or (_22685_, _22684_, _22619_);
  and (_22686_, _22685_, _01347_);
  and (_22687_, _22686_, _22683_);
  or (_22688_, _22687_, _22605_);
  and (_43212_, _22688_, _42618_);
  and (_22689_, _01351_, \oc8051_golden_model_1.TL0 [2]);
  and (_22691_, _11804_, \oc8051_golden_model_1.TL0 [2]);
  nor (_22692_, _11804_, _07776_);
  or (_22693_, _22692_, _22691_);
  or (_22694_, _22693_, _07215_);
  and (_22695_, _14770_, _07919_);
  or (_22696_, _22695_, _22691_);
  and (_22697_, _22696_, _06341_);
  and (_22698_, _07142_, \oc8051_golden_model_1.TL0 [2]);
  and (_22699_, _07919_, \oc8051_golden_model_1.ACC [2]);
  or (_22700_, _22699_, _22691_);
  and (_22702_, _22700_, _07141_);
  or (_22703_, _22702_, _22698_);
  and (_22704_, _22703_, _07151_);
  or (_22705_, _22704_, _06461_);
  or (_22706_, _22705_, _22697_);
  or (_22707_, _22693_, _07166_);
  and (_22708_, _22707_, _06465_);
  and (_22709_, _22708_, _22706_);
  and (_22710_, _22700_, _06464_);
  or (_22711_, _22710_, _10080_);
  or (_22713_, _22711_, _22709_);
  and (_22714_, _22713_, _22694_);
  or (_22715_, _22714_, _07460_);
  and (_22716_, _09450_, _07919_);
  or (_22717_, _22691_, _07208_);
  or (_22718_, _22717_, _22716_);
  and (_22719_, _22718_, _22715_);
  or (_22720_, _22719_, _10094_);
  and (_22721_, _14859_, _07919_);
  or (_22722_, _22691_, _05982_);
  or (_22724_, _22722_, _22721_);
  and (_22725_, _22724_, _06219_);
  and (_22726_, _22725_, _22720_);
  and (_22727_, _07919_, _08973_);
  or (_22728_, _22727_, _22691_);
  and (_22729_, _22728_, _06218_);
  or (_22730_, _22729_, _06369_);
  or (_22731_, _22730_, _22726_);
  and (_22732_, _14751_, _07919_);
  or (_22733_, _22732_, _22691_);
  or (_22735_, _22733_, _07237_);
  and (_22736_, _22735_, _07240_);
  and (_22737_, _22736_, _22731_);
  and (_22738_, _11259_, _07919_);
  or (_22739_, _22738_, _22691_);
  and (_22740_, _22739_, _06536_);
  or (_22741_, _22740_, _22737_);
  and (_22742_, _22741_, _07242_);
  or (_22743_, _22691_, _08440_);
  and (_22744_, _22728_, _06375_);
  and (_22746_, _22744_, _22743_);
  or (_22747_, _22746_, _22742_);
  and (_22748_, _22747_, _07234_);
  and (_22749_, _22700_, _06545_);
  and (_22750_, _22749_, _22743_);
  or (_22751_, _22750_, _06366_);
  or (_22752_, _22751_, _22748_);
  and (_22753_, _14748_, _07919_);
  or (_22754_, _22691_, _09056_);
  or (_22755_, _22754_, _22753_);
  and (_22757_, _22755_, _09061_);
  and (_22758_, _22757_, _22752_);
  nor (_22759_, _11258_, _11804_);
  or (_22760_, _22759_, _22691_);
  and (_22761_, _22760_, _06528_);
  or (_22762_, _22761_, _22758_);
  and (_22763_, _22762_, _06926_);
  and (_22764_, _22696_, _06568_);
  or (_22765_, _22764_, _06278_);
  or (_22766_, _22765_, _22763_);
  and (_22768_, _14926_, _07919_);
  or (_22769_, _22691_, _06279_);
  or (_22770_, _22769_, _22768_);
  and (_22771_, _22770_, _01347_);
  and (_22772_, _22771_, _22766_);
  or (_22773_, _22772_, _22689_);
  and (_43213_, _22773_, _42618_);
  and (_22774_, _01351_, \oc8051_golden_model_1.TL0 [3]);
  and (_22775_, _11804_, \oc8051_golden_model_1.TL0 [3]);
  and (_22776_, _14953_, _07919_);
  or (_22778_, _22776_, _22775_);
  or (_22779_, _22778_, _07151_);
  and (_22780_, _07919_, \oc8051_golden_model_1.ACC [3]);
  or (_22781_, _22780_, _22775_);
  and (_22782_, _22781_, _07141_);
  and (_22783_, _07142_, \oc8051_golden_model_1.TL0 [3]);
  or (_22784_, _22783_, _06341_);
  or (_22785_, _22784_, _22782_);
  and (_22786_, _22785_, _07166_);
  and (_22787_, _22786_, _22779_);
  nor (_22789_, _11804_, _07594_);
  or (_22790_, _22789_, _22775_);
  and (_22791_, _22790_, _06461_);
  or (_22792_, _22791_, _22787_);
  and (_22793_, _22792_, _06465_);
  and (_22794_, _22781_, _06464_);
  or (_22795_, _22794_, _10080_);
  or (_22796_, _22795_, _22793_);
  or (_22797_, _22790_, _07215_);
  and (_22798_, _22797_, _22796_);
  or (_22800_, _22798_, _07460_);
  and (_22801_, _09449_, _07919_);
  or (_22802_, _22775_, _07208_);
  or (_22803_, _22802_, _22801_);
  and (_22804_, _22803_, _05982_);
  and (_22805_, _22804_, _22800_);
  and (_22806_, _15048_, _07919_);
  or (_22807_, _22806_, _22775_);
  and (_22808_, _22807_, _10094_);
  or (_22809_, _22808_, _06218_);
  or (_22811_, _22809_, _22805_);
  and (_22812_, _07919_, _08930_);
  or (_22813_, _22812_, _22775_);
  or (_22814_, _22813_, _06219_);
  and (_22815_, _22814_, _22811_);
  or (_22816_, _22815_, _06369_);
  and (_22817_, _14943_, _07919_);
  or (_22818_, _22817_, _22775_);
  or (_22819_, _22818_, _07237_);
  and (_22820_, _22819_, _07240_);
  and (_22822_, _22820_, _22816_);
  and (_22823_, _12577_, _07919_);
  or (_22824_, _22823_, _22775_);
  and (_22825_, _22824_, _06536_);
  or (_22826_, _22825_, _22822_);
  and (_22827_, _22826_, _07242_);
  or (_22828_, _22775_, _08292_);
  and (_22829_, _22813_, _06375_);
  and (_22830_, _22829_, _22828_);
  or (_22831_, _22830_, _22827_);
  and (_22832_, _22831_, _07234_);
  and (_22833_, _22781_, _06545_);
  and (_22834_, _22833_, _22828_);
  or (_22835_, _22834_, _06366_);
  or (_22836_, _22835_, _22832_);
  and (_22837_, _14940_, _07919_);
  or (_22838_, _22775_, _09056_);
  or (_22839_, _22838_, _22837_);
  and (_22840_, _22839_, _09061_);
  and (_22841_, _22840_, _22836_);
  nor (_22844_, _11256_, _11804_);
  or (_22845_, _22844_, _22775_);
  and (_22846_, _22845_, _06528_);
  or (_22847_, _22846_, _22841_);
  and (_22848_, _22847_, _06926_);
  and (_22849_, _22778_, _06568_);
  or (_22850_, _22849_, _06278_);
  or (_22851_, _22850_, _22848_);
  and (_22852_, _15128_, _07919_);
  or (_22853_, _22775_, _06279_);
  or (_22855_, _22853_, _22852_);
  and (_22856_, _22855_, _01347_);
  and (_22857_, _22856_, _22851_);
  or (_22858_, _22857_, _22774_);
  and (_43214_, _22858_, _42618_);
  and (_22859_, _01351_, \oc8051_golden_model_1.TL0 [4]);
  and (_22860_, _11804_, \oc8051_golden_model_1.TL0 [4]);
  nor (_22861_, _08541_, _11804_);
  or (_22862_, _22861_, _22860_);
  or (_22863_, _22862_, _07215_);
  and (_22865_, _15162_, _07919_);
  or (_22866_, _22865_, _22860_);
  or (_22867_, _22866_, _07151_);
  and (_22868_, _07919_, \oc8051_golden_model_1.ACC [4]);
  or (_22869_, _22868_, _22860_);
  and (_22870_, _22869_, _07141_);
  and (_22871_, _07142_, \oc8051_golden_model_1.TL0 [4]);
  or (_22872_, _22871_, _06341_);
  or (_22873_, _22872_, _22870_);
  and (_22874_, _22873_, _07166_);
  and (_22876_, _22874_, _22867_);
  and (_22877_, _22862_, _06461_);
  or (_22878_, _22877_, _22876_);
  and (_22879_, _22878_, _06465_);
  and (_22880_, _22869_, _06464_);
  or (_22881_, _22880_, _10080_);
  or (_22882_, _22881_, _22879_);
  and (_22883_, _22882_, _22863_);
  or (_22884_, _22883_, _07460_);
  and (_22885_, _09448_, _07919_);
  or (_22887_, _22860_, _07208_);
  or (_22888_, _22887_, _22885_);
  and (_22889_, _22888_, _22884_);
  or (_22890_, _22889_, _10094_);
  and (_22891_, _15254_, _07919_);
  or (_22892_, _22860_, _05982_);
  or (_22893_, _22892_, _22891_);
  and (_22894_, _22893_, _06219_);
  and (_22895_, _22894_, _22890_);
  and (_22896_, _08959_, _07919_);
  or (_22898_, _22896_, _22860_);
  and (_22899_, _22898_, _06218_);
  or (_22900_, _22899_, _06369_);
  or (_22901_, _22900_, _22895_);
  and (_22902_, _15269_, _07919_);
  or (_22903_, _22902_, _22860_);
  or (_22904_, _22903_, _07237_);
  and (_22905_, _22904_, _07240_);
  and (_22906_, _22905_, _22901_);
  and (_22907_, _11254_, _07919_);
  or (_22909_, _22907_, _22860_);
  and (_22910_, _22909_, _06536_);
  or (_22911_, _22910_, _22906_);
  and (_22912_, _22911_, _07242_);
  or (_22913_, _22860_, _08544_);
  and (_22914_, _22898_, _06375_);
  and (_22915_, _22914_, _22913_);
  or (_22916_, _22915_, _22912_);
  and (_22917_, _22916_, _07234_);
  and (_22918_, _22869_, _06545_);
  and (_22920_, _22918_, _22913_);
  or (_22921_, _22920_, _06366_);
  or (_22922_, _22921_, _22917_);
  and (_22923_, _15266_, _07919_);
  or (_22924_, _22860_, _09056_);
  or (_22925_, _22924_, _22923_);
  and (_22926_, _22925_, _09061_);
  and (_22927_, _22926_, _22922_);
  nor (_22928_, _11253_, _11804_);
  or (_22929_, _22928_, _22860_);
  and (_22931_, _22929_, _06528_);
  or (_22932_, _22931_, _22927_);
  and (_22933_, _22932_, _06926_);
  and (_22934_, _22866_, _06568_);
  or (_22935_, _22934_, _06278_);
  or (_22936_, _22935_, _22933_);
  and (_22937_, _15329_, _07919_);
  or (_22938_, _22860_, _06279_);
  or (_22939_, _22938_, _22937_);
  and (_22940_, _22939_, _01347_);
  and (_22942_, _22940_, _22936_);
  or (_22943_, _22942_, _22859_);
  and (_43215_, _22943_, _42618_);
  and (_22944_, _01351_, \oc8051_golden_model_1.TL0 [5]);
  and (_22945_, _11804_, \oc8051_golden_model_1.TL0 [5]);
  nor (_22946_, _08244_, _11804_);
  or (_22947_, _22946_, _22945_);
  or (_22948_, _22947_, _07215_);
  and (_22949_, _15358_, _07919_);
  or (_22950_, _22949_, _22945_);
  or (_22952_, _22950_, _07151_);
  and (_22953_, _07919_, \oc8051_golden_model_1.ACC [5]);
  or (_22954_, _22953_, _22945_);
  and (_22955_, _22954_, _07141_);
  and (_22956_, _07142_, \oc8051_golden_model_1.TL0 [5]);
  or (_22957_, _22956_, _06341_);
  or (_22958_, _22957_, _22955_);
  and (_22959_, _22958_, _07166_);
  and (_22960_, _22959_, _22952_);
  and (_22961_, _22947_, _06461_);
  or (_22963_, _22961_, _22960_);
  and (_22964_, _22963_, _06465_);
  and (_22965_, _22954_, _06464_);
  or (_22966_, _22965_, _10080_);
  or (_22967_, _22966_, _22964_);
  and (_22968_, _22967_, _22948_);
  or (_22969_, _22968_, _07460_);
  and (_22970_, _09447_, _07919_);
  or (_22971_, _22945_, _07208_);
  or (_22972_, _22971_, _22970_);
  and (_22974_, _22972_, _05982_);
  and (_22975_, _22974_, _22969_);
  and (_22976_, _15459_, _07919_);
  or (_22977_, _22976_, _22945_);
  and (_22978_, _22977_, _10094_);
  or (_22979_, _22978_, _06218_);
  or (_22980_, _22979_, _22975_);
  and (_22981_, _08946_, _07919_);
  or (_22982_, _22981_, _22945_);
  or (_22983_, _22982_, _06219_);
  and (_22985_, _22983_, _22980_);
  or (_22986_, _22985_, _06369_);
  and (_22987_, _15353_, _07919_);
  or (_22988_, _22987_, _22945_);
  or (_22989_, _22988_, _07237_);
  and (_22990_, _22989_, _07240_);
  and (_22991_, _22990_, _22986_);
  and (_22992_, _11250_, _07919_);
  or (_22993_, _22992_, _22945_);
  and (_22994_, _22993_, _06536_);
  or (_22996_, _22994_, _22991_);
  and (_22997_, _22996_, _07242_);
  or (_22998_, _22945_, _08247_);
  and (_22999_, _22982_, _06375_);
  and (_23000_, _22999_, _22998_);
  or (_23001_, _23000_, _22997_);
  and (_23002_, _23001_, _07234_);
  and (_23003_, _22954_, _06545_);
  and (_23004_, _23003_, _22998_);
  or (_23005_, _23004_, _06366_);
  or (_23007_, _23005_, _23002_);
  and (_23008_, _15350_, _07919_);
  or (_23009_, _22945_, _09056_);
  or (_23010_, _23009_, _23008_);
  and (_23011_, _23010_, _09061_);
  and (_23012_, _23011_, _23007_);
  nor (_23013_, _11249_, _11804_);
  or (_23014_, _23013_, _22945_);
  and (_23015_, _23014_, _06528_);
  or (_23016_, _23015_, _23012_);
  and (_23018_, _23016_, _06926_);
  and (_23019_, _22950_, _06568_);
  or (_23020_, _23019_, _06278_);
  or (_23021_, _23020_, _23018_);
  and (_23022_, _15532_, _07919_);
  or (_23023_, _22945_, _06279_);
  or (_23024_, _23023_, _23022_);
  and (_23025_, _23024_, _01347_);
  and (_23026_, _23025_, _23021_);
  or (_23027_, _23026_, _22944_);
  and (_43216_, _23027_, _42618_);
  and (_23029_, _01351_, \oc8051_golden_model_1.TL0 [6]);
  and (_23030_, _11804_, \oc8051_golden_model_1.TL0 [6]);
  nor (_23031_, _08142_, _11804_);
  or (_23032_, _23031_, _23030_);
  or (_23033_, _23032_, _07215_);
  and (_23034_, _15554_, _07919_);
  or (_23035_, _23034_, _23030_);
  or (_23036_, _23035_, _07151_);
  and (_23037_, _07919_, \oc8051_golden_model_1.ACC [6]);
  or (_23039_, _23037_, _23030_);
  and (_23040_, _23039_, _07141_);
  and (_23041_, _07142_, \oc8051_golden_model_1.TL0 [6]);
  or (_23042_, _23041_, _06341_);
  or (_23043_, _23042_, _23040_);
  and (_23044_, _23043_, _07166_);
  and (_23045_, _23044_, _23036_);
  and (_23046_, _23032_, _06461_);
  or (_23047_, _23046_, _23045_);
  and (_23048_, _23047_, _06465_);
  and (_23050_, _23039_, _06464_);
  or (_23051_, _23050_, _10080_);
  or (_23052_, _23051_, _23048_);
  and (_23053_, _23052_, _23033_);
  or (_23054_, _23053_, _07460_);
  and (_23055_, _09446_, _07919_);
  or (_23056_, _23030_, _07208_);
  or (_23057_, _23056_, _23055_);
  and (_23058_, _23057_, _05982_);
  and (_23059_, _23058_, _23054_);
  and (_23061_, _15657_, _07919_);
  or (_23062_, _23061_, _23030_);
  and (_23063_, _23062_, _10094_);
  or (_23064_, _23063_, _06218_);
  or (_23065_, _23064_, _23059_);
  and (_23066_, _15664_, _07919_);
  or (_23067_, _23066_, _23030_);
  or (_23068_, _23067_, _06219_);
  and (_23069_, _23068_, _23065_);
  or (_23070_, _23069_, _06369_);
  and (_23072_, _15549_, _07919_);
  or (_23073_, _23072_, _23030_);
  or (_23074_, _23073_, _07237_);
  and (_23075_, _23074_, _07240_);
  and (_23076_, _23075_, _23070_);
  and (_23077_, _11247_, _07919_);
  or (_23078_, _23077_, _23030_);
  and (_23079_, _23078_, _06536_);
  or (_23080_, _23079_, _23076_);
  and (_23081_, _23080_, _07242_);
  or (_23083_, _23030_, _08145_);
  and (_23084_, _23067_, _06375_);
  and (_23085_, _23084_, _23083_);
  or (_23086_, _23085_, _23081_);
  and (_23087_, _23086_, _07234_);
  and (_23088_, _23039_, _06545_);
  and (_23089_, _23088_, _23083_);
  or (_23090_, _23089_, _06366_);
  or (_23091_, _23090_, _23087_);
  and (_23092_, _15546_, _07919_);
  or (_23093_, _23030_, _09056_);
  or (_23094_, _23093_, _23092_);
  and (_23095_, _23094_, _09061_);
  and (_23096_, _23095_, _23091_);
  nor (_23097_, _11246_, _11804_);
  or (_23098_, _23097_, _23030_);
  and (_23099_, _23098_, _06528_);
  or (_23100_, _23099_, _23096_);
  and (_23101_, _23100_, _06926_);
  and (_23102_, _23035_, _06568_);
  or (_23105_, _23102_, _06278_);
  or (_23106_, _23105_, _23101_);
  and (_23107_, _15734_, _07919_);
  or (_23108_, _23030_, _06279_);
  or (_23109_, _23108_, _23107_);
  and (_23110_, _23109_, _01347_);
  and (_23111_, _23110_, _23106_);
  or (_23112_, _23111_, _23029_);
  and (_43217_, _23112_, _42618_);
  not (_23113_, \oc8051_golden_model_1.TCON [0]);
  nor (_23115_, _01347_, _23113_);
  nand (_23116_, _11263_, _07928_);
  nor (_23117_, _07928_, _23113_);
  nor (_23118_, _23117_, _07234_);
  nand (_23119_, _23118_, _23116_);
  and (_23120_, _07928_, _07133_);
  or (_23121_, _23120_, _23117_);
  or (_23122_, _23121_, _07215_);
  nor (_23123_, _08390_, _11882_);
  or (_23124_, _23123_, _23117_);
  or (_23126_, _23124_, _07151_);
  and (_23127_, _07928_, \oc8051_golden_model_1.ACC [0]);
  or (_23128_, _23127_, _23117_);
  and (_23129_, _23128_, _07141_);
  nor (_23130_, _07141_, _23113_);
  or (_23131_, _23130_, _06341_);
  or (_23132_, _23131_, _23129_);
  and (_23133_, _23132_, _06273_);
  and (_23134_, _23133_, _23126_);
  nor (_23135_, _08616_, _23113_);
  and (_23137_, _14382_, _08616_);
  or (_23138_, _23137_, _23135_);
  and (_23139_, _23138_, _06272_);
  or (_23140_, _23139_, _23134_);
  and (_23141_, _23140_, _07166_);
  and (_23142_, _23121_, _06461_);
  or (_23143_, _23142_, _06464_);
  or (_23144_, _23143_, _23141_);
  or (_23145_, _23128_, _06465_);
  and (_23146_, _23145_, _06269_);
  and (_23148_, _23146_, _23144_);
  and (_23149_, _23117_, _06268_);
  or (_23150_, _23149_, _06261_);
  or (_23151_, _23150_, _23148_);
  or (_23152_, _23124_, _06262_);
  and (_23153_, _23152_, _06258_);
  and (_23154_, _23153_, _23151_);
  and (_23155_, _14413_, _08616_);
  or (_23156_, _23155_, _23135_);
  and (_23157_, _23156_, _06257_);
  or (_23159_, _23157_, _10080_);
  or (_23160_, _23159_, _23154_);
  and (_23161_, _23160_, _23122_);
  or (_23162_, _23161_, _07460_);
  and (_23163_, _09392_, _07928_);
  or (_23164_, _23117_, _07208_);
  or (_23165_, _23164_, _23163_);
  and (_23166_, _23165_, _23162_);
  or (_23167_, _23166_, _10094_);
  and (_23168_, _14467_, _07928_);
  or (_23170_, _23117_, _05982_);
  or (_23171_, _23170_, _23168_);
  and (_23172_, _23171_, _06219_);
  and (_23173_, _23172_, _23167_);
  and (_23174_, _07928_, _08954_);
  or (_23175_, _23174_, _23117_);
  and (_23176_, _23175_, _06218_);
  or (_23177_, _23176_, _06369_);
  or (_23178_, _23177_, _23173_);
  and (_23179_, _14366_, _07928_);
  or (_23181_, _23179_, _23117_);
  or (_23182_, _23181_, _07237_);
  and (_23183_, _23182_, _07240_);
  and (_23184_, _23183_, _23178_);
  nor (_23185_, _12580_, _11882_);
  or (_23186_, _23185_, _23117_);
  and (_23187_, _23116_, _06536_);
  and (_23188_, _23187_, _23186_);
  or (_23189_, _23188_, _23184_);
  and (_23190_, _23189_, _07242_);
  nand (_23192_, _23175_, _06375_);
  nor (_23193_, _23192_, _23123_);
  or (_23194_, _23193_, _06545_);
  or (_23195_, _23194_, _23190_);
  and (_23196_, _23195_, _23119_);
  or (_23197_, _23196_, _06366_);
  and (_23198_, _14363_, _07928_);
  or (_23199_, _23117_, _09056_);
  or (_23200_, _23199_, _23198_);
  and (_23201_, _23200_, _09061_);
  and (_23203_, _23201_, _23197_);
  and (_23204_, _23186_, _06528_);
  or (_23205_, _23204_, _06568_);
  or (_23206_, _23205_, _23203_);
  or (_23207_, _23124_, _06926_);
  and (_23208_, _23207_, _23206_);
  or (_23209_, _23208_, _05927_);
  or (_23210_, _23117_, _05928_);
  and (_23211_, _23210_, _23209_);
  or (_23212_, _23211_, _06278_);
  or (_23214_, _23124_, _06279_);
  and (_23215_, _23214_, _01347_);
  and (_23216_, _23215_, _23212_);
  or (_23217_, _23216_, _23115_);
  and (_43219_, _23217_, _42618_);
  not (_23218_, \oc8051_golden_model_1.TCON [1]);
  nor (_23219_, _01347_, _23218_);
  nor (_23220_, _07928_, _23218_);
  nor (_23221_, _11261_, _11882_);
  or (_23222_, _23221_, _23220_);
  or (_23224_, _23222_, _09061_);
  nor (_23225_, _11882_, _07357_);
  or (_23226_, _23225_, _23220_);
  or (_23227_, _23226_, _07166_);
  or (_23228_, _07928_, \oc8051_golden_model_1.TCON [1]);
  and (_23229_, _14562_, _07928_);
  not (_23230_, _23229_);
  and (_23231_, _23230_, _23228_);
  or (_23232_, _23231_, _07151_);
  and (_23233_, _07928_, \oc8051_golden_model_1.ACC [1]);
  or (_23235_, _23233_, _23220_);
  and (_23236_, _23235_, _07141_);
  nor (_23237_, _07141_, _23218_);
  or (_23238_, _23237_, _06341_);
  or (_23239_, _23238_, _23236_);
  and (_23240_, _23239_, _06273_);
  and (_23241_, _23240_, _23232_);
  nor (_23242_, _08616_, _23218_);
  and (_23243_, _14557_, _08616_);
  or (_23244_, _23243_, _23242_);
  and (_23246_, _23244_, _06272_);
  or (_23247_, _23246_, _06461_);
  or (_23248_, _23247_, _23241_);
  and (_23249_, _23248_, _23227_);
  or (_23250_, _23249_, _06464_);
  or (_23251_, _23235_, _06465_);
  and (_23252_, _23251_, _06269_);
  and (_23253_, _23252_, _23250_);
  and (_23254_, _14560_, _08616_);
  or (_23255_, _23254_, _23242_);
  and (_23257_, _23255_, _06268_);
  or (_23258_, _23257_, _06261_);
  or (_23259_, _23258_, _23253_);
  and (_23260_, _23243_, _14556_);
  or (_23261_, _23242_, _06262_);
  or (_23262_, _23261_, _23260_);
  and (_23263_, _23262_, _06258_);
  and (_23264_, _23263_, _23259_);
  or (_23265_, _23242_, _14597_);
  and (_23266_, _23265_, _06257_);
  and (_23268_, _23266_, _23244_);
  or (_23269_, _23268_, _10080_);
  or (_23270_, _23269_, _23264_);
  or (_23271_, _23226_, _07215_);
  and (_23272_, _23271_, _23270_);
  or (_23273_, _23272_, _07460_);
  and (_23274_, _09451_, _07928_);
  or (_23275_, _23220_, _07208_);
  or (_23276_, _23275_, _23274_);
  and (_23277_, _23276_, _05982_);
  and (_23279_, _23277_, _23273_);
  and (_23280_, _14653_, _07928_);
  or (_23281_, _23280_, _23220_);
  and (_23282_, _23281_, _10094_);
  or (_23283_, _23282_, _23279_);
  and (_23284_, _23283_, _06219_);
  nand (_23285_, _07928_, _07038_);
  and (_23286_, _23228_, _06218_);
  and (_23287_, _23286_, _23285_);
  or (_23288_, _23287_, _23284_);
  and (_23290_, _23288_, _07237_);
  or (_23291_, _14668_, _11882_);
  and (_23292_, _23228_, _06369_);
  and (_23293_, _23292_, _23291_);
  or (_23294_, _23293_, _06536_);
  or (_23295_, _23294_, _23290_);
  nand (_23296_, _11260_, _07928_);
  and (_23297_, _23296_, _23222_);
  or (_23298_, _23297_, _07240_);
  and (_23299_, _23298_, _07242_);
  and (_23301_, _23299_, _23295_);
  or (_23302_, _14666_, _11882_);
  and (_23303_, _23228_, _06375_);
  and (_23304_, _23303_, _23302_);
  or (_23305_, _23304_, _06545_);
  or (_23306_, _23305_, _23301_);
  nor (_23307_, _23220_, _07234_);
  nand (_23308_, _23307_, _23296_);
  and (_23309_, _23308_, _09056_);
  and (_23310_, _23309_, _23306_);
  or (_23312_, _23285_, _08341_);
  and (_23313_, _23228_, _06366_);
  and (_23314_, _23313_, _23312_);
  or (_23315_, _23314_, _06528_);
  or (_23316_, _23315_, _23310_);
  and (_23317_, _23316_, _23224_);
  or (_23318_, _23317_, _06568_);
  or (_23319_, _23231_, _06926_);
  and (_23320_, _23319_, _05928_);
  and (_23321_, _23320_, _23318_);
  and (_23323_, _23255_, _05927_);
  or (_23324_, _23323_, _06278_);
  or (_23325_, _23324_, _23321_);
  or (_23326_, _23220_, _06279_);
  or (_23327_, _23326_, _23229_);
  and (_23328_, _23327_, _01347_);
  and (_23329_, _23328_, _23325_);
  or (_23330_, _23329_, _23219_);
  and (_43220_, _23330_, _42618_);
  and (_23331_, _01351_, \oc8051_golden_model_1.TCON [2]);
  and (_23333_, _11882_, \oc8051_golden_model_1.TCON [2]);
  nor (_23334_, _11882_, _07776_);
  or (_23335_, _23334_, _23333_);
  or (_23336_, _23335_, _07215_);
  or (_23337_, _23335_, _07166_);
  and (_23338_, _14770_, _07928_);
  or (_23339_, _23338_, _23333_);
  or (_23340_, _23339_, _07151_);
  and (_23341_, _07928_, \oc8051_golden_model_1.ACC [2]);
  or (_23342_, _23341_, _23333_);
  and (_23344_, _23342_, _07141_);
  and (_23345_, _07142_, \oc8051_golden_model_1.TCON [2]);
  or (_23346_, _23345_, _06341_);
  or (_23347_, _23346_, _23344_);
  and (_23348_, _23347_, _06273_);
  and (_23349_, _23348_, _23340_);
  and (_23350_, _11890_, \oc8051_golden_model_1.TCON [2]);
  and (_23351_, _14774_, _08616_);
  or (_23352_, _23351_, _23350_);
  and (_23353_, _23352_, _06272_);
  or (_23355_, _23353_, _06461_);
  or (_23356_, _23355_, _23349_);
  and (_23357_, _23356_, _23337_);
  or (_23358_, _23357_, _06464_);
  or (_23359_, _23342_, _06465_);
  and (_23360_, _23359_, _06269_);
  and (_23361_, _23360_, _23358_);
  and (_23362_, _14756_, _08616_);
  or (_23363_, _23362_, _23350_);
  and (_23364_, _23363_, _06268_);
  or (_23366_, _23364_, _06261_);
  or (_23367_, _23366_, _23361_);
  and (_23368_, _23351_, _14789_);
  or (_23369_, _23350_, _06262_);
  or (_23370_, _23369_, _23368_);
  and (_23371_, _23370_, _06258_);
  and (_23372_, _23371_, _23367_);
  and (_23373_, _14804_, _08616_);
  or (_23374_, _23373_, _23350_);
  and (_23375_, _23374_, _06257_);
  or (_23376_, _23375_, _10080_);
  or (_23377_, _23376_, _23372_);
  and (_23378_, _23377_, _23336_);
  or (_23379_, _23378_, _07460_);
  and (_23380_, _09450_, _07928_);
  or (_23381_, _23333_, _07208_);
  or (_23382_, _23381_, _23380_);
  and (_23383_, _23382_, _05982_);
  and (_23384_, _23383_, _23379_);
  and (_23385_, _14859_, _07928_);
  or (_23388_, _23385_, _23333_);
  and (_23389_, _23388_, _10094_);
  or (_23390_, _23389_, _06218_);
  or (_23391_, _23390_, _23384_);
  and (_23392_, _07928_, _08973_);
  or (_23393_, _23392_, _23333_);
  or (_23394_, _23393_, _06219_);
  and (_23395_, _23394_, _23391_);
  or (_23396_, _23395_, _06369_);
  and (_23397_, _14751_, _07928_);
  or (_23399_, _23397_, _23333_);
  or (_23400_, _23399_, _07237_);
  and (_23401_, _23400_, _07240_);
  and (_23402_, _23401_, _23396_);
  and (_23403_, _11259_, _07928_);
  or (_23404_, _23403_, _23333_);
  and (_23405_, _23404_, _06536_);
  or (_23406_, _23405_, _23402_);
  and (_23407_, _23406_, _07242_);
  or (_23408_, _23333_, _08440_);
  and (_23410_, _23393_, _06375_);
  and (_23411_, _23410_, _23408_);
  or (_23412_, _23411_, _23407_);
  and (_23413_, _23412_, _07234_);
  and (_23414_, _23342_, _06545_);
  and (_23415_, _23414_, _23408_);
  or (_23416_, _23415_, _06366_);
  or (_23417_, _23416_, _23413_);
  and (_23418_, _14748_, _07928_);
  or (_23419_, _23333_, _09056_);
  or (_23421_, _23419_, _23418_);
  and (_23422_, _23421_, _09061_);
  and (_23423_, _23422_, _23417_);
  nor (_23424_, _11258_, _11882_);
  or (_23425_, _23424_, _23333_);
  and (_23426_, _23425_, _06528_);
  or (_23427_, _23426_, _06568_);
  or (_23428_, _23427_, _23423_);
  or (_23429_, _23339_, _06926_);
  and (_23430_, _23429_, _05928_);
  and (_23432_, _23430_, _23428_);
  and (_23433_, _23363_, _05927_);
  or (_23434_, _23433_, _06278_);
  or (_23435_, _23434_, _23432_);
  and (_23436_, _14926_, _07928_);
  or (_23437_, _23333_, _06279_);
  or (_23438_, _23437_, _23436_);
  and (_23439_, _23438_, _01347_);
  and (_23440_, _23439_, _23435_);
  or (_23441_, _23440_, _23331_);
  and (_43221_, _23441_, _42618_);
  and (_23443_, _01351_, \oc8051_golden_model_1.TCON [3]);
  and (_23444_, _11882_, \oc8051_golden_model_1.TCON [3]);
  nor (_23445_, _11882_, _07594_);
  or (_23446_, _23445_, _23444_);
  or (_23447_, _23446_, _07215_);
  and (_23448_, _14953_, _07928_);
  or (_23449_, _23448_, _23444_);
  or (_23450_, _23449_, _07151_);
  and (_23451_, _07928_, \oc8051_golden_model_1.ACC [3]);
  or (_23453_, _23451_, _23444_);
  and (_23454_, _23453_, _07141_);
  and (_23455_, _07142_, \oc8051_golden_model_1.TCON [3]);
  or (_23456_, _23455_, _06341_);
  or (_23457_, _23456_, _23454_);
  and (_23458_, _23457_, _06273_);
  and (_23459_, _23458_, _23450_);
  and (_23460_, _11890_, \oc8051_golden_model_1.TCON [3]);
  and (_23461_, _14950_, _08616_);
  or (_23462_, _23461_, _23460_);
  and (_23464_, _23462_, _06272_);
  or (_23465_, _23464_, _06461_);
  or (_23466_, _23465_, _23459_);
  or (_23467_, _23446_, _07166_);
  and (_23468_, _23467_, _23466_);
  or (_23469_, _23468_, _06464_);
  or (_23470_, _23453_, _06465_);
  and (_23471_, _23470_, _06269_);
  and (_23472_, _23471_, _23469_);
  and (_23473_, _14948_, _08616_);
  or (_23475_, _23473_, _23460_);
  and (_23476_, _23475_, _06268_);
  or (_23477_, _23476_, _06261_);
  or (_23478_, _23477_, _23472_);
  or (_23479_, _23460_, _14979_);
  and (_23480_, _23479_, _23462_);
  or (_23481_, _23480_, _06262_);
  and (_23482_, _23481_, _06258_);
  and (_23483_, _23482_, _23478_);
  or (_23484_, _23460_, _14992_);
  and (_23486_, _23484_, _06257_);
  and (_23487_, _23486_, _23462_);
  or (_23488_, _23487_, _10080_);
  or (_23489_, _23488_, _23483_);
  and (_23490_, _23489_, _23447_);
  or (_23491_, _23490_, _07460_);
  and (_23492_, _09449_, _07928_);
  or (_23493_, _23444_, _07208_);
  or (_23494_, _23493_, _23492_);
  and (_23495_, _23494_, _05982_);
  and (_23497_, _23495_, _23491_);
  and (_23498_, _15048_, _07928_);
  or (_23499_, _23498_, _23444_);
  and (_23500_, _23499_, _10094_);
  or (_23501_, _23500_, _06218_);
  or (_23502_, _23501_, _23497_);
  and (_23503_, _07928_, _08930_);
  or (_23504_, _23503_, _23444_);
  or (_23505_, _23504_, _06219_);
  and (_23506_, _23505_, _23502_);
  or (_23508_, _23506_, _06369_);
  and (_23509_, _14943_, _07928_);
  or (_23510_, _23509_, _23444_);
  or (_23511_, _23510_, _07237_);
  and (_23512_, _23511_, _07240_);
  and (_23513_, _23512_, _23508_);
  and (_23514_, _12577_, _07928_);
  or (_23515_, _23514_, _23444_);
  and (_23516_, _23515_, _06536_);
  or (_23517_, _23516_, _23513_);
  and (_23519_, _23517_, _07242_);
  or (_23520_, _23444_, _08292_);
  and (_23521_, _23504_, _06375_);
  and (_23522_, _23521_, _23520_);
  or (_23523_, _23522_, _23519_);
  and (_23524_, _23523_, _07234_);
  and (_23525_, _23453_, _06545_);
  and (_23526_, _23525_, _23520_);
  or (_23527_, _23526_, _06366_);
  or (_23528_, _23527_, _23524_);
  and (_23530_, _14940_, _07928_);
  or (_23531_, _23444_, _09056_);
  or (_23532_, _23531_, _23530_);
  and (_23533_, _23532_, _09061_);
  and (_23534_, _23533_, _23528_);
  nor (_23535_, _11256_, _11882_);
  or (_23536_, _23535_, _23444_);
  and (_23537_, _23536_, _06528_);
  or (_23538_, _23537_, _06568_);
  or (_23539_, _23538_, _23534_);
  or (_23541_, _23449_, _06926_);
  and (_23542_, _23541_, _05928_);
  and (_23543_, _23542_, _23539_);
  and (_23544_, _23475_, _05927_);
  or (_23545_, _23544_, _06278_);
  or (_23546_, _23545_, _23543_);
  and (_23547_, _15128_, _07928_);
  or (_23548_, _23444_, _06279_);
  or (_23549_, _23548_, _23547_);
  and (_23550_, _23549_, _01347_);
  and (_23552_, _23550_, _23546_);
  or (_23553_, _23552_, _23443_);
  and (_43223_, _23553_, _42618_);
  and (_23554_, _01351_, \oc8051_golden_model_1.TCON [4]);
  and (_23555_, _11882_, \oc8051_golden_model_1.TCON [4]);
  nor (_23556_, _08541_, _11882_);
  or (_23557_, _23556_, _23555_);
  or (_23558_, _23557_, _07215_);
  and (_23559_, _11890_, \oc8051_golden_model_1.TCON [4]);
  and (_23560_, _15176_, _08616_);
  or (_23562_, _23560_, _23559_);
  and (_23563_, _23562_, _06268_);
  and (_23564_, _15162_, _07928_);
  or (_23565_, _23564_, _23555_);
  or (_23566_, _23565_, _07151_);
  and (_23567_, _07928_, \oc8051_golden_model_1.ACC [4]);
  or (_23568_, _23567_, _23555_);
  and (_23569_, _23568_, _07141_);
  and (_23570_, _07142_, \oc8051_golden_model_1.TCON [4]);
  or (_23571_, _23570_, _06341_);
  or (_23573_, _23571_, _23569_);
  and (_23574_, _23573_, _06273_);
  and (_23575_, _23574_, _23566_);
  and (_23576_, _15166_, _08616_);
  or (_23577_, _23576_, _23559_);
  and (_23578_, _23577_, _06272_);
  or (_23579_, _23578_, _06461_);
  or (_23580_, _23579_, _23575_);
  or (_23581_, _23557_, _07166_);
  and (_23582_, _23581_, _23580_);
  or (_23584_, _23582_, _06464_);
  or (_23585_, _23568_, _06465_);
  and (_23586_, _23585_, _06269_);
  and (_23587_, _23586_, _23584_);
  or (_23588_, _23587_, _23563_);
  and (_23589_, _23588_, _06262_);
  or (_23590_, _23559_, _15183_);
  and (_23591_, _23590_, _06261_);
  and (_23592_, _23591_, _23577_);
  or (_23593_, _23592_, _23589_);
  and (_23595_, _23593_, _06258_);
  and (_23596_, _15200_, _08616_);
  or (_23597_, _23596_, _23559_);
  and (_23598_, _23597_, _06257_);
  or (_23599_, _23598_, _10080_);
  or (_23600_, _23599_, _23595_);
  and (_23601_, _23600_, _23558_);
  or (_23602_, _23601_, _07460_);
  and (_23603_, _09448_, _07928_);
  or (_23604_, _23555_, _07208_);
  or (_23605_, _23604_, _23603_);
  and (_23606_, _23605_, _05982_);
  and (_23607_, _23606_, _23602_);
  and (_23608_, _15254_, _07928_);
  or (_23609_, _23608_, _23555_);
  and (_23610_, _23609_, _10094_);
  or (_23611_, _23610_, _06218_);
  or (_23612_, _23611_, _23607_);
  and (_23613_, _08959_, _07928_);
  or (_23614_, _23613_, _23555_);
  or (_23616_, _23614_, _06219_);
  and (_23617_, _23616_, _23612_);
  or (_23618_, _23617_, _06369_);
  and (_23619_, _15269_, _07928_);
  or (_23620_, _23619_, _23555_);
  or (_23621_, _23620_, _07237_);
  and (_23622_, _23621_, _07240_);
  and (_23623_, _23622_, _23618_);
  and (_23624_, _11254_, _07928_);
  or (_23625_, _23624_, _23555_);
  and (_23627_, _23625_, _06536_);
  or (_23628_, _23627_, _23623_);
  and (_23629_, _23628_, _07242_);
  or (_23630_, _23555_, _08544_);
  and (_23631_, _23614_, _06375_);
  and (_23632_, _23631_, _23630_);
  or (_23633_, _23632_, _23629_);
  and (_23634_, _23633_, _07234_);
  and (_23635_, _23568_, _06545_);
  and (_23636_, _23635_, _23630_);
  or (_23638_, _23636_, _06366_);
  or (_23639_, _23638_, _23634_);
  and (_23640_, _15266_, _07928_);
  or (_23641_, _23555_, _09056_);
  or (_23642_, _23641_, _23640_);
  and (_23643_, _23642_, _09061_);
  and (_23644_, _23643_, _23639_);
  nor (_23645_, _11253_, _11882_);
  or (_23646_, _23645_, _23555_);
  and (_23647_, _23646_, _06528_);
  or (_23648_, _23647_, _06568_);
  or (_23649_, _23648_, _23644_);
  or (_23650_, _23565_, _06926_);
  and (_23651_, _23650_, _05928_);
  and (_23652_, _23651_, _23649_);
  and (_23653_, _23562_, _05927_);
  or (_23654_, _23653_, _06278_);
  or (_23655_, _23654_, _23652_);
  and (_23656_, _15329_, _07928_);
  or (_23657_, _23555_, _06279_);
  or (_23659_, _23657_, _23656_);
  and (_23660_, _23659_, _01347_);
  and (_23661_, _23660_, _23655_);
  or (_23662_, _23661_, _23554_);
  and (_43224_, _23662_, _42618_);
  and (_23663_, _01351_, \oc8051_golden_model_1.TCON [5]);
  and (_23664_, _11882_, \oc8051_golden_model_1.TCON [5]);
  and (_23665_, _15358_, _07928_);
  or (_23666_, _23665_, _23664_);
  or (_23667_, _23666_, _07151_);
  and (_23668_, _07928_, \oc8051_golden_model_1.ACC [5]);
  or (_23669_, _23668_, _23664_);
  and (_23670_, _23669_, _07141_);
  and (_23671_, _07142_, \oc8051_golden_model_1.TCON [5]);
  or (_23672_, _23671_, _06341_);
  or (_23673_, _23672_, _23670_);
  and (_23674_, _23673_, _06273_);
  and (_23675_, _23674_, _23667_);
  and (_23676_, _11890_, \oc8051_golden_model_1.TCON [5]);
  and (_23677_, _15372_, _08616_);
  or (_23679_, _23677_, _23676_);
  and (_23680_, _23679_, _06272_);
  or (_23681_, _23680_, _06461_);
  or (_23682_, _23681_, _23675_);
  nor (_23683_, _08244_, _11882_);
  or (_23684_, _23683_, _23664_);
  or (_23685_, _23684_, _07166_);
  and (_23686_, _23685_, _23682_);
  or (_23687_, _23686_, _06464_);
  or (_23688_, _23669_, _06465_);
  and (_23690_, _23688_, _06269_);
  and (_23691_, _23690_, _23687_);
  and (_23692_, _15355_, _08616_);
  or (_23693_, _23692_, _23676_);
  and (_23694_, _23693_, _06268_);
  or (_23695_, _23694_, _06261_);
  or (_23696_, _23695_, _23691_);
  or (_23697_, _23676_, _15387_);
  and (_23698_, _23697_, _23679_);
  or (_23699_, _23698_, _06262_);
  and (_23700_, _23699_, _06258_);
  and (_23701_, _23700_, _23696_);
  or (_23702_, _23676_, _15403_);
  and (_23703_, _23702_, _06257_);
  and (_23704_, _23703_, _23679_);
  or (_23705_, _23704_, _10080_);
  or (_23706_, _23705_, _23701_);
  or (_23707_, _23684_, _07215_);
  and (_23708_, _23707_, _23706_);
  or (_23709_, _23708_, _07460_);
  and (_23711_, _09447_, _07928_);
  or (_23712_, _23664_, _07208_);
  or (_23713_, _23712_, _23711_);
  and (_23714_, _23713_, _05982_);
  and (_23715_, _23714_, _23709_);
  and (_23716_, _15459_, _07928_);
  or (_23717_, _23716_, _23664_);
  and (_23718_, _23717_, _10094_);
  or (_23719_, _23718_, _06218_);
  or (_23720_, _23719_, _23715_);
  and (_23722_, _08946_, _07928_);
  or (_23723_, _23722_, _23664_);
  or (_23724_, _23723_, _06219_);
  and (_23725_, _23724_, _23720_);
  or (_23726_, _23725_, _06369_);
  and (_23727_, _15353_, _07928_);
  or (_23728_, _23727_, _23664_);
  or (_23729_, _23728_, _07237_);
  and (_23730_, _23729_, _07240_);
  and (_23731_, _23730_, _23726_);
  and (_23732_, _11250_, _07928_);
  or (_23733_, _23732_, _23664_);
  and (_23734_, _23733_, _06536_);
  or (_23735_, _23734_, _23731_);
  and (_23736_, _23735_, _07242_);
  or (_23737_, _23664_, _08247_);
  and (_23738_, _23723_, _06375_);
  and (_23739_, _23738_, _23737_);
  or (_23740_, _23739_, _23736_);
  and (_23741_, _23740_, _07234_);
  and (_23743_, _23669_, _06545_);
  and (_23744_, _23743_, _23737_);
  or (_23745_, _23744_, _06366_);
  or (_23746_, _23745_, _23741_);
  and (_23747_, _15350_, _07928_);
  or (_23748_, _23664_, _09056_);
  or (_23749_, _23748_, _23747_);
  and (_23750_, _23749_, _09061_);
  and (_23751_, _23750_, _23746_);
  nor (_23752_, _11249_, _11882_);
  or (_23754_, _23752_, _23664_);
  and (_23755_, _23754_, _06528_);
  or (_23756_, _23755_, _06568_);
  or (_23757_, _23756_, _23751_);
  or (_23758_, _23666_, _06926_);
  and (_23759_, _23758_, _05928_);
  and (_23760_, _23759_, _23757_);
  and (_23761_, _23693_, _05927_);
  or (_23762_, _23761_, _06278_);
  or (_23763_, _23762_, _23760_);
  and (_23764_, _15532_, _07928_);
  or (_23765_, _23664_, _06279_);
  or (_23766_, _23765_, _23764_);
  and (_23767_, _23766_, _01347_);
  and (_23768_, _23767_, _23763_);
  or (_23769_, _23768_, _23663_);
  and (_43225_, _23769_, _42618_);
  and (_23770_, _01351_, \oc8051_golden_model_1.TCON [6]);
  and (_23771_, _11882_, \oc8051_golden_model_1.TCON [6]);
  and (_23772_, _15554_, _07928_);
  or (_23774_, _23772_, _23771_);
  or (_23775_, _23774_, _07151_);
  and (_23776_, _07928_, \oc8051_golden_model_1.ACC [6]);
  or (_23777_, _23776_, _23771_);
  and (_23778_, _23777_, _07141_);
  and (_23779_, _07142_, \oc8051_golden_model_1.TCON [6]);
  or (_23780_, _23779_, _06341_);
  or (_23781_, _23780_, _23778_);
  and (_23782_, _23781_, _06273_);
  and (_23783_, _23782_, _23775_);
  and (_23785_, _11890_, \oc8051_golden_model_1.TCON [6]);
  and (_23786_, _15570_, _08616_);
  or (_23787_, _23786_, _23785_);
  and (_23788_, _23787_, _06272_);
  or (_23789_, _23788_, _06461_);
  or (_23790_, _23789_, _23783_);
  nor (_23791_, _08142_, _11882_);
  or (_23792_, _23791_, _23771_);
  or (_23793_, _23792_, _07166_);
  and (_23794_, _23793_, _23790_);
  or (_23795_, _23794_, _06464_);
  or (_23796_, _23777_, _06465_);
  and (_23797_, _23796_, _06269_);
  and (_23798_, _23797_, _23795_);
  and (_23799_, _15551_, _08616_);
  or (_23800_, _23799_, _23785_);
  and (_23801_, _23800_, _06268_);
  or (_23802_, _23801_, _06261_);
  or (_23803_, _23802_, _23798_);
  or (_23804_, _23785_, _15585_);
  and (_23805_, _23804_, _23787_);
  or (_23806_, _23805_, _06262_);
  and (_23807_, _23806_, _06258_);
  and (_23808_, _23807_, _23803_);
  and (_23809_, _15602_, _08616_);
  or (_23810_, _23809_, _23785_);
  and (_23811_, _23810_, _06257_);
  or (_23812_, _23811_, _10080_);
  or (_23813_, _23812_, _23808_);
  or (_23814_, _23792_, _07215_);
  and (_23817_, _23814_, _23813_);
  or (_23818_, _23817_, _07460_);
  and (_23819_, _09446_, _07928_);
  or (_23820_, _23771_, _07208_);
  or (_23821_, _23820_, _23819_);
  and (_23822_, _23821_, _05982_);
  and (_23823_, _23822_, _23818_);
  and (_23824_, _15657_, _07928_);
  or (_23825_, _23824_, _23771_);
  and (_23826_, _23825_, _10094_);
  or (_23827_, _23826_, _06218_);
  or (_23828_, _23827_, _23823_);
  and (_23829_, _15664_, _07928_);
  or (_23830_, _23829_, _23771_);
  or (_23831_, _23830_, _06219_);
  and (_23832_, _23831_, _23828_);
  or (_23833_, _23832_, _06369_);
  and (_23834_, _15549_, _07928_);
  or (_23835_, _23834_, _23771_);
  or (_23836_, _23835_, _07237_);
  and (_23838_, _23836_, _07240_);
  and (_23839_, _23838_, _23833_);
  and (_23840_, _11247_, _07928_);
  or (_23841_, _23840_, _23771_);
  and (_23842_, _23841_, _06536_);
  or (_23843_, _23842_, _23839_);
  and (_23844_, _23843_, _07242_);
  or (_23845_, _23771_, _08145_);
  and (_23846_, _23830_, _06375_);
  and (_23847_, _23846_, _23845_);
  or (_23849_, _23847_, _23844_);
  and (_23850_, _23849_, _07234_);
  and (_23851_, _23777_, _06545_);
  and (_23852_, _23851_, _23845_);
  or (_23853_, _23852_, _06366_);
  or (_23854_, _23853_, _23850_);
  and (_23855_, _15546_, _07928_);
  or (_23856_, _23771_, _09056_);
  or (_23857_, _23856_, _23855_);
  and (_23858_, _23857_, _09061_);
  and (_23859_, _23858_, _23854_);
  nor (_23860_, _11246_, _11882_);
  or (_23861_, _23860_, _23771_);
  and (_23862_, _23861_, _06528_);
  or (_23863_, _23862_, _06568_);
  or (_23864_, _23863_, _23859_);
  or (_23865_, _23774_, _06926_);
  and (_23866_, _23865_, _05928_);
  and (_23867_, _23866_, _23864_);
  and (_23868_, _23800_, _05927_);
  or (_23870_, _23868_, _06278_);
  or (_23871_, _23870_, _23867_);
  and (_23872_, _15734_, _07928_);
  or (_23873_, _23771_, _06279_);
  or (_23874_, _23873_, _23872_);
  and (_23875_, _23874_, _01347_);
  and (_23876_, _23875_, _23871_);
  or (_23877_, _23876_, _23770_);
  and (_43226_, _23877_, _42618_);
  and (_23878_, _01351_, \oc8051_golden_model_1.TH1 [0]);
  and (_23880_, _07910_, \oc8051_golden_model_1.ACC [0]);
  and (_23881_, _23880_, _08390_);
  and (_23882_, _11985_, \oc8051_golden_model_1.TH1 [0]);
  or (_23883_, _23882_, _07234_);
  or (_23884_, _23883_, _23881_);
  and (_23885_, _07910_, _07133_);
  or (_23886_, _23885_, _23882_);
  or (_23887_, _23886_, _07215_);
  nor (_23888_, _08390_, _11985_);
  or (_23889_, _23888_, _23882_);
  or (_23890_, _23889_, _07151_);
  or (_23891_, _23882_, _23880_);
  and (_23892_, _23891_, _07141_);
  and (_23893_, _07142_, \oc8051_golden_model_1.TH1 [0]);
  or (_23894_, _23893_, _06341_);
  or (_23895_, _23894_, _23892_);
  and (_23896_, _23895_, _07166_);
  and (_23897_, _23896_, _23890_);
  and (_23898_, _23886_, _06461_);
  or (_23899_, _23898_, _23897_);
  and (_23901_, _23899_, _06465_);
  and (_23902_, _23891_, _06464_);
  or (_23903_, _23902_, _10080_);
  or (_23904_, _23903_, _23901_);
  and (_23905_, _23904_, _23887_);
  or (_23906_, _23905_, _07460_);
  and (_23907_, _09392_, _07910_);
  or (_23908_, _23882_, _07208_);
  or (_23909_, _23908_, _23907_);
  and (_23910_, _23909_, _23906_);
  or (_23912_, _23910_, _10094_);
  and (_23913_, _14467_, _07910_);
  or (_23914_, _23882_, _05982_);
  or (_23915_, _23914_, _23913_);
  and (_23916_, _23915_, _06219_);
  and (_23917_, _23916_, _23912_);
  and (_23918_, _07910_, _08954_);
  or (_23919_, _23918_, _23882_);
  and (_23920_, _23919_, _06218_);
  or (_23921_, _23920_, _06369_);
  or (_23922_, _23921_, _23917_);
  and (_23923_, _14366_, _07910_);
  or (_23924_, _23923_, _23882_);
  or (_23925_, _23924_, _07237_);
  and (_23926_, _23925_, _07240_);
  and (_23927_, _23926_, _23922_);
  nor (_23928_, _12580_, _11985_);
  or (_23929_, _23928_, _23882_);
  nor (_23930_, _23881_, _07240_);
  and (_23931_, _23930_, _23929_);
  or (_23933_, _23931_, _23927_);
  and (_23934_, _23933_, _07242_);
  nand (_23935_, _23919_, _06375_);
  nor (_23936_, _23935_, _23888_);
  or (_23937_, _23936_, _06545_);
  or (_23938_, _23937_, _23934_);
  and (_23939_, _23938_, _23884_);
  or (_23940_, _23939_, _06366_);
  and (_23941_, _14363_, _07910_);
  or (_23942_, _23882_, _09056_);
  or (_23944_, _23942_, _23941_);
  and (_23945_, _23944_, _09061_);
  and (_23946_, _23945_, _23940_);
  and (_23947_, _23929_, _06528_);
  or (_23948_, _23947_, _19502_);
  or (_23949_, _23948_, _23946_);
  or (_23950_, _23889_, _06661_);
  and (_23951_, _23950_, _01347_);
  and (_23952_, _23951_, _23949_);
  or (_23953_, _23952_, _23878_);
  and (_43228_, _23953_, _42618_);
  and (_23954_, _01351_, \oc8051_golden_model_1.TH1 [1]);
  nand (_23955_, _07910_, _07038_);
  or (_23956_, _07910_, \oc8051_golden_model_1.TH1 [1]);
  and (_23957_, _23956_, _06218_);
  and (_23958_, _23957_, _23955_);
  and (_23959_, _11985_, \oc8051_golden_model_1.TH1 [1]);
  nor (_23960_, _11985_, _07357_);
  or (_23961_, _23960_, _23959_);
  or (_23962_, _23961_, _07215_);
  and (_23964_, _14562_, _07910_);
  not (_23965_, _23964_);
  and (_23966_, _23965_, _23956_);
  or (_23967_, _23966_, _07151_);
  and (_23968_, _07910_, \oc8051_golden_model_1.ACC [1]);
  or (_23969_, _23968_, _23959_);
  and (_23970_, _23969_, _07141_);
  and (_23971_, _07142_, \oc8051_golden_model_1.TH1 [1]);
  or (_23972_, _23971_, _06341_);
  or (_23973_, _23972_, _23970_);
  and (_23975_, _23973_, _07166_);
  and (_23976_, _23975_, _23967_);
  and (_23977_, _23961_, _06461_);
  or (_23978_, _23977_, _23976_);
  and (_23979_, _23978_, _06465_);
  and (_23980_, _23969_, _06464_);
  or (_23981_, _23980_, _10080_);
  or (_23982_, _23981_, _23979_);
  and (_23983_, _23982_, _23962_);
  or (_23984_, _23983_, _07460_);
  and (_23985_, _09451_, _07910_);
  or (_23986_, _23959_, _07208_);
  or (_23987_, _23986_, _23985_);
  and (_23988_, _23987_, _05982_);
  and (_23989_, _23988_, _23984_);
  or (_23990_, _14653_, _11985_);
  and (_23991_, _23956_, _10094_);
  and (_23992_, _23991_, _23990_);
  or (_23993_, _23992_, _23989_);
  and (_23994_, _23993_, _06219_);
  or (_23996_, _23994_, _23958_);
  and (_23997_, _23996_, _07237_);
  or (_23998_, _14668_, _11985_);
  and (_23999_, _23956_, _06369_);
  and (_24000_, _23999_, _23998_);
  or (_24001_, _24000_, _06536_);
  or (_24002_, _24001_, _23997_);
  and (_24003_, _11262_, _07910_);
  or (_24004_, _24003_, _23959_);
  or (_24005_, _24004_, _07240_);
  and (_24007_, _24005_, _07242_);
  and (_24008_, _24007_, _24002_);
  or (_24009_, _14666_, _11985_);
  and (_24010_, _23956_, _06375_);
  and (_24011_, _24010_, _24009_);
  or (_24012_, _24011_, _06545_);
  or (_24013_, _24012_, _24008_);
  and (_24014_, _23968_, _08341_);
  or (_24015_, _23959_, _07234_);
  or (_24016_, _24015_, _24014_);
  and (_24018_, _24016_, _09056_);
  and (_24019_, _24018_, _24013_);
  or (_24020_, _23955_, _08341_);
  and (_24021_, _23956_, _06366_);
  and (_24022_, _24021_, _24020_);
  or (_24023_, _24022_, _06528_);
  or (_24024_, _24023_, _24019_);
  nor (_24025_, _11261_, _11985_);
  or (_24026_, _24025_, _23959_);
  or (_24027_, _24026_, _09061_);
  and (_24028_, _24027_, _06926_);
  and (_24029_, _24028_, _24024_);
  and (_24030_, _23966_, _06568_);
  or (_24031_, _24030_, _06278_);
  or (_24032_, _24031_, _24029_);
  or (_24033_, _23959_, _06279_);
  or (_24034_, _24033_, _23964_);
  and (_24035_, _24034_, _01347_);
  and (_24036_, _24035_, _24032_);
  or (_24037_, _24036_, _23954_);
  and (_43229_, _24037_, _42618_);
  and (_24039_, _01351_, \oc8051_golden_model_1.TH1 [2]);
  and (_24040_, _11985_, \oc8051_golden_model_1.TH1 [2]);
  and (_24041_, _09450_, _07910_);
  or (_24042_, _24041_, _24040_);
  and (_24043_, _24042_, _07460_);
  and (_24044_, _14770_, _07910_);
  or (_24045_, _24044_, _24040_);
  or (_24046_, _24045_, _07151_);
  and (_24047_, _07910_, \oc8051_golden_model_1.ACC [2]);
  or (_24049_, _24047_, _24040_);
  and (_24050_, _24049_, _07141_);
  and (_24051_, _07142_, \oc8051_golden_model_1.TH1 [2]);
  or (_24052_, _24051_, _06341_);
  or (_24053_, _24052_, _24050_);
  and (_24054_, _24053_, _07166_);
  and (_24055_, _24054_, _24046_);
  nor (_24056_, _11985_, _07776_);
  or (_24057_, _24056_, _24040_);
  and (_24058_, _24057_, _06461_);
  or (_24059_, _24058_, _24055_);
  and (_24060_, _24059_, _06465_);
  and (_24061_, _24049_, _06464_);
  or (_24062_, _24061_, _10080_);
  or (_24063_, _24062_, _24060_);
  or (_24064_, _24057_, _07215_);
  and (_24065_, _24064_, _07208_);
  and (_24066_, _24065_, _24063_);
  or (_24067_, _24066_, _10094_);
  or (_24068_, _24067_, _24043_);
  and (_24070_, _14859_, _07910_);
  or (_24071_, _24040_, _05982_);
  or (_24072_, _24071_, _24070_);
  and (_24073_, _24072_, _06219_);
  and (_24074_, _24073_, _24068_);
  and (_24075_, _07910_, _08973_);
  or (_24076_, _24075_, _24040_);
  and (_24077_, _24076_, _06218_);
  or (_24078_, _24077_, _06369_);
  or (_24079_, _24078_, _24074_);
  and (_24081_, _14751_, _07910_);
  or (_24082_, _24081_, _24040_);
  or (_24083_, _24082_, _07237_);
  and (_24084_, _24083_, _07240_);
  and (_24085_, _24084_, _24079_);
  and (_24086_, _11259_, _07910_);
  or (_24087_, _24086_, _24040_);
  and (_24088_, _24087_, _06536_);
  or (_24089_, _24088_, _24085_);
  and (_24090_, _24089_, _07242_);
  or (_24092_, _24040_, _08440_);
  and (_24093_, _24076_, _06375_);
  and (_24094_, _24093_, _24092_);
  or (_24095_, _24094_, _24090_);
  and (_24096_, _24095_, _07234_);
  and (_24097_, _24049_, _06545_);
  and (_24098_, _24097_, _24092_);
  or (_24099_, _24098_, _06366_);
  or (_24100_, _24099_, _24096_);
  and (_24101_, _14748_, _07910_);
  or (_24102_, _24040_, _09056_);
  or (_24103_, _24102_, _24101_);
  and (_24104_, _24103_, _09061_);
  and (_24105_, _24104_, _24100_);
  nor (_24106_, _11258_, _11985_);
  or (_24107_, _24106_, _24040_);
  and (_24108_, _24107_, _06528_);
  or (_24109_, _24108_, _24105_);
  and (_24110_, _24109_, _06926_);
  and (_24111_, _24045_, _06568_);
  or (_24113_, _24111_, _06278_);
  or (_24114_, _24113_, _24110_);
  and (_24115_, _14926_, _07910_);
  or (_24116_, _24040_, _06279_);
  or (_24117_, _24116_, _24115_);
  and (_24118_, _24117_, _01347_);
  and (_24119_, _24118_, _24114_);
  or (_24120_, _24119_, _24039_);
  and (_43230_, _24120_, _42618_);
  and (_24121_, _01351_, \oc8051_golden_model_1.TH1 [3]);
  and (_24123_, _11985_, \oc8051_golden_model_1.TH1 [3]);
  and (_24124_, _14953_, _07910_);
  or (_24125_, _24124_, _24123_);
  or (_24126_, _24125_, _07151_);
  and (_24127_, _07910_, \oc8051_golden_model_1.ACC [3]);
  or (_24128_, _24127_, _24123_);
  and (_24129_, _24128_, _07141_);
  and (_24130_, _07142_, \oc8051_golden_model_1.TH1 [3]);
  or (_24131_, _24130_, _06341_);
  or (_24132_, _24131_, _24129_);
  and (_24133_, _24132_, _07166_);
  and (_24134_, _24133_, _24126_);
  nor (_24135_, _11985_, _07594_);
  or (_24136_, _24135_, _24123_);
  and (_24137_, _24136_, _06461_);
  or (_24138_, _24137_, _24134_);
  and (_24139_, _24138_, _06465_);
  and (_24140_, _24128_, _06464_);
  or (_24141_, _24140_, _10080_);
  or (_24142_, _24141_, _24139_);
  or (_24144_, _24136_, _07215_);
  and (_24145_, _24144_, _24142_);
  or (_24146_, _24145_, _07460_);
  and (_24147_, _09449_, _07910_);
  or (_24148_, _24123_, _07208_);
  or (_24149_, _24148_, _24147_);
  and (_24150_, _24149_, _05982_);
  and (_24151_, _24150_, _24146_);
  and (_24152_, _15048_, _07910_);
  or (_24153_, _24152_, _24123_);
  and (_24155_, _24153_, _10094_);
  or (_24156_, _24155_, _06218_);
  or (_24157_, _24156_, _24151_);
  and (_24158_, _07910_, _08930_);
  or (_24159_, _24158_, _24123_);
  or (_24160_, _24159_, _06219_);
  and (_24161_, _24160_, _24157_);
  or (_24162_, _24161_, _06369_);
  and (_24163_, _14943_, _07910_);
  or (_24164_, _24163_, _24123_);
  or (_24166_, _24164_, _07237_);
  and (_24167_, _24166_, _07240_);
  and (_24168_, _24167_, _24162_);
  and (_24169_, _12577_, _07910_);
  or (_24170_, _24169_, _24123_);
  and (_24171_, _24170_, _06536_);
  or (_24172_, _24171_, _24168_);
  and (_24173_, _24172_, _07242_);
  or (_24174_, _24123_, _08292_);
  and (_24175_, _24159_, _06375_);
  and (_24177_, _24175_, _24174_);
  or (_24178_, _24177_, _24173_);
  and (_24179_, _24178_, _07234_);
  and (_24180_, _24128_, _06545_);
  and (_24181_, _24180_, _24174_);
  or (_24182_, _24181_, _06366_);
  or (_24183_, _24182_, _24179_);
  and (_24184_, _14940_, _07910_);
  or (_24185_, _24123_, _09056_);
  or (_24186_, _24185_, _24184_);
  and (_24188_, _24186_, _09061_);
  and (_24189_, _24188_, _24183_);
  nor (_24190_, _11256_, _11985_);
  or (_24191_, _24190_, _24123_);
  and (_24192_, _24191_, _06528_);
  or (_24193_, _24192_, _24189_);
  and (_24194_, _24193_, _06926_);
  and (_24195_, _24125_, _06568_);
  or (_24196_, _24195_, _06278_);
  or (_24197_, _24196_, _24194_);
  and (_24199_, _15128_, _07910_);
  or (_24200_, _24123_, _06279_);
  or (_24201_, _24200_, _24199_);
  and (_24202_, _24201_, _01347_);
  and (_24203_, _24202_, _24197_);
  or (_24204_, _24203_, _24121_);
  and (_43231_, _24204_, _42618_);
  and (_24205_, _01351_, \oc8051_golden_model_1.TH1 [4]);
  and (_24206_, _11985_, \oc8051_golden_model_1.TH1 [4]);
  nor (_24207_, _08541_, _11985_);
  or (_24209_, _24207_, _24206_);
  or (_24210_, _24209_, _07215_);
  and (_24211_, _15162_, _07910_);
  or (_24212_, _24211_, _24206_);
  or (_24213_, _24212_, _07151_);
  and (_24214_, _07910_, \oc8051_golden_model_1.ACC [4]);
  or (_24215_, _24214_, _24206_);
  and (_24216_, _24215_, _07141_);
  and (_24217_, _07142_, \oc8051_golden_model_1.TH1 [4]);
  or (_24218_, _24217_, _06341_);
  or (_24220_, _24218_, _24216_);
  and (_24221_, _24220_, _07166_);
  and (_24222_, _24221_, _24213_);
  and (_24223_, _24209_, _06461_);
  or (_24224_, _24223_, _24222_);
  and (_24225_, _24224_, _06465_);
  and (_24226_, _24215_, _06464_);
  or (_24227_, _24226_, _10080_);
  or (_24228_, _24227_, _24225_);
  and (_24229_, _24228_, _24210_);
  or (_24231_, _24229_, _07460_);
  and (_24232_, _09448_, _07910_);
  or (_24233_, _24206_, _07208_);
  or (_24234_, _24233_, _24232_);
  and (_24235_, _24234_, _24231_);
  or (_24236_, _24235_, _10094_);
  and (_24237_, _15254_, _07910_);
  or (_24238_, _24206_, _05982_);
  or (_24239_, _24238_, _24237_);
  and (_24240_, _24239_, _06219_);
  and (_24241_, _24240_, _24236_);
  and (_24242_, _08959_, _07910_);
  or (_24243_, _24242_, _24206_);
  and (_24244_, _24243_, _06218_);
  or (_24245_, _24244_, _06369_);
  or (_24246_, _24245_, _24241_);
  and (_24247_, _15269_, _07910_);
  or (_24248_, _24247_, _24206_);
  or (_24249_, _24248_, _07237_);
  and (_24250_, _24249_, _07240_);
  and (_24251_, _24250_, _24246_);
  and (_24252_, _11254_, _07910_);
  or (_24253_, _24252_, _24206_);
  and (_24254_, _24253_, _06536_);
  or (_24255_, _24254_, _24251_);
  and (_24256_, _24255_, _07242_);
  or (_24257_, _24206_, _08544_);
  and (_24258_, _24243_, _06375_);
  and (_24259_, _24258_, _24257_);
  or (_24260_, _24259_, _24256_);
  and (_24262_, _24260_, _07234_);
  and (_24263_, _24215_, _06545_);
  and (_24264_, _24263_, _24257_);
  or (_24265_, _24264_, _06366_);
  or (_24266_, _24265_, _24262_);
  and (_24267_, _15266_, _07910_);
  or (_24268_, _24206_, _09056_);
  or (_24269_, _24268_, _24267_);
  and (_24270_, _24269_, _09061_);
  and (_24271_, _24270_, _24266_);
  nor (_24273_, _11253_, _11985_);
  or (_24274_, _24273_, _24206_);
  and (_24275_, _24274_, _06528_);
  or (_24276_, _24275_, _24271_);
  and (_24277_, _24276_, _06926_);
  and (_24278_, _24212_, _06568_);
  or (_24279_, _24278_, _06278_);
  or (_24280_, _24279_, _24277_);
  and (_24281_, _15329_, _07910_);
  or (_24282_, _24206_, _06279_);
  or (_24285_, _24282_, _24281_);
  and (_24286_, _24285_, _01347_);
  and (_24287_, _24286_, _24280_);
  or (_24288_, _24287_, _24205_);
  and (_43232_, _24288_, _42618_);
  and (_24289_, _01351_, \oc8051_golden_model_1.TH1 [5]);
  and (_24290_, _11985_, \oc8051_golden_model_1.TH1 [5]);
  nor (_24291_, _08244_, _11985_);
  or (_24292_, _24291_, _24290_);
  or (_24293_, _24292_, _07215_);
  and (_24295_, _15358_, _07910_);
  or (_24296_, _24295_, _24290_);
  or (_24297_, _24296_, _07151_);
  and (_24298_, _07910_, \oc8051_golden_model_1.ACC [5]);
  or (_24299_, _24298_, _24290_);
  and (_24300_, _24299_, _07141_);
  and (_24301_, _07142_, \oc8051_golden_model_1.TH1 [5]);
  or (_24302_, _24301_, _06341_);
  or (_24303_, _24302_, _24300_);
  and (_24304_, _24303_, _07166_);
  and (_24306_, _24304_, _24297_);
  and (_24307_, _24292_, _06461_);
  or (_24308_, _24307_, _24306_);
  and (_24309_, _24308_, _06465_);
  and (_24310_, _24299_, _06464_);
  or (_24311_, _24310_, _10080_);
  or (_24312_, _24311_, _24309_);
  and (_24313_, _24312_, _24293_);
  or (_24314_, _24313_, _07460_);
  and (_24315_, _09447_, _07910_);
  or (_24317_, _24290_, _07208_);
  or (_24318_, _24317_, _24315_);
  and (_24319_, _24318_, _05982_);
  and (_24320_, _24319_, _24314_);
  and (_24321_, _15459_, _07910_);
  or (_24322_, _24321_, _24290_);
  and (_24323_, _24322_, _10094_);
  or (_24324_, _24323_, _06218_);
  or (_24325_, _24324_, _24320_);
  and (_24326_, _08946_, _07910_);
  or (_24328_, _24326_, _24290_);
  or (_24329_, _24328_, _06219_);
  and (_24330_, _24329_, _24325_);
  or (_24331_, _24330_, _06369_);
  and (_24332_, _15353_, _07910_);
  or (_24333_, _24332_, _24290_);
  or (_24334_, _24333_, _07237_);
  and (_24335_, _24334_, _07240_);
  and (_24336_, _24335_, _24331_);
  and (_24337_, _11250_, _07910_);
  or (_24339_, _24337_, _24290_);
  and (_24340_, _24339_, _06536_);
  or (_24341_, _24340_, _24336_);
  and (_24342_, _24341_, _07242_);
  or (_24343_, _24290_, _08247_);
  and (_24344_, _24328_, _06375_);
  and (_24345_, _24344_, _24343_);
  or (_24346_, _24345_, _24342_);
  and (_24347_, _24346_, _07234_);
  and (_24348_, _24299_, _06545_);
  and (_24350_, _24348_, _24343_);
  or (_24351_, _24350_, _06366_);
  or (_24352_, _24351_, _24347_);
  and (_24353_, _15350_, _07910_);
  or (_24354_, _24290_, _09056_);
  or (_24355_, _24354_, _24353_);
  and (_24356_, _24355_, _09061_);
  and (_24357_, _24356_, _24352_);
  nor (_24358_, _11249_, _11985_);
  or (_24359_, _24358_, _24290_);
  and (_24361_, _24359_, _06528_);
  or (_24362_, _24361_, _24357_);
  and (_24363_, _24362_, _06926_);
  and (_24364_, _24296_, _06568_);
  or (_24365_, _24364_, _06278_);
  or (_24366_, _24365_, _24363_);
  and (_24367_, _15532_, _07910_);
  or (_24368_, _24290_, _06279_);
  or (_24369_, _24368_, _24367_);
  and (_24370_, _24369_, _01347_);
  and (_24372_, _24370_, _24366_);
  or (_24373_, _24372_, _24289_);
  and (_43233_, _24373_, _42618_);
  and (_24374_, _01351_, \oc8051_golden_model_1.TH1 [6]);
  and (_24375_, _11985_, \oc8051_golden_model_1.TH1 [6]);
  and (_24376_, _15554_, _07910_);
  or (_24377_, _24376_, _24375_);
  or (_24378_, _24377_, _07151_);
  and (_24379_, _07910_, \oc8051_golden_model_1.ACC [6]);
  or (_24380_, _24379_, _24375_);
  and (_24382_, _24380_, _07141_);
  and (_24383_, _07142_, \oc8051_golden_model_1.TH1 [6]);
  or (_24384_, _24383_, _06341_);
  or (_24385_, _24384_, _24382_);
  and (_24386_, _24385_, _07166_);
  and (_24387_, _24386_, _24378_);
  nor (_24388_, _08142_, _11985_);
  or (_24389_, _24388_, _24375_);
  and (_24390_, _24389_, _06461_);
  or (_24391_, _24390_, _24387_);
  and (_24393_, _24391_, _06465_);
  and (_24394_, _24380_, _06464_);
  or (_24395_, _24394_, _10080_);
  or (_24396_, _24395_, _24393_);
  or (_24397_, _24389_, _07215_);
  and (_24398_, _24397_, _24396_);
  or (_24399_, _24398_, _07460_);
  and (_24400_, _09446_, _07910_);
  or (_24401_, _24375_, _07208_);
  or (_24402_, _24401_, _24400_);
  and (_24404_, _24402_, _05982_);
  and (_24405_, _24404_, _24399_);
  and (_24406_, _15657_, _07910_);
  or (_24407_, _24406_, _24375_);
  and (_24408_, _24407_, _10094_);
  or (_24409_, _24408_, _06218_);
  or (_24410_, _24409_, _24405_);
  and (_24411_, _15664_, _07910_);
  or (_24412_, _24411_, _24375_);
  or (_24413_, _24412_, _06219_);
  and (_24415_, _24413_, _24410_);
  or (_24416_, _24415_, _06369_);
  and (_24417_, _15549_, _07910_);
  or (_24418_, _24417_, _24375_);
  or (_24419_, _24418_, _07237_);
  and (_24420_, _24419_, _07240_);
  and (_24421_, _24420_, _24416_);
  and (_24422_, _11247_, _07910_);
  or (_24423_, _24422_, _24375_);
  and (_24424_, _24423_, _06536_);
  or (_24426_, _24424_, _24421_);
  and (_24427_, _24426_, _07242_);
  or (_24428_, _24375_, _08145_);
  and (_24429_, _24412_, _06375_);
  and (_24430_, _24429_, _24428_);
  or (_24431_, _24430_, _24427_);
  and (_24432_, _24431_, _07234_);
  and (_24433_, _24380_, _06545_);
  and (_24434_, _24433_, _24428_);
  or (_24435_, _24434_, _06366_);
  or (_24437_, _24435_, _24432_);
  and (_24438_, _15546_, _07910_);
  or (_24439_, _24375_, _09056_);
  or (_24440_, _24439_, _24438_);
  and (_24441_, _24440_, _09061_);
  and (_24442_, _24441_, _24437_);
  nor (_24443_, _11246_, _11985_);
  or (_24444_, _24443_, _24375_);
  and (_24445_, _24444_, _06528_);
  or (_24446_, _24445_, _24442_);
  and (_24448_, _24446_, _06926_);
  and (_24449_, _24377_, _06568_);
  or (_24450_, _24449_, _06278_);
  or (_24451_, _24450_, _24448_);
  and (_24452_, _15734_, _07910_);
  or (_24453_, _24375_, _06279_);
  or (_24454_, _24453_, _24452_);
  and (_24455_, _24454_, _01347_);
  and (_24456_, _24455_, _24451_);
  or (_24457_, _24456_, _24374_);
  and (_43234_, _24457_, _42618_);
  and (_24459_, _01351_, \oc8051_golden_model_1.TH0 [0]);
  and (_24460_, _07922_, \oc8051_golden_model_1.ACC [0]);
  and (_24461_, _24460_, _08390_);
  and (_24462_, _12063_, \oc8051_golden_model_1.TH0 [0]);
  or (_24463_, _24462_, _07234_);
  or (_24464_, _24463_, _24461_);
  or (_24465_, _24462_, _24460_);
  and (_24466_, _24465_, _06464_);
  or (_24467_, _24466_, _10080_);
  nor (_24469_, _08390_, _12063_);
  or (_24470_, _24469_, _24462_);
  and (_24471_, _24470_, _06341_);
  and (_24472_, _07142_, \oc8051_golden_model_1.TH0 [0]);
  and (_24473_, _24465_, _07141_);
  or (_24474_, _24473_, _24472_);
  and (_24475_, _24474_, _07151_);
  or (_24476_, _24475_, _06461_);
  or (_24477_, _24476_, _24471_);
  and (_24478_, _24477_, _06465_);
  or (_24480_, _24478_, _24467_);
  and (_24481_, _07922_, _07133_);
  or (_24482_, _24462_, _22611_);
  or (_24483_, _24482_, _24481_);
  and (_24484_, _24483_, _24480_);
  or (_24485_, _24484_, _07460_);
  and (_24486_, _09392_, _07922_);
  or (_24487_, _24462_, _07208_);
  or (_24488_, _24487_, _24486_);
  and (_24489_, _24488_, _24485_);
  or (_24491_, _24489_, _10094_);
  and (_24492_, _14467_, _07922_);
  or (_24493_, _24462_, _05982_);
  or (_24494_, _24493_, _24492_);
  and (_24495_, _24494_, _06219_);
  and (_24496_, _24495_, _24491_);
  and (_24497_, _07922_, _08954_);
  or (_24498_, _24497_, _24462_);
  and (_24499_, _24498_, _06218_);
  or (_24500_, _24499_, _06369_);
  or (_24502_, _24500_, _24496_);
  and (_24503_, _14366_, _07922_);
  or (_24504_, _24503_, _24462_);
  or (_24505_, _24504_, _07237_);
  and (_24506_, _24505_, _07240_);
  and (_24507_, _24506_, _24502_);
  nor (_24508_, _12580_, _12063_);
  or (_24509_, _24508_, _24462_);
  nor (_24510_, _24461_, _07240_);
  and (_24511_, _24510_, _24509_);
  or (_24512_, _24511_, _24507_);
  and (_24513_, _24512_, _07242_);
  nand (_24514_, _24498_, _06375_);
  nor (_24515_, _24514_, _24469_);
  or (_24516_, _24515_, _06545_);
  or (_24517_, _24516_, _24513_);
  and (_24518_, _24517_, _24464_);
  or (_24519_, _24518_, _06366_);
  and (_24520_, _14363_, _07922_);
  or (_24521_, _24462_, _09056_);
  or (_24524_, _24521_, _24520_);
  and (_24525_, _24524_, _09061_);
  and (_24526_, _24525_, _24519_);
  and (_24527_, _24509_, _06528_);
  or (_24528_, _24527_, _19502_);
  or (_24529_, _24528_, _24526_);
  or (_24530_, _24470_, _06661_);
  and (_24531_, _24530_, _01347_);
  and (_24532_, _24531_, _24529_);
  or (_24533_, _24532_, _24459_);
  and (_43236_, _24533_, _42618_);
  not (_24535_, \oc8051_golden_model_1.TH0 [1]);
  nor (_24536_, _01347_, _24535_);
  nor (_24537_, _07922_, _24535_);
  nor (_24538_, _12063_, _07357_);
  or (_24539_, _24538_, _24537_);
  or (_24540_, _24539_, _07215_);
  or (_24541_, _07922_, \oc8051_golden_model_1.TH0 [1]);
  and (_24542_, _14562_, _07922_);
  not (_24543_, _24542_);
  and (_24545_, _24543_, _24541_);
  or (_24546_, _24545_, _07151_);
  and (_24547_, _07922_, \oc8051_golden_model_1.ACC [1]);
  or (_24548_, _24547_, _24537_);
  and (_24549_, _24548_, _07141_);
  nor (_24550_, _07141_, _24535_);
  or (_24551_, _24550_, _06341_);
  or (_24552_, _24551_, _24549_);
  and (_24553_, _24552_, _07166_);
  and (_24554_, _24553_, _24546_);
  and (_24556_, _24539_, _06461_);
  or (_24557_, _24556_, _24554_);
  and (_24558_, _24557_, _06465_);
  and (_24559_, _24548_, _06464_);
  or (_24560_, _24559_, _10080_);
  or (_24561_, _24560_, _24558_);
  and (_24562_, _24561_, _24540_);
  or (_24563_, _24562_, _07460_);
  and (_24564_, _09451_, _07922_);
  or (_24565_, _24537_, _07208_);
  or (_24567_, _24565_, _24564_);
  and (_24568_, _24567_, _05982_);
  and (_24569_, _24568_, _24563_);
  or (_24570_, _14653_, _12063_);
  and (_24571_, _24541_, _10094_);
  and (_24572_, _24571_, _24570_);
  or (_24573_, _24572_, _24569_);
  and (_24574_, _24573_, _06219_);
  nand (_24575_, _07922_, _07038_);
  and (_24576_, _24541_, _06218_);
  and (_24578_, _24576_, _24575_);
  or (_24579_, _24578_, _24574_);
  and (_24580_, _24579_, _07237_);
  or (_24581_, _14668_, _12063_);
  and (_24582_, _24541_, _06369_);
  and (_24583_, _24582_, _24581_);
  or (_24584_, _24583_, _06536_);
  or (_24585_, _24584_, _24580_);
  nor (_24586_, _11261_, _12063_);
  or (_24587_, _24586_, _24537_);
  nand (_24589_, _11260_, _07922_);
  and (_24590_, _24589_, _24587_);
  or (_24591_, _24590_, _07240_);
  and (_24592_, _24591_, _07242_);
  and (_24593_, _24592_, _24585_);
  or (_24594_, _14666_, _12063_);
  and (_24595_, _24541_, _06375_);
  and (_24596_, _24595_, _24594_);
  or (_24597_, _24596_, _06545_);
  or (_24598_, _24597_, _24593_);
  nor (_24600_, _24537_, _07234_);
  nand (_24601_, _24600_, _24589_);
  and (_24602_, _24601_, _09056_);
  and (_24603_, _24602_, _24598_);
  or (_24604_, _24575_, _08341_);
  and (_24605_, _24541_, _06366_);
  and (_24606_, _24605_, _24604_);
  or (_24607_, _24606_, _06528_);
  or (_24608_, _24607_, _24603_);
  or (_24609_, _24587_, _09061_);
  and (_24611_, _24609_, _06926_);
  and (_24612_, _24611_, _24608_);
  and (_24613_, _24545_, _06568_);
  or (_24614_, _24613_, _06278_);
  or (_24615_, _24614_, _24612_);
  or (_24616_, _24537_, _06279_);
  or (_24617_, _24616_, _24542_);
  and (_24618_, _24617_, _01347_);
  and (_24619_, _24618_, _24615_);
  or (_24620_, _24619_, _24536_);
  and (_43237_, _24620_, _42618_);
  and (_24622_, _01351_, \oc8051_golden_model_1.TH0 [2]);
  and (_24623_, _12063_, \oc8051_golden_model_1.TH0 [2]);
  and (_24624_, _09450_, _07922_);
  or (_24625_, _24624_, _24623_);
  and (_24626_, _24625_, _07460_);
  and (_24627_, _14770_, _07922_);
  or (_24628_, _24627_, _24623_);
  or (_24629_, _24628_, _07151_);
  and (_24630_, _07922_, \oc8051_golden_model_1.ACC [2]);
  or (_24632_, _24630_, _24623_);
  and (_24633_, _24632_, _07141_);
  and (_24634_, _07142_, \oc8051_golden_model_1.TH0 [2]);
  or (_24635_, _24634_, _06341_);
  or (_24636_, _24635_, _24633_);
  and (_24637_, _24636_, _07166_);
  and (_24638_, _24637_, _24629_);
  nor (_24639_, _12063_, _07776_);
  or (_24640_, _24639_, _24623_);
  and (_24641_, _24640_, _06461_);
  or (_24643_, _24641_, _24638_);
  and (_24644_, _24643_, _06465_);
  and (_24645_, _24632_, _06464_);
  or (_24646_, _24645_, _10080_);
  or (_24647_, _24646_, _24644_);
  or (_24648_, _24640_, _07215_);
  and (_24649_, _24648_, _07208_);
  and (_24650_, _24649_, _24647_);
  or (_24651_, _24650_, _10094_);
  or (_24652_, _24651_, _24626_);
  and (_24654_, _14859_, _07922_);
  or (_24655_, _24623_, _05982_);
  or (_24656_, _24655_, _24654_);
  and (_24657_, _24656_, _06219_);
  and (_24658_, _24657_, _24652_);
  and (_24659_, _07922_, _08973_);
  or (_24660_, _24659_, _24623_);
  and (_24661_, _24660_, _06218_);
  or (_24662_, _24661_, _06369_);
  or (_24663_, _24662_, _24658_);
  and (_24665_, _14751_, _07922_);
  or (_24666_, _24665_, _24623_);
  or (_24667_, _24666_, _07237_);
  and (_24668_, _24667_, _07240_);
  and (_24669_, _24668_, _24663_);
  and (_24670_, _11259_, _07922_);
  or (_24671_, _24670_, _24623_);
  and (_24672_, _24671_, _06536_);
  or (_24673_, _24672_, _24669_);
  and (_24674_, _24673_, _07242_);
  or (_24676_, _24623_, _08440_);
  and (_24677_, _24660_, _06375_);
  and (_24678_, _24677_, _24676_);
  or (_24679_, _24678_, _24674_);
  and (_24680_, _24679_, _07234_);
  and (_24681_, _24632_, _06545_);
  and (_24682_, _24681_, _24676_);
  or (_24683_, _24682_, _06366_);
  or (_24684_, _24683_, _24680_);
  and (_24685_, _14748_, _07922_);
  or (_24687_, _24623_, _09056_);
  or (_24688_, _24687_, _24685_);
  and (_24689_, _24688_, _09061_);
  and (_24690_, _24689_, _24684_);
  nor (_24691_, _11258_, _12063_);
  or (_24692_, _24691_, _24623_);
  and (_24693_, _24692_, _06528_);
  or (_24694_, _24693_, _24690_);
  and (_24695_, _24694_, _06926_);
  and (_24696_, _24628_, _06568_);
  or (_24698_, _24696_, _06278_);
  or (_24699_, _24698_, _24695_);
  and (_24700_, _14926_, _07922_);
  or (_24701_, _24623_, _06279_);
  or (_24702_, _24701_, _24700_);
  and (_24703_, _24702_, _01347_);
  and (_24704_, _24703_, _24699_);
  or (_24705_, _24704_, _24622_);
  and (_43238_, _24705_, _42618_);
  and (_24706_, _01351_, \oc8051_golden_model_1.TH0 [3]);
  and (_24708_, _12063_, \oc8051_golden_model_1.TH0 [3]);
  and (_24709_, _14953_, _07922_);
  or (_24710_, _24709_, _24708_);
  or (_24711_, _24710_, _07151_);
  and (_24712_, _07922_, \oc8051_golden_model_1.ACC [3]);
  or (_24713_, _24712_, _24708_);
  and (_24714_, _24713_, _07141_);
  and (_24715_, _07142_, \oc8051_golden_model_1.TH0 [3]);
  or (_24716_, _24715_, _06341_);
  or (_24717_, _24716_, _24714_);
  and (_24719_, _24717_, _07166_);
  and (_24720_, _24719_, _24711_);
  nor (_24721_, _12063_, _07594_);
  or (_24722_, _24721_, _24708_);
  and (_24723_, _24722_, _06461_);
  or (_24724_, _24723_, _24720_);
  and (_24725_, _24724_, _06465_);
  and (_24726_, _24713_, _06464_);
  or (_24727_, _24726_, _10080_);
  or (_24728_, _24727_, _24725_);
  or (_24730_, _24722_, _07215_);
  and (_24731_, _24730_, _24728_);
  or (_24732_, _24731_, _07460_);
  and (_24733_, _09449_, _07922_);
  or (_24734_, _24708_, _07208_);
  or (_24735_, _24734_, _24733_);
  and (_24736_, _24735_, _05982_);
  and (_24737_, _24736_, _24732_);
  and (_24738_, _15048_, _07922_);
  or (_24739_, _24738_, _24708_);
  and (_24741_, _24739_, _10094_);
  or (_24742_, _24741_, _06218_);
  or (_24743_, _24742_, _24737_);
  and (_24744_, _07922_, _08930_);
  or (_24745_, _24744_, _24708_);
  or (_24746_, _24745_, _06219_);
  and (_24747_, _24746_, _24743_);
  or (_24748_, _24747_, _06369_);
  and (_24749_, _14943_, _07922_);
  or (_24750_, _24749_, _24708_);
  or (_24752_, _24750_, _07237_);
  and (_24753_, _24752_, _07240_);
  and (_24754_, _24753_, _24748_);
  and (_24755_, _12577_, _07922_);
  or (_24756_, _24755_, _24708_);
  and (_24757_, _24756_, _06536_);
  or (_24758_, _24757_, _24754_);
  and (_24759_, _24758_, _07242_);
  or (_24760_, _24708_, _08292_);
  and (_24761_, _24745_, _06375_);
  and (_24763_, _24761_, _24760_);
  or (_24764_, _24763_, _24759_);
  and (_24765_, _24764_, _07234_);
  and (_24766_, _24713_, _06545_);
  and (_24767_, _24766_, _24760_);
  or (_24768_, _24767_, _06366_);
  or (_24769_, _24768_, _24765_);
  and (_24770_, _14940_, _07922_);
  or (_24771_, _24708_, _09056_);
  or (_24772_, _24771_, _24770_);
  and (_24774_, _24772_, _09061_);
  and (_24775_, _24774_, _24769_);
  nor (_24776_, _11256_, _12063_);
  or (_24777_, _24776_, _24708_);
  and (_24778_, _24777_, _06528_);
  or (_24779_, _24778_, _24775_);
  and (_24780_, _24779_, _06926_);
  and (_24781_, _24710_, _06568_);
  or (_24782_, _24781_, _06278_);
  or (_24783_, _24782_, _24780_);
  and (_24785_, _15128_, _07922_);
  or (_24786_, _24708_, _06279_);
  or (_24787_, _24786_, _24785_);
  and (_24788_, _24787_, _01347_);
  and (_24789_, _24788_, _24783_);
  or (_24790_, _24789_, _24706_);
  and (_43239_, _24790_, _42618_);
  and (_24791_, _01351_, \oc8051_golden_model_1.TH0 [4]);
  and (_24792_, _12063_, \oc8051_golden_model_1.TH0 [4]);
  and (_24793_, _15162_, _07922_);
  or (_24795_, _24793_, _24792_);
  or (_24796_, _24795_, _07151_);
  and (_24797_, _07922_, \oc8051_golden_model_1.ACC [4]);
  or (_24798_, _24797_, _24792_);
  and (_24799_, _24798_, _07141_);
  and (_24800_, _07142_, \oc8051_golden_model_1.TH0 [4]);
  or (_24801_, _24800_, _06341_);
  or (_24802_, _24801_, _24799_);
  and (_24803_, _24802_, _07166_);
  and (_24804_, _24803_, _24796_);
  nor (_24806_, _08541_, _12063_);
  or (_24807_, _24806_, _24792_);
  and (_24808_, _24807_, _06461_);
  or (_24809_, _24808_, _24804_);
  and (_24810_, _24809_, _06465_);
  and (_24811_, _24798_, _06464_);
  or (_24812_, _24811_, _10080_);
  or (_24813_, _24812_, _24810_);
  or (_24814_, _24807_, _07215_);
  and (_24815_, _24814_, _24813_);
  or (_24817_, _24815_, _07460_);
  and (_24818_, _09448_, _07922_);
  or (_24819_, _24792_, _07208_);
  or (_24820_, _24819_, _24818_);
  and (_24821_, _24820_, _24817_);
  or (_24822_, _24821_, _10094_);
  and (_24823_, _15254_, _07922_);
  or (_24824_, _24792_, _05982_);
  or (_24825_, _24824_, _24823_);
  and (_24826_, _24825_, _06219_);
  and (_24828_, _24826_, _24822_);
  and (_24829_, _08959_, _07922_);
  or (_24830_, _24829_, _24792_);
  and (_24831_, _24830_, _06218_);
  or (_24832_, _24831_, _06369_);
  or (_24833_, _24832_, _24828_);
  and (_24834_, _15269_, _07922_);
  or (_24835_, _24834_, _24792_);
  or (_24836_, _24835_, _07237_);
  and (_24837_, _24836_, _07240_);
  and (_24839_, _24837_, _24833_);
  and (_24840_, _11254_, _07922_);
  or (_24841_, _24840_, _24792_);
  and (_24842_, _24841_, _06536_);
  or (_24843_, _24842_, _24839_);
  and (_24844_, _24843_, _07242_);
  or (_24845_, _24792_, _08544_);
  and (_24846_, _24830_, _06375_);
  and (_24847_, _24846_, _24845_);
  or (_24848_, _24847_, _24844_);
  and (_24850_, _24848_, _07234_);
  and (_24851_, _24798_, _06545_);
  and (_24852_, _24851_, _24845_);
  or (_24853_, _24852_, _06366_);
  or (_24854_, _24853_, _24850_);
  and (_24855_, _15266_, _07922_);
  or (_24856_, _24792_, _09056_);
  or (_24857_, _24856_, _24855_);
  and (_24858_, _24857_, _09061_);
  and (_24859_, _24858_, _24854_);
  nor (_24861_, _11253_, _12063_);
  or (_24862_, _24861_, _24792_);
  and (_24863_, _24862_, _06528_);
  or (_24864_, _24863_, _24859_);
  and (_24865_, _24864_, _06926_);
  and (_24866_, _24795_, _06568_);
  or (_24867_, _24866_, _06278_);
  or (_24868_, _24867_, _24865_);
  and (_24869_, _15329_, _07922_);
  or (_24870_, _24792_, _06279_);
  or (_24872_, _24870_, _24869_);
  and (_24873_, _24872_, _01347_);
  and (_24874_, _24873_, _24868_);
  or (_24875_, _24874_, _24791_);
  and (_43240_, _24875_, _42618_);
  and (_24876_, _01351_, \oc8051_golden_model_1.TH0 [5]);
  and (_24877_, _12063_, \oc8051_golden_model_1.TH0 [5]);
  nor (_24878_, _08244_, _12063_);
  or (_24879_, _24878_, _24877_);
  or (_24880_, _24879_, _07215_);
  and (_24882_, _15358_, _07922_);
  or (_24883_, _24882_, _24877_);
  or (_24884_, _24883_, _07151_);
  and (_24885_, _07922_, \oc8051_golden_model_1.ACC [5]);
  or (_24886_, _24885_, _24877_);
  and (_24887_, _24886_, _07141_);
  and (_24888_, _07142_, \oc8051_golden_model_1.TH0 [5]);
  or (_24889_, _24888_, _06341_);
  or (_24890_, _24889_, _24887_);
  and (_24891_, _24890_, _07166_);
  and (_24893_, _24891_, _24884_);
  and (_24894_, _24879_, _06461_);
  or (_24895_, _24894_, _24893_);
  and (_24896_, _24895_, _06465_);
  and (_24897_, _24886_, _06464_);
  or (_24898_, _24897_, _10080_);
  or (_24899_, _24898_, _24896_);
  and (_24900_, _24899_, _24880_);
  or (_24901_, _24900_, _07460_);
  and (_24902_, _09447_, _07922_);
  or (_24904_, _24877_, _07208_);
  or (_24905_, _24904_, _24902_);
  and (_24906_, _24905_, _05982_);
  and (_24907_, _24906_, _24901_);
  and (_24908_, _15459_, _07922_);
  or (_24909_, _24908_, _24877_);
  and (_24910_, _24909_, _10094_);
  or (_24911_, _24910_, _06218_);
  or (_24912_, _24911_, _24907_);
  and (_24913_, _08946_, _07922_);
  or (_24915_, _24913_, _24877_);
  or (_24916_, _24915_, _06219_);
  and (_24917_, _24916_, _24912_);
  or (_24918_, _24917_, _06369_);
  and (_24919_, _15353_, _07922_);
  or (_24920_, _24919_, _24877_);
  or (_24921_, _24920_, _07237_);
  and (_24922_, _24921_, _07240_);
  and (_24923_, _24922_, _24918_);
  and (_24924_, _11250_, _07922_);
  or (_24926_, _24924_, _24877_);
  and (_24927_, _24926_, _06536_);
  or (_24928_, _24927_, _24923_);
  and (_24929_, _24928_, _07242_);
  or (_24930_, _24877_, _08247_);
  and (_24931_, _24915_, _06375_);
  and (_24932_, _24931_, _24930_);
  or (_24933_, _24932_, _24929_);
  and (_24934_, _24933_, _07234_);
  and (_24935_, _24886_, _06545_);
  and (_24937_, _24935_, _24930_);
  or (_24938_, _24937_, _06366_);
  or (_24939_, _24938_, _24934_);
  and (_24940_, _15350_, _07922_);
  or (_24941_, _24877_, _09056_);
  or (_24942_, _24941_, _24940_);
  and (_24943_, _24942_, _09061_);
  and (_24944_, _24943_, _24939_);
  nor (_24945_, _11249_, _12063_);
  or (_24946_, _24945_, _24877_);
  and (_24948_, _24946_, _06528_);
  or (_24949_, _24948_, _24944_);
  and (_24950_, _24949_, _06926_);
  and (_24951_, _24883_, _06568_);
  or (_24952_, _24951_, _06278_);
  or (_24953_, _24952_, _24950_);
  and (_24954_, _15532_, _07922_);
  or (_24955_, _24877_, _06279_);
  or (_24956_, _24955_, _24954_);
  and (_24957_, _24956_, _01347_);
  and (_24959_, _24957_, _24953_);
  or (_24960_, _24959_, _24876_);
  and (_43242_, _24960_, _42618_);
  and (_24961_, _01351_, \oc8051_golden_model_1.TH0 [6]);
  and (_24962_, _12063_, \oc8051_golden_model_1.TH0 [6]);
  nor (_24963_, _08142_, _12063_);
  or (_24964_, _24963_, _24962_);
  or (_24965_, _24964_, _07215_);
  and (_24966_, _15554_, _07922_);
  or (_24967_, _24966_, _24962_);
  or (_24969_, _24967_, _07151_);
  and (_24970_, _07922_, \oc8051_golden_model_1.ACC [6]);
  or (_24971_, _24970_, _24962_);
  and (_24972_, _24971_, _07141_);
  and (_24973_, _07142_, \oc8051_golden_model_1.TH0 [6]);
  or (_24974_, _24973_, _06341_);
  or (_24975_, _24974_, _24972_);
  and (_24976_, _24975_, _07166_);
  and (_24977_, _24976_, _24969_);
  and (_24978_, _24964_, _06461_);
  or (_24980_, _24978_, _24977_);
  and (_24981_, _24980_, _06465_);
  and (_24982_, _24971_, _06464_);
  or (_24983_, _24982_, _10080_);
  or (_24984_, _24983_, _24981_);
  and (_24985_, _24984_, _24965_);
  or (_24986_, _24985_, _07460_);
  and (_24987_, _09446_, _07922_);
  or (_24988_, _24962_, _07208_);
  or (_24989_, _24988_, _24987_);
  and (_24991_, _24989_, _05982_);
  and (_24992_, _24991_, _24986_);
  and (_24993_, _15657_, _07922_);
  or (_24994_, _24993_, _24962_);
  and (_24995_, _24994_, _10094_);
  or (_24996_, _24995_, _06218_);
  or (_24997_, _24996_, _24992_);
  and (_24998_, _15664_, _07922_);
  or (_24999_, _24998_, _24962_);
  or (_25000_, _24999_, _06219_);
  and (_25002_, _25000_, _24997_);
  or (_25003_, _25002_, _06369_);
  and (_25004_, _15549_, _07922_);
  or (_25005_, _25004_, _24962_);
  or (_25006_, _25005_, _07237_);
  and (_25007_, _25006_, _07240_);
  and (_25008_, _25007_, _25003_);
  and (_25009_, _11247_, _07922_);
  or (_25010_, _25009_, _24962_);
  and (_25011_, _25010_, _06536_);
  or (_25013_, _25011_, _25008_);
  and (_25014_, _25013_, _07242_);
  or (_25015_, _24962_, _08145_);
  and (_25016_, _24999_, _06375_);
  and (_25017_, _25016_, _25015_);
  or (_25018_, _25017_, _25014_);
  and (_25019_, _25018_, _07234_);
  and (_25020_, _24971_, _06545_);
  and (_25021_, _25020_, _25015_);
  or (_25022_, _25021_, _06366_);
  or (_25024_, _25022_, _25019_);
  and (_25025_, _15546_, _07922_);
  or (_25026_, _24962_, _09056_);
  or (_25027_, _25026_, _25025_);
  and (_25028_, _25027_, _09061_);
  and (_25029_, _25028_, _25024_);
  nor (_25030_, _11246_, _12063_);
  or (_25031_, _25030_, _24962_);
  and (_25032_, _25031_, _06528_);
  or (_25033_, _25032_, _25029_);
  and (_25035_, _25033_, _06926_);
  and (_25036_, _24967_, _06568_);
  or (_25037_, _25036_, _06278_);
  or (_25038_, _25037_, _25035_);
  and (_25039_, _15734_, _07922_);
  or (_25040_, _24962_, _06279_);
  or (_25041_, _25040_, _25039_);
  and (_25042_, _25041_, _01347_);
  and (_25043_, _25042_, _25038_);
  or (_25044_, _25043_, _24961_);
  and (_43243_, _25044_, _42618_);
  and (_25046_, _13052_, _12141_);
  nor (_25047_, _25046_, _05630_);
  and (_25048_, _13030_, _13037_);
  nor (_25049_, _25048_, _05630_);
  and (_25050_, _12151_, _11285_);
  nor (_25051_, _25050_, _05630_);
  and (_25052_, _10559_, \oc8051_golden_model_1.PC [0]);
  nor (_25053_, _10559_, \oc8051_golden_model_1.PC [0]);
  nor (_25054_, _25053_, _25052_);
  and (_25055_, _25054_, _12800_);
  not (_25056_, _12800_);
  and (_25057_, _12162_, _09056_);
  nor (_25058_, _25057_, _05630_);
  and (_25059_, _10979_, _07242_);
  nor (_25060_, _25059_, _05630_);
  not (_25061_, _12755_);
  and (_25062_, _12169_, _07237_);
  nor (_25063_, _25062_, _05630_);
  not (_25064_, _12733_);
  and (_25067_, _06218_, _05630_);
  nor (_25068_, _06872_, _06007_);
  and (_25069_, _12587_, _05630_);
  and (_25070_, _06872_, \oc8051_golden_model_1.PC [0]);
  nor (_25071_, _25070_, _12251_);
  not (_25072_, _25071_);
  nor (_25073_, _25072_, _12587_);
  nor (_25074_, _25073_, _25069_);
  nor (_25075_, _25074_, _06774_);
  and (_25076_, _12333_, _05630_);
  not (_25078_, _25076_);
  and (_25079_, _25071_, _12335_);
  nor (_25080_, _25079_, _12177_);
  and (_25081_, _25080_, _25078_);
  nor (_25082_, _06872_, _06013_);
  and (_25083_, _12513_, _05630_);
  nor (_25084_, _12513_, _05630_);
  nor (_25085_, _25084_, _25083_);
  and (_25086_, _25085_, _07504_);
  nor (_25087_, _06872_, _07504_);
  or (_25089_, _25087_, _12516_);
  nor (_25090_, _25089_, _25086_);
  nor (_25091_, _12512_, _05630_);
  nor (_25092_, _25091_, _25090_);
  nor (_25093_, _25092_, _12387_);
  and (_25094_, _12507_, \oc8051_golden_model_1.PC [0]);
  and (_25095_, _06251_, _05630_);
  nor (_25096_, _25095_, _12458_);
  and (_25097_, _25096_, _12393_);
  or (_25098_, _25097_, _25094_);
  nor (_25100_, _25098_, _08654_);
  nor (_25101_, _25100_, _25093_);
  nor (_25102_, _25101_, _07154_);
  and (_25103_, _07154_, \oc8051_golden_model_1.PC [0]);
  nor (_25104_, _25103_, _06341_);
  not (_25105_, _25104_);
  nor (_25106_, _25105_, _25102_);
  not (_25107_, _25106_);
  and (_25108_, _25072_, _12534_);
  and (_25109_, _12536_, \oc8051_golden_model_1.PC [0]);
  or (_25111_, _25109_, _07151_);
  nor (_25112_, _25111_, _25108_);
  nor (_25113_, _25112_, _12542_);
  and (_25114_, _25113_, _25107_);
  nor (_25115_, _12541_, _05630_);
  nor (_25116_, _25115_, _07611_);
  not (_25117_, _25116_);
  nor (_25118_, _25117_, _25114_);
  nor (_25119_, _06872_, _06010_);
  and (_25120_, _12560_, _12550_);
  not (_25122_, _25120_);
  nor (_25123_, _25122_, _25119_);
  not (_25124_, _25123_);
  nor (_25125_, _25124_, _25118_);
  nor (_25126_, _25120_, _05630_);
  nor (_25127_, _25126_, _12563_);
  not (_25128_, _25127_);
  nor (_25129_, _25128_, _25125_);
  or (_25130_, _25129_, _12379_);
  nor (_25131_, _25130_, _25082_);
  and (_25133_, _12371_, _05630_);
  not (_25134_, _25133_);
  nor (_25135_, _25072_, _12371_);
  nor (_25136_, _25135_, _12378_);
  and (_25137_, _25136_, _25134_);
  nor (_25138_, _25137_, _25131_);
  nor (_25139_, _25138_, _06347_);
  nor (_25140_, _25139_, _06480_);
  not (_25141_, _25140_);
  nor (_25142_, _25141_, _25081_);
  nor (_25144_, _25142_, _25075_);
  nor (_25145_, _25144_, _06371_);
  and (_25146_, _12604_, _05630_);
  nor (_25147_, _25072_, _12604_);
  or (_25148_, _25147_, _25146_);
  and (_25149_, _25148_, _06371_);
  or (_25150_, _25149_, _25145_);
  and (_25151_, _25150_, _12175_);
  and (_25152_, _12174_, _05630_);
  or (_25153_, _25152_, _25151_);
  and (_25155_, _25153_, _06007_);
  or (_25156_, _25155_, _12631_);
  nor (_25157_, _25156_, _25068_);
  not (_25158_, _06020_);
  nor (_25159_, _12630_, _05630_);
  nor (_25160_, _25159_, _25158_);
  not (_25161_, _25160_);
  nor (_25162_, _25161_, _25157_);
  nor (_25163_, _06872_, _06020_);
  and (_25164_, _12639_, _05984_);
  not (_25166_, _25164_);
  nor (_25167_, _25166_, _25163_);
  not (_25168_, _25167_);
  nor (_25169_, _25168_, _25162_);
  nor (_25170_, _25164_, _05630_);
  nor (_25171_, _25170_, _06254_);
  not (_25172_, _25171_);
  nor (_25173_, _25172_, _25169_);
  nor (_25174_, _06872_, _05978_);
  nor (_25175_, _06373_, _10094_);
  and (_25177_, _25175_, _12172_);
  not (_25178_, _25177_);
  nor (_25179_, _25178_, _25174_);
  not (_25180_, _25179_);
  nor (_25181_, _25180_, _25173_);
  nor (_25182_, _25177_, _05630_);
  nor (_25183_, _25182_, _12668_);
  not (_25184_, _25183_);
  nor (_25185_, _25184_, _25181_);
  nor (_25186_, _06872_, _05946_);
  or (_25188_, _25186_, _12674_);
  or (_25189_, _25188_, _25185_);
  or (_25190_, _25096_, _12679_);
  and (_25191_, _25190_, _25189_);
  and (_25192_, _25191_, _06219_);
  or (_25193_, _25192_, _25067_);
  and (_25194_, _25193_, _12691_);
  and (_25195_, _12690_, _06090_);
  or (_25196_, _25195_, _25194_);
  and (_25197_, _25196_, _05952_);
  nor (_25199_, _06872_, _05952_);
  or (_25200_, _25199_, _25197_);
  and (_25201_, _25200_, _25064_);
  not (_25202_, _25062_);
  nor (_25203_, _25096_, _11342_);
  and (_25204_, _11342_, _05630_);
  nor (_25205_, _25204_, _25064_);
  not (_25206_, _25205_);
  nor (_25207_, _25206_, _25203_);
  nor (_25208_, _25207_, _25202_);
  not (_25210_, _25208_);
  nor (_25211_, _25210_, _25201_);
  nor (_25212_, _25211_, _25063_);
  and (_25213_, _25212_, _05955_);
  nor (_25214_, _06872_, _05955_);
  or (_25215_, _25214_, _25213_);
  and (_25216_, _25215_, _25061_);
  not (_25217_, _25059_);
  nor (_25218_, _11342_, _05630_);
  and (_25219_, _25096_, _11342_);
  or (_25221_, _25219_, _25218_);
  and (_25222_, _25221_, _12755_);
  nor (_25223_, _25222_, _25217_);
  not (_25224_, _25223_);
  nor (_25225_, _25224_, _25216_);
  nor (_25226_, _25225_, _25060_);
  and (_25227_, _25226_, _05961_);
  nor (_25228_, _06872_, _05961_);
  or (_25229_, _25228_, _25227_);
  and (_25230_, _25229_, _12782_);
  not (_25232_, _25057_);
  and (_25233_, \oc8051_golden_model_1.PSW [7], \oc8051_golden_model_1.PC [0]);
  and (_25234_, _25096_, _10558_);
  or (_25235_, _25234_, _25233_);
  and (_25236_, _25235_, _12776_);
  nor (_25237_, _25236_, _25232_);
  not (_25238_, _25237_);
  nor (_25239_, _25238_, _25230_);
  nor (_25240_, _25239_, _25058_);
  and (_25241_, _25240_, _05966_);
  nor (_25243_, _06872_, _05966_);
  or (_25244_, _25243_, _25241_);
  and (_25245_, _25244_, _25056_);
  and (_25246_, _12154_, _11126_);
  not (_25247_, _25246_);
  or (_25248_, _25247_, _25245_);
  nor (_25249_, _25248_, _25055_);
  nor (_25250_, _25246_, _05630_);
  nor (_25251_, _25250_, _06551_);
  not (_25252_, _25251_);
  nor (_25254_, _25252_, _25249_);
  and (_25255_, _09392_, _06551_);
  or (_25256_, _25255_, _25254_);
  and (_25257_, _25256_, _05959_);
  nor (_25258_, _06872_, _05959_);
  or (_25259_, _25258_, _25257_);
  and (_25260_, _25259_, _06558_);
  and (_25261_, _25072_, _13004_);
  nor (_25262_, _13004_, _05630_);
  or (_25263_, _25262_, _06558_);
  or (_25265_, _25263_, _25261_);
  and (_25266_, _25265_, _25050_);
  not (_25267_, _25266_);
  nor (_25268_, _25267_, _25260_);
  nor (_25269_, _25268_, _25051_);
  and (_25270_, _25269_, _06282_);
  and (_25271_, _09392_, _06281_);
  or (_25272_, _25271_, _25270_);
  and (_25273_, _25272_, _05964_);
  nor (_25274_, _06872_, _05964_);
  nor (_25276_, _25274_, _25273_);
  nor (_25277_, _25276_, _06362_);
  not (_25278_, _25048_);
  and (_25279_, _13004_, \oc8051_golden_model_1.PC [0]);
  nor (_25280_, _25071_, _13004_);
  nor (_25281_, _25280_, _25279_);
  and (_25282_, _25281_, _06362_);
  nor (_25283_, _25282_, _25278_);
  not (_25284_, _25283_);
  nor (_25285_, _25284_, _25277_);
  nor (_25287_, _25285_, _25049_);
  nor (_25288_, _25287_, _07695_);
  and (_25289_, _07695_, _06872_);
  nor (_25290_, _25289_, _05927_);
  not (_25291_, _25290_);
  or (_25292_, _25291_, _25288_);
  not (_25293_, _25046_);
  and (_25294_, _25281_, _05927_);
  nor (_25295_, _25294_, _25293_);
  and (_25296_, _25295_, _25292_);
  or (_25298_, _25296_, _25047_);
  nor (_25299_, _06379_, _05939_);
  nand (_25300_, _25299_, _25298_);
  not (_25301_, _25299_);
  and (_25302_, _25301_, _06872_);
  nor (_25303_, _25302_, _13068_);
  and (_25304_, _25303_, _25300_);
  and (_25305_, _13068_, _05630_);
  or (_25306_, _25305_, _25304_);
  or (_25307_, _25306_, _01351_);
  or (_25309_, _01347_, \oc8051_golden_model_1.PC [0]);
  and (_25310_, _25309_, _42618_);
  and (_43245_, _25310_, _25307_);
  and (_25311_, _06278_, _05597_);
  nor (_25312_, _13037_, _06111_);
  nor (_25313_, _08568_, _06111_);
  nor (_25314_, _12151_, _06111_);
  nor (_25315_, _12154_, _06111_);
  nor (_25316_, _12157_, _06111_);
  nor (_25317_, _10979_, _06111_);
  nor (_25318_, _12169_, _06111_);
  nor (_25319_, _09030_, _05597_);
  nor (_25320_, _12639_, _06111_);
  and (_25321_, _12621_, _12616_);
  and (_25322_, _25321_, _12620_);
  nor (_25323_, _25322_, _05597_);
  and (_25324_, _12174_, _06043_);
  and (_25325_, _12371_, _06043_);
  nor (_25326_, _12253_, _12251_);
  nor (_25327_, _25326_, _12254_);
  not (_25330_, _25327_);
  nor (_25331_, _25330_, _12371_);
  or (_25332_, _25331_, _25325_);
  nor (_25333_, _25332_, _12378_);
  nor (_25334_, _12560_, _06111_);
  and (_25335_, _10759_, _06784_);
  nor (_25336_, _25335_, _06111_);
  and (_25337_, _10754_, _06043_);
  nor (_25338_, _07038_, _07504_);
  and (_25339_, _07486_, \oc8051_golden_model_1.PC [0]);
  nor (_25341_, _25339_, _07141_);
  nor (_25342_, _25341_, \oc8051_golden_model_1.PC [1]);
  and (_25343_, _25341_, \oc8051_golden_model_1.PC [1]);
  nor (_25344_, _25343_, _25342_);
  and (_25345_, _25344_, _06782_);
  and (_25346_, _06781_, _06043_);
  nor (_25347_, _25346_, _25345_);
  and (_25348_, _25347_, _07504_);
  nor (_25349_, _25348_, _10754_);
  not (_25350_, _25349_);
  nor (_25352_, _25350_, _25338_);
  nor (_25353_, _25352_, _25337_);
  not (_25354_, _25335_);
  nor (_25355_, _25354_, _25353_);
  or (_25356_, _25355_, _10768_);
  nor (_25357_, _25356_, _25336_);
  nor (_25358_, _06043_, _06015_);
  nor (_25359_, _25358_, _12387_);
  not (_25360_, _25359_);
  nor (_25361_, _25360_, _25357_);
  or (_25363_, _12393_, \oc8051_golden_model_1.PC [1]);
  and (_25364_, _12389_, _12391_);
  and (_25365_, _08554_, _08553_);
  nand (_25366_, _25365_, _25364_);
  nor (_25367_, _12460_, _12458_);
  nor (_25368_, _25367_, _12461_);
  nand (_25369_, _25368_, _25366_);
  and (_25370_, _25369_, _12387_);
  and (_25371_, _25370_, _25363_);
  or (_25372_, _25371_, _25361_);
  nand (_25374_, _25372_, _07155_);
  and (_25375_, _07154_, _06043_);
  nor (_25376_, _25375_, _06341_);
  nand (_25377_, _25376_, _25374_);
  or (_25378_, _25327_, _12536_);
  or (_25379_, _12534_, _06043_);
  and (_25380_, _25379_, _06341_);
  nand (_25381_, _25380_, _25378_);
  and (_25382_, _25381_, _12541_);
  nand (_25383_, _25382_, _25377_);
  nor (_25385_, _12541_, _06111_);
  nor (_25386_, _25385_, _06272_);
  nand (_25387_, _25386_, _25383_);
  and (_25388_, _06272_, _05597_);
  nor (_25389_, _25388_, _07611_);
  nand (_25390_, _25389_, _25387_);
  and (_25391_, _07038_, _07611_);
  nor (_25392_, _25391_, _06461_);
  nand (_25393_, _25392_, _25390_);
  and (_25394_, _06461_, _05597_);
  nor (_25396_, _25394_, _12551_);
  nand (_25397_, _25396_, _25393_);
  nor (_25398_, _12550_, _06111_);
  nor (_25399_, _25398_, _06464_);
  nand (_25400_, _25399_, _25397_);
  not (_25401_, _12560_);
  and (_25402_, _06464_, _05597_);
  nor (_25403_, _25402_, _25401_);
  and (_25404_, _25403_, _25400_);
  or (_25405_, _25404_, _25334_);
  nand (_25407_, _25405_, _06269_);
  and (_25408_, _06268_, \oc8051_golden_model_1.PC [1]);
  nor (_25409_, _25408_, _12563_);
  and (_25410_, _25409_, _25407_);
  nor (_25411_, _07038_, _06013_);
  or (_25412_, _25411_, _25410_);
  nand (_25413_, _25412_, _07303_);
  and (_25414_, _06267_, _05597_);
  nor (_25415_, _25414_, _12379_);
  and (_25416_, _25415_, _25413_);
  or (_25418_, _25416_, _25333_);
  nand (_25419_, _25418_, _12177_);
  or (_25420_, _25330_, _12333_);
  or (_25421_, _12335_, _06111_);
  and (_25422_, _25421_, _06347_);
  nand (_25423_, _25422_, _25420_);
  and (_25424_, _25423_, _06774_);
  nand (_25425_, _25424_, _25419_);
  and (_25426_, _12587_, _06111_);
  nor (_25427_, _25327_, _12587_);
  or (_25429_, _25427_, _06774_);
  or (_25430_, _25429_, _25426_);
  nand (_25431_, _25430_, _25425_);
  nand (_25432_, _25431_, _12176_);
  and (_25433_, _12604_, _06043_);
  nor (_25434_, _25330_, _12604_);
  or (_25435_, _25434_, _25433_);
  and (_25436_, _25435_, _06371_);
  nor (_25437_, _25436_, _12174_);
  and (_25438_, _25437_, _25432_);
  or (_25440_, _25438_, _25324_);
  nand (_25441_, _25440_, _06262_);
  and (_25442_, _06261_, \oc8051_golden_model_1.PC [1]);
  nor (_25443_, _25442_, _12613_);
  nand (_25444_, _25443_, _25441_);
  not (_25445_, _25322_);
  nor (_25446_, _07038_, _06007_);
  nor (_25447_, _25446_, _25445_);
  and (_25448_, _25447_, _25444_);
  or (_25449_, _25448_, _25323_);
  nand (_25451_, _25449_, _12630_);
  nor (_25452_, _12630_, _06111_);
  nor (_25453_, _25452_, _06505_);
  nand (_25454_, _25453_, _25451_);
  and (_25455_, _06505_, _05597_);
  nor (_25456_, _25455_, _25158_);
  nand (_25457_, _25456_, _25454_);
  and (_25458_, _07038_, _25158_);
  nor (_25459_, _25458_, _06504_);
  nand (_25460_, _25459_, _25457_);
  not (_25462_, _17307_);
  and (_25463_, _10588_, _14204_);
  and (_25464_, _06504_, _05597_);
  not (_25465_, _25464_);
  and (_25466_, _25465_, _17311_);
  and (_25467_, _25466_, _25463_);
  and (_25468_, _25467_, _25462_);
  and (_25469_, _25468_, _25460_);
  or (_25470_, _25469_, _25320_);
  nand (_25471_, _25470_, _12643_);
  nor (_25473_, _12643_, _05597_);
  nor (_25474_, _25473_, _10515_);
  nand (_25475_, _25474_, _25471_);
  nor (_25476_, _06043_, _05984_);
  nor (_25477_, _25476_, _06257_);
  and (_25478_, _25477_, _25475_);
  and (_25479_, _06257_, \oc8051_golden_model_1.PC [1]);
  or (_25480_, _25479_, _25478_);
  nand (_25481_, _25480_, _05978_);
  and (_25482_, _07038_, _06254_);
  nor (_25484_, _25482_, _06373_);
  nand (_25485_, _25484_, _25481_);
  and (_25486_, _06373_, _06043_);
  nor (_25487_, _25486_, _12659_);
  nand (_25488_, _25487_, _25485_);
  nor (_25489_, _07216_, _05597_);
  nor (_25490_, _25489_, _10094_);
  nand (_25491_, _25490_, _25488_);
  not (_25492_, _12172_);
  nor (_25493_, _06111_, _05982_);
  nor (_25495_, _25493_, _25492_);
  nand (_25496_, _25495_, _25491_);
  nor (_25497_, _12172_, _06111_);
  nor (_25498_, _25497_, _06323_);
  nand (_25499_, _25498_, _25496_);
  and (_25500_, _06323_, _05597_);
  nor (_25501_, _25500_, _12668_);
  nand (_25502_, _25501_, _25499_);
  and (_25503_, _07038_, _12668_);
  nor (_25504_, _25503_, _12674_);
  nand (_25506_, _25504_, _25502_);
  and (_25507_, _25368_, _12674_);
  nor (_25508_, _25507_, _09031_);
  and (_25509_, _25508_, _25506_);
  or (_25510_, _25509_, _25319_);
  nand (_25511_, _25510_, _06219_);
  and (_25512_, _06218_, _06111_);
  nor (_25513_, _25512_, _10929_);
  nand (_25514_, _25513_, _25511_);
  and (_25515_, _10929_, _05597_);
  nor (_25517_, _25515_, _12690_);
  nand (_25518_, _25517_, _25514_);
  and (_25519_, _12690_, _06109_);
  nor (_25520_, _25519_, _06322_);
  nand (_25521_, _25520_, _25518_);
  and (_25522_, _06322_, _05597_);
  nor (_25523_, _25522_, _06217_);
  nand (_25524_, _25523_, _25521_);
  and (_25525_, _07038_, _06217_);
  nor (_25526_, _25525_, _12733_);
  nand (_25528_, _25526_, _25524_);
  and (_25529_, _11342_, _05597_);
  and (_25530_, _25368_, _12759_);
  or (_25531_, _25530_, _25529_);
  and (_25532_, _25531_, _12733_);
  nor (_25533_, _25532_, _12737_);
  and (_25534_, _25533_, _25528_);
  or (_25535_, _25534_, _25318_);
  nand (_25536_, _25535_, _12166_);
  nor (_25537_, _12166_, _05597_);
  nor (_25539_, _25537_, _06369_);
  nand (_25540_, _25539_, _25536_);
  and (_25541_, _06369_, _06043_);
  nor (_25542_, _25541_, _06536_);
  and (_25543_, _25542_, _25540_);
  and (_25544_, _06536_, \oc8051_golden_model_1.PC [1]);
  or (_25545_, _25544_, _25543_);
  nand (_25546_, _25545_, _05955_);
  and (_25547_, _07038_, _12750_);
  nor (_25548_, _25547_, _12755_);
  nand (_25550_, _25548_, _25546_);
  nor (_25551_, _25368_, _12759_);
  nor (_25552_, _11342_, _05597_);
  nor (_25553_, _25552_, _25061_);
  not (_25554_, _25553_);
  nor (_25555_, _25554_, _25551_);
  nor (_25556_, _25555_, _10980_);
  and (_25557_, _25556_, _25550_);
  or (_25558_, _25557_, _25317_);
  nand (_25559_, _25558_, _12164_);
  nor (_25561_, _12164_, _05597_);
  nor (_25562_, _25561_, _06375_);
  nand (_25563_, _25562_, _25559_);
  and (_25564_, _06375_, _06043_);
  nor (_25565_, _25564_, _06545_);
  and (_25566_, _25565_, _25563_);
  and (_25567_, _06545_, \oc8051_golden_model_1.PC [1]);
  or (_25568_, _25567_, _25566_);
  nand (_25569_, _25568_, _05961_);
  and (_25570_, _07038_, _07233_);
  nor (_25572_, _25570_, _12776_);
  nand (_25573_, _25572_, _25569_);
  nor (_25574_, _25368_, \oc8051_golden_model_1.PSW [7]);
  and (_25575_, \oc8051_golden_model_1.PSW [7], \oc8051_golden_model_1.PC [1]);
  nor (_25576_, _25575_, _12782_);
  not (_25577_, _25576_);
  nor (_25578_, _25577_, _25574_);
  nor (_25579_, _25578_, _17507_);
  and (_25580_, _25579_, _25573_);
  nor (_25581_, _25580_, _25316_);
  or (_25583_, _25581_, _12160_);
  and (_25584_, _12160_, _06043_);
  nor (_25585_, _25584_, _11011_);
  nand (_25586_, _25585_, _25583_);
  and (_25587_, _11011_, _06111_);
  nor (_25588_, _25587_, _11023_);
  nand (_25589_, _25588_, _25586_);
  nor (_25590_, _11022_, _05597_);
  nor (_25591_, _25590_, _06366_);
  nand (_25592_, _25591_, _25589_);
  and (_25594_, _06366_, _06043_);
  nor (_25595_, _25594_, _06528_);
  and (_25596_, _25595_, _25592_);
  and (_25597_, _06528_, \oc8051_golden_model_1.PC [1]);
  or (_25598_, _25597_, _25596_);
  nand (_25599_, _25598_, _05966_);
  and (_25600_, _07038_, _12795_);
  nor (_25601_, _25600_, _12800_);
  nand (_25602_, _25601_, _25599_);
  nor (_25603_, \oc8051_golden_model_1.PSW [7], \oc8051_golden_model_1.PC [1]);
  and (_25605_, _25368_, \oc8051_golden_model_1.PSW [7]);
  or (_25606_, _25605_, _25603_);
  and (_25607_, _25606_, _12800_);
  nor (_25608_, _25607_, _12804_);
  and (_25609_, _25608_, _25602_);
  or (_25610_, _25609_, _25315_);
  nand (_25611_, _25610_, _12153_);
  nor (_25612_, _12153_, _05597_);
  nor (_25613_, _25612_, _11125_);
  nand (_25614_, _25613_, _25611_);
  and (_25616_, _11125_, _06111_);
  nor (_25617_, _25616_, _06551_);
  and (_25618_, _25617_, _25614_);
  and (_25619_, _09347_, _06551_);
  or (_25620_, _25619_, _25618_);
  nand (_25621_, _25620_, _05959_);
  and (_25622_, _07038_, _07253_);
  nor (_25623_, _25622_, _06365_);
  nand (_25624_, _25623_, _25621_);
  not (_25625_, _12151_);
  and (_25626_, _25330_, _13004_);
  not (_25627_, _25626_);
  nor (_25628_, _13004_, _06043_);
  nor (_25629_, _25628_, _06558_);
  and (_25630_, _25629_, _25627_);
  nor (_25631_, _25630_, _25625_);
  and (_25632_, _25631_, _25624_);
  or (_25633_, _25632_, _25314_);
  nand (_25634_, _25633_, _13012_);
  nor (_25635_, _13012_, _05597_);
  nor (_25638_, _25635_, _11284_);
  nand (_25639_, _25638_, _25634_);
  and (_25640_, _11284_, _06111_);
  nor (_25641_, _25640_, _06281_);
  and (_25642_, _25641_, _25639_);
  and (_25643_, _09347_, _06281_);
  or (_25644_, _25643_, _25642_);
  nand (_25645_, _25644_, _05964_);
  not (_25646_, _05964_);
  and (_25647_, _07038_, _25646_);
  nor (_25649_, _25647_, _06362_);
  nand (_25650_, _25649_, _25645_);
  and (_25651_, _13004_, _06111_);
  nor (_25652_, _25327_, _13004_);
  nor (_25653_, _25652_, _25651_);
  and (_25654_, _25653_, _06362_);
  nor (_25655_, _25654_, _15693_);
  and (_25656_, _25655_, _25650_);
  nor (_25657_, _25656_, _25313_);
  nor (_25658_, _07482_, _06567_);
  or (_25660_, _25658_, _25657_);
  and (_25661_, _25658_, _06043_);
  nor (_25662_, _25661_, _06568_);
  nand (_25663_, _25662_, _25660_);
  and (_25664_, _06568_, _05597_);
  nor (_25665_, _25664_, _13038_);
  and (_25666_, _25665_, _25663_);
  or (_25667_, _25666_, _25312_);
  nand (_25668_, _25667_, _07271_);
  and (_25669_, _07695_, _07038_);
  nor (_25671_, _25669_, _05927_);
  nand (_25672_, _25671_, _25668_);
  and (_25673_, _25653_, _05927_);
  nor (_25674_, _25673_, _15111_);
  nand (_25675_, _25674_, _25672_);
  nor (_25676_, _15107_, _06111_);
  nor (_25677_, _25676_, _15115_);
  nand (_25678_, _25677_, _25675_);
  and (_25679_, _15115_, _06111_);
  nor (_25680_, _25679_, _07281_);
  nand (_25682_, _25680_, _25678_);
  and (_25683_, _07281_, _06043_);
  nor (_25684_, _25683_, _06278_);
  and (_25685_, _25684_, _25682_);
  or (_25686_, _25685_, _25311_);
  nand (_25687_, _25686_, _12141_);
  nor (_25688_, _12141_, _06043_);
  nor (_25689_, _25688_, _25301_);
  nand (_25690_, _25689_, _25687_);
  and (_25691_, _25301_, _07038_);
  nor (_25693_, _25691_, _13068_);
  and (_25694_, _25693_, _25690_);
  and (_25695_, _13068_, _06111_);
  or (_25696_, _25695_, _25694_);
  or (_25697_, _25696_, _01351_);
  or (_25698_, _01347_, \oc8051_golden_model_1.PC [1]);
  and (_25699_, _25698_, _42618_);
  and (_43246_, _25699_, _25697_);
  and (_25700_, _13068_, _06040_);
  and (_25701_, _06278_, _06079_);
  and (_25703_, _06568_, _06079_);
  nor (_25704_, _12151_, _06040_);
  nor (_25705_, _12154_, _06040_);
  nor (_25706_, _12162_, _06040_);
  nor (_25707_, _10979_, _06040_);
  nor (_25708_, _12169_, _06040_);
  and (_25709_, _06332_, _06321_);
  nor (_25710_, _06699_, _05951_);
  nand (_25711_, _25710_, _06079_);
  and (_25712_, _07214_, _06085_);
  nor (_25714_, _25322_, _06079_);
  and (_25715_, _12174_, _06074_);
  and (_25716_, _12258_, _12255_);
  nor (_25717_, _25716_, _12259_);
  not (_25718_, _25717_);
  and (_25719_, _25718_, _12335_);
  and (_25720_, _12333_, _12248_);
  or (_25721_, _25720_, _25719_);
  and (_25722_, _25721_, _06347_);
  or (_25723_, _12393_, _06085_);
  and (_25725_, _12465_, _12462_);
  nor (_25726_, _25725_, _12466_);
  nand (_25727_, _25726_, _12393_);
  and (_25728_, _25727_, _12387_);
  and (_25729_, _25728_, _25723_);
  or (_25730_, _07504_, _06697_);
  nor (_25731_, _07486_, \oc8051_golden_model_1.PC [2]);
  or (_25732_, _25731_, _07141_);
  nand (_25733_, _07141_, _06079_);
  and (_25734_, _25733_, _06782_);
  and (_25736_, _25734_, _25732_);
  nor (_25737_, _12513_, _06040_);
  or (_25738_, _25737_, _06758_);
  or (_25739_, _25738_, _25736_);
  and (_25740_, _25739_, _12512_);
  and (_25741_, _25740_, _25730_);
  nor (_25742_, _12512_, _06040_);
  or (_25743_, _25742_, _25741_);
  and (_25744_, _25743_, _08654_);
  or (_25745_, _25744_, _25729_);
  and (_25747_, _25745_, _07155_);
  and (_25748_, _07154_, _06074_);
  or (_25749_, _25748_, _06341_);
  or (_25750_, _25749_, _25747_);
  and (_25751_, _25718_, _12534_);
  and (_25752_, _12536_, _12248_);
  or (_25753_, _25752_, _07151_);
  or (_25754_, _25753_, _25751_);
  and (_25755_, _25754_, _12541_);
  and (_25756_, _25755_, _25750_);
  nor (_25758_, _12541_, _06040_);
  or (_25759_, _25758_, _06272_);
  or (_25760_, _25759_, _25756_);
  nand (_25761_, _06272_, _06079_);
  and (_25762_, _25761_, _06010_);
  and (_25763_, _25762_, _25760_);
  and (_25764_, _06697_, _07611_);
  or (_25765_, _25764_, _06461_);
  or (_25766_, _25765_, _25763_);
  nand (_25767_, _06461_, _06079_);
  and (_25769_, _25767_, _12550_);
  and (_25770_, _25769_, _25766_);
  nor (_25771_, _12550_, _06040_);
  or (_25772_, _25771_, _06464_);
  or (_25773_, _25772_, _25770_);
  nand (_25774_, _06464_, _06079_);
  and (_25775_, _25774_, _12560_);
  and (_25776_, _25775_, _25773_);
  nor (_25777_, _12560_, _06040_);
  or (_25778_, _25777_, _06268_);
  or (_25780_, _25778_, _25776_);
  nand (_25781_, _06268_, _06079_);
  and (_25782_, _25781_, _06013_);
  and (_25783_, _25782_, _25780_);
  and (_25784_, _06697_, _12563_);
  or (_25785_, _25784_, _06267_);
  or (_25786_, _25785_, _25783_);
  nand (_25787_, _06267_, _06079_);
  and (_25788_, _25787_, _12378_);
  and (_25789_, _25788_, _25786_);
  nand (_25791_, _12371_, _12247_);
  or (_25792_, _25718_, _12371_);
  and (_25793_, _25792_, _12379_);
  and (_25794_, _25793_, _25791_);
  or (_25795_, _25794_, _25789_);
  and (_25796_, _25795_, _12177_);
  or (_25797_, _25796_, _25722_);
  and (_25798_, _25797_, _06774_);
  or (_25799_, _25718_, _12587_);
  nand (_25800_, _12587_, _12247_);
  and (_25802_, _25800_, _06480_);
  and (_25803_, _25802_, _25799_);
  or (_25804_, _25803_, _06371_);
  or (_25805_, _25804_, _25798_);
  nor (_25806_, _25717_, _12604_);
  and (_25807_, _12604_, _12248_);
  or (_25808_, _25807_, _12176_);
  or (_25809_, _25808_, _25806_);
  and (_25810_, _25809_, _12175_);
  and (_25811_, _25810_, _25805_);
  or (_25813_, _25811_, _25715_);
  and (_25814_, _25813_, _06262_);
  and (_25815_, _06261_, _06085_);
  or (_25816_, _25815_, _12613_);
  or (_25817_, _25816_, _25814_);
  or (_25818_, _06697_, _06007_);
  and (_25819_, _25818_, _25322_);
  and (_25820_, _25819_, _25817_);
  or (_25821_, _25820_, _25714_);
  and (_25822_, _25821_, _12630_);
  nor (_25824_, _12630_, _06040_);
  or (_25825_, _25824_, _06505_);
  or (_25826_, _25825_, _25822_);
  nand (_25827_, _06505_, _06079_);
  and (_25828_, _25827_, _06020_);
  and (_25829_, _25828_, _25826_);
  and (_25830_, _06697_, _25158_);
  or (_25831_, _25830_, _06504_);
  or (_25832_, _25831_, _25829_);
  nand (_25833_, _06504_, _06079_);
  and (_25835_, _25833_, _12639_);
  and (_25836_, _25835_, _25832_);
  nor (_25837_, _12639_, _06040_);
  or (_25838_, _25837_, _25836_);
  and (_25839_, _25838_, _12643_);
  nor (_25840_, _12643_, _06079_);
  or (_25841_, _25840_, _10515_);
  or (_25842_, _25841_, _25839_);
  or (_25843_, _06074_, _05984_);
  and (_25844_, _25843_, _06258_);
  and (_25846_, _25844_, _25842_);
  and (_25847_, _06257_, _06085_);
  or (_25848_, _25847_, _25846_);
  and (_25849_, _25848_, _05978_);
  and (_25850_, _06697_, _06254_);
  or (_25851_, _25850_, _06373_);
  or (_25852_, _25851_, _25849_);
  nor (_25853_, _07461_, _06759_);
  nand (_25854_, _12247_, _06373_);
  nand (_25855_, _25854_, _25853_);
  nor (_25857_, _25855_, _07455_);
  and (_25858_, _25857_, _25852_);
  nor (_25859_, _25858_, _25712_);
  nor (_25860_, _07482_, _05945_);
  nor (_25861_, _25860_, _25859_);
  and (_25862_, _25860_, _06085_);
  or (_25863_, _25862_, _10094_);
  or (_25864_, _25863_, _25861_);
  or (_25865_, _12248_, _05982_);
  and (_25866_, _25865_, _12172_);
  and (_25868_, _25866_, _25864_);
  nor (_25869_, _12172_, _06040_);
  or (_25870_, _25869_, _06323_);
  or (_25871_, _25870_, _25868_);
  nand (_25872_, _06323_, _06079_);
  and (_25873_, _25872_, _05946_);
  and (_25874_, _25873_, _25871_);
  and (_25875_, _06697_, _12668_);
  or (_25876_, _25875_, _25874_);
  and (_25877_, _25876_, _12679_);
  nor (_25879_, _25726_, _12679_);
  or (_25880_, _25879_, _25710_);
  or (_25881_, _25880_, _25877_);
  and (_25882_, _25881_, _25711_);
  or (_25883_, _25882_, _25709_);
  nand (_25884_, _25709_, _06079_);
  and (_25885_, _25884_, _09029_);
  and (_25886_, _25885_, _25883_);
  nor (_25887_, _09029_, _06079_);
  or (_25888_, _25887_, _06218_);
  or (_25890_, _25888_, _25886_);
  and (_25891_, _12247_, _06218_);
  nor (_25892_, _25891_, _10929_);
  and (_25893_, _25892_, _25890_);
  and (_25894_, _10929_, _06085_);
  or (_25895_, _25894_, _25893_);
  nand (_25896_, _25895_, _12691_);
  and (_25897_, _12690_, _06071_);
  nor (_25898_, _25897_, _06322_);
  nand (_25899_, _25898_, _25896_);
  and (_25901_, _06322_, _06079_);
  nor (_25902_, _25901_, _06217_);
  nand (_25903_, _25902_, _25899_);
  and (_25904_, _06697_, _06217_);
  nor (_25905_, _25904_, _12733_);
  nand (_25906_, _25905_, _25903_);
  nor (_25907_, _25726_, _11342_);
  and (_25908_, _11342_, _06085_);
  nor (_25909_, _25908_, _25064_);
  not (_25910_, _25909_);
  nor (_25912_, _25910_, _25907_);
  nor (_25913_, _25912_, _12737_);
  and (_25914_, _25913_, _25906_);
  or (_25915_, _25914_, _25708_);
  nand (_25916_, _25915_, _12166_);
  nor (_25917_, _12166_, _06079_);
  nor (_25918_, _25917_, _06369_);
  nand (_25919_, _25918_, _25916_);
  and (_25920_, _12247_, _06369_);
  nor (_25921_, _25920_, _06536_);
  and (_25923_, _25921_, _25919_);
  and (_25924_, _06536_, _06085_);
  or (_25925_, _25924_, _25923_);
  nand (_25926_, _25925_, _05955_);
  and (_25927_, _06697_, _12750_);
  nor (_25928_, _25927_, _12755_);
  nand (_25929_, _25928_, _25926_);
  nor (_25930_, _11342_, _06085_);
  and (_25931_, _25726_, _11342_);
  or (_25932_, _25931_, _25930_);
  and (_25934_, _25932_, _12755_);
  nor (_25935_, _25934_, _10980_);
  and (_25936_, _25935_, _25929_);
  or (_25937_, _25936_, _25707_);
  nand (_25938_, _25937_, _12164_);
  nor (_25939_, _12164_, _06079_);
  nor (_25940_, _25939_, _06375_);
  nand (_25941_, _25940_, _25938_);
  and (_25942_, _12247_, _06375_);
  nor (_25943_, _25942_, _06545_);
  and (_25945_, _25943_, _25941_);
  and (_25946_, _06545_, _06085_);
  or (_25947_, _25946_, _25945_);
  nand (_25948_, _25947_, _05961_);
  and (_25949_, _06697_, _07233_);
  nor (_25950_, _25949_, _12776_);
  nand (_25951_, _25950_, _25948_);
  nor (_25952_, _25726_, \oc8051_golden_model_1.PSW [7]);
  nor (_25953_, _06079_, _10558_);
  nor (_25954_, _25953_, _12782_);
  not (_25955_, _25954_);
  nor (_25956_, _25955_, _25952_);
  nor (_25957_, _25956_, _12780_);
  and (_25958_, _25957_, _25951_);
  or (_25959_, _25958_, _25706_);
  nand (_25960_, _25959_, _11022_);
  nor (_25961_, _11022_, _06079_);
  nor (_25962_, _25961_, _06366_);
  nand (_25963_, _25962_, _25960_);
  and (_25964_, _12247_, _06366_);
  nor (_25967_, _25964_, _06528_);
  and (_25968_, _25967_, _25963_);
  and (_25969_, _06528_, _06085_);
  or (_25970_, _25969_, _25968_);
  nand (_25971_, _25970_, _05966_);
  and (_25972_, _06697_, _12795_);
  nor (_25973_, _25972_, _12800_);
  nand (_25974_, _25973_, _25971_);
  nor (_25975_, _25726_, _10558_);
  nor (_25976_, _06079_, \oc8051_golden_model_1.PSW [7]);
  nor (_25978_, _25976_, _25056_);
  not (_25979_, _25978_);
  nor (_25980_, _25979_, _25975_);
  nor (_25981_, _25980_, _12804_);
  and (_25982_, _25981_, _25974_);
  or (_25983_, _25982_, _25705_);
  nand (_25984_, _25983_, _12153_);
  nor (_25985_, _12153_, _06079_);
  nor (_25986_, _25985_, _11125_);
  nand (_25987_, _25986_, _25984_);
  and (_25989_, _11125_, _06040_);
  nor (_25990_, _25989_, _06551_);
  and (_25991_, _25990_, _25987_);
  and (_25992_, _09302_, _06551_);
  or (_25993_, _25992_, _25991_);
  nand (_25994_, _25993_, _05959_);
  and (_25995_, _06697_, _07253_);
  nor (_25996_, _25995_, _06365_);
  nand (_25997_, _25996_, _25994_);
  nor (_25998_, _12247_, _13004_);
  and (_26000_, _25718_, _13004_);
  or (_26001_, _26000_, _06558_);
  or (_26002_, _26001_, _25998_);
  and (_26003_, _26002_, _12151_);
  and (_26004_, _26003_, _25997_);
  or (_26005_, _26004_, _25704_);
  nand (_26006_, _26005_, _13012_);
  nor (_26007_, _13012_, _06079_);
  nor (_26008_, _26007_, _11284_);
  nand (_26009_, _26008_, _26006_);
  and (_26011_, _11284_, _06040_);
  nor (_26012_, _26011_, _06281_);
  and (_26013_, _26012_, _26009_);
  and (_26014_, _09302_, _06281_);
  or (_26015_, _26014_, _26013_);
  nand (_26016_, _26015_, _05964_);
  and (_26017_, _06697_, _25646_);
  nor (_26018_, _26017_, _06362_);
  nand (_26019_, _26018_, _26016_);
  nor (_26020_, _25717_, _13004_);
  and (_26022_, _12248_, _13004_);
  nor (_26023_, _26022_, _26020_);
  and (_26024_, _26023_, _06362_);
  nor (_26025_, _26024_, _13031_);
  nand (_26026_, _26025_, _26019_);
  nor (_26027_, _13030_, _06040_);
  nor (_26028_, _26027_, _06568_);
  and (_26029_, _26028_, _26026_);
  or (_26030_, _26029_, _25703_);
  nand (_26031_, _26030_, _13037_);
  nor (_26033_, _13037_, _06074_);
  nor (_26034_, _26033_, _07695_);
  nand (_26035_, _26034_, _26031_);
  and (_26036_, _07695_, _06697_);
  nor (_26037_, _26036_, _05927_);
  nand (_26038_, _26037_, _26035_);
  and (_26039_, _26023_, _05927_);
  nor (_26040_, _26039_, _13053_);
  nand (_26041_, _26040_, _26038_);
  nor (_26042_, _13052_, _06040_);
  nor (_26044_, _26042_, _06278_);
  and (_26045_, _26044_, _26041_);
  or (_26046_, _26045_, _25701_);
  nand (_26047_, _26046_, _12141_);
  nor (_26048_, _12141_, _06074_);
  nor (_26049_, _26048_, _25301_);
  nand (_26050_, _26049_, _26047_);
  and (_26051_, _25301_, _06697_);
  nor (_26052_, _26051_, _13068_);
  and (_26053_, _26052_, _26050_);
  or (_26055_, _26053_, _25700_);
  or (_26056_, _26055_, _01351_);
  or (_26057_, _01347_, \oc8051_golden_model_1.PC [2]);
  and (_26058_, _26057_, _42618_);
  and (_43247_, _26058_, _26056_);
  and (_26059_, _13068_, _06028_);
  and (_26060_, _06278_, _05932_);
  and (_26061_, _06568_, _05932_);
  nor (_26062_, _12151_, _06028_);
  nor (_26063_, _12154_, _06028_);
  nor (_26065_, _12162_, _06028_);
  nor (_26066_, _10979_, _06028_);
  nor (_26067_, _12169_, _06028_);
  nor (_26068_, _09030_, _05932_);
  nor (_26069_, _25322_, _05932_);
  and (_26070_, _12174_, _06027_);
  or (_26071_, _12534_, _12242_);
  or (_26072_, _12245_, _12244_);
  and (_26073_, _26072_, _12260_);
  nor (_26074_, _26072_, _12260_);
  nor (_26076_, _26074_, _26073_);
  or (_26077_, _26076_, _12536_);
  and (_26078_, _26077_, _26071_);
  or (_26079_, _26078_, _07151_);
  and (_26080_, _12507_, _05932_);
  or (_26081_, _12455_, _12454_);
  and (_26082_, _26081_, _12467_);
  nor (_26083_, _26081_, _12467_);
  nor (_26084_, _26083_, _26082_);
  and (_26085_, _26084_, _12393_);
  nor (_26087_, _26085_, _26080_);
  nand (_26088_, _26087_, _12387_);
  nor (_26089_, _12512_, _06028_);
  nor (_26090_, _07486_, \oc8051_golden_model_1.PC [3]);
  nor (_26091_, _26090_, _07141_);
  and (_26092_, _07141_, _05932_);
  nor (_26093_, _26092_, _06781_);
  not (_26094_, _26093_);
  nor (_26095_, _26094_, _26091_);
  not (_26096_, _26095_);
  nor (_26098_, _12513_, _06028_);
  nor (_26099_, _26098_, _06758_);
  and (_26100_, _26099_, _26096_);
  nor (_26101_, _07504_, _06452_);
  or (_26102_, _26101_, _12516_);
  nor (_26103_, _26102_, _26100_);
  nor (_26104_, _26103_, _26089_);
  nor (_26105_, _26104_, _12387_);
  nor (_26106_, _26105_, _07154_);
  and (_26107_, _26106_, _26088_);
  and (_26109_, _07154_, _06028_);
  or (_26110_, _26109_, _06341_);
  or (_26111_, _26110_, _26107_);
  nand (_26112_, _26111_, _26079_);
  nand (_26113_, _26112_, _12541_);
  nor (_26114_, _12541_, _06028_);
  nor (_26115_, _26114_, _06272_);
  nand (_26116_, _26115_, _26113_);
  and (_26117_, _06272_, _05932_);
  nor (_26118_, _26117_, _07611_);
  nand (_26120_, _26118_, _26116_);
  and (_26121_, _06452_, _07611_);
  nor (_26122_, _26121_, _06461_);
  nand (_26123_, _26122_, _26120_);
  and (_26124_, _06461_, _05932_);
  nor (_26125_, _26124_, _12551_);
  nand (_26126_, _26125_, _26123_);
  nor (_26127_, _12550_, _06028_);
  nor (_26128_, _26127_, _06464_);
  nand (_26129_, _26128_, _26126_);
  and (_26131_, _06464_, _05932_);
  nor (_26132_, _26131_, _25401_);
  nand (_26133_, _26132_, _26129_);
  nor (_26134_, _12560_, _06028_);
  nor (_26135_, _26134_, _06268_);
  nand (_26136_, _26135_, _26133_);
  and (_26137_, _06268_, _05932_);
  nor (_26138_, _26137_, _12563_);
  nand (_26139_, _26138_, _26136_);
  and (_26140_, _06452_, _12563_);
  nor (_26142_, _26140_, _06267_);
  nand (_26143_, _26142_, _26139_);
  and (_26144_, _06267_, _05932_);
  nor (_26145_, _26144_, _12379_);
  nand (_26146_, _26145_, _26143_);
  and (_26147_, _12371_, _12242_);
  not (_26148_, _26076_);
  nor (_26149_, _26148_, _12371_);
  or (_26150_, _26149_, _12378_);
  nor (_26151_, _26150_, _26147_);
  nor (_26153_, _26151_, _06347_);
  nand (_26154_, _26153_, _26146_);
  or (_26155_, _26148_, _12333_);
  or (_26156_, _12335_, _12243_);
  nand (_26157_, _26156_, _26155_);
  nand (_26158_, _26157_, _06347_);
  and (_26159_, _26158_, _06774_);
  nand (_26160_, _26159_, _26154_);
  and (_26161_, _12587_, _12242_);
  not (_26162_, _26161_);
  nor (_26164_, _26148_, _12587_);
  nor (_26165_, _26164_, _06774_);
  and (_26166_, _26165_, _26162_);
  nor (_26167_, _26166_, _06371_);
  nand (_26168_, _26167_, _26160_);
  and (_26169_, _12604_, _12243_);
  nor (_26170_, _26076_, _12604_);
  or (_26171_, _26170_, _12176_);
  nor (_26172_, _26171_, _26169_);
  nor (_26173_, _26172_, _12174_);
  and (_26175_, _26173_, _26168_);
  or (_26176_, _26175_, _26070_);
  nand (_26177_, _26176_, _06262_);
  and (_26178_, _06261_, _06033_);
  nor (_26179_, _26178_, _12613_);
  nand (_26180_, _26179_, _26177_);
  nor (_26181_, _06452_, _06007_);
  nor (_26182_, _26181_, _25445_);
  and (_26183_, _26182_, _26180_);
  or (_26184_, _26183_, _26069_);
  nand (_26186_, _26184_, _12630_);
  nor (_26187_, _12630_, _06028_);
  nor (_26188_, _26187_, _06505_);
  nand (_26189_, _26188_, _26186_);
  and (_26190_, _06505_, _05932_);
  nor (_26191_, _26190_, _25158_);
  nand (_26192_, _26191_, _26189_);
  and (_26193_, _06452_, _25158_);
  nor (_26194_, _26193_, _06504_);
  nand (_26195_, _26194_, _26192_);
  not (_26197_, _12639_);
  and (_26198_, _06504_, _05932_);
  nor (_26199_, _26198_, _26197_);
  and (_26200_, _26199_, _26195_);
  nor (_26201_, _12639_, _06028_);
  or (_26202_, _26201_, _26200_);
  nand (_26203_, _26202_, _12643_);
  nor (_26204_, _12643_, _05932_);
  nor (_26205_, _26204_, _10515_);
  nand (_26206_, _26205_, _26203_);
  nor (_26208_, _05984_, _06027_);
  nor (_26209_, _26208_, _06257_);
  and (_26210_, _26209_, _26206_);
  and (_26211_, _06257_, _06033_);
  or (_26212_, _26211_, _26210_);
  nand (_26213_, _26212_, _05978_);
  and (_26214_, _06452_, _06254_);
  nor (_26215_, _26214_, _06373_);
  nand (_26216_, _26215_, _26213_);
  and (_26217_, _12242_, _06373_);
  nor (_26219_, _26217_, _12659_);
  nand (_26220_, _26219_, _26216_);
  nor (_26221_, _07216_, _05932_);
  nor (_26222_, _26221_, _10094_);
  nand (_26223_, _26222_, _26220_);
  nor (_26224_, _12243_, _05982_);
  nor (_26225_, _26224_, _25492_);
  nand (_26226_, _26225_, _26223_);
  nor (_26227_, _12172_, _06028_);
  nor (_26228_, _26227_, _06323_);
  nand (_26230_, _26228_, _26226_);
  and (_26231_, _06323_, _05932_);
  nor (_26232_, _26231_, _12668_);
  nand (_26233_, _26232_, _26230_);
  and (_26234_, _06452_, _12668_);
  nor (_26235_, _26234_, _12674_);
  nand (_26236_, _26235_, _26233_);
  and (_26237_, _26084_, _12674_);
  nor (_26238_, _26237_, _09031_);
  and (_26239_, _26238_, _26236_);
  or (_26241_, _26239_, _26068_);
  nand (_26242_, _26241_, _06219_);
  and (_26243_, _12243_, _06218_);
  nor (_26244_, _26243_, _10929_);
  nand (_26245_, _26244_, _26242_);
  and (_26246_, _10929_, _05932_);
  nor (_26247_, _26246_, _12690_);
  nand (_26248_, _26247_, _26245_);
  and (_26249_, _12690_, _06004_);
  nor (_26250_, _26249_, _06322_);
  and (_26252_, _26250_, _26248_);
  and (_26253_, _06322_, _05932_);
  or (_26254_, _26253_, _06217_);
  or (_26255_, _26254_, _26252_);
  and (_26256_, _06452_, _06217_);
  nor (_26257_, _26256_, _12733_);
  nand (_26258_, _26257_, _26255_);
  and (_26259_, _11342_, _05932_);
  and (_26260_, _26084_, _12759_);
  or (_26261_, _26260_, _26259_);
  and (_26263_, _26261_, _12733_);
  nor (_26264_, _26263_, _12737_);
  and (_26265_, _26264_, _26258_);
  or (_26266_, _26265_, _26067_);
  nand (_26267_, _26266_, _12166_);
  nor (_26268_, _12166_, _05932_);
  nor (_26269_, _26268_, _06369_);
  and (_26270_, _26269_, _26267_);
  and (_26271_, _12242_, _06369_);
  or (_26272_, _26271_, _06536_);
  nor (_26274_, _26272_, _26270_);
  and (_26275_, _06536_, _06033_);
  or (_26276_, _26275_, _26274_);
  nand (_26277_, _26276_, _05955_);
  and (_26278_, _06452_, _12750_);
  nor (_26279_, _26278_, _12755_);
  nand (_26280_, _26279_, _26277_);
  nor (_26281_, _11342_, _06033_);
  and (_26282_, _26084_, _11342_);
  or (_26283_, _26282_, _26281_);
  and (_26285_, _26283_, _12755_);
  nor (_26286_, _26285_, _10980_);
  and (_26287_, _26286_, _26280_);
  or (_26288_, _26287_, _26066_);
  nand (_26289_, _26288_, _12164_);
  nor (_26290_, _12164_, _05932_);
  nor (_26291_, _26290_, _06375_);
  nand (_26292_, _26291_, _26289_);
  and (_26293_, _12242_, _06375_);
  nor (_26294_, _26293_, _06545_);
  and (_26296_, _26294_, _26292_);
  and (_26297_, _06545_, _06033_);
  or (_26298_, _26297_, _26296_);
  nand (_26299_, _26298_, _05961_);
  and (_26300_, _06452_, _07233_);
  nor (_26301_, _26300_, _12776_);
  nand (_26302_, _26301_, _26299_);
  nor (_26303_, _26084_, \oc8051_golden_model_1.PSW [7]);
  nor (_26304_, _05932_, _10558_);
  nor (_26305_, _26304_, _12782_);
  not (_26307_, _26305_);
  nor (_26308_, _26307_, _26303_);
  nor (_26309_, _26308_, _12780_);
  and (_26310_, _26309_, _26302_);
  or (_26311_, _26310_, _26065_);
  nand (_26312_, _26311_, _11022_);
  nor (_26313_, _11022_, _05932_);
  nor (_26314_, _26313_, _06366_);
  and (_26315_, _26314_, _26312_);
  and (_26316_, _12242_, _06366_);
  or (_26318_, _26316_, _06528_);
  nor (_26319_, _26318_, _26315_);
  and (_26320_, _06528_, _06033_);
  or (_26321_, _26320_, _26319_);
  nand (_26322_, _26321_, _05966_);
  and (_26323_, _06452_, _12795_);
  nor (_26324_, _26323_, _12800_);
  nand (_26325_, _26324_, _26322_);
  and (_26326_, _05932_, _10558_);
  and (_26327_, _26084_, \oc8051_golden_model_1.PSW [7]);
  or (_26329_, _26327_, _26326_);
  and (_26330_, _26329_, _12800_);
  nor (_26331_, _26330_, _12804_);
  and (_26332_, _26331_, _26325_);
  or (_26333_, _26332_, _26063_);
  nand (_26334_, _26333_, _12153_);
  nor (_26335_, _12153_, _05932_);
  nor (_26336_, _26335_, _11125_);
  nand (_26337_, _26336_, _26334_);
  and (_26338_, _11125_, _06028_);
  nor (_26340_, _26338_, _06551_);
  and (_26341_, _26340_, _26337_);
  and (_26342_, _09257_, _06551_);
  or (_26343_, _26342_, _26341_);
  nand (_26344_, _26343_, _05959_);
  and (_26345_, _06452_, _07253_);
  nor (_26346_, _26345_, _06365_);
  nand (_26347_, _26346_, _26344_);
  and (_26348_, _26148_, _13004_);
  nor (_26349_, _12242_, _13004_);
  or (_26351_, _26349_, _06558_);
  or (_26352_, _26351_, _26348_);
  and (_26353_, _26352_, _12151_);
  and (_26354_, _26353_, _26347_);
  or (_26355_, _26354_, _26062_);
  nand (_26356_, _26355_, _13012_);
  nor (_26357_, _13012_, _05932_);
  nor (_26358_, _26357_, _11284_);
  nand (_26359_, _26358_, _26356_);
  and (_26360_, _11284_, _06028_);
  nor (_26362_, _26360_, _06281_);
  and (_26363_, _26362_, _26359_);
  and (_26364_, _09257_, _06281_);
  or (_26365_, _26364_, _26363_);
  nand (_26366_, _26365_, _05964_);
  and (_26367_, _06452_, _25646_);
  nor (_26368_, _26367_, _06362_);
  nand (_26369_, _26368_, _26366_);
  nor (_26370_, _26076_, _13004_);
  and (_26371_, _12243_, _13004_);
  nor (_26373_, _26371_, _26370_);
  and (_26374_, _26373_, _06362_);
  nor (_26375_, _26374_, _13031_);
  nand (_26376_, _26375_, _26369_);
  nor (_26377_, _13030_, _06028_);
  nor (_26378_, _26377_, _06568_);
  and (_26379_, _26378_, _26376_);
  or (_26380_, _26379_, _26061_);
  nand (_26381_, _26380_, _13037_);
  nor (_26382_, _13037_, _06027_);
  nor (_26384_, _26382_, _07695_);
  nand (_26385_, _26384_, _26381_);
  and (_26386_, _07695_, _06452_);
  nor (_26387_, _26386_, _05927_);
  nand (_26388_, _26387_, _26385_);
  and (_26389_, _26373_, _05927_);
  nor (_26390_, _26389_, _13053_);
  nand (_26391_, _26390_, _26388_);
  nor (_26392_, _13052_, _06028_);
  nor (_26393_, _26392_, _06278_);
  and (_26395_, _26393_, _26391_);
  or (_26396_, _26395_, _26060_);
  nand (_26397_, _26396_, _12141_);
  nor (_26398_, _12141_, _06027_);
  nor (_26399_, _26398_, _25301_);
  nand (_26400_, _26399_, _26397_);
  and (_26401_, _25301_, _06452_);
  nor (_26402_, _26401_, _13068_);
  and (_26403_, _26402_, _26400_);
  or (_26404_, _26403_, _26059_);
  or (_26406_, _26404_, _01351_);
  or (_26407_, _01347_, \oc8051_golden_model_1.PC [3]);
  and (_26408_, _26407_, _42618_);
  and (_43249_, _26408_, _26406_);
  and (_26409_, _08892_, _07695_);
  and (_26410_, _12451_, _10558_);
  and (_26411_, _12472_, _12469_);
  nor (_26412_, _26411_, _12473_);
  and (_26413_, _26412_, \oc8051_golden_model_1.PSW [7]);
  or (_26414_, _26413_, _26410_);
  and (_26416_, _26414_, _12800_);
  nor (_26417_, _12452_, _11342_);
  and (_26418_, _26412_, _11342_);
  or (_26419_, _26418_, _26417_);
  and (_26420_, _26419_, _12755_);
  and (_26421_, _12451_, _11342_);
  and (_26422_, _26412_, _12759_);
  or (_26423_, _26422_, _26421_);
  and (_26424_, _26423_, _12733_);
  nor (_26425_, _12451_, _09030_);
  and (_26427_, _12452_, _06257_);
  not (_26428_, \oc8051_golden_model_1.PC [4]);
  nor (_26429_, _05616_, _26428_);
  and (_26430_, _05616_, _26428_);
  nor (_26431_, _26430_, _26429_);
  not (_26432_, _26431_);
  and (_26433_, _26432_, _12174_);
  and (_26434_, _12452_, _06268_);
  nor (_26435_, _26431_, _12550_);
  nand (_26436_, _26412_, _25366_);
  or (_26437_, _12393_, _12452_);
  and (_26438_, _26437_, _26436_);
  and (_26439_, _26438_, _12387_);
  nor (_26440_, _26432_, _12512_);
  and (_26441_, _08892_, _06758_);
  or (_26442_, _07486_, _26428_);
  and (_26443_, _26442_, _07142_);
  and (_26444_, _12452_, _07141_);
  or (_26445_, _26444_, _06781_);
  or (_26446_, _26445_, _26443_);
  or (_26448_, _26432_, _12513_);
  and (_26449_, _26448_, _07504_);
  and (_26450_, _26449_, _26446_);
  nor (_26451_, _26450_, _12516_);
  not (_26452_, _26451_);
  nor (_26453_, _26452_, _26441_);
  or (_26454_, _26453_, _12387_);
  nor (_26455_, _26454_, _26440_);
  or (_26456_, _26455_, _26439_);
  nand (_26457_, _26456_, _07155_);
  and (_26459_, _26432_, _07154_);
  nor (_26460_, _26459_, _06341_);
  nand (_26461_, _26460_, _26457_);
  or (_26462_, _12534_, _12238_);
  and (_26463_, _12265_, _12262_);
  nor (_26464_, _26463_, _12266_);
  or (_26465_, _26464_, _12536_);
  and (_26466_, _26465_, _06341_);
  nand (_26467_, _26466_, _26462_);
  and (_26468_, _26467_, _12541_);
  and (_26469_, _26468_, _26461_);
  nor (_26470_, _26431_, _12541_);
  or (_26471_, _26470_, _26469_);
  nand (_26472_, _26471_, _06273_);
  and (_26473_, _12452_, _06272_);
  nor (_26474_, _26473_, _07611_);
  and (_26475_, _26474_, _26472_);
  nor (_26476_, _08892_, _06010_);
  or (_26477_, _26476_, _06461_);
  nor (_26478_, _26477_, _26475_);
  and (_26479_, _12452_, _06461_);
  or (_26480_, _26479_, _26478_);
  and (_26481_, _26480_, _12550_);
  or (_26482_, _26481_, _26435_);
  nand (_26483_, _26482_, _06465_);
  and (_26484_, _12452_, _06464_);
  nor (_26485_, _26484_, _25401_);
  nand (_26486_, _26485_, _26483_);
  nor (_26487_, _26432_, _12560_);
  nor (_26488_, _26487_, _06268_);
  and (_26489_, _26488_, _26486_);
  or (_26490_, _26489_, _26434_);
  nand (_26491_, _26490_, _06013_);
  and (_26492_, _08892_, _12563_);
  nor (_26493_, _26492_, _06267_);
  nand (_26494_, _26493_, _26491_);
  and (_26495_, _12451_, _06267_);
  nor (_26496_, _26495_, _12379_);
  and (_26497_, _26496_, _26494_);
  and (_26498_, _12371_, _12238_);
  not (_26499_, _26464_);
  nor (_26500_, _26499_, _12371_);
  or (_26501_, _26500_, _12378_);
  nor (_26502_, _26501_, _26498_);
  nor (_26503_, _26502_, _26497_);
  or (_26504_, _26503_, _06347_);
  and (_26505_, _26464_, _12335_);
  and (_26506_, _12333_, _12238_);
  or (_26507_, _26506_, _12177_);
  or (_26508_, _26507_, _26505_);
  nand (_26509_, _26508_, _26504_);
  or (_26510_, _26509_, _06480_);
  nor (_26511_, _26499_, _12587_);
  and (_26512_, _12587_, _12238_);
  nor (_26513_, _26512_, _26511_);
  or (_26514_, _26513_, _06774_);
  and (_26515_, _26514_, _26510_);
  or (_26516_, _26515_, _06371_);
  and (_26517_, _12604_, _12238_);
  not (_26518_, _12604_);
  and (_26520_, _26464_, _26518_);
  or (_26521_, _26520_, _26517_);
  and (_26522_, _26521_, _06371_);
  nor (_26523_, _26522_, _12174_);
  and (_26524_, _26523_, _26516_);
  or (_26525_, _26524_, _26433_);
  nand (_26526_, _26525_, _06262_);
  and (_26527_, _12452_, _06261_);
  nor (_26528_, _26527_, _12613_);
  nand (_26529_, _26528_, _26526_);
  nor (_26531_, _08892_, _06007_);
  nor (_26532_, _26531_, _25445_);
  nand (_26533_, _26532_, _26529_);
  nor (_26534_, _25322_, _12451_);
  nor (_26535_, _26534_, _12631_);
  nand (_26536_, _26535_, _26533_);
  nor (_26537_, _26432_, _12630_);
  nor (_26538_, _26537_, _06505_);
  nand (_26539_, _26538_, _26536_);
  and (_26540_, _12452_, _06505_);
  nor (_26541_, _26540_, _25158_);
  and (_26542_, _26541_, _26539_);
  nor (_26543_, _08892_, _06020_);
  or (_26544_, _26543_, _06504_);
  or (_26545_, _26544_, _26542_);
  and (_26546_, _12452_, _06504_);
  nor (_26547_, _26546_, _26197_);
  nand (_26548_, _26547_, _26545_);
  nor (_26549_, _26432_, _12639_);
  nor (_26550_, _26549_, _12644_);
  nand (_26552_, _26550_, _26548_);
  nor (_26553_, _12451_, _12643_);
  nor (_26554_, _26553_, _10515_);
  nand (_26555_, _26554_, _26552_);
  nor (_26556_, _26432_, _05984_);
  nor (_26557_, _26556_, _06257_);
  and (_26558_, _26557_, _26555_);
  or (_26559_, _26558_, _26427_);
  nand (_26560_, _26559_, _05978_);
  and (_26561_, _08892_, _06254_);
  nor (_26563_, _26561_, _06373_);
  nand (_26564_, _26563_, _26560_);
  and (_26565_, _12238_, _06373_);
  nor (_26566_, _26565_, _12659_);
  nand (_26567_, _26566_, _26564_);
  nor (_26568_, _12451_, _07216_);
  nor (_26569_, _26568_, _10094_);
  and (_26570_, _26569_, _26567_);
  nor (_26571_, _12239_, _05982_);
  nor (_26572_, _26571_, _26570_);
  nand (_26574_, _26572_, _12172_);
  nor (_26575_, _26431_, _12172_);
  nor (_26576_, _26575_, _06323_);
  nand (_26577_, _26576_, _26574_);
  and (_26578_, _12451_, _06323_);
  nor (_26579_, _26578_, _12668_);
  nand (_26580_, _26579_, _26577_);
  and (_26581_, _08892_, _12668_);
  nor (_26582_, _26581_, _12674_);
  nand (_26583_, _26582_, _26580_);
  and (_26585_, _26412_, _12674_);
  nor (_26586_, _26585_, _09031_);
  and (_26587_, _26586_, _26583_);
  or (_26588_, _26587_, _26425_);
  nand (_26589_, _26588_, _06219_);
  and (_26590_, _12239_, _06218_);
  nor (_26591_, _26590_, _10929_);
  nand (_26592_, _26591_, _26589_);
  and (_26593_, _12451_, _10929_);
  nor (_26594_, _26593_, _12690_);
  nand (_26595_, _26594_, _26592_);
  and (_26596_, _12709_, _12706_);
  nor (_26597_, _26596_, _12710_);
  nor (_26598_, _26597_, _12691_);
  nor (_26599_, _26598_, _06322_);
  nand (_26600_, _26599_, _26595_);
  and (_26601_, _12451_, _06322_);
  nor (_26602_, _26601_, _06217_);
  nand (_26603_, _26602_, _26600_);
  and (_26604_, _08892_, _06217_);
  nor (_26606_, _26604_, _12733_);
  and (_26607_, _26606_, _26603_);
  or (_26608_, _26607_, _26424_);
  nand (_26609_, _26608_, _12169_);
  not (_26610_, _12166_);
  nor (_26611_, _26432_, _12169_);
  nor (_26612_, _26611_, _26610_);
  nand (_26613_, _26612_, _26609_);
  nor (_26614_, _12451_, _12166_);
  nor (_26615_, _26614_, _06369_);
  nand (_26617_, _26615_, _26613_);
  and (_26618_, _12238_, _06369_);
  nor (_26619_, _26618_, _06536_);
  and (_26620_, _26619_, _26617_);
  and (_26621_, _12452_, _06536_);
  or (_26622_, _26621_, _26620_);
  nand (_26623_, _26622_, _05955_);
  and (_26624_, _08892_, _12750_);
  nor (_26625_, _26624_, _12755_);
  and (_26626_, _26625_, _26623_);
  or (_26628_, _26626_, _26420_);
  nand (_26629_, _26628_, _10979_);
  not (_26630_, _12164_);
  nor (_26631_, _26432_, _10979_);
  nor (_26632_, _26631_, _26630_);
  nand (_26633_, _26632_, _26629_);
  nor (_26634_, _12164_, _12451_);
  nor (_26635_, _26634_, _06375_);
  nand (_26636_, _26635_, _26633_);
  and (_26637_, _12238_, _06375_);
  nor (_26639_, _26637_, _06545_);
  and (_26640_, _26639_, _26636_);
  and (_26641_, _12452_, _06545_);
  or (_26642_, _26641_, _26640_);
  nand (_26643_, _26642_, _05961_);
  and (_26644_, _08892_, _07233_);
  nor (_26645_, _26644_, _12776_);
  and (_26646_, _26645_, _26643_);
  and (_26647_, _12451_, \oc8051_golden_model_1.PSW [7]);
  and (_26648_, _26412_, _10558_);
  or (_26650_, _26648_, _26647_);
  and (_26651_, _26650_, _12776_);
  or (_26652_, _26651_, _26646_);
  nand (_26653_, _26652_, _12162_);
  nor (_26654_, _26432_, _12162_);
  nor (_26655_, _26654_, _11023_);
  nand (_26656_, _26655_, _26653_);
  nor (_26657_, _12451_, _11022_);
  nor (_26658_, _26657_, _06366_);
  nand (_26659_, _26658_, _26656_);
  and (_26660_, _12238_, _06366_);
  nor (_26661_, _26660_, _06528_);
  and (_26662_, _26661_, _26659_);
  and (_26663_, _12452_, _06528_);
  or (_26664_, _26663_, _26662_);
  nand (_26665_, _26664_, _05966_);
  and (_26666_, _08892_, _12795_);
  nor (_26667_, _26666_, _12800_);
  and (_26668_, _26667_, _26665_);
  or (_26669_, _26668_, _26416_);
  nand (_26671_, _26669_, _12154_);
  nor (_26672_, _26432_, _12154_);
  nor (_26673_, _26672_, _14297_);
  nand (_26674_, _26673_, _26671_);
  nor (_26675_, _12451_, _12153_);
  nor (_26676_, _26675_, _11125_);
  nand (_26677_, _26676_, _26674_);
  and (_26678_, _26431_, _11125_);
  nor (_26679_, _26678_, _06551_);
  and (_26680_, _26679_, _26677_);
  and (_26682_, _09212_, _06551_);
  or (_26683_, _26682_, _26680_);
  nand (_26684_, _26683_, _05959_);
  and (_26685_, _08892_, _07253_);
  nor (_26686_, _26685_, _06365_);
  and (_26687_, _26686_, _26684_);
  nor (_26688_, _12239_, _13004_);
  and (_26689_, _26464_, _13004_);
  nor (_26690_, _26689_, _26688_);
  nor (_26691_, _26690_, _06558_);
  or (_26693_, _26691_, _26687_);
  nand (_26694_, _26693_, _12151_);
  nor (_26695_, _26432_, _12151_);
  nor (_26696_, _26695_, _19056_);
  nand (_26697_, _26696_, _26694_);
  nor (_26698_, _13012_, _12451_);
  nor (_26699_, _26698_, _11284_);
  nand (_26700_, _26699_, _26697_);
  and (_26701_, _26431_, _11284_);
  nor (_26702_, _26701_, _06281_);
  nand (_26704_, _26702_, _26700_);
  and (_26705_, _09212_, _06281_);
  nor (_26706_, _26705_, _25646_);
  nand (_26707_, _26706_, _26704_);
  nor (_26708_, _08892_, _05964_);
  nor (_26709_, _26708_, _06362_);
  nand (_26710_, _26709_, _26707_);
  and (_26711_, _12239_, _13004_);
  nor (_26712_, _26464_, _13004_);
  nor (_26713_, _26712_, _26711_);
  nor (_26715_, _26713_, _06921_);
  nor (_26716_, _26715_, _13031_);
  nand (_26717_, _26716_, _26710_);
  nor (_26718_, _26432_, _13030_);
  nor (_26719_, _26718_, _06568_);
  nand (_26720_, _26719_, _26717_);
  and (_26721_, _12452_, _06568_);
  nor (_26722_, _26721_, _13038_);
  nand (_26723_, _26722_, _26720_);
  nor (_26724_, _26432_, _13037_);
  nor (_26725_, _26724_, _07695_);
  and (_26726_, _26725_, _26723_);
  or (_26727_, _26726_, _26409_);
  nand (_26728_, _26727_, _05928_);
  nor (_26729_, _26713_, _05928_);
  nor (_26730_, _26729_, _13053_);
  nand (_26731_, _26730_, _26728_);
  nor (_26732_, _26432_, _13052_);
  nor (_26733_, _26732_, _06278_);
  nand (_26734_, _26733_, _26731_);
  and (_26736_, _12452_, _06278_);
  nor (_26737_, _26736_, _13059_);
  nand (_26738_, _26737_, _26734_);
  nor (_26739_, _26432_, _12141_);
  nor (_26740_, _26739_, _25301_);
  nand (_26741_, _26740_, _26738_);
  and (_26742_, _25301_, _08892_);
  nor (_26743_, _26742_, _13068_);
  and (_26744_, _26743_, _26741_);
  and (_26745_, _26431_, _13068_);
  or (_26747_, _26745_, _26744_);
  or (_26748_, _26747_, _01351_);
  or (_26749_, _01347_, \oc8051_golden_model_1.PC [4]);
  and (_26750_, _26749_, _42618_);
  and (_43250_, _26750_, _26748_);
  and (_26751_, _12446_, _06278_);
  and (_26752_, _12446_, _06568_);
  nor (_26753_, \oc8051_golden_model_1.PC [5], \oc8051_golden_model_1.PC [0]);
  nor (_26754_, _12446_, _05630_);
  nor (_26755_, _26754_, _26753_);
  nor (_26757_, _26755_, _12151_);
  nor (_26758_, _26755_, _12154_);
  nor (_26759_, _26755_, _12162_);
  nor (_26760_, _26755_, _10979_);
  nor (_26761_, _26755_, _12169_);
  nor (_26762_, _12446_, _09030_);
  nor (_26763_, _25322_, _12446_);
  not (_26764_, _26755_);
  and (_26765_, _26764_, _12174_);
  or (_26766_, _12534_, _12233_);
  or (_26768_, _12236_, _12235_);
  not (_26769_, _26768_);
  nor (_26770_, _26769_, _12267_);
  and (_26771_, _26769_, _12267_);
  nor (_26772_, _26771_, _26770_);
  not (_26773_, _26772_);
  or (_26774_, _26773_, _12536_);
  and (_26775_, _26774_, _26766_);
  or (_26776_, _26775_, _07151_);
  and (_26777_, _12507_, _12446_);
  or (_26779_, _12448_, _12449_);
  and (_26780_, _26779_, _12474_);
  nor (_26781_, _26779_, _12474_);
  nor (_26782_, _26781_, _26780_);
  and (_26783_, _26782_, _12393_);
  nor (_26784_, _26783_, _26777_);
  nand (_26785_, _26784_, _12387_);
  nor (_26786_, _07486_, \oc8051_golden_model_1.PC [5]);
  nor (_26787_, _26786_, _07141_);
  and (_26788_, _12446_, _07141_);
  nor (_26789_, _26788_, _06781_);
  not (_26790_, _26789_);
  nor (_26791_, _26790_, _26787_);
  not (_26792_, _26791_);
  nor (_26793_, _26755_, _12513_);
  nor (_26794_, _26793_, _06758_);
  and (_26795_, _26794_, _26792_);
  nor (_26796_, _08926_, _07504_);
  or (_26797_, _26796_, _12516_);
  nor (_26798_, _26797_, _26795_);
  nor (_26800_, _26755_, _12512_);
  nor (_26801_, _26800_, _26798_);
  nor (_26802_, _26801_, _12387_);
  nor (_26803_, _26802_, _07154_);
  and (_26804_, _26803_, _26785_);
  and (_26805_, _26755_, _07154_);
  or (_26806_, _26805_, _06341_);
  or (_26807_, _26806_, _26804_);
  nand (_26808_, _26807_, _26776_);
  nand (_26809_, _26808_, _12541_);
  nor (_26811_, _26755_, _12541_);
  nor (_26812_, _26811_, _06272_);
  nand (_26813_, _26812_, _26809_);
  and (_26814_, _12446_, _06272_);
  nor (_26815_, _26814_, _07611_);
  nand (_26816_, _26815_, _26813_);
  and (_26817_, _08926_, _07611_);
  nor (_26818_, _26817_, _06461_);
  nand (_26819_, _26818_, _26816_);
  and (_26820_, _12446_, _06461_);
  nor (_26822_, _26820_, _12551_);
  nand (_26823_, _26822_, _26819_);
  nor (_26824_, _26755_, _12550_);
  nor (_26825_, _26824_, _06464_);
  nand (_26826_, _26825_, _26823_);
  and (_26827_, _12446_, _06464_);
  nor (_26828_, _26827_, _25401_);
  nand (_26829_, _26828_, _26826_);
  nor (_26830_, _26755_, _12560_);
  nor (_26831_, _26830_, _06268_);
  nand (_26833_, _26831_, _26829_);
  and (_26834_, _12446_, _06268_);
  nor (_26835_, _26834_, _12563_);
  nand (_26836_, _26835_, _26833_);
  and (_26837_, _08926_, _12563_);
  nor (_26838_, _26837_, _06267_);
  nand (_26839_, _26838_, _26836_);
  and (_26840_, _12446_, _06267_);
  nor (_26841_, _26840_, _12379_);
  nand (_26842_, _26841_, _26839_);
  and (_26844_, _12371_, _12233_);
  nor (_26845_, _26772_, _12371_);
  or (_26846_, _26845_, _26844_);
  nor (_26847_, _26846_, _12378_);
  nor (_26848_, _26847_, _06347_);
  nand (_26849_, _26848_, _26842_);
  or (_26850_, _26772_, _12333_);
  or (_26851_, _12335_, _12234_);
  nand (_26852_, _26851_, _26850_);
  nand (_26853_, _26852_, _06347_);
  and (_26854_, _26853_, _06774_);
  nand (_26855_, _26854_, _26849_);
  nor (_26856_, _26772_, _12587_);
  not (_26857_, _26856_);
  and (_26858_, _12587_, _12233_);
  nor (_26859_, _26858_, _06774_);
  and (_26860_, _26859_, _26857_);
  nor (_26861_, _26860_, _06371_);
  nand (_26862_, _26861_, _26855_);
  and (_26863_, _12604_, _12234_);
  and (_26865_, _26772_, _26518_);
  or (_26866_, _26865_, _12176_);
  nor (_26867_, _26866_, _26863_);
  nor (_26868_, _26867_, _12174_);
  and (_26869_, _26868_, _26862_);
  or (_26870_, _26869_, _26765_);
  nand (_26871_, _26870_, _06262_);
  and (_26872_, _12447_, _06261_);
  nor (_26873_, _26872_, _12613_);
  nand (_26874_, _26873_, _26871_);
  nor (_26876_, _08926_, _06007_);
  nor (_26877_, _26876_, _25445_);
  and (_26878_, _26877_, _26874_);
  or (_26879_, _26878_, _26763_);
  nand (_26880_, _26879_, _12630_);
  nor (_26881_, _26755_, _12630_);
  nor (_26882_, _26881_, _06505_);
  nand (_26883_, _26882_, _26880_);
  and (_26884_, _12446_, _06505_);
  nor (_26885_, _26884_, _25158_);
  nand (_26887_, _26885_, _26883_);
  and (_26888_, _08926_, _25158_);
  nor (_26889_, _26888_, _06504_);
  nand (_26890_, _26889_, _26887_);
  and (_26891_, _12446_, _06504_);
  nor (_26892_, _26891_, _26197_);
  and (_26893_, _26892_, _26890_);
  nor (_26894_, _26755_, _12639_);
  or (_26895_, _26894_, _26893_);
  nand (_26896_, _26895_, _12643_);
  nor (_26898_, _12446_, _12643_);
  nor (_26899_, _26898_, _10515_);
  nand (_26900_, _26899_, _26896_);
  nor (_26901_, _26764_, _05984_);
  nor (_26902_, _26901_, _06257_);
  and (_26903_, _26902_, _26900_);
  and (_26904_, _12447_, _06257_);
  or (_26905_, _26904_, _26903_);
  nand (_26906_, _26905_, _05978_);
  and (_26907_, _08926_, _06254_);
  nor (_26909_, _26907_, _06373_);
  nand (_26910_, _26909_, _26906_);
  and (_26911_, _12233_, _06373_);
  nor (_26912_, _26911_, _12659_);
  nand (_26913_, _26912_, _26910_);
  nor (_26914_, _12446_, _07216_);
  nor (_26915_, _26914_, _10094_);
  nand (_26916_, _26915_, _26913_);
  nor (_26917_, _12234_, _05982_);
  nor (_26918_, _26917_, _25492_);
  nand (_26920_, _26918_, _26916_);
  nor (_26921_, _26755_, _12172_);
  nor (_26922_, _26921_, _06323_);
  nand (_26923_, _26922_, _26920_);
  and (_26924_, _12446_, _06323_);
  nor (_26925_, _26924_, _12668_);
  nand (_26926_, _26925_, _26923_);
  and (_26927_, _08926_, _12668_);
  nor (_26928_, _26927_, _12674_);
  nand (_26929_, _26928_, _26926_);
  and (_26931_, _26782_, _12674_);
  nor (_26932_, _26931_, _09031_);
  and (_26933_, _26932_, _26929_);
  or (_26934_, _26933_, _26762_);
  nand (_26935_, _26934_, _06219_);
  and (_26936_, _12234_, _06218_);
  nor (_26937_, _26936_, _10929_);
  nand (_26938_, _26937_, _26935_);
  and (_26939_, _12446_, _10929_);
  nor (_26940_, _26939_, _12690_);
  nand (_26941_, _26940_, _26938_);
  and (_26942_, _12711_, _12704_);
  nor (_26943_, _26942_, _12712_);
  nor (_26944_, _26943_, _12691_);
  nor (_26945_, _26944_, _06322_);
  nand (_26946_, _26945_, _26941_);
  and (_26947_, _12446_, _06322_);
  nor (_26948_, _26947_, _06217_);
  nand (_26949_, _26948_, _26946_);
  and (_26950_, _08926_, _06217_);
  nor (_26952_, _26950_, _12733_);
  nand (_26953_, _26952_, _26949_);
  and (_26954_, _12446_, _11342_);
  and (_26955_, _26782_, _12759_);
  or (_26956_, _26955_, _26954_);
  and (_26957_, _26956_, _12733_);
  nor (_26958_, _26957_, _12737_);
  and (_26959_, _26958_, _26953_);
  or (_26960_, _26959_, _26761_);
  nand (_26961_, _26960_, _12166_);
  nor (_26963_, _12446_, _12166_);
  nor (_26964_, _26963_, _06369_);
  nand (_26965_, _26964_, _26961_);
  and (_26966_, _12233_, _06369_);
  nor (_26967_, _26966_, _06536_);
  and (_26968_, _26967_, _26965_);
  and (_26969_, _12447_, _06536_);
  or (_26970_, _26969_, _26968_);
  nand (_26971_, _26970_, _05955_);
  and (_26972_, _08926_, _12750_);
  nor (_26974_, _26972_, _12755_);
  nand (_26975_, _26974_, _26971_);
  nor (_26976_, _12447_, _11342_);
  and (_26977_, _26782_, _11342_);
  or (_26978_, _26977_, _26976_);
  and (_26979_, _26978_, _12755_);
  nor (_26980_, _26979_, _10980_);
  and (_26981_, _26980_, _26975_);
  or (_26982_, _26981_, _26760_);
  nand (_26983_, _26982_, _12164_);
  nor (_26985_, _12164_, _12446_);
  nor (_26986_, _26985_, _06375_);
  nand (_26987_, _26986_, _26983_);
  and (_26988_, _12233_, _06375_);
  nor (_26989_, _26988_, _06545_);
  and (_26990_, _26989_, _26987_);
  and (_26991_, _12447_, _06545_);
  or (_26992_, _26991_, _26990_);
  nand (_26993_, _26992_, _05961_);
  and (_26994_, _08926_, _07233_);
  nor (_26996_, _26994_, _12776_);
  nand (_26997_, _26996_, _26993_);
  nor (_26998_, _26782_, \oc8051_golden_model_1.PSW [7]);
  nor (_26999_, _12446_, _10558_);
  nor (_27000_, _26999_, _12782_);
  not (_27001_, _27000_);
  nor (_27002_, _27001_, _26998_);
  nor (_27003_, _27002_, _12780_);
  and (_27004_, _27003_, _26997_);
  or (_27005_, _27004_, _26759_);
  nand (_27006_, _27005_, _11022_);
  nor (_27007_, _12446_, _11022_);
  nor (_27008_, _27007_, _06366_);
  nand (_27009_, _27008_, _27006_);
  and (_27010_, _12233_, _06366_);
  nor (_27011_, _27010_, _06528_);
  and (_27012_, _27011_, _27009_);
  and (_27013_, _12447_, _06528_);
  or (_27014_, _27013_, _27012_);
  nand (_27015_, _27014_, _05966_);
  and (_27017_, _08926_, _12795_);
  nor (_27018_, _27017_, _12800_);
  nand (_27019_, _27018_, _27015_);
  and (_27020_, _12446_, _10558_);
  and (_27021_, _26782_, \oc8051_golden_model_1.PSW [7]);
  or (_27022_, _27021_, _27020_);
  and (_27023_, _27022_, _12800_);
  nor (_27024_, _27023_, _12804_);
  and (_27025_, _27024_, _27019_);
  or (_27026_, _27025_, _26758_);
  nand (_27028_, _27026_, _12153_);
  nor (_27029_, _12446_, _12153_);
  nor (_27030_, _27029_, _11125_);
  nand (_27031_, _27030_, _27028_);
  and (_27032_, _26755_, _11125_);
  nor (_27033_, _27032_, _06551_);
  and (_27034_, _27033_, _27031_);
  and (_27035_, _09167_, _06551_);
  or (_27036_, _27035_, _27034_);
  nand (_27037_, _27036_, _05959_);
  and (_27039_, _08926_, _07253_);
  nor (_27040_, _27039_, _06365_);
  nand (_27041_, _27040_, _27037_);
  and (_27042_, _26772_, _13004_);
  nor (_27043_, _12233_, _13004_);
  or (_27044_, _27043_, _06558_);
  or (_27045_, _27044_, _27042_);
  and (_27046_, _27045_, _12151_);
  and (_27047_, _27046_, _27041_);
  or (_27048_, _27047_, _26757_);
  nand (_27050_, _27048_, _13012_);
  nor (_27051_, _13012_, _12446_);
  nor (_27052_, _27051_, _11284_);
  nand (_27053_, _27052_, _27050_);
  and (_27054_, _26755_, _11284_);
  nor (_27055_, _27054_, _06281_);
  and (_27056_, _27055_, _27053_);
  and (_27057_, _09167_, _06281_);
  or (_27058_, _27057_, _27056_);
  nand (_27059_, _27058_, _05964_);
  and (_27061_, _08926_, _25646_);
  nor (_27062_, _27061_, _06362_);
  nand (_27063_, _27062_, _27059_);
  and (_27064_, _12234_, _13004_);
  nor (_27065_, _26773_, _13004_);
  nor (_27066_, _27065_, _27064_);
  and (_27067_, _27066_, _06362_);
  nor (_27068_, _27067_, _13031_);
  nand (_27069_, _27068_, _27063_);
  nor (_27070_, _26755_, _13030_);
  nor (_27072_, _27070_, _06568_);
  and (_27073_, _27072_, _27069_);
  or (_27074_, _27073_, _26752_);
  nand (_27075_, _27074_, _13037_);
  nor (_27076_, _26764_, _13037_);
  nor (_27077_, _27076_, _07695_);
  nand (_27078_, _27077_, _27075_);
  and (_27079_, _08926_, _07695_);
  nor (_27080_, _27079_, _05927_);
  nand (_27081_, _27080_, _27078_);
  and (_27083_, _27066_, _05927_);
  nor (_27084_, _27083_, _13053_);
  nand (_27085_, _27084_, _27081_);
  nor (_27086_, _26755_, _13052_);
  nor (_27087_, _27086_, _06278_);
  and (_27088_, _27087_, _27085_);
  or (_27089_, _27088_, _26751_);
  nand (_27090_, _27089_, _12141_);
  nor (_27091_, _26764_, _12141_);
  nor (_27092_, _27091_, _25301_);
  nand (_27094_, _27092_, _27090_);
  and (_27095_, _25301_, _08926_);
  nor (_27096_, _27095_, _13068_);
  and (_27097_, _27096_, _27094_);
  and (_27098_, _26755_, _13068_);
  or (_27099_, _27098_, _27097_);
  or (_27100_, _27099_, _01351_);
  or (_27101_, _01347_, \oc8051_golden_model_1.PC [5]);
  and (_27102_, _27101_, _42618_);
  and (_43251_, _27102_, _27100_);
  and (_27104_, _08657_, _12142_);
  and (_27105_, _08656_, _12142_);
  nor (_27106_, _27105_, \oc8051_golden_model_1.PC [6]);
  nor (_27107_, _27106_, _27104_);
  and (_27108_, _27107_, _13068_);
  and (_27109_, _08857_, _07695_);
  not (_27110_, _27107_);
  and (_27111_, _27110_, _11284_);
  and (_27112_, _12226_, _06366_);
  and (_27113_, _12226_, _06375_);
  and (_27115_, _12226_, _06369_);
  nor (_27116_, _25322_, _12439_);
  and (_27117_, _27110_, _12174_);
  and (_27118_, _12333_, _12226_);
  and (_27119_, _12269_, _12230_);
  nor (_27120_, _27119_, _12270_);
  not (_27121_, _27120_);
  and (_27122_, _27121_, _12335_);
  nor (_27123_, _27122_, _27118_);
  nor (_27124_, _27123_, _12177_);
  and (_27126_, _12440_, _06268_);
  nor (_27127_, _27107_, _12550_);
  or (_27128_, _27120_, _12536_);
  or (_27129_, _12534_, _12225_);
  and (_27130_, _27129_, _06341_);
  nand (_27131_, _27130_, _27128_);
  and (_27132_, _12507_, _12439_);
  nor (_27133_, _12476_, _12443_);
  nor (_27134_, _27133_, _12477_);
  and (_27135_, _27134_, _12393_);
  nor (_27137_, _27135_, _27132_);
  nand (_27138_, _27137_, _12387_);
  and (_27139_, _08857_, _06758_);
  and (_27140_, _12440_, _07141_);
  nor (_27141_, _27140_, _06781_);
  and (_27142_, _07487_, \oc8051_golden_model_1.PC [6]);
  or (_27143_, _27142_, _07141_);
  and (_27144_, _27143_, _27141_);
  nor (_27145_, _27110_, _12513_);
  or (_27146_, _27145_, _06758_);
  nor (_27148_, _27146_, _27144_);
  nor (_27149_, _27148_, _12516_);
  not (_27150_, _27149_);
  nor (_27151_, _27150_, _27139_);
  nor (_27152_, _27110_, _12512_);
  nor (_27153_, _27152_, _12387_);
  not (_27154_, _27153_);
  nor (_27155_, _27154_, _27151_);
  not (_27156_, _27155_);
  nor (_27157_, _07154_, _06341_);
  and (_27159_, _27157_, _27156_);
  nand (_27160_, _27159_, _27138_);
  nand (_27161_, _27160_, _27131_);
  and (_27162_, _27161_, _12541_);
  or (_27163_, _12542_, _07154_);
  and (_27164_, _27163_, _27107_);
  or (_27165_, _27164_, _06272_);
  or (_27166_, _27165_, _27162_);
  and (_27167_, _12440_, _06272_);
  nor (_27168_, _27167_, _07611_);
  and (_27170_, _27168_, _27166_);
  nor (_27171_, _08857_, _06010_);
  or (_27172_, _27171_, _06461_);
  nor (_27173_, _27172_, _27170_);
  and (_27174_, _12440_, _06461_);
  or (_27175_, _27174_, _27173_);
  and (_27176_, _27175_, _12550_);
  or (_27177_, _27176_, _27127_);
  nand (_27178_, _27177_, _06465_);
  and (_27179_, _12440_, _06464_);
  nor (_27181_, _27179_, _25401_);
  nand (_27182_, _27181_, _27178_);
  nor (_27183_, _27110_, _12560_);
  nor (_27184_, _27183_, _06268_);
  and (_27185_, _27184_, _27182_);
  or (_27186_, _27185_, _27126_);
  nand (_27187_, _27186_, _06013_);
  and (_27188_, _08857_, _12563_);
  nor (_27189_, _27188_, _06267_);
  nand (_27190_, _27189_, _27187_);
  and (_27192_, _12439_, _06267_);
  nor (_27193_, _27192_, _12379_);
  and (_27194_, _27193_, _27190_);
  and (_27195_, _12371_, _12225_);
  nor (_27196_, _27121_, _12371_);
  or (_27197_, _27196_, _12378_);
  nor (_27198_, _27197_, _27195_);
  or (_27199_, _27198_, _27194_);
  and (_27200_, _27199_, _12177_);
  nor (_27201_, _27200_, _27124_);
  or (_27203_, _27201_, _06480_);
  nor (_27204_, _27121_, _12587_);
  and (_27205_, _12587_, _12225_);
  or (_27206_, _27205_, _06774_);
  or (_27207_, _27206_, _27204_);
  and (_27208_, _27207_, _12176_);
  nand (_27209_, _27208_, _27203_);
  and (_27210_, _12604_, _12225_);
  and (_27211_, _27120_, _26518_);
  or (_27212_, _27211_, _27210_);
  and (_27214_, _27212_, _06371_);
  nor (_27215_, _27214_, _12174_);
  and (_27216_, _27215_, _27209_);
  or (_27217_, _27216_, _27117_);
  nand (_27218_, _27217_, _06262_);
  and (_27219_, _12440_, _06261_);
  nor (_27220_, _27219_, _12613_);
  nand (_27221_, _27220_, _27218_);
  nor (_27222_, _08857_, _06007_);
  nor (_27223_, _27222_, _25445_);
  and (_27225_, _27223_, _27221_);
  or (_27226_, _27225_, _27116_);
  nand (_27227_, _27226_, _12630_);
  nor (_27228_, _27107_, _12630_);
  nor (_27229_, _27228_, _06505_);
  nand (_27230_, _27229_, _27227_);
  and (_27231_, _12439_, _06505_);
  nor (_27232_, _27231_, _25158_);
  nand (_27233_, _27232_, _27230_);
  and (_27234_, _08857_, _25158_);
  nor (_27235_, _27234_, _06504_);
  nand (_27236_, _27235_, _27233_);
  and (_27237_, _12439_, _06504_);
  nor (_27238_, _27237_, _26197_);
  nand (_27239_, _27238_, _27236_);
  nor (_27240_, _27107_, _12639_);
  nor (_27241_, _27240_, _12644_);
  nand (_27242_, _27241_, _27239_);
  nor (_27243_, _12440_, _12643_);
  nor (_27244_, _27243_, _10515_);
  and (_27247_, _27244_, _27242_);
  nor (_27248_, _27107_, _05984_);
  or (_27249_, _27248_, _27247_);
  nand (_27250_, _27249_, _06258_);
  and (_27251_, _12440_, _06257_);
  nor (_27252_, _27251_, _06254_);
  nand (_27253_, _27252_, _27250_);
  nor (_27254_, _08857_, _05978_);
  nor (_27255_, _27254_, _06373_);
  nand (_27256_, _27255_, _27253_);
  and (_27258_, _12226_, _06373_);
  nor (_27259_, _27258_, _12659_);
  nand (_27260_, _27259_, _27256_);
  nor (_27261_, _12440_, _07216_);
  nor (_27262_, _27261_, _10094_);
  nand (_27263_, _27262_, _27260_);
  nor (_27264_, _12225_, _05982_);
  nor (_27265_, _27264_, _25492_);
  nand (_27266_, _27265_, _27263_);
  nor (_27267_, _27110_, _12172_);
  nor (_27269_, _27267_, _06323_);
  nand (_27270_, _27269_, _27266_);
  and (_27271_, _12440_, _06323_);
  nor (_27272_, _27271_, _12668_);
  nand (_27273_, _27272_, _27270_);
  nor (_27274_, _08857_, _05946_);
  nor (_27275_, _27274_, _12674_);
  nand (_27276_, _27275_, _27273_);
  nor (_27277_, _27134_, _12679_);
  nor (_27278_, _27277_, _09031_);
  nand (_27280_, _27278_, _27276_);
  nor (_27281_, _12440_, _09030_);
  nor (_27282_, _27281_, _06218_);
  nand (_27283_, _27282_, _27280_);
  and (_27284_, _12226_, _06218_);
  nor (_27285_, _27284_, _10929_);
  nand (_27286_, _27285_, _27283_);
  and (_27287_, _12439_, _10929_);
  nor (_27288_, _27287_, _12690_);
  nand (_27289_, _27288_, _27286_);
  and (_27291_, _12713_, _12700_);
  nor (_27292_, _27291_, _12714_);
  nor (_27293_, _27292_, _12691_);
  nor (_27294_, _27293_, _06322_);
  nand (_27295_, _27294_, _27289_);
  and (_27296_, _12439_, _06322_);
  nor (_27297_, _27296_, _06217_);
  nand (_27298_, _27297_, _27295_);
  and (_27299_, _08857_, _06217_);
  nor (_27300_, _27299_, _12733_);
  nand (_27302_, _27300_, _27298_);
  and (_27303_, _12439_, _11342_);
  and (_27304_, _27134_, _12759_);
  or (_27305_, _27304_, _27303_);
  and (_27306_, _27305_, _12733_);
  nor (_27307_, _27306_, _12737_);
  nand (_27308_, _27307_, _27302_);
  nor (_27309_, _27107_, _12169_);
  nor (_27310_, _27309_, _26610_);
  nand (_27311_, _27310_, _27308_);
  nor (_27313_, _12440_, _12166_);
  nor (_27314_, _27313_, _06369_);
  and (_27315_, _27314_, _27311_);
  or (_27316_, _27315_, _27115_);
  nand (_27317_, _27316_, _07240_);
  and (_27318_, _12440_, _06536_);
  nor (_27319_, _27318_, _12750_);
  and (_27320_, _27319_, _27317_);
  nor (_27321_, _08857_, _05955_);
  or (_27322_, _27321_, _27320_);
  nand (_27324_, _27322_, _25061_);
  nor (_27325_, _12440_, _11342_);
  and (_27326_, _27134_, _11342_);
  or (_27327_, _27326_, _27325_);
  and (_27328_, _27327_, _12755_);
  nor (_27329_, _27328_, _10980_);
  nand (_27330_, _27329_, _27324_);
  nor (_27331_, _27107_, _10979_);
  nor (_27332_, _27331_, _26630_);
  nand (_27333_, _27332_, _27330_);
  nor (_27335_, _12164_, _12440_);
  nor (_27336_, _27335_, _06375_);
  and (_27337_, _27336_, _27333_);
  or (_27338_, _27337_, _27113_);
  nand (_27339_, _27338_, _07234_);
  and (_27340_, _12440_, _06545_);
  nor (_27341_, _27340_, _07233_);
  and (_27342_, _27341_, _27339_);
  nor (_27343_, _08857_, _05961_);
  or (_27344_, _27343_, _27342_);
  nand (_27346_, _27344_, _12782_);
  nor (_27347_, _27134_, \oc8051_golden_model_1.PSW [7]);
  nor (_27348_, _12439_, _10558_);
  nor (_27349_, _27348_, _12782_);
  not (_27350_, _27349_);
  nor (_27351_, _27350_, _27347_);
  nor (_27352_, _27351_, _12780_);
  nand (_27353_, _27352_, _27346_);
  nor (_27354_, _27107_, _12162_);
  nor (_27355_, _27354_, _11023_);
  nand (_27357_, _27355_, _27353_);
  nor (_27358_, _12440_, _11022_);
  nor (_27359_, _27358_, _06366_);
  and (_27360_, _27359_, _27357_);
  or (_27361_, _27360_, _27112_);
  nand (_27362_, _27361_, _09061_);
  and (_27363_, _12440_, _06528_);
  nor (_27364_, _27363_, _12795_);
  and (_27365_, _27364_, _27362_);
  nor (_27366_, _08857_, _05966_);
  or (_27368_, _27366_, _27365_);
  nand (_27369_, _27368_, _25056_);
  and (_27370_, _12439_, _10558_);
  and (_27371_, _27134_, \oc8051_golden_model_1.PSW [7]);
  or (_27372_, _27371_, _27370_);
  and (_27373_, _27372_, _12800_);
  nor (_27374_, _27373_, _12804_);
  nand (_27375_, _27374_, _27369_);
  nor (_27376_, _27107_, _12154_);
  nor (_27377_, _27376_, _14297_);
  nand (_27379_, _27377_, _27375_);
  nor (_27380_, _12440_, _12153_);
  nor (_27381_, _27380_, _11125_);
  nand (_27382_, _27381_, _27379_);
  and (_27383_, _27110_, _11125_);
  nor (_27384_, _27383_, _06551_);
  nand (_27385_, _27384_, _27382_);
  and (_27386_, _09446_, _06551_);
  nor (_27387_, _27386_, _07253_);
  nand (_27388_, _27387_, _27385_);
  and (_27390_, _08857_, _07253_);
  nor (_27391_, _27390_, _06365_);
  nand (_27392_, _27391_, _27388_);
  nor (_27393_, _12225_, _13004_);
  and (_27394_, _27121_, _13004_);
  or (_27395_, _27394_, _06558_);
  or (_27396_, _27395_, _27393_);
  and (_27397_, _27396_, _12151_);
  nand (_27398_, _27397_, _27392_);
  nor (_27399_, _27107_, _12151_);
  nor (_27401_, _27399_, _19056_);
  nand (_27402_, _27401_, _27398_);
  nor (_27403_, _13012_, _12440_);
  nor (_27404_, _27403_, _11284_);
  and (_27405_, _27404_, _27402_);
  or (_27406_, _27405_, _27111_);
  nand (_27407_, _27406_, _06282_);
  and (_27408_, _09122_, _06281_);
  nor (_27409_, _27408_, _25646_);
  nand (_27410_, _27409_, _27407_);
  nor (_27412_, _08857_, _05964_);
  nor (_27413_, _27412_, _06362_);
  and (_27414_, _27413_, _27410_);
  nor (_27415_, _27120_, _13004_);
  and (_27416_, _12226_, _13004_);
  nor (_27417_, _27416_, _27415_);
  nor (_27418_, _27417_, _06921_);
  or (_27419_, _27418_, _27414_);
  and (_27420_, _27419_, _13030_);
  nor (_27421_, _27107_, _13030_);
  or (_27423_, _27421_, _27420_);
  nand (_27424_, _27423_, _06926_);
  and (_27425_, _12440_, _06568_);
  nor (_27426_, _27425_, _13038_);
  nand (_27427_, _27426_, _27424_);
  nor (_27428_, _27110_, _13037_);
  nor (_27429_, _27428_, _07695_);
  and (_27430_, _27429_, _27427_);
  or (_27431_, _27430_, _27109_);
  nand (_27432_, _27431_, _05928_);
  nor (_27434_, _27417_, _05928_);
  nor (_27435_, _27434_, _13053_);
  nand (_27436_, _27435_, _27432_);
  nor (_27437_, _27110_, _13052_);
  nor (_27438_, _27437_, _06278_);
  nand (_27439_, _27438_, _27436_);
  and (_27440_, _12440_, _06278_);
  nor (_27441_, _27440_, _13059_);
  nand (_27442_, _27441_, _27439_);
  nor (_27443_, _27110_, _12141_);
  nor (_27445_, _27443_, _25301_);
  nand (_27446_, _27445_, _27442_);
  and (_27447_, _25301_, _08857_);
  nor (_27448_, _27447_, _13068_);
  and (_27449_, _27448_, _27446_);
  or (_27450_, _27449_, _27108_);
  or (_27451_, _27450_, _01351_);
  or (_27452_, _01347_, \oc8051_golden_model_1.PC [6]);
  and (_27453_, _27452_, _42618_);
  and (_43252_, _27453_, _27451_);
  and (_27455_, _08661_, _06278_);
  and (_27456_, _27104_, \oc8051_golden_model_1.PC [7]);
  nor (_27457_, _27104_, \oc8051_golden_model_1.PC [7]);
  nor (_27458_, _27457_, _27456_);
  nor (_27459_, _27458_, _12151_);
  nor (_27460_, _27458_, _12154_);
  nor (_27461_, _27458_, _12162_);
  nor (_27462_, _27458_, _10979_);
  nor (_27463_, _27458_, _12169_);
  nor (_27464_, _09030_, _08661_);
  nor (_27466_, _27458_, _12639_);
  nor (_27467_, _25322_, _08661_);
  or (_27468_, _12534_, _09415_);
  or (_27469_, _12221_, _12222_);
  and (_27470_, _27469_, _12271_);
  nor (_27471_, _27469_, _12271_);
  nor (_27472_, _27471_, _27470_);
  or (_27473_, _27472_, _12536_);
  and (_27474_, _27473_, _27468_);
  or (_27475_, _27474_, _07151_);
  and (_27477_, _12507_, _08661_);
  and (_27478_, _12478_, _12436_);
  nor (_27479_, _27478_, _12479_);
  and (_27480_, _27479_, _12393_);
  nor (_27481_, _27480_, _27477_);
  nand (_27482_, _27481_, _12387_);
  nor (_27483_, _07486_, \oc8051_golden_model_1.PC [7]);
  nor (_27484_, _27483_, _07141_);
  and (_27485_, _08661_, _07141_);
  nor (_27486_, _27485_, _06781_);
  not (_27488_, _27486_);
  nor (_27489_, _27488_, _27484_);
  not (_27490_, _27489_);
  nor (_27491_, _27458_, _12513_);
  nor (_27492_, _27491_, _06758_);
  and (_27493_, _27492_, _27490_);
  nor (_27494_, _08608_, _07504_);
  or (_27495_, _27494_, _12516_);
  nor (_27496_, _27495_, _27493_);
  nor (_27497_, _27458_, _12512_);
  nor (_27499_, _27497_, _27496_);
  nor (_27500_, _27499_, _12387_);
  nor (_27501_, _27500_, _07154_);
  and (_27502_, _27501_, _27482_);
  and (_27503_, _27458_, _07154_);
  or (_27504_, _27503_, _06341_);
  or (_27505_, _27504_, _27502_);
  nand (_27506_, _27505_, _27475_);
  nand (_27507_, _27506_, _12541_);
  nor (_27508_, _27458_, _12541_);
  nor (_27510_, _27508_, _06272_);
  nand (_27511_, _27510_, _27507_);
  and (_27512_, _08661_, _06272_);
  nor (_27513_, _27512_, _07611_);
  nand (_27514_, _27513_, _27511_);
  and (_27515_, _08608_, _07611_);
  nor (_27516_, _27515_, _06461_);
  nand (_27517_, _27516_, _27514_);
  and (_27518_, _08661_, _06461_);
  nor (_27519_, _27518_, _12551_);
  nand (_27521_, _27519_, _27517_);
  nor (_27522_, _27458_, _12550_);
  nor (_27523_, _27522_, _06464_);
  nand (_27524_, _27523_, _27521_);
  and (_27525_, _08661_, _06464_);
  nor (_27526_, _27525_, _25401_);
  nand (_27527_, _27526_, _27524_);
  nor (_27528_, _27458_, _12560_);
  nor (_27529_, _27528_, _06268_);
  nand (_27530_, _27529_, _27527_);
  and (_27532_, _08661_, _06268_);
  nor (_27533_, _27532_, _12563_);
  nand (_27534_, _27533_, _27530_);
  and (_27535_, _08608_, _12563_);
  nor (_27536_, _27535_, _06267_);
  nand (_27537_, _27536_, _27534_);
  and (_27538_, _08661_, _06267_);
  nor (_27539_, _27538_, _12379_);
  nand (_27540_, _27539_, _27537_);
  and (_27541_, _12371_, _09415_);
  not (_27543_, _27472_);
  nor (_27544_, _27543_, _12371_);
  or (_27545_, _27544_, _12378_);
  nor (_27546_, _27545_, _27541_);
  nor (_27547_, _27546_, _06347_);
  nand (_27548_, _27547_, _27540_);
  or (_27549_, _27543_, _12333_);
  or (_27550_, _12335_, _09416_);
  nand (_27551_, _27550_, _27549_);
  nand (_27552_, _27551_, _06347_);
  and (_27554_, _27552_, _06774_);
  and (_27555_, _27554_, _27548_);
  and (_27556_, _12587_, _09415_);
  nor (_27557_, _27543_, _12587_);
  or (_27558_, _27557_, _06774_);
  nor (_27559_, _27558_, _27556_);
  or (_27560_, _27559_, _06371_);
  or (_27561_, _27560_, _27555_);
  nand (_27562_, _12604_, _09415_);
  nand (_27563_, _27472_, _26518_);
  and (_27565_, _27563_, _27562_);
  or (_27566_, _27565_, _12176_);
  and (_27567_, _27566_, _27561_);
  or (_27568_, _27567_, _12174_);
  nand (_27569_, _27458_, _12174_);
  and (_27570_, _27569_, _27568_);
  nand (_27571_, _27570_, _06262_);
  and (_27572_, _08794_, _06261_);
  nor (_27573_, _27572_, _12613_);
  nand (_27574_, _27573_, _27571_);
  nor (_27576_, _08608_, _06007_);
  nor (_27577_, _27576_, _25445_);
  and (_27578_, _27577_, _27574_);
  or (_27579_, _27578_, _27467_);
  nand (_27580_, _27579_, _12630_);
  nor (_27581_, _27458_, _12630_);
  nor (_27582_, _27581_, _06505_);
  nand (_27583_, _27582_, _27580_);
  and (_27584_, _08661_, _06505_);
  nor (_27585_, _27584_, _25158_);
  nand (_27587_, _27585_, _27583_);
  and (_27588_, _08608_, _25158_);
  nor (_27589_, _27588_, _06504_);
  nand (_27590_, _27589_, _27587_);
  and (_27591_, _08661_, _06504_);
  nor (_27592_, _27591_, _26197_);
  and (_27593_, _27592_, _27590_);
  or (_27594_, _27593_, _27466_);
  nand (_27595_, _27594_, _12643_);
  nor (_27596_, _12643_, _08661_);
  nor (_27598_, _27596_, _10515_);
  nand (_27599_, _27598_, _27595_);
  not (_27600_, _27458_);
  nor (_27601_, _27600_, _05984_);
  nor (_27602_, _27601_, _06257_);
  and (_27603_, _27602_, _27599_);
  and (_27604_, _08794_, _06257_);
  or (_27605_, _27604_, _27603_);
  nand (_27606_, _27605_, _05978_);
  and (_27607_, _08608_, _06254_);
  nor (_27609_, _27607_, _06373_);
  nand (_27610_, _27609_, _27606_);
  and (_27611_, _09415_, _06373_);
  nor (_27612_, _27611_, _12659_);
  nand (_27613_, _27612_, _27610_);
  nor (_27614_, _08661_, _07216_);
  nor (_27615_, _27614_, _10094_);
  nand (_27616_, _27615_, _27613_);
  nor (_27617_, _09416_, _05982_);
  nor (_27618_, _27617_, _25492_);
  nand (_27620_, _27618_, _27616_);
  nor (_27621_, _27458_, _12172_);
  nor (_27622_, _27621_, _06323_);
  nand (_27623_, _27622_, _27620_);
  and (_27624_, _08661_, _06323_);
  nor (_27625_, _27624_, _12668_);
  nand (_27626_, _27625_, _27623_);
  and (_27627_, _08608_, _12668_);
  nor (_27628_, _27627_, _12674_);
  nand (_27629_, _27628_, _27626_);
  and (_27631_, _27479_, _12674_);
  nor (_27632_, _27631_, _09031_);
  and (_27633_, _27632_, _27629_);
  or (_27634_, _27633_, _27464_);
  nand (_27635_, _27634_, _06219_);
  and (_27636_, _09416_, _06218_);
  nor (_27637_, _27636_, _10929_);
  nand (_27638_, _27637_, _27635_);
  and (_27639_, _10929_, _08661_);
  nor (_27640_, _27639_, _12690_);
  nand (_27642_, _27640_, _27638_);
  or (_27643_, _12695_, _12694_);
  not (_27644_, _27643_);
  and (_27645_, _27644_, _12715_);
  nor (_27646_, _27644_, _12715_);
  nor (_27647_, _27646_, _27645_);
  and (_27648_, _27647_, _12690_);
  nor (_27649_, _27648_, _06322_);
  nand (_27650_, _27649_, _27642_);
  and (_27651_, _08661_, _06322_);
  nor (_27653_, _27651_, _06217_);
  nand (_27654_, _27653_, _27650_);
  and (_27655_, _08608_, _06217_);
  nor (_27656_, _27655_, _12733_);
  nand (_27657_, _27656_, _27654_);
  and (_27658_, _11342_, _08661_);
  and (_27659_, _27479_, _12759_);
  or (_27660_, _27659_, _27658_);
  and (_27661_, _27660_, _12733_);
  nor (_27662_, _27661_, _12737_);
  and (_27664_, _27662_, _27657_);
  or (_27665_, _27664_, _27463_);
  nand (_27666_, _27665_, _12166_);
  nor (_27667_, _12166_, _08661_);
  nor (_27668_, _27667_, _06369_);
  nand (_27669_, _27668_, _27666_);
  and (_27670_, _09415_, _06369_);
  nor (_27671_, _27670_, _06536_);
  and (_27672_, _27671_, _27669_);
  and (_27673_, _08794_, _06536_);
  or (_27675_, _27673_, _27672_);
  nand (_27676_, _27675_, _05955_);
  and (_27677_, _08608_, _12750_);
  nor (_27678_, _27677_, _12755_);
  nand (_27679_, _27678_, _27676_);
  nor (_27680_, _11342_, _08794_);
  and (_27681_, _27479_, _11342_);
  or (_27682_, _27681_, _27680_);
  and (_27683_, _27682_, _12755_);
  nor (_27684_, _27683_, _10980_);
  and (_27686_, _27684_, _27679_);
  or (_27687_, _27686_, _27462_);
  nand (_27688_, _27687_, _12164_);
  nor (_27689_, _12164_, _08661_);
  nor (_27690_, _27689_, _06375_);
  nand (_27691_, _27690_, _27688_);
  and (_27692_, _09415_, _06375_);
  nor (_27693_, _27692_, _06545_);
  and (_27694_, _27693_, _27691_);
  and (_27695_, _08794_, _06545_);
  or (_27697_, _27695_, _27694_);
  nand (_27698_, _27697_, _05961_);
  and (_27699_, _08608_, _07233_);
  nor (_27700_, _27699_, _12776_);
  nand (_27701_, _27700_, _27698_);
  nor (_27702_, _27479_, \oc8051_golden_model_1.PSW [7]);
  nor (_27703_, _08661_, _10558_);
  nor (_27704_, _27703_, _12782_);
  not (_27705_, _27704_);
  nor (_27706_, _27705_, _27702_);
  nor (_27708_, _27706_, _12780_);
  and (_27709_, _27708_, _27701_);
  or (_27710_, _27709_, _27461_);
  nand (_27711_, _27710_, _11022_);
  nor (_27712_, _11022_, _08661_);
  nor (_27713_, _27712_, _06366_);
  nand (_27714_, _27713_, _27711_);
  and (_27715_, _09415_, _06366_);
  nor (_27716_, _27715_, _06528_);
  and (_27717_, _27716_, _27714_);
  and (_27719_, _08794_, _06528_);
  or (_27720_, _27719_, _27717_);
  nand (_27721_, _27720_, _05966_);
  and (_27722_, _08608_, _12795_);
  nor (_27723_, _27722_, _12800_);
  nand (_27724_, _27723_, _27721_);
  and (_27725_, _08661_, _10558_);
  and (_27726_, _27479_, \oc8051_golden_model_1.PSW [7]);
  or (_27727_, _27726_, _27725_);
  and (_27728_, _27727_, _12800_);
  nor (_27730_, _27728_, _12804_);
  and (_27731_, _27730_, _27724_);
  or (_27732_, _27731_, _27460_);
  nand (_27733_, _27732_, _12153_);
  nor (_27734_, _12153_, _08661_);
  nor (_27735_, _27734_, _11125_);
  nand (_27736_, _27735_, _27733_);
  and (_27737_, _27458_, _11125_);
  nor (_27738_, _27737_, _06551_);
  and (_27739_, _27738_, _27736_);
  nor (_27741_, _08755_, _06716_);
  or (_27742_, _27741_, _27739_);
  nand (_27743_, _27742_, _05959_);
  and (_27744_, _08608_, _07253_);
  nor (_27745_, _27744_, _06365_);
  nand (_27746_, _27745_, _27743_);
  and (_27747_, _27543_, _13004_);
  nor (_27748_, _09415_, _13004_);
  or (_27749_, _27748_, _06558_);
  or (_27750_, _27749_, _27747_);
  and (_27752_, _27750_, _12151_);
  and (_27753_, _27752_, _27746_);
  or (_27754_, _27753_, _27459_);
  nand (_27755_, _27754_, _13012_);
  nor (_27756_, _13012_, _08661_);
  nor (_27757_, _27756_, _11284_);
  nand (_27758_, _27757_, _27755_);
  and (_27759_, _27458_, _11284_);
  nor (_27760_, _27759_, _06281_);
  and (_27761_, _27760_, _27758_);
  nor (_27763_, _08755_, _06282_);
  or (_27764_, _27763_, _27761_);
  nand (_27765_, _27764_, _05964_);
  and (_27766_, _08608_, _25646_);
  nor (_27767_, _27766_, _06362_);
  nand (_27768_, _27767_, _27765_);
  and (_27769_, _09416_, _13004_);
  nor (_27770_, _27472_, _13004_);
  nor (_27771_, _27770_, _27769_);
  and (_27772_, _27771_, _06362_);
  nor (_27774_, _27772_, _13031_);
  nand (_27775_, _27774_, _27768_);
  nor (_27776_, _27458_, _13030_);
  nor (_27777_, _27776_, _06568_);
  nand (_27778_, _27777_, _27775_);
  and (_27779_, _08661_, _06568_);
  nor (_27780_, _27779_, _13038_);
  and (_27781_, _27780_, _27778_);
  nor (_27782_, _27458_, _13037_);
  or (_27783_, _27782_, _27781_);
  nand (_27785_, _27783_, _07271_);
  and (_27786_, _08608_, _07695_);
  nor (_27787_, _27786_, _05927_);
  nand (_27788_, _27787_, _27785_);
  and (_27789_, _27771_, _05927_);
  nor (_27790_, _27789_, _13053_);
  nand (_27791_, _27790_, _27788_);
  nor (_27792_, _27458_, _13052_);
  nor (_27793_, _27792_, _06278_);
  and (_27794_, _27793_, _27791_);
  or (_27796_, _27794_, _27455_);
  nand (_27797_, _27796_, _12141_);
  nor (_27798_, _27600_, _12141_);
  nor (_27799_, _27798_, _25301_);
  nand (_27800_, _27799_, _27797_);
  and (_27801_, _25301_, _08608_);
  nor (_27802_, _27801_, _13068_);
  and (_27803_, _27802_, _27800_);
  and (_27804_, _27458_, _13068_);
  or (_27805_, _27804_, _27803_);
  or (_27807_, _27805_, _01351_);
  or (_27808_, _01347_, \oc8051_golden_model_1.PC [7]);
  and (_27809_, _27808_, _42618_);
  and (_43253_, _27809_, _27807_);
  nor (_27810_, _12140_, _06251_);
  nor (_27811_, _14508_, _06251_);
  and (_27812_, _27456_, \oc8051_golden_model_1.PC [8]);
  nor (_27813_, _27456_, \oc8051_golden_model_1.PC [8]);
  nor (_27814_, _27813_, _27812_);
  nor (_27815_, _27814_, _12151_);
  nor (_27817_, _27814_, _12154_);
  nor (_27818_, _27814_, _12162_);
  nor (_27819_, _27814_, _10979_);
  and (_27820_, _12275_, _06369_);
  nor (_27821_, _27814_, _12169_);
  nor (_27822_, _12431_, _09030_);
  and (_27823_, _12431_, _06323_);
  nor (_27824_, _25322_, _12431_);
  and (_27825_, _12431_, _06268_);
  or (_27826_, _06461_, _07611_);
  nand (_27828_, _12431_, _06272_);
  and (_27829_, _12536_, _12276_);
  nor (_27830_, _12279_, _12273_);
  nor (_27831_, _27830_, _12280_);
  not (_27832_, _27831_);
  and (_27833_, _27832_, _12534_);
  or (_27834_, _27833_, _27829_);
  and (_27835_, _27834_, _06341_);
  not (_27836_, _12431_);
  or (_27837_, _12393_, _27836_);
  and (_27839_, _12483_, _12480_);
  nor (_27840_, _27839_, _12484_);
  nand (_27841_, _27840_, _12393_);
  and (_27842_, _27841_, _27837_);
  and (_27843_, _27842_, _12387_);
  nand (_27844_, _12431_, _07141_);
  nand (_27845_, _07142_, \oc8051_golden_model_1.PC [8]);
  or (_27846_, _27845_, _07486_);
  and (_27847_, _27846_, _27844_);
  or (_27848_, _27847_, _06781_);
  and (_27850_, _27848_, _07504_);
  or (_27851_, _27850_, _12516_);
  not (_27852_, _27814_);
  or (_27853_, _27852_, _12514_);
  and (_27854_, _27853_, _08654_);
  and (_27855_, _27854_, _27851_);
  or (_27856_, _27855_, _07154_);
  or (_27857_, _27856_, _27843_);
  nand (_27858_, _27814_, _07154_);
  and (_27859_, _27858_, _07151_);
  and (_27861_, _27859_, _27857_);
  or (_27862_, _27861_, _27835_);
  and (_27863_, _27862_, _12541_);
  nor (_27864_, _27814_, _12541_);
  or (_27865_, _27864_, _06272_);
  or (_27866_, _27865_, _27863_);
  and (_27867_, _27866_, _27828_);
  nor (_27868_, _27867_, _27826_);
  and (_27869_, _12431_, _06461_);
  nor (_27870_, _27869_, _12551_);
  not (_27871_, _27870_);
  nor (_27872_, _27871_, _27868_);
  nor (_27873_, _27814_, _12550_);
  nor (_27874_, _27873_, _06464_);
  not (_27875_, _27874_);
  nor (_27876_, _27875_, _27872_);
  and (_27877_, _12431_, _06464_);
  nor (_27878_, _27877_, _25401_);
  not (_27879_, _27878_);
  or (_27880_, _27879_, _27876_);
  nor (_27883_, _27814_, _12560_);
  nor (_27884_, _27883_, _06268_);
  and (_27885_, _27884_, _27880_);
  or (_27886_, _27885_, _27825_);
  nand (_27887_, _27886_, _12564_);
  and (_27888_, _12431_, _06267_);
  nor (_27889_, _27888_, _12379_);
  nand (_27890_, _27889_, _27887_);
  and (_27891_, _12371_, _12275_);
  nor (_27892_, _27832_, _12371_);
  or (_27894_, _27892_, _27891_);
  nor (_27895_, _27894_, _12378_);
  nor (_27896_, _27895_, _06347_);
  nand (_27897_, _27896_, _27890_);
  and (_27898_, _27831_, _12335_);
  and (_27899_, _12333_, _12275_);
  nor (_27900_, _27899_, _27898_);
  nor (_27901_, _27900_, _12177_);
  nor (_27902_, _27901_, _06480_);
  nand (_27903_, _27902_, _27897_);
  and (_27905_, _12587_, _12275_);
  not (_27906_, _27905_);
  nor (_27907_, _27832_, _12587_);
  nor (_27908_, _27907_, _06774_);
  and (_27909_, _27908_, _27906_);
  nor (_27910_, _27909_, _06371_);
  nand (_27911_, _27910_, _27903_);
  and (_27912_, _12604_, _12275_);
  and (_27913_, _27831_, _26518_);
  or (_27914_, _27913_, _27912_);
  and (_27916_, _27914_, _06371_);
  nor (_27917_, _27916_, _12174_);
  nand (_27918_, _27917_, _27911_);
  and (_27919_, _27852_, _12174_);
  nor (_27920_, _27919_, _06261_);
  nand (_27921_, _27920_, _27918_);
  and (_27922_, _12431_, _06261_);
  not (_27923_, _27922_);
  and (_27924_, _25322_, _06007_);
  and (_27925_, _27924_, _27923_);
  and (_27927_, _27925_, _27921_);
  or (_27928_, _27927_, _27824_);
  nand (_27929_, _27928_, _12630_);
  nor (_27930_, _27814_, _12630_);
  nor (_27931_, _27930_, _06505_);
  nand (_27932_, _27931_, _27929_);
  and (_27933_, _12431_, _06505_);
  nor (_27934_, _27933_, _25158_);
  nand (_27935_, _27934_, _27932_);
  nand (_27936_, _27935_, _14057_);
  and (_27938_, _12431_, _06504_);
  nor (_27939_, _27938_, _26197_);
  and (_27940_, _27939_, _27936_);
  nor (_27941_, _27814_, _12639_);
  or (_27942_, _27941_, _27940_);
  nand (_27943_, _27942_, _12643_);
  nor (_27944_, _12431_, _12643_);
  nor (_27945_, _27944_, _10515_);
  nand (_27946_, _27945_, _27943_);
  nor (_27947_, _27852_, _05984_);
  nor (_27949_, _27947_, _06257_);
  nand (_27950_, _27949_, _27946_);
  nor (_27951_, _06373_, _06254_);
  not (_27952_, _27951_);
  and (_27953_, _27836_, _06257_);
  nor (_27954_, _27953_, _27952_);
  nand (_27955_, _27954_, _27950_);
  and (_27956_, _12275_, _06373_);
  nor (_27957_, _27956_, _12659_);
  nand (_27958_, _27957_, _27955_);
  nor (_27960_, _12431_, _07216_);
  nor (_27961_, _27960_, _10094_);
  nand (_27962_, _27961_, _27958_);
  nor (_27963_, _12276_, _05982_);
  nor (_27964_, _27963_, _25492_);
  nand (_27965_, _27964_, _27962_);
  nor (_27966_, _27814_, _12172_);
  nor (_27967_, _27966_, _06323_);
  and (_27968_, _27967_, _27965_);
  or (_27969_, _27968_, _27823_);
  nor (_27971_, _12674_, _12668_);
  nand (_27972_, _27971_, _27969_);
  and (_27973_, _27840_, _12674_);
  nor (_27974_, _27973_, _09031_);
  and (_27975_, _27974_, _27972_);
  or (_27976_, _27975_, _27822_);
  nand (_27977_, _27976_, _06219_);
  and (_27978_, _12276_, _06218_);
  nor (_27979_, _27978_, _10929_);
  nand (_27980_, _27979_, _27977_);
  and (_27982_, _12431_, _10929_);
  nor (_27983_, _27982_, _12690_);
  nand (_27984_, _27983_, _27980_);
  and (_27985_, _12717_, _12693_);
  nor (_27986_, _27985_, _12718_);
  nor (_27987_, _27986_, _12691_);
  nor (_27988_, _27987_, _06322_);
  nand (_27989_, _27988_, _27984_);
  and (_27990_, _12431_, _06322_);
  nor (_27991_, _27990_, _06217_);
  nand (_27993_, _27991_, _27989_);
  nand (_27994_, _27993_, _25064_);
  and (_27995_, _12431_, _11342_);
  and (_27996_, _27840_, _12759_);
  or (_27997_, _27996_, _27995_);
  and (_27998_, _27997_, _12733_);
  nor (_27999_, _27998_, _12737_);
  and (_28000_, _27999_, _27994_);
  or (_28001_, _28000_, _27821_);
  nand (_28002_, _28001_, _12166_);
  nor (_28004_, _12431_, _12166_);
  nor (_28005_, _28004_, _06369_);
  and (_28006_, _28005_, _28002_);
  or (_28007_, _28006_, _27820_);
  nand (_28008_, _28007_, _07240_);
  and (_28009_, _12431_, _06536_);
  nor (_28010_, _28009_, _12750_);
  nand (_28011_, _28010_, _28008_);
  nand (_28012_, _28011_, _25061_);
  nor (_28013_, _27836_, _11342_);
  and (_28015_, _27840_, _11342_);
  or (_28016_, _28015_, _28013_);
  and (_28017_, _28016_, _12755_);
  nor (_28018_, _28017_, _10980_);
  and (_28019_, _28018_, _28012_);
  or (_28020_, _28019_, _27819_);
  nand (_28021_, _28020_, _12164_);
  nor (_28022_, _12164_, _12431_);
  nor (_28023_, _28022_, _06375_);
  nand (_28024_, _28023_, _28021_);
  and (_28026_, _12275_, _06375_);
  nor (_28027_, _28026_, _06545_);
  nand (_28028_, _28027_, _28024_);
  nor (_28029_, _12776_, _07233_);
  and (_28030_, _27836_, _06545_);
  not (_28031_, _28030_);
  and (_28032_, _28031_, _28029_);
  nand (_28033_, _28032_, _28028_);
  nor (_28034_, _27840_, \oc8051_golden_model_1.PSW [7]);
  nor (_28035_, _12431_, _10558_);
  nor (_28037_, _28035_, _12782_);
  not (_28038_, _28037_);
  nor (_28039_, _28038_, _28034_);
  nor (_28040_, _28039_, _12780_);
  and (_28041_, _28040_, _28033_);
  or (_28042_, _28041_, _27818_);
  nand (_28043_, _28042_, _11022_);
  nor (_28044_, _12431_, _11022_);
  nor (_28045_, _28044_, _06366_);
  nand (_28046_, _28045_, _28043_);
  and (_28048_, _12275_, _06366_);
  nor (_28049_, _28048_, _06528_);
  nand (_28050_, _28049_, _28046_);
  nor (_28051_, _12800_, _12795_);
  and (_28052_, _27836_, _06528_);
  not (_28053_, _28052_);
  and (_28054_, _28053_, _28051_);
  nand (_28055_, _28054_, _28050_);
  and (_28056_, _12431_, _10558_);
  and (_28057_, _27840_, \oc8051_golden_model_1.PSW [7]);
  or (_28059_, _28057_, _28056_);
  and (_28060_, _28059_, _12800_);
  nor (_28061_, _28060_, _12804_);
  and (_28062_, _28061_, _28055_);
  or (_28063_, _28062_, _27817_);
  nand (_28064_, _28063_, _12153_);
  nor (_28065_, _12431_, _12153_);
  nor (_28066_, _28065_, _11125_);
  and (_28067_, _28066_, _28064_);
  and (_28068_, _27814_, _11125_);
  or (_28070_, _28068_, _28067_);
  nand (_28071_, _28070_, _06716_);
  and (_28072_, _07133_, _06551_);
  nor (_28073_, _28072_, _07253_);
  nand (_28074_, _28073_, _28071_);
  nand (_28075_, _28074_, _06558_);
  and (_28076_, _27832_, _13004_);
  nor (_28077_, _12275_, _13004_);
  or (_28078_, _28077_, _06558_);
  or (_28079_, _28078_, _28076_);
  and (_28081_, _28079_, _12151_);
  and (_28082_, _28081_, _28075_);
  or (_28083_, _28082_, _27815_);
  nand (_28084_, _28083_, _13012_);
  nor (_28085_, _13012_, _12431_);
  nor (_28086_, _28085_, _11284_);
  and (_28087_, _28086_, _28084_);
  and (_28088_, _27814_, _11284_);
  or (_28089_, _28088_, _28087_);
  nand (_28090_, _28089_, _06282_);
  and (_28092_, _07133_, _06281_);
  nor (_28093_, _28092_, _25646_);
  nand (_28094_, _28093_, _28090_);
  nand (_28095_, _28094_, _06921_);
  and (_28096_, _12276_, _13004_);
  nor (_28097_, _27831_, _13004_);
  nor (_28098_, _28097_, _28096_);
  and (_28099_, _28098_, _06362_);
  nor (_28100_, _28099_, _13031_);
  nand (_28101_, _28100_, _28095_);
  nor (_28103_, _27814_, _13030_);
  nor (_28104_, _28103_, _06568_);
  nand (_28105_, _28104_, _28101_);
  and (_28106_, _12431_, _06568_);
  nor (_28107_, _28106_, _13038_);
  nand (_28108_, _28107_, _28105_);
  nor (_28109_, _27814_, _13037_);
  nor (_28110_, _28109_, _06361_);
  and (_28111_, _28110_, _28108_);
  or (_28112_, _28111_, _27811_);
  nor (_28114_, _05940_, _05927_);
  nand (_28115_, _28114_, _28112_);
  and (_28116_, _28098_, _05927_);
  nor (_28117_, _28116_, _13053_);
  nand (_28118_, _28117_, _28115_);
  nor (_28119_, _27814_, _13052_);
  nor (_28120_, _28119_, _06278_);
  nand (_28121_, _28120_, _28118_);
  and (_28122_, _12431_, _06278_);
  nor (_28123_, _28122_, _13059_);
  nand (_28125_, _28123_, _28121_);
  nor (_28126_, _27814_, _12141_);
  nor (_28127_, _28126_, _06379_);
  and (_28128_, _28127_, _28125_);
  or (_28129_, _28128_, _27810_);
  nor (_28130_, _13068_, _05939_);
  and (_28131_, _28130_, _28129_);
  and (_28132_, _27814_, _13068_);
  or (_28133_, _28132_, _28131_);
  or (_28134_, _28133_, _01351_);
  or (_28136_, _01347_, \oc8051_golden_model_1.PC [8]);
  and (_28137_, _28136_, _42618_);
  and (_43254_, _28137_, _28134_);
  nor (_28138_, _07004_, _12140_);
  nor (_28139_, _07004_, _14508_);
  and (_28140_, _27812_, \oc8051_golden_model_1.PC [9]);
  nor (_28141_, _27812_, \oc8051_golden_model_1.PC [9]);
  nor (_28142_, _28141_, _28140_);
  nor (_28143_, _28142_, _12151_);
  nor (_28144_, _28142_, _12154_);
  and (_28146_, _12216_, _06366_);
  nor (_28147_, _28142_, _12162_);
  and (_28148_, _12216_, _06375_);
  nor (_28149_, _28142_, _10979_);
  and (_28150_, _12216_, _06369_);
  nor (_28151_, _28142_, _12169_);
  nor (_28152_, _12426_, _09030_);
  and (_28153_, _12426_, _06323_);
  and (_28154_, _12426_, _06504_);
  nor (_28155_, _06504_, _25158_);
  not (_28157_, _28142_);
  and (_28158_, _28157_, _12174_);
  nor (_28159_, _12280_, _12277_);
  and (_28160_, _28159_, _12220_);
  nor (_28161_, _28159_, _12220_);
  nor (_28162_, _28161_, _28160_);
  and (_28163_, _28162_, _12335_);
  and (_28164_, _12333_, _12217_);
  nor (_28165_, _28164_, _28163_);
  nor (_28166_, _28165_, _12177_);
  nand (_28168_, _12426_, _07141_);
  nand (_28169_, _07142_, \oc8051_golden_model_1.PC [9]);
  or (_28170_, _28169_, _07486_);
  and (_28171_, _28170_, _28168_);
  or (_28172_, _28171_, _06781_);
  and (_28173_, _28172_, _07504_);
  or (_28174_, _28173_, _12516_);
  or (_28175_, _28157_, _12514_);
  and (_28176_, _28175_, _08654_);
  and (_28177_, _28176_, _28174_);
  and (_28178_, _12507_, _12426_);
  or (_28179_, _12427_, _12428_);
  not (_28180_, _28179_);
  nor (_28181_, _28180_, _12485_);
  and (_28182_, _28180_, _12485_);
  nor (_28183_, _28182_, _28181_);
  nor (_28184_, _28183_, _12507_);
  nor (_28185_, _28184_, _28178_);
  and (_28186_, _28185_, _12387_);
  or (_28187_, _28186_, _28177_);
  nand (_28190_, _28187_, _07155_);
  and (_28191_, _28157_, _07154_);
  nor (_28192_, _28191_, _06341_);
  and (_28193_, _28192_, _28190_);
  and (_28194_, _28162_, _12534_);
  and (_28195_, _12536_, _12217_);
  or (_28196_, _28195_, _07151_);
  nor (_28197_, _28196_, _28194_);
  or (_28198_, _28197_, _12542_);
  or (_28199_, _28198_, _28193_);
  nor (_28201_, _28142_, _12541_);
  nor (_28202_, _28201_, _06272_);
  nand (_28203_, _28202_, _28199_);
  and (_28204_, _12426_, _06272_);
  nor (_28205_, _28204_, _07611_);
  nand (_28206_, _28205_, _28203_);
  nand (_28207_, _28206_, _07166_);
  and (_28208_, _12426_, _06461_);
  nor (_28209_, _28208_, _12551_);
  nand (_28210_, _28209_, _28207_);
  nor (_28212_, _28142_, _12550_);
  nor (_28213_, _28212_, _06464_);
  nand (_28214_, _28213_, _28210_);
  and (_28215_, _12426_, _06464_);
  nor (_28216_, _28215_, _25401_);
  nand (_28217_, _28216_, _28214_);
  nor (_28218_, _28142_, _12560_);
  nor (_28219_, _28218_, _06268_);
  nand (_28220_, _28219_, _28217_);
  and (_28221_, _12426_, _06268_);
  nor (_28223_, _28221_, _12563_);
  nand (_28224_, _28223_, _28220_);
  nand (_28225_, _28224_, _07303_);
  and (_28226_, _12426_, _06267_);
  nor (_28227_, _28226_, _12379_);
  and (_28228_, _28227_, _28225_);
  and (_28229_, _12371_, _12216_);
  nor (_28230_, _28162_, _12371_);
  or (_28231_, _28230_, _12378_);
  nor (_28232_, _28231_, _28229_);
  or (_28234_, _28232_, _28228_);
  and (_28235_, _28234_, _12177_);
  or (_28236_, _28235_, _28166_);
  or (_28237_, _28236_, _06480_);
  nor (_28238_, _28162_, _12587_);
  and (_28239_, _12587_, _12216_);
  nor (_28240_, _28239_, _28238_);
  or (_28241_, _28240_, _06774_);
  and (_28242_, _28241_, _28237_);
  or (_28243_, _28242_, _06371_);
  and (_28245_, _12604_, _12216_);
  nor (_28246_, _28162_, _12604_);
  or (_28247_, _28246_, _28245_);
  and (_28248_, _28247_, _06371_);
  nor (_28249_, _28248_, _12174_);
  and (_28250_, _28249_, _28243_);
  or (_28251_, _28250_, _28158_);
  nand (_28252_, _28251_, _06262_);
  not (_28253_, _12426_);
  and (_28254_, _28253_, _06261_);
  not (_28256_, _28254_);
  and (_28257_, _28256_, _27924_);
  nand (_28258_, _28257_, _28252_);
  nor (_28259_, _25322_, _28253_);
  nor (_28260_, _28259_, _12631_);
  nand (_28261_, _28260_, _28258_);
  nor (_28262_, _28142_, _12630_);
  nor (_28263_, _28262_, _06505_);
  and (_28264_, _28263_, _28261_);
  and (_28265_, _12426_, _06505_);
  or (_28267_, _28265_, _28264_);
  and (_28268_, _28267_, _28155_);
  or (_28269_, _28268_, _28154_);
  nand (_28270_, _28269_, _12639_);
  nor (_28271_, _28157_, _12639_);
  nor (_28272_, _28271_, _12644_);
  nand (_28273_, _28272_, _28270_);
  nor (_28274_, _12426_, _12643_);
  nor (_28275_, _28274_, _10515_);
  nand (_28276_, _28275_, _28273_);
  nor (_28278_, _28157_, _05984_);
  nor (_28279_, _28278_, _06257_);
  nand (_28280_, _28279_, _28276_);
  and (_28281_, _28253_, _06257_);
  nor (_28282_, _28281_, _27952_);
  nand (_28283_, _28282_, _28280_);
  and (_28284_, _12216_, _06373_);
  nor (_28285_, _28284_, _12659_);
  nand (_28286_, _28285_, _28283_);
  nor (_28287_, _12426_, _07216_);
  nor (_28289_, _28287_, _10094_);
  nand (_28290_, _28289_, _28286_);
  nor (_28291_, _12217_, _05982_);
  nor (_28292_, _28291_, _25492_);
  nand (_28293_, _28292_, _28290_);
  nor (_28294_, _28142_, _12172_);
  nor (_28295_, _28294_, _06323_);
  and (_28296_, _28295_, _28293_);
  or (_28297_, _28296_, _28153_);
  nand (_28298_, _28297_, _27971_);
  nor (_28300_, _28183_, _12679_);
  nor (_28301_, _28300_, _09031_);
  and (_28302_, _28301_, _28298_);
  or (_28303_, _28302_, _28152_);
  nand (_28304_, _28303_, _06219_);
  and (_28305_, _12217_, _06218_);
  nor (_28306_, _28305_, _10929_);
  nand (_28307_, _28306_, _28304_);
  and (_28308_, _12426_, _10929_);
  nor (_28309_, _28308_, _12690_);
  nand (_28311_, _28309_, _28307_);
  nor (_28312_, _12718_, \oc8051_golden_model_1.DPH [1]);
  nor (_28313_, _28312_, _12719_);
  nor (_28314_, _28313_, _12691_);
  nor (_28315_, _28314_, _06322_);
  nand (_28316_, _28315_, _28311_);
  and (_28317_, _12426_, _06322_);
  nor (_28318_, _28317_, _06217_);
  nand (_28319_, _28318_, _28316_);
  nand (_28320_, _28319_, _25064_);
  and (_28322_, _12426_, _11342_);
  nor (_28323_, _28183_, _11342_);
  or (_28324_, _28323_, _28322_);
  and (_28325_, _28324_, _12733_);
  nor (_28326_, _28325_, _12737_);
  and (_28327_, _28326_, _28320_);
  or (_28328_, _28327_, _28151_);
  nand (_28329_, _28328_, _12166_);
  nor (_28330_, _12426_, _12166_);
  nor (_28331_, _28330_, _06369_);
  and (_28333_, _28331_, _28329_);
  or (_28334_, _28333_, _28150_);
  nand (_28335_, _28334_, _07240_);
  and (_28336_, _12426_, _06536_);
  nor (_28337_, _28336_, _12750_);
  nand (_28338_, _28337_, _28335_);
  nand (_28339_, _28338_, _25061_);
  and (_28340_, _28183_, _11342_);
  nor (_28341_, _12426_, _11342_);
  nor (_28342_, _28341_, _25061_);
  not (_28344_, _28342_);
  nor (_28345_, _28344_, _28340_);
  nor (_28346_, _28345_, _10980_);
  and (_28347_, _28346_, _28339_);
  or (_28348_, _28347_, _28149_);
  nand (_28349_, _28348_, _12164_);
  nor (_28350_, _12164_, _12426_);
  nor (_28351_, _28350_, _06375_);
  and (_28352_, _28351_, _28349_);
  or (_28353_, _28352_, _28148_);
  nand (_28355_, _28353_, _07234_);
  and (_28356_, _12426_, _06545_);
  nor (_28357_, _28356_, _07233_);
  nand (_28358_, _28357_, _28355_);
  nand (_28359_, _28358_, _12782_);
  and (_28360_, _12426_, \oc8051_golden_model_1.PSW [7]);
  nor (_28361_, _28183_, \oc8051_golden_model_1.PSW [7]);
  or (_28362_, _28361_, _28360_);
  and (_28363_, _28362_, _12776_);
  nor (_28364_, _28363_, _12780_);
  and (_28366_, _28364_, _28359_);
  or (_28367_, _28366_, _28147_);
  nand (_28368_, _28367_, _11022_);
  nor (_28369_, _12426_, _11022_);
  nor (_28370_, _28369_, _06366_);
  and (_28371_, _28370_, _28368_);
  or (_28372_, _28371_, _28146_);
  nand (_28373_, _28372_, _09061_);
  and (_28374_, _12426_, _06528_);
  nor (_28375_, _28374_, _12795_);
  nand (_28377_, _28375_, _28373_);
  nand (_28378_, _28377_, _25056_);
  and (_28379_, _12426_, _10558_);
  nor (_28380_, _28183_, _10558_);
  or (_28381_, _28380_, _28379_);
  and (_28382_, _28381_, _12800_);
  nor (_28383_, _28382_, _12804_);
  and (_28384_, _28383_, _28378_);
  or (_28385_, _28384_, _28144_);
  nand (_28386_, _28385_, _12153_);
  nor (_28388_, _12426_, _12153_);
  nor (_28389_, _28388_, _11125_);
  nand (_28390_, _28389_, _28386_);
  and (_28391_, _28142_, _11125_);
  nor (_28392_, _28391_, _06551_);
  nand (_28393_, _28392_, _28390_);
  nor (_28394_, _06365_, _07253_);
  not (_28395_, _28394_);
  and (_28396_, _07357_, _06551_);
  nor (_28397_, _28396_, _28395_);
  nand (_28399_, _28397_, _28393_);
  nor (_28400_, _12216_, _13004_);
  and (_28401_, _28162_, _13004_);
  or (_28402_, _28401_, _06558_);
  or (_28403_, _28402_, _28400_);
  and (_28404_, _28403_, _12151_);
  and (_28405_, _28404_, _28399_);
  or (_28406_, _28405_, _28143_);
  nand (_28407_, _28406_, _13012_);
  nor (_28408_, _13012_, _12426_);
  nor (_28410_, _28408_, _11284_);
  nand (_28411_, _28410_, _28407_);
  and (_28412_, _28142_, _11284_);
  nor (_28413_, _28412_, _06281_);
  nand (_28414_, _28413_, _28411_);
  nor (_28415_, _06362_, _25646_);
  not (_28416_, _28415_);
  and (_28417_, _07357_, _06281_);
  nor (_28418_, _28417_, _28416_);
  nand (_28419_, _28418_, _28414_);
  and (_28421_, _12216_, _13004_);
  nor (_28422_, _28162_, _13004_);
  or (_28423_, _28422_, _28421_);
  and (_28424_, _28423_, _06362_);
  nor (_28425_, _28424_, _13031_);
  nand (_28426_, _28425_, _28419_);
  nor (_28427_, _28142_, _13030_);
  nor (_28428_, _28427_, _06568_);
  nand (_28429_, _28428_, _28426_);
  and (_28430_, _12426_, _06568_);
  nor (_28432_, _28430_, _13038_);
  nand (_28433_, _28432_, _28429_);
  nor (_28434_, _28142_, _13037_);
  nor (_28435_, _28434_, _06361_);
  and (_28436_, _28435_, _28433_);
  or (_28437_, _28436_, _28139_);
  nand (_28438_, _28437_, _28114_);
  and (_28439_, _28423_, _05927_);
  nor (_28440_, _28439_, _13053_);
  nand (_28441_, _28440_, _28438_);
  nor (_28443_, _28142_, _13052_);
  nor (_28444_, _28443_, _06278_);
  nand (_28445_, _28444_, _28441_);
  and (_28446_, _12426_, _06278_);
  nor (_28447_, _28446_, _13059_);
  nand (_28448_, _28447_, _28445_);
  nor (_28449_, _28142_, _12141_);
  nor (_28450_, _28449_, _06379_);
  and (_28451_, _28450_, _28448_);
  or (_28452_, _28451_, _28138_);
  and (_28454_, _28452_, _28130_);
  and (_28455_, _28142_, _13068_);
  or (_28456_, _28455_, _28454_);
  or (_28457_, _28456_, _01351_);
  or (_28458_, _01347_, \oc8051_golden_model_1.PC [9]);
  and (_28459_, _28458_, _42618_);
  and (_43255_, _28459_, _28457_);
  nand (_28460_, _12203_, _06366_);
  nand (_28461_, _12203_, _06375_);
  nand (_28462_, _12203_, _06369_);
  nand (_28464_, _07412_, _05925_);
  and (_28465_, _28140_, \oc8051_golden_model_1.PC [10]);
  nor (_28466_, _28140_, \oc8051_golden_model_1.PC [10]);
  nor (_28467_, _28466_, _28465_);
  and (_28468_, _28467_, _25492_);
  and (_28469_, _28467_, _25401_);
  or (_28470_, _28467_, _12550_);
  and (_28471_, _28467_, _27163_);
  nor (_28472_, _12284_, _12281_);
  not (_28473_, _28472_);
  and (_28475_, _28473_, _12213_);
  nor (_28476_, _28473_, _12213_);
  nor (_28477_, _28476_, _28475_);
  or (_28478_, _28477_, _12536_);
  or (_28479_, _12534_, _12202_);
  and (_28480_, _28479_, _06341_);
  and (_28481_, _28480_, _28478_);
  and (_28482_, _12507_, _12421_);
  nor (_28483_, _12488_, _12424_);
  nor (_28484_, _28483_, _12489_);
  and (_28486_, _28484_, _12393_);
  or (_28487_, _28486_, _28482_);
  or (_28488_, _28487_, _08654_);
  and (_28489_, _12421_, _07141_);
  nand (_28490_, _07142_, \oc8051_golden_model_1.PC [10]);
  nor (_28491_, _28490_, _07486_);
  or (_28492_, _28491_, _28489_);
  and (_28493_, _28492_, _06782_);
  or (_28494_, _28493_, _06758_);
  and (_28495_, _28494_, _12512_);
  not (_28497_, _12514_);
  and (_28498_, _28467_, _28497_);
  or (_28499_, _28498_, _12387_);
  or (_28500_, _28499_, _28495_);
  and (_28501_, _28500_, _27157_);
  and (_28502_, _28501_, _28488_);
  or (_28503_, _28502_, _28481_);
  and (_28504_, _28503_, _12541_);
  or (_28505_, _28504_, _28471_);
  and (_28506_, _28505_, _06466_);
  and (_28508_, _12421_, _06467_);
  nor (_28509_, _28508_, _07611_);
  nand (_28510_, _28509_, _12550_);
  or (_28511_, _28510_, _28506_);
  and (_28512_, _28511_, _28470_);
  or (_28513_, _28512_, _06464_);
  or (_28514_, _12421_, _06465_);
  and (_28515_, _28514_, _12560_);
  and (_28516_, _28515_, _28513_);
  or (_28517_, _28516_, _28469_);
  and (_28519_, _28517_, _06269_);
  and (_28520_, _12421_, _06268_);
  or (_28521_, _28520_, _12563_);
  or (_28522_, _28521_, _28519_);
  and (_28523_, _28522_, _07303_);
  nand (_28524_, _12421_, _06267_);
  nand (_28525_, _28524_, _12378_);
  or (_28526_, _28525_, _28523_);
  or (_28527_, _28477_, _12371_);
  nand (_28528_, _12371_, _12203_);
  and (_28529_, _28528_, _28527_);
  or (_28530_, _28529_, _12378_);
  and (_28531_, _28530_, _12177_);
  and (_28532_, _28531_, _28526_);
  and (_28533_, _28477_, _12335_);
  and (_28534_, _12333_, _12202_);
  or (_28535_, _28534_, _28533_);
  and (_28536_, _28535_, _06347_);
  or (_28537_, _28536_, _06480_);
  or (_28538_, _28537_, _28532_);
  and (_28541_, _12587_, _12202_);
  not (_28542_, _12587_);
  and (_28543_, _28477_, _28542_);
  or (_28544_, _28543_, _06774_);
  or (_28545_, _28544_, _28541_);
  and (_28546_, _28545_, _12176_);
  and (_28547_, _28546_, _28538_);
  or (_28548_, _28477_, _12604_);
  nand (_28549_, _12604_, _12203_);
  and (_28550_, _28549_, _06371_);
  and (_28552_, _28550_, _28548_);
  or (_28553_, _28552_, _12174_);
  or (_28554_, _28553_, _28547_);
  or (_28555_, _28467_, _12175_);
  and (_28556_, _25322_, _06262_);
  and (_28557_, _28556_, _28555_);
  and (_28558_, _28557_, _28554_);
  not (_28559_, _12421_);
  nor (_28560_, _28556_, _28559_);
  nand (_28561_, _12630_, _06007_);
  or (_28563_, _28561_, _28560_);
  or (_28564_, _28563_, _28558_);
  or (_28565_, _28467_, _12630_);
  and (_28566_, _28565_, _14058_);
  and (_28567_, _28566_, _28564_);
  or (_28568_, _28567_, _25158_);
  and (_28569_, _28568_, _14057_);
  or (_28570_, _28559_, _06506_);
  nand (_28571_, _28570_, _12639_);
  or (_28572_, _28571_, _28569_);
  or (_28574_, _28467_, _12639_);
  and (_28575_, _28574_, _12643_);
  and (_28576_, _28575_, _28572_);
  nor (_28577_, _28559_, _12643_);
  or (_28578_, _28577_, _10515_);
  or (_28579_, _28578_, _28576_);
  or (_28580_, _28467_, _05984_);
  and (_28581_, _28580_, _06258_);
  and (_28582_, _28581_, _28579_);
  nand (_28583_, _12421_, _06257_);
  nand (_28585_, _28583_, _27951_);
  or (_28586_, _28585_, _28582_);
  nand (_28587_, _12203_, _06373_);
  and (_28588_, _28587_, _07216_);
  and (_28589_, _28588_, _28586_);
  nor (_28590_, _28559_, _07216_);
  or (_28591_, _28590_, _10094_);
  or (_28592_, _28591_, _28589_);
  or (_28593_, _12202_, _05982_);
  and (_28594_, _28593_, _12172_);
  and (_28596_, _28594_, _28592_);
  nor (_28597_, _28596_, _28468_);
  nor (_28598_, _28597_, _06323_);
  nand (_28599_, _12421_, _06323_);
  nand (_28600_, _28599_, _27971_);
  or (_28601_, _28600_, _28598_);
  or (_28602_, _28484_, _12679_);
  and (_28603_, _28602_, _09030_);
  and (_28604_, _28603_, _28601_);
  nor (_28605_, _28559_, _09030_);
  or (_28607_, _28605_, _06218_);
  or (_28608_, _28607_, _28604_);
  and (_28609_, _12203_, _06218_);
  nor (_28610_, _28609_, _10929_);
  and (_28611_, _28610_, _28608_);
  and (_28612_, _12421_, _10929_);
  or (_28613_, _28612_, _12690_);
  or (_28614_, _28613_, _28611_);
  nor (_28615_, _12719_, \oc8051_golden_model_1.DPH [2]);
  nor (_28616_, _28615_, _12720_);
  or (_28618_, _28616_, _12691_);
  and (_28619_, _28618_, _06881_);
  and (_28620_, _28619_, _28614_);
  and (_28621_, _12421_, _06322_);
  or (_28622_, _28621_, _28620_);
  and (_28623_, _28622_, _28464_);
  or (_28624_, _28484_, _11342_);
  or (_28625_, _12421_, _12759_);
  and (_28626_, _28625_, _12733_);
  and (_28627_, _28626_, _28624_);
  or (_28629_, _28627_, _12737_);
  or (_28630_, _28629_, _28623_);
  or (_28631_, _28467_, _12169_);
  and (_28632_, _28631_, _12166_);
  and (_28633_, _28632_, _28630_);
  nor (_28634_, _28559_, _12166_);
  or (_28635_, _28634_, _06369_);
  or (_28636_, _28635_, _28633_);
  and (_28637_, _28636_, _28462_);
  or (_28638_, _28637_, _06536_);
  nand (_28640_, _28559_, _06536_);
  nor (_28641_, _12755_, _12750_);
  and (_28642_, _28641_, _28640_);
  and (_28643_, _28642_, _28638_);
  or (_28644_, _28484_, _12759_);
  or (_28645_, _12421_, _11342_);
  and (_28646_, _28645_, _12755_);
  and (_28647_, _28646_, _28644_);
  or (_28648_, _28647_, _10980_);
  or (_28649_, _28648_, _28643_);
  or (_28651_, _28467_, _10979_);
  and (_28652_, _28651_, _12164_);
  and (_28653_, _28652_, _28649_);
  nor (_28654_, _12164_, _28559_);
  or (_28655_, _28654_, _06375_);
  or (_28656_, _28655_, _28653_);
  and (_28657_, _28656_, _28461_);
  or (_28658_, _28657_, _06545_);
  nand (_28659_, _28559_, _06545_);
  and (_28660_, _28659_, _28029_);
  and (_28662_, _28660_, _28658_);
  or (_28663_, _28484_, \oc8051_golden_model_1.PSW [7]);
  or (_28664_, _12421_, _10558_);
  and (_28665_, _28664_, _12776_);
  and (_28666_, _28665_, _28663_);
  or (_28667_, _28666_, _12780_);
  or (_28668_, _28667_, _28662_);
  or (_28669_, _28467_, _12162_);
  and (_28670_, _28669_, _11022_);
  and (_28671_, _28670_, _28668_);
  nor (_28673_, _28559_, _11022_);
  or (_28674_, _28673_, _06366_);
  or (_28675_, _28674_, _28671_);
  and (_28676_, _28675_, _28460_);
  or (_28677_, _28676_, _06528_);
  nand (_28678_, _28559_, _06528_);
  and (_28679_, _28678_, _28051_);
  and (_28680_, _28679_, _28677_);
  or (_28681_, _28484_, _10558_);
  or (_28682_, _12421_, \oc8051_golden_model_1.PSW [7]);
  and (_28684_, _28682_, _12800_);
  and (_28685_, _28684_, _28681_);
  or (_28686_, _28685_, _12804_);
  or (_28687_, _28686_, _28680_);
  or (_28688_, _28467_, _12154_);
  and (_28689_, _28688_, _12153_);
  and (_28690_, _28689_, _28687_);
  nor (_28691_, _28559_, _12153_);
  or (_28692_, _28691_, _11125_);
  or (_28693_, _28692_, _28690_);
  or (_28695_, _28467_, _11126_);
  and (_28696_, _28695_, _28693_);
  or (_28697_, _28696_, _06551_);
  nand (_28698_, _07776_, _06551_);
  and (_28699_, _28698_, _28394_);
  and (_28700_, _28699_, _28697_);
  not (_28701_, _13004_);
  or (_28702_, _28477_, _28701_);
  or (_28703_, _12202_, _13004_);
  and (_28704_, _28703_, _06365_);
  and (_28706_, _28704_, _28702_);
  or (_28707_, _28706_, _25625_);
  or (_28708_, _28707_, _28700_);
  or (_28709_, _28467_, _12151_);
  and (_28710_, _28709_, _13012_);
  and (_28711_, _28710_, _28708_);
  nor (_28712_, _13012_, _28559_);
  or (_28713_, _28712_, _11284_);
  or (_28714_, _28713_, _28711_);
  or (_28715_, _28467_, _11285_);
  and (_28717_, _28715_, _28714_);
  or (_28718_, _28717_, _06281_);
  nand (_28719_, _07776_, _06281_);
  and (_28720_, _28719_, _28415_);
  and (_28721_, _28720_, _28718_);
  or (_28722_, _28477_, _13004_);
  nand (_28723_, _12203_, _13004_);
  and (_28724_, _28723_, _28722_);
  and (_28725_, _28724_, _06362_);
  or (_28726_, _28725_, _13031_);
  or (_28728_, _28726_, _28721_);
  or (_28729_, _28467_, _13030_);
  and (_28730_, _28729_, _28728_);
  or (_28731_, _28730_, _06568_);
  nand (_28732_, _28559_, _06568_);
  and (_28733_, _28732_, _13037_);
  and (_28734_, _28733_, _28731_);
  and (_28735_, _28467_, _13038_);
  or (_28736_, _28735_, _06361_);
  or (_28737_, _28736_, _28734_);
  nand (_28739_, _06656_, _06361_);
  and (_28740_, _28739_, _28114_);
  and (_28741_, _28740_, _28737_);
  and (_28742_, _28724_, _05927_);
  or (_28743_, _28742_, _13053_);
  or (_28744_, _28743_, _28741_);
  or (_28745_, _28467_, _13052_);
  and (_28746_, _28745_, _28744_);
  or (_28747_, _28746_, _06278_);
  nand (_28748_, _28559_, _06278_);
  and (_28750_, _28748_, _12141_);
  and (_28751_, _28750_, _28747_);
  and (_28752_, _28467_, _13059_);
  or (_28753_, _28752_, _06379_);
  or (_28754_, _28753_, _28751_);
  nand (_28755_, _06656_, _06379_);
  and (_28756_, _28755_, _28130_);
  and (_28757_, _28756_, _28754_);
  and (_28758_, _28467_, _13068_);
  or (_28759_, _28758_, _28757_);
  or (_28761_, _28759_, _01351_);
  or (_28762_, _01347_, \oc8051_golden_model_1.PC [10]);
  and (_28763_, _28762_, _42618_);
  and (_43256_, _28763_, _28761_);
  and (_28764_, _28465_, \oc8051_golden_model_1.PC [11]);
  nor (_28765_, _28465_, \oc8051_golden_model_1.PC [11]);
  nor (_28766_, _28765_, _28764_);
  or (_28767_, _28766_, _12151_);
  or (_28768_, _28766_, _12162_);
  or (_28769_, _28766_, _10979_);
  or (_28771_, _28766_, _12169_);
  or (_28772_, _12417_, _09030_);
  nor (_28773_, _12208_, _05982_);
  and (_28774_, _12333_, _12207_);
  nor (_28775_, _28475_, _12204_);
  and (_28776_, _28775_, _12211_);
  nor (_28777_, _28775_, _12211_);
  or (_28778_, _28777_, _28776_);
  and (_28779_, _28778_, _12335_);
  or (_28780_, _28779_, _12177_);
  or (_28782_, _28780_, _28774_);
  nand (_28783_, _12371_, _12208_);
  or (_28784_, _28778_, _12371_);
  and (_28785_, _28784_, _12379_);
  and (_28786_, _28785_, _28783_);
  and (_28787_, _12417_, _06464_);
  or (_28788_, _12545_, _12417_);
  or (_28789_, _12534_, _12207_);
  or (_28790_, _28778_, _12536_);
  and (_28791_, _28790_, _06341_);
  and (_28793_, _28791_, _28789_);
  or (_28794_, _12418_, _12419_);
  nand (_28795_, _28794_, _12490_);
  or (_28796_, _28794_, _12490_);
  and (_28797_, _28796_, _28795_);
  and (_28798_, _28797_, _25366_);
  or (_28799_, _28798_, _08654_);
  and (_28800_, _12507_, _12417_);
  or (_28801_, _28800_, _28799_);
  or (_28802_, _12517_, _12417_);
  nor (_28804_, _06781_, _07141_);
  nor (_28805_, _06758_, \oc8051_golden_model_1.PC [11]);
  nand (_28806_, _28805_, _28804_);
  or (_28807_, _28806_, _07486_);
  nand (_28808_, _28807_, _28802_);
  nand (_28809_, _28808_, _12512_);
  or (_28810_, _28766_, _12514_);
  and (_28811_, _28810_, _28809_);
  or (_28812_, _28811_, _12387_);
  and (_28813_, _28812_, _27157_);
  and (_28815_, _28813_, _28801_);
  or (_28816_, _28815_, _28793_);
  and (_28817_, _28816_, _12541_);
  and (_28818_, _28766_, _27163_);
  or (_28819_, _28818_, _12546_);
  or (_28820_, _28819_, _28817_);
  and (_28821_, _28820_, _28788_);
  or (_28822_, _28821_, _12551_);
  or (_28823_, _28766_, _12550_);
  and (_28824_, _28823_, _06465_);
  and (_28826_, _28824_, _28822_);
  or (_28827_, _28826_, _28787_);
  and (_28828_, _28827_, _12560_);
  and (_28829_, _28766_, _25401_);
  or (_28830_, _28829_, _12566_);
  or (_28831_, _28830_, _28828_);
  or (_28832_, _12565_, _12417_);
  and (_28833_, _28832_, _12378_);
  and (_28834_, _28833_, _28831_);
  or (_28835_, _28834_, _28786_);
  or (_28837_, _28835_, _06347_);
  and (_28838_, _28837_, _06774_);
  and (_28839_, _28838_, _28782_);
  and (_28840_, _28778_, _28542_);
  and (_28841_, _12587_, _12207_);
  or (_28842_, _28841_, _28840_);
  and (_28843_, _28842_, _06480_);
  or (_28844_, _28843_, _28839_);
  and (_28845_, _28844_, _12176_);
  or (_28846_, _28778_, _12604_);
  nand (_28848_, _12604_, _12208_);
  and (_28849_, _28848_, _06371_);
  and (_28850_, _28849_, _28846_);
  or (_28851_, _28850_, _28845_);
  and (_28852_, _28851_, _12175_);
  nand (_28853_, _28766_, _12174_);
  nand (_28854_, _28853_, _12623_);
  or (_28855_, _28854_, _28852_);
  or (_28856_, _12623_, _12417_);
  and (_28857_, _28856_, _12630_);
  and (_28859_, _28857_, _28855_);
  and (_28860_, _28766_, _12631_);
  or (_28861_, _28860_, _12636_);
  or (_28862_, _28861_, _28859_);
  or (_28863_, _12635_, _12417_);
  and (_28864_, _28863_, _12639_);
  and (_28865_, _28864_, _28862_);
  and (_28866_, _28766_, _26197_);
  or (_28867_, _28866_, _12644_);
  or (_28868_, _28867_, _28865_);
  or (_28870_, _12417_, _12643_);
  and (_28871_, _28870_, _05984_);
  and (_28872_, _28871_, _28868_);
  nand (_28873_, _28766_, _10515_);
  nand (_28874_, _28873_, _12652_);
  or (_28875_, _28874_, _28872_);
  or (_28876_, _12652_, _12417_);
  and (_28877_, _28876_, _06374_);
  and (_28878_, _28877_, _28875_);
  nand (_28879_, _12207_, _06373_);
  nand (_28881_, _28879_, _07216_);
  or (_28882_, _28881_, _28878_);
  or (_28883_, _12417_, _07216_);
  and (_28884_, _28883_, _05982_);
  and (_28885_, _28884_, _28882_);
  or (_28886_, _28885_, _28773_);
  and (_28887_, _28886_, _12172_);
  and (_28888_, _28766_, _25492_);
  or (_28889_, _28888_, _12670_);
  or (_28890_, _28889_, _28887_);
  or (_28892_, _12669_, _12417_);
  and (_28893_, _28892_, _12679_);
  and (_28894_, _28893_, _28890_);
  and (_28895_, _28797_, _12674_);
  or (_28896_, _28895_, _09031_);
  or (_28897_, _28896_, _28894_);
  and (_28898_, _28897_, _28772_);
  or (_28899_, _28898_, _06218_);
  and (_28900_, _12208_, _06218_);
  nor (_28901_, _28900_, _10929_);
  and (_28902_, _28901_, _28899_);
  and (_28903_, _12417_, _10929_);
  or (_28904_, _28903_, _28902_);
  and (_28905_, _28904_, _12691_);
  or (_28906_, _12720_, \oc8051_golden_model_1.DPH [3]);
  nor (_28907_, _12721_, _12691_);
  and (_28908_, _28907_, _28906_);
  or (_28909_, _28908_, _12730_);
  or (_28910_, _28909_, _28905_);
  or (_28911_, _12729_, _12417_);
  and (_28914_, _28911_, _25064_);
  and (_28915_, _28914_, _28910_);
  or (_28916_, _28797_, _11342_);
  or (_28917_, _12417_, _12759_);
  and (_28918_, _28917_, _12733_);
  and (_28919_, _28918_, _28916_);
  or (_28920_, _28919_, _12737_);
  or (_28921_, _28920_, _28915_);
  and (_28922_, _28921_, _28771_);
  or (_28923_, _28922_, _26610_);
  or (_28925_, _12417_, _12166_);
  and (_28926_, _28925_, _07237_);
  and (_28927_, _28926_, _28923_);
  nand (_28928_, _12207_, _06369_);
  nand (_28929_, _28928_, _12751_);
  or (_28930_, _28929_, _28927_);
  or (_28931_, _12751_, _12417_);
  and (_28932_, _28931_, _25061_);
  and (_28933_, _28932_, _28930_);
  or (_28934_, _28797_, _12759_);
  or (_28936_, _12417_, _11342_);
  and (_28937_, _28936_, _12755_);
  and (_28938_, _28937_, _28934_);
  or (_28939_, _28938_, _10980_);
  or (_28940_, _28939_, _28933_);
  and (_28941_, _28940_, _28769_);
  or (_28942_, _28941_, _26630_);
  or (_28943_, _12164_, _12417_);
  and (_28944_, _28943_, _07242_);
  and (_28945_, _28944_, _28942_);
  nand (_28947_, _12207_, _06375_);
  nand (_28948_, _28947_, _12772_);
  or (_28949_, _28948_, _28945_);
  or (_28950_, _12772_, _12417_);
  and (_28951_, _28950_, _12782_);
  and (_28952_, _28951_, _28949_);
  or (_28953_, _28797_, \oc8051_golden_model_1.PSW [7]);
  or (_28954_, _12417_, _10558_);
  and (_28955_, _28954_, _12776_);
  and (_28956_, _28955_, _28953_);
  or (_28958_, _28956_, _12780_);
  or (_28959_, _28958_, _28952_);
  and (_28960_, _28959_, _28768_);
  or (_28961_, _28960_, _11023_);
  or (_28962_, _12417_, _11022_);
  and (_28963_, _28962_, _09056_);
  and (_28964_, _28963_, _28961_);
  nand (_28965_, _12207_, _06366_);
  nand (_28966_, _28965_, _12796_);
  or (_28967_, _28966_, _28964_);
  or (_28969_, _12796_, _12417_);
  and (_28970_, _28969_, _25056_);
  and (_28971_, _28970_, _28967_);
  or (_28972_, _28797_, _10558_);
  or (_28973_, _12417_, \oc8051_golden_model_1.PSW [7]);
  and (_28974_, _28973_, _12800_);
  and (_28975_, _28974_, _28972_);
  or (_28976_, _28975_, _28971_);
  and (_28977_, _28976_, _12154_);
  and (_28978_, _28766_, _12804_);
  or (_28980_, _28978_, _14297_);
  or (_28981_, _28980_, _28977_);
  or (_28982_, _12417_, _12153_);
  and (_28983_, _28982_, _11126_);
  and (_28984_, _28983_, _28981_);
  and (_28985_, _28766_, _11125_);
  or (_28986_, _28985_, _06551_);
  or (_28987_, _28986_, _28984_);
  nand (_28988_, _07594_, _06551_);
  and (_28989_, _28988_, _28987_);
  or (_28991_, _28989_, _07253_);
  nor (_28992_, _12417_, _05959_);
  nor (_28993_, _28992_, _06365_);
  and (_28994_, _28993_, _28991_);
  or (_28995_, _28778_, _28701_);
  or (_28996_, _12207_, _13004_);
  and (_28997_, _28996_, _06365_);
  and (_28998_, _28997_, _28995_);
  or (_28999_, _28998_, _25625_);
  or (_29000_, _28999_, _28994_);
  and (_29002_, _29000_, _28767_);
  or (_29003_, _29002_, _19056_);
  or (_29004_, _13012_, _12417_);
  and (_29005_, _29004_, _11285_);
  and (_29006_, _29005_, _29003_);
  and (_29007_, _28766_, _11284_);
  or (_29008_, _29007_, _06281_);
  or (_29009_, _29008_, _29006_);
  nand (_29010_, _07594_, _06281_);
  and (_29011_, _29010_, _29009_);
  or (_29013_, _29011_, _25646_);
  nor (_29014_, _12417_, _05964_);
  nor (_29015_, _29014_, _06362_);
  and (_29016_, _29015_, _29013_);
  or (_29017_, _28778_, _13004_);
  nand (_29018_, _12208_, _13004_);
  and (_29019_, _29018_, _29017_);
  and (_29020_, _29019_, _06362_);
  or (_29021_, _29020_, _13031_);
  or (_29022_, _29021_, _29016_);
  or (_29024_, _28766_, _13030_);
  and (_29025_, _29024_, _06926_);
  and (_29026_, _29025_, _29022_);
  nand (_29027_, _12417_, _06568_);
  nand (_29028_, _29027_, _13037_);
  or (_29029_, _29028_, _29026_);
  or (_29030_, _28766_, _13037_);
  and (_29031_, _29030_, _14508_);
  and (_29032_, _29031_, _29029_);
  nor (_29033_, _14508_, _06213_);
  or (_29035_, _29033_, _05940_);
  or (_29036_, _29035_, _29032_);
  or (_29037_, _12417_, _14710_);
  and (_29038_, _29037_, _05928_);
  and (_29039_, _29038_, _29036_);
  and (_29040_, _29019_, _05927_);
  or (_29041_, _29040_, _13053_);
  or (_29042_, _29041_, _29039_);
  or (_29043_, _28766_, _13052_);
  and (_29044_, _29043_, _06279_);
  and (_29046_, _29044_, _29042_);
  nand (_29047_, _12417_, _06278_);
  nand (_29048_, _29047_, _12141_);
  or (_29049_, _29048_, _29046_);
  or (_29050_, _28766_, _12141_);
  and (_29051_, _29050_, _12140_);
  and (_29052_, _29051_, _29049_);
  nor (_29053_, _12140_, _06213_);
  or (_29054_, _29053_, _05939_);
  or (_29055_, _29054_, _29052_);
  not (_29057_, _13068_);
  not (_29058_, _05939_);
  or (_29059_, _12417_, _29058_);
  and (_29060_, _29059_, _29057_);
  and (_29061_, _29060_, _29055_);
  and (_29062_, _28766_, _13068_);
  or (_29063_, _29062_, _29061_);
  or (_29064_, _29063_, _01351_);
  or (_29065_, _01347_, \oc8051_golden_model_1.PC [11]);
  and (_29066_, _29065_, _42618_);
  and (_43257_, _29066_, _29064_);
  and (_29068_, _06968_, _06379_);
  or (_29069_, _29068_, _05939_);
  and (_29070_, _28764_, \oc8051_golden_model_1.PC [12]);
  nor (_29071_, _28764_, \oc8051_golden_model_1.PC [12]);
  nor (_29072_, _29071_, _29070_);
  not (_29073_, _29072_);
  and (_29074_, _29073_, _11284_);
  not (_29075_, _12414_);
  nor (_29076_, _12796_, _29075_);
  nor (_29078_, _12772_, _29075_);
  nor (_29079_, _12751_, _29075_);
  and (_29080_, _12291_, _12288_);
  nor (_29081_, _29080_, _12292_);
  or (_29082_, _29081_, _12333_);
  or (_29083_, _12335_, _12198_);
  and (_29084_, _29083_, _06347_);
  nand (_29085_, _29084_, _29082_);
  nand (_29086_, _12371_, _12198_);
  not (_29087_, _29081_);
  or (_29089_, _29087_, _12371_);
  and (_29090_, _29089_, _12379_);
  and (_29091_, _29090_, _29086_);
  or (_29092_, _29087_, _12536_);
  or (_29093_, _12534_, _12199_);
  nand (_29094_, _29093_, _29092_);
  nand (_29095_, _29094_, _06341_);
  and (_29096_, _12507_, _12414_);
  nor (_29097_, _12494_, _12492_);
  nor (_29098_, _29097_, _12495_);
  and (_29100_, _29098_, _12393_);
  nor (_29101_, _29100_, _29096_);
  nand (_29102_, _29101_, _12387_);
  nor (_29103_, _29073_, _12514_);
  not (_29104_, _29103_);
  nor (_29105_, _12517_, _29075_);
  and (_29106_, _28804_, _07504_);
  and (_29107_, _07487_, \oc8051_golden_model_1.PC [12]);
  and (_29108_, _29107_, _29106_);
  nor (_29109_, _29108_, _29105_);
  nor (_29111_, _29109_, _12516_);
  nor (_29112_, _29111_, _12387_);
  and (_29113_, _29112_, _29104_);
  not (_29114_, _29113_);
  and (_29115_, _29114_, _27157_);
  nand (_29116_, _29115_, _29102_);
  nand (_29117_, _29116_, _29095_);
  and (_29118_, _29117_, _12541_);
  and (_29119_, _29072_, _27163_);
  or (_29120_, _29119_, _12546_);
  or (_29122_, _29120_, _29118_);
  nor (_29123_, _12545_, _12414_);
  nor (_29124_, _29123_, _12551_);
  and (_29125_, _29124_, _29122_);
  nor (_29126_, _29073_, _12550_);
  or (_29127_, _29126_, _06464_);
  nor (_29128_, _29127_, _29125_);
  and (_29129_, _29075_, _06464_);
  or (_29130_, _29129_, _29128_);
  nand (_29131_, _29130_, _12560_);
  nor (_29133_, _29072_, _12560_);
  nor (_29134_, _29133_, _12566_);
  and (_29135_, _29134_, _29131_);
  nor (_29136_, _12565_, _29075_);
  or (_29137_, _29136_, _12379_);
  nor (_29138_, _29137_, _29135_);
  or (_29139_, _29138_, _06347_);
  or (_29140_, _29139_, _29091_);
  and (_29141_, _29140_, _29085_);
  nand (_29142_, _29141_, _06774_);
  nor (_29144_, _29087_, _12587_);
  and (_29145_, _12587_, _12198_);
  or (_29146_, _29145_, _29144_);
  nor (_29147_, _29146_, _06774_);
  nor (_29148_, _29147_, _06371_);
  nand (_29149_, _29148_, _29142_);
  and (_29150_, _12604_, _12198_);
  and (_29151_, _29081_, _26518_);
  or (_29152_, _29151_, _29150_);
  and (_29153_, _29152_, _06371_);
  nor (_29155_, _29153_, _12174_);
  and (_29156_, _29155_, _29149_);
  and (_29157_, _29073_, _12174_);
  or (_29158_, _29157_, _29156_);
  and (_29159_, _29158_, _12623_);
  nor (_29160_, _12623_, _12414_);
  or (_29161_, _29160_, _29159_);
  nand (_29162_, _29161_, _12630_);
  nor (_29163_, _29072_, _12630_);
  nor (_29164_, _29163_, _12636_);
  nand (_29166_, _29164_, _29162_);
  nor (_29167_, _12635_, _29075_);
  nor (_29168_, _29167_, _26197_);
  nand (_29169_, _29168_, _29166_);
  nor (_29170_, _29072_, _12639_);
  nor (_29171_, _29170_, _12644_);
  nand (_29172_, _29171_, _29169_);
  nor (_29173_, _29075_, _12643_);
  nor (_29174_, _29173_, _10515_);
  nand (_29175_, _29174_, _29172_);
  nor (_29177_, _29072_, _05984_);
  nor (_29178_, _29177_, _12653_);
  nand (_29179_, _29178_, _29175_);
  nor (_29180_, _12652_, _29075_);
  nor (_29181_, _29180_, _06373_);
  nand (_29182_, _29181_, _29179_);
  and (_29183_, _12199_, _06373_);
  nor (_29184_, _29183_, _12659_);
  nand (_29185_, _29184_, _29182_);
  nor (_29186_, _29075_, _07216_);
  nor (_29188_, _29186_, _10094_);
  nand (_29189_, _29188_, _29185_);
  nor (_29190_, _12198_, _05982_);
  nor (_29191_, _29190_, _25492_);
  nand (_29192_, _29191_, _29189_);
  nor (_29193_, _29073_, _12172_);
  nor (_29194_, _29193_, _12670_);
  nand (_29195_, _29194_, _29192_);
  nor (_29196_, _12669_, _12414_);
  nor (_29197_, _29196_, _12674_);
  and (_29199_, _29197_, _29195_);
  and (_29200_, _29098_, _12674_);
  nor (_29201_, _29200_, _29199_);
  or (_29202_, _29201_, _09031_);
  or (_29203_, _29075_, _09030_);
  and (_29204_, _29203_, _06219_);
  nand (_29205_, _29204_, _29202_);
  and (_29206_, _12199_, _06218_);
  nor (_29207_, _29206_, _10929_);
  nand (_29208_, _29207_, _29205_);
  and (_29210_, _12414_, _10929_);
  nor (_29211_, _29210_, _12690_);
  and (_29212_, _29211_, _29208_);
  nor (_29213_, _12721_, \oc8051_golden_model_1.DPH [4]);
  nor (_29214_, _29213_, _12722_);
  nor (_29215_, _29214_, _12691_);
  or (_29216_, _29215_, _29212_);
  nand (_29217_, _29216_, _12729_);
  nor (_29218_, _12729_, _12414_);
  nor (_29219_, _29218_, _12733_);
  nand (_29221_, _29219_, _29217_);
  nor (_29222_, _29098_, _11342_);
  nor (_29223_, _12414_, _12759_);
  nor (_29224_, _29223_, _25064_);
  not (_29225_, _29224_);
  nor (_29226_, _29225_, _29222_);
  nor (_29227_, _29226_, _12737_);
  nand (_29228_, _29227_, _29221_);
  nor (_29229_, _29072_, _12169_);
  nor (_29230_, _29229_, _26610_);
  nand (_29232_, _29230_, _29228_);
  nor (_29233_, _29075_, _12166_);
  nor (_29234_, _29233_, _06369_);
  nand (_29235_, _29234_, _29232_);
  and (_29236_, _12199_, _06369_);
  nor (_29237_, _29236_, _12752_);
  and (_29238_, _29237_, _29235_);
  or (_29239_, _29238_, _29079_);
  nand (_29240_, _29239_, _25061_);
  and (_29241_, _12414_, _12759_);
  and (_29243_, _29098_, _11342_);
  or (_29244_, _29243_, _29241_);
  and (_29245_, _29244_, _12755_);
  nor (_29246_, _29245_, _10980_);
  nand (_29247_, _29246_, _29240_);
  nor (_29248_, _29072_, _10979_);
  nor (_29249_, _29248_, _26630_);
  nand (_29250_, _29249_, _29247_);
  nor (_29251_, _12164_, _29075_);
  nor (_29252_, _29251_, _06375_);
  nand (_29254_, _29252_, _29250_);
  and (_29255_, _12199_, _06375_);
  nor (_29256_, _29255_, _12773_);
  and (_29257_, _29256_, _29254_);
  or (_29258_, _29257_, _29078_);
  nand (_29259_, _29258_, _12782_);
  and (_29260_, _12414_, \oc8051_golden_model_1.PSW [7]);
  and (_29261_, _29098_, _10558_);
  or (_29262_, _29261_, _29260_);
  and (_29263_, _29262_, _12776_);
  nor (_29265_, _29263_, _12780_);
  nand (_29266_, _29265_, _29259_);
  nor (_29267_, _29072_, _12162_);
  nor (_29268_, _29267_, _11023_);
  nand (_29269_, _29268_, _29266_);
  nor (_29270_, _29075_, _11022_);
  nor (_29271_, _29270_, _06366_);
  nand (_29272_, _29271_, _29269_);
  and (_29273_, _12199_, _06366_);
  nor (_29274_, _29273_, _12797_);
  and (_29276_, _29274_, _29272_);
  or (_29277_, _29276_, _29076_);
  nand (_29278_, _29277_, _25056_);
  and (_29279_, _12414_, _10558_);
  and (_29280_, _29098_, \oc8051_golden_model_1.PSW [7]);
  or (_29281_, _29280_, _29279_);
  and (_29282_, _29281_, _12800_);
  nor (_29283_, _29282_, _12804_);
  nand (_29284_, _29283_, _29278_);
  nor (_29285_, _29072_, _12154_);
  nor (_29287_, _29285_, _14297_);
  nand (_29288_, _29287_, _29284_);
  nor (_29289_, _29075_, _12153_);
  nor (_29290_, _29289_, _11125_);
  nand (_29291_, _29290_, _29288_);
  and (_29292_, _29073_, _11125_);
  nor (_29293_, _29292_, _06551_);
  and (_29294_, _29293_, _29291_);
  nor (_29295_, _08541_, _06716_);
  or (_29296_, _29295_, _07253_);
  or (_29298_, _29296_, _29294_);
  nor (_29299_, _12414_, _05959_);
  nor (_29300_, _29299_, _06365_);
  nand (_29301_, _29300_, _29298_);
  and (_29302_, _29087_, _13004_);
  nor (_29303_, _12198_, _13004_);
  or (_29304_, _29303_, _06558_);
  or (_29305_, _29304_, _29302_);
  and (_29306_, _29305_, _12151_);
  nand (_29307_, _29306_, _29301_);
  nor (_29309_, _29072_, _12151_);
  nor (_29310_, _29309_, _19056_);
  nand (_29311_, _29310_, _29307_);
  nor (_29312_, _13012_, _29075_);
  nor (_29313_, _29312_, _11284_);
  and (_29314_, _29313_, _29311_);
  or (_29315_, _29314_, _29074_);
  nand (_29316_, _29315_, _06282_);
  and (_29317_, _08541_, _06281_);
  nor (_29318_, _29317_, _25646_);
  and (_29320_, _29318_, _29316_);
  nor (_29321_, _29075_, _05964_);
  or (_29322_, _29321_, _06362_);
  nor (_29323_, _29322_, _29320_);
  nor (_29324_, _29081_, _13004_);
  and (_29325_, _12199_, _13004_);
  nor (_29326_, _29325_, _29324_);
  nor (_29327_, _29326_, _06921_);
  or (_29328_, _29327_, _29323_);
  and (_29329_, _29328_, _13030_);
  nor (_29331_, _29072_, _13030_);
  or (_29332_, _29331_, _29329_);
  nand (_29333_, _29332_, _06926_);
  and (_29334_, _29075_, _06568_);
  nor (_29335_, _29334_, _13038_);
  nand (_29336_, _29335_, _29333_);
  nor (_29337_, _29073_, _13037_);
  nor (_29338_, _29337_, _06361_);
  nand (_29339_, _29338_, _29336_);
  and (_29340_, _06968_, _06361_);
  nor (_29342_, _29340_, _05940_);
  nand (_29343_, _29342_, _29339_);
  and (_29344_, _12414_, _05940_);
  nor (_29345_, _29344_, _05927_);
  nand (_29346_, _29345_, _29343_);
  nor (_29347_, _29326_, _05928_);
  nor (_29348_, _29347_, _13053_);
  nand (_29349_, _29348_, _29346_);
  nor (_29350_, _29073_, _13052_);
  nor (_29351_, _29350_, _06278_);
  nand (_29353_, _29351_, _29349_);
  and (_29354_, _29075_, _06278_);
  nor (_29355_, _29354_, _13059_);
  nand (_29356_, _29355_, _29353_);
  nor (_29357_, _29073_, _12141_);
  nor (_29358_, _29357_, _06379_);
  and (_29359_, _29358_, _29356_);
  or (_29360_, _29359_, _29069_);
  and (_29361_, _12414_, _05939_);
  nor (_29362_, _29361_, _13068_);
  and (_29364_, _29362_, _29360_);
  and (_29365_, _29073_, _13068_);
  nor (_29366_, _29365_, _29364_);
  or (_29367_, _29366_, _01351_);
  or (_29368_, _01347_, \oc8051_golden_model_1.PC [12]);
  and (_29369_, _29368_, _42618_);
  and (_43258_, _29369_, _29367_);
  and (_29370_, _29070_, \oc8051_golden_model_1.PC [13]);
  nor (_29371_, _29070_, \oc8051_golden_model_1.PC [13]);
  nor (_29372_, _29371_, _29370_);
  or (_29374_, _29372_, _12151_);
  or (_29375_, _29372_, _12154_);
  or (_29376_, _29372_, _12162_);
  or (_29377_, _29372_, _10979_);
  or (_29378_, _29372_, _12169_);
  or (_29379_, _12409_, _09030_);
  nor (_29380_, _12194_, _05982_);
  or (_29381_, _12196_, _12195_);
  not (_29382_, _29381_);
  nor (_29383_, _29382_, _12293_);
  and (_29385_, _29382_, _12293_);
  or (_29386_, _29385_, _29383_);
  or (_29387_, _29386_, _12587_);
  nand (_29388_, _12587_, _12194_);
  and (_29389_, _29388_, _06480_);
  and (_29390_, _29389_, _29387_);
  and (_29391_, _12333_, _12193_);
  and (_29392_, _29386_, _12335_);
  or (_29393_, _29392_, _12177_);
  or (_29394_, _29393_, _29391_);
  nand (_29396_, _12371_, _12194_);
  or (_29397_, _29386_, _12371_);
  and (_29398_, _29397_, _12379_);
  and (_29399_, _29398_, _29396_);
  and (_29400_, _12409_, _06464_);
  or (_29401_, _12545_, _12409_);
  or (_29402_, _29386_, _12536_);
  or (_29403_, _12534_, _12193_);
  and (_29404_, _29403_, _06341_);
  and (_29405_, _29404_, _29402_);
  or (_29407_, _12410_, _12411_);
  not (_29408_, _29407_);
  nor (_29409_, _29408_, _12496_);
  and (_29410_, _29408_, _12496_);
  or (_29411_, _29410_, _29409_);
  and (_29412_, _29411_, _25366_);
  or (_29413_, _29412_, _08654_);
  and (_29414_, _12507_, _12409_);
  or (_29415_, _29414_, _29413_);
  or (_29416_, _29372_, _12514_);
  or (_29418_, _12517_, _12409_);
  nor (_29419_, _07486_, \oc8051_golden_model_1.PC [13]);
  nand (_29420_, _29419_, _29106_);
  and (_29421_, _29420_, _29418_);
  or (_29422_, _29421_, _12516_);
  and (_29423_, _29422_, _29416_);
  or (_29424_, _29423_, _12387_);
  and (_29425_, _29424_, _27157_);
  and (_29426_, _29425_, _29415_);
  or (_29427_, _29426_, _29405_);
  and (_29428_, _29427_, _12541_);
  and (_29429_, _29372_, _27163_);
  or (_29430_, _29429_, _12546_);
  or (_29431_, _29430_, _29428_);
  and (_29432_, _29431_, _29401_);
  or (_29433_, _29432_, _12551_);
  or (_29434_, _29372_, _12550_);
  and (_29435_, _29434_, _06465_);
  and (_29436_, _29435_, _29433_);
  or (_29437_, _29436_, _29400_);
  and (_29440_, _29437_, _12560_);
  and (_29441_, _29372_, _25401_);
  or (_29442_, _29441_, _12566_);
  or (_29443_, _29442_, _29440_);
  or (_29444_, _12565_, _12409_);
  and (_29445_, _29444_, _12378_);
  and (_29446_, _29445_, _29443_);
  or (_29447_, _29446_, _29399_);
  or (_29448_, _29447_, _06347_);
  and (_29449_, _29448_, _06774_);
  and (_29451_, _29449_, _29394_);
  or (_29452_, _29451_, _29390_);
  and (_29453_, _29452_, _12176_);
  or (_29454_, _29386_, _12604_);
  nand (_29455_, _12604_, _12194_);
  and (_29456_, _29455_, _06371_);
  and (_29457_, _29456_, _29454_);
  or (_29458_, _29457_, _29453_);
  and (_29459_, _29458_, _12175_);
  nand (_29460_, _29372_, _12174_);
  nand (_29462_, _29460_, _12623_);
  or (_29463_, _29462_, _29459_);
  or (_29464_, _12623_, _12409_);
  and (_29465_, _29464_, _12630_);
  and (_29466_, _29465_, _29463_);
  and (_29467_, _29372_, _12631_);
  or (_29468_, _29467_, _12636_);
  or (_29469_, _29468_, _29466_);
  or (_29470_, _12635_, _12409_);
  and (_29471_, _29470_, _12639_);
  and (_29473_, _29471_, _29469_);
  and (_29474_, _29372_, _26197_);
  or (_29475_, _29474_, _12644_);
  or (_29476_, _29475_, _29473_);
  or (_29477_, _12409_, _12643_);
  and (_29478_, _29477_, _05984_);
  and (_29479_, _29478_, _29476_);
  nand (_29480_, _29372_, _10515_);
  nand (_29481_, _29480_, _12652_);
  or (_29482_, _29481_, _29479_);
  or (_29484_, _12652_, _12409_);
  and (_29485_, _29484_, _06374_);
  and (_29486_, _29485_, _29482_);
  nand (_29487_, _12193_, _06373_);
  nand (_29488_, _29487_, _07216_);
  or (_29489_, _29488_, _29486_);
  or (_29490_, _12409_, _07216_);
  and (_29491_, _29490_, _05982_);
  and (_29492_, _29491_, _29489_);
  or (_29493_, _29492_, _29380_);
  and (_29495_, _29493_, _12172_);
  and (_29496_, _29372_, _25492_);
  or (_29497_, _29496_, _12670_);
  or (_29498_, _29497_, _29495_);
  or (_29499_, _12669_, _12409_);
  and (_29500_, _29499_, _12679_);
  and (_29501_, _29500_, _29498_);
  and (_29502_, _29411_, _12674_);
  or (_29503_, _29502_, _09031_);
  or (_29504_, _29503_, _29501_);
  and (_29506_, _29504_, _29379_);
  or (_29507_, _29506_, _06218_);
  and (_29508_, _12194_, _06218_);
  nor (_29509_, _29508_, _10929_);
  and (_29510_, _29509_, _29507_);
  and (_29511_, _12409_, _10929_);
  or (_29512_, _29511_, _29510_);
  and (_29513_, _29512_, _12691_);
  or (_29514_, _12722_, \oc8051_golden_model_1.DPH [5]);
  nor (_29515_, _12723_, _12691_);
  and (_29517_, _29515_, _29514_);
  or (_29518_, _29517_, _12730_);
  or (_29519_, _29518_, _29513_);
  or (_29520_, _12729_, _12409_);
  and (_29521_, _29520_, _25064_);
  and (_29522_, _29521_, _29519_);
  or (_29523_, _29411_, _11342_);
  or (_29524_, _12409_, _12759_);
  and (_29525_, _29524_, _12733_);
  and (_29526_, _29525_, _29523_);
  or (_29528_, _29526_, _12737_);
  or (_29529_, _29528_, _29522_);
  and (_29530_, _29529_, _29378_);
  or (_29531_, _29530_, _26610_);
  or (_29532_, _12409_, _12166_);
  and (_29533_, _29532_, _07237_);
  and (_29534_, _29533_, _29531_);
  nand (_29535_, _12193_, _06369_);
  nand (_29536_, _29535_, _12751_);
  or (_29537_, _29536_, _29534_);
  or (_29539_, _12751_, _12409_);
  and (_29540_, _29539_, _25061_);
  and (_29541_, _29540_, _29537_);
  or (_29542_, _29411_, _12759_);
  or (_29543_, _12409_, _11342_);
  and (_29544_, _29543_, _12755_);
  and (_29545_, _29544_, _29542_);
  or (_29546_, _29545_, _10980_);
  or (_29547_, _29546_, _29541_);
  and (_29548_, _29547_, _29377_);
  or (_29550_, _29548_, _26630_);
  or (_29551_, _12164_, _12409_);
  and (_29552_, _29551_, _07242_);
  and (_29553_, _29552_, _29550_);
  nand (_29554_, _12193_, _06375_);
  nand (_29555_, _29554_, _12772_);
  or (_29556_, _29555_, _29553_);
  or (_29557_, _12772_, _12409_);
  and (_29558_, _29557_, _12782_);
  and (_29559_, _29558_, _29556_);
  or (_29561_, _29411_, \oc8051_golden_model_1.PSW [7]);
  or (_29562_, _12409_, _10558_);
  and (_29563_, _29562_, _12776_);
  and (_29564_, _29563_, _29561_);
  or (_29565_, _29564_, _12780_);
  or (_29566_, _29565_, _29559_);
  and (_29567_, _29566_, _29376_);
  or (_29568_, _29567_, _11023_);
  or (_29569_, _12409_, _11022_);
  and (_29570_, _29569_, _09056_);
  and (_29572_, _29570_, _29568_);
  nand (_29573_, _12193_, _06366_);
  nand (_29574_, _29573_, _12796_);
  or (_29575_, _29574_, _29572_);
  or (_29576_, _12796_, _12409_);
  and (_29577_, _29576_, _25056_);
  and (_29578_, _29577_, _29575_);
  or (_29579_, _29411_, _10558_);
  or (_29580_, _12409_, \oc8051_golden_model_1.PSW [7]);
  and (_29581_, _29580_, _12800_);
  and (_29583_, _29581_, _29579_);
  or (_29584_, _29583_, _12804_);
  or (_29585_, _29584_, _29578_);
  and (_29586_, _29585_, _29375_);
  or (_29587_, _29586_, _14297_);
  or (_29588_, _12409_, _12153_);
  and (_29589_, _29588_, _11126_);
  and (_29590_, _29589_, _29587_);
  and (_29591_, _29372_, _11125_);
  or (_29592_, _29591_, _06551_);
  or (_29594_, _29592_, _29590_);
  nand (_29595_, _08244_, _06551_);
  and (_29596_, _29595_, _29594_);
  or (_29597_, _29596_, _07253_);
  nor (_29598_, _12409_, _05959_);
  nor (_29599_, _29598_, _06365_);
  and (_29600_, _29599_, _29597_);
  or (_29601_, _29386_, _28701_);
  or (_29602_, _12193_, _13004_);
  and (_29603_, _29602_, _06365_);
  and (_29605_, _29603_, _29601_);
  or (_29606_, _29605_, _25625_);
  or (_29607_, _29606_, _29600_);
  and (_29608_, _29607_, _29374_);
  or (_29609_, _29608_, _19056_);
  or (_29610_, _13012_, _12409_);
  and (_29611_, _29610_, _11285_);
  and (_29612_, _29611_, _29609_);
  and (_29613_, _29372_, _11284_);
  or (_29614_, _29613_, _06281_);
  or (_29616_, _29614_, _29612_);
  nand (_29617_, _08244_, _06281_);
  and (_29618_, _29617_, _29616_);
  or (_29619_, _29618_, _25646_);
  nor (_29620_, _12409_, _05964_);
  nor (_29621_, _29620_, _06362_);
  and (_29622_, _29621_, _29619_);
  or (_29623_, _29386_, _13004_);
  nand (_29624_, _12194_, _13004_);
  and (_29625_, _29624_, _29623_);
  and (_29627_, _29625_, _06362_);
  or (_29628_, _29627_, _13031_);
  or (_29629_, _29628_, _29622_);
  or (_29630_, _29372_, _13030_);
  and (_29631_, _29630_, _06926_);
  and (_29632_, _29631_, _29629_);
  nand (_29633_, _12409_, _06568_);
  nand (_29634_, _29633_, _13037_);
  or (_29635_, _29634_, _29632_);
  or (_29636_, _29372_, _13037_);
  and (_29638_, _29636_, _14508_);
  and (_29639_, _29638_, _29635_);
  nor (_29640_, _06611_, _14508_);
  or (_29641_, _29640_, _05940_);
  or (_29642_, _29641_, _29639_);
  or (_29643_, _12409_, _14710_);
  and (_29644_, _29643_, _05928_);
  and (_29645_, _29644_, _29642_);
  and (_29646_, _29625_, _05927_);
  or (_29647_, _29646_, _13053_);
  or (_29649_, _29647_, _29645_);
  or (_29650_, _29372_, _13052_);
  and (_29651_, _29650_, _06279_);
  and (_29652_, _29651_, _29649_);
  nand (_29653_, _12409_, _06278_);
  nand (_29654_, _29653_, _12141_);
  or (_29655_, _29654_, _29652_);
  or (_29656_, _29372_, _12141_);
  and (_29657_, _29656_, _12140_);
  and (_29658_, _29657_, _29655_);
  nor (_29660_, _06611_, _12140_);
  or (_29661_, _29660_, _05939_);
  or (_29662_, _29661_, _29658_);
  or (_29663_, _12409_, _29058_);
  and (_29664_, _29663_, _29057_);
  and (_29665_, _29664_, _29662_);
  and (_29666_, _29372_, _13068_);
  or (_29667_, _29666_, _29665_);
  or (_29668_, _29667_, _01351_);
  or (_29669_, _01347_, \oc8051_golden_model_1.PC [13]);
  and (_29671_, _29669_, _42618_);
  and (_43260_, _29671_, _29668_);
  and (_29672_, _29370_, \oc8051_golden_model_1.PC [14]);
  nor (_29673_, _29370_, \oc8051_golden_model_1.PC [14]);
  nor (_29674_, _29673_, _29672_);
  nor (_29675_, _29674_, _11285_);
  not (_29676_, _12403_);
  nor (_29677_, _12796_, _29676_);
  nor (_29678_, _12772_, _29676_);
  nor (_29679_, _12751_, _29676_);
  nor (_29681_, _12729_, _29676_);
  and (_29682_, _12295_, _12191_);
  nor (_29683_, _29682_, _12296_);
  not (_29684_, _29683_);
  nand (_29685_, _29684_, _12335_);
  or (_29686_, _12335_, _12186_);
  and (_29687_, _29686_, _06347_);
  nand (_29688_, _29687_, _29685_);
  not (_29689_, _29674_);
  nor (_29690_, _29689_, _12560_);
  nor (_29692_, _29674_, _12550_);
  or (_29693_, _29683_, _12536_);
  or (_29694_, _12534_, _12186_);
  and (_29695_, _29694_, _29693_);
  nor (_29696_, _29695_, _07151_);
  or (_29697_, _12393_, _29676_);
  and (_29698_, _12498_, _12407_);
  nor (_29699_, _29698_, _12499_);
  nand (_29700_, _29699_, _25366_);
  and (_29701_, _29700_, _12387_);
  nand (_29702_, _29701_, _29697_);
  nor (_29703_, _29689_, _12514_);
  not (_29704_, _29703_);
  nor (_29705_, _12517_, _29676_);
  and (_29706_, _07487_, \oc8051_golden_model_1.PC [14]);
  and (_29707_, _29706_, _29106_);
  nor (_29708_, _29707_, _29705_);
  nor (_29709_, _29708_, _12516_);
  nor (_29710_, _29709_, _12387_);
  and (_29711_, _29710_, _29704_);
  nor (_29714_, _29711_, _07154_);
  nand (_29715_, _29714_, _29702_);
  and (_29716_, _29674_, _07154_);
  nor (_29717_, _29716_, _06341_);
  and (_29718_, _29717_, _29715_);
  or (_29719_, _29718_, _29696_);
  nand (_29720_, _29719_, _12541_);
  nor (_29721_, _29674_, _12541_);
  nor (_29722_, _29721_, _12546_);
  and (_29723_, _29722_, _29720_);
  nor (_29725_, _12545_, _29676_);
  nor (_29726_, _29725_, _29723_);
  and (_29727_, _29726_, _12550_);
  or (_29728_, _29727_, _29692_);
  nand (_29729_, _29728_, _06465_);
  nor (_29730_, _12403_, _06465_);
  nor (_29731_, _29730_, _25401_);
  and (_29732_, _29731_, _29729_);
  or (_29733_, _29732_, _29690_);
  nand (_29734_, _29733_, _12565_);
  nor (_29736_, _12565_, _29676_);
  nor (_29737_, _29736_, _12379_);
  and (_29738_, _29737_, _29734_);
  and (_29739_, _12371_, _12186_);
  nor (_29740_, _29684_, _12371_);
  or (_29741_, _29740_, _12378_);
  nor (_29742_, _29741_, _29739_);
  or (_29743_, _29742_, _06347_);
  or (_29744_, _29743_, _29738_);
  and (_29745_, _29744_, _29688_);
  nand (_29747_, _29745_, _06774_);
  and (_29748_, _12587_, _12186_);
  nor (_29749_, _29684_, _12587_);
  or (_29750_, _29749_, _29748_);
  nor (_29751_, _29750_, _06774_);
  nor (_29752_, _29751_, _06371_);
  nand (_29753_, _29752_, _29747_);
  and (_29754_, _12604_, _12186_);
  and (_29755_, _29683_, _26518_);
  or (_29756_, _29755_, _29754_);
  and (_29758_, _29756_, _06371_);
  nor (_29759_, _29758_, _12174_);
  and (_29760_, _29759_, _29753_);
  nor (_29761_, _29674_, _12175_);
  or (_29762_, _29761_, _29760_);
  and (_29763_, _29762_, _12623_);
  nor (_29764_, _12623_, _12403_);
  or (_29765_, _29764_, _29763_);
  nand (_29766_, _29765_, _12630_);
  nor (_29767_, _29674_, _12630_);
  nor (_29769_, _29767_, _12636_);
  nand (_29770_, _29769_, _29766_);
  nor (_29771_, _12635_, _29676_);
  nor (_29772_, _29771_, _26197_);
  nand (_29773_, _29772_, _29770_);
  nor (_29774_, _29674_, _12639_);
  nor (_29775_, _29774_, _12644_);
  nand (_29776_, _29775_, _29773_);
  nor (_29777_, _29676_, _12643_);
  nor (_29778_, _29777_, _10515_);
  nand (_29780_, _29778_, _29776_);
  nor (_29781_, _29674_, _05984_);
  nor (_29782_, _29781_, _12653_);
  nand (_29783_, _29782_, _29780_);
  nor (_29784_, _12652_, _29676_);
  nor (_29785_, _29784_, _06373_);
  nand (_29786_, _29785_, _29783_);
  nor (_29787_, _12186_, _06374_);
  nor (_29788_, _29787_, _12659_);
  nand (_29789_, _29788_, _29786_);
  nor (_29791_, _29676_, _07216_);
  nor (_29792_, _29791_, _10094_);
  nand (_29793_, _29792_, _29789_);
  nor (_29794_, _12186_, _05982_);
  nor (_29795_, _29794_, _25492_);
  nand (_29796_, _29795_, _29793_);
  nor (_29797_, _29689_, _12172_);
  nor (_29798_, _29797_, _12670_);
  nand (_29799_, _29798_, _29796_);
  nor (_29800_, _12669_, _12403_);
  nor (_29802_, _29800_, _12674_);
  and (_29803_, _29802_, _29799_);
  and (_29804_, _29699_, _12674_);
  nor (_29805_, _29804_, _29803_);
  or (_29806_, _29805_, _09031_);
  or (_29807_, _29676_, _09030_);
  and (_29808_, _29807_, _06219_);
  nand (_29809_, _29808_, _29806_);
  nor (_29810_, _12186_, _06219_);
  nor (_29811_, _29810_, _10929_);
  nand (_29813_, _29811_, _29809_);
  and (_29814_, _12403_, _10929_);
  nor (_29815_, _29814_, _12690_);
  nand (_29816_, _29815_, _29813_);
  nor (_29817_, _12723_, \oc8051_golden_model_1.DPH [6]);
  nor (_29818_, _29817_, _12724_);
  nor (_29819_, _29818_, _12691_);
  nor (_29820_, _29819_, _12730_);
  and (_29821_, _29820_, _29816_);
  or (_29822_, _29821_, _29681_);
  nand (_29824_, _29822_, _25064_);
  and (_29825_, _12403_, _11342_);
  and (_29826_, _29699_, _12759_);
  or (_29827_, _29826_, _29825_);
  and (_29828_, _29827_, _12733_);
  nor (_29829_, _29828_, _12737_);
  nand (_29830_, _29829_, _29824_);
  nor (_29831_, _29674_, _12169_);
  nor (_29832_, _29831_, _26610_);
  nand (_29833_, _29832_, _29830_);
  nor (_29835_, _29676_, _12166_);
  nor (_29836_, _29835_, _06369_);
  nand (_29837_, _29836_, _29833_);
  nor (_29838_, _12186_, _07237_);
  nor (_29839_, _29838_, _12752_);
  and (_29840_, _29839_, _29837_);
  or (_29841_, _29840_, _29679_);
  nand (_29842_, _29841_, _25061_);
  and (_29843_, _12403_, _12759_);
  and (_29844_, _29699_, _11342_);
  or (_29846_, _29844_, _29843_);
  and (_29847_, _29846_, _12755_);
  nor (_29848_, _29847_, _10980_);
  nand (_29849_, _29848_, _29842_);
  nor (_29850_, _29674_, _10979_);
  nor (_29851_, _29850_, _26630_);
  nand (_29852_, _29851_, _29849_);
  nor (_29853_, _12164_, _29676_);
  nor (_29854_, _29853_, _06375_);
  nand (_29855_, _29854_, _29852_);
  nor (_29857_, _12186_, _07242_);
  nor (_29858_, _29857_, _12773_);
  and (_29859_, _29858_, _29855_);
  or (_29860_, _29859_, _29678_);
  nand (_29861_, _29860_, _12782_);
  and (_29862_, _12403_, \oc8051_golden_model_1.PSW [7]);
  and (_29863_, _29699_, _10558_);
  or (_29864_, _29863_, _29862_);
  and (_29865_, _29864_, _12776_);
  nor (_29866_, _29865_, _12780_);
  nand (_29868_, _29866_, _29861_);
  nor (_29869_, _29674_, _12162_);
  nor (_29870_, _29869_, _11023_);
  nand (_29871_, _29870_, _29868_);
  nor (_29872_, _29676_, _11022_);
  nor (_29873_, _29872_, _06366_);
  nand (_29874_, _29873_, _29871_);
  nor (_29875_, _12186_, _09056_);
  nor (_29876_, _29875_, _12797_);
  and (_29877_, _29876_, _29874_);
  or (_29879_, _29877_, _29677_);
  nand (_29880_, _29879_, _25056_);
  and (_29881_, _12403_, _10558_);
  and (_29882_, _29699_, \oc8051_golden_model_1.PSW [7]);
  or (_29883_, _29882_, _29881_);
  and (_29884_, _29883_, _12800_);
  nor (_29885_, _29884_, _12804_);
  nand (_29886_, _29885_, _29880_);
  nor (_29887_, _29674_, _12154_);
  nor (_29888_, _29887_, _14297_);
  nand (_29890_, _29888_, _29886_);
  nor (_29891_, _29676_, _12153_);
  nor (_29892_, _29891_, _11125_);
  nand (_29893_, _29892_, _29890_);
  nor (_29894_, _29674_, _11126_);
  nor (_29895_, _29894_, _06551_);
  nand (_29896_, _29895_, _29893_);
  nor (_29897_, _08142_, _06716_);
  nor (_29898_, _29897_, _07253_);
  nand (_29899_, _29898_, _29896_);
  nor (_29901_, _12403_, _05959_);
  nor (_29902_, _29901_, _06365_);
  nand (_29903_, _29902_, _29899_);
  and (_29904_, _29684_, _13004_);
  nor (_29905_, _12186_, _13004_);
  or (_29906_, _29905_, _06558_);
  or (_29907_, _29906_, _29904_);
  and (_29908_, _29907_, _12151_);
  nand (_29909_, _29908_, _29903_);
  nor (_29910_, _29674_, _12151_);
  nor (_29912_, _29910_, _19056_);
  nand (_29913_, _29912_, _29909_);
  nor (_29914_, _13012_, _29676_);
  nor (_29915_, _29914_, _11284_);
  and (_29916_, _29915_, _29913_);
  or (_29917_, _29916_, _29675_);
  nand (_29918_, _29917_, _06282_);
  and (_29919_, _08142_, _06281_);
  nor (_29920_, _29919_, _25646_);
  nand (_29921_, _29920_, _29918_);
  and (_29923_, _12403_, _25646_);
  nor (_29924_, _29923_, _06362_);
  and (_29925_, _29924_, _29921_);
  and (_29926_, _12187_, _13004_);
  nor (_29927_, _29683_, _13004_);
  nor (_29928_, _29927_, _29926_);
  nor (_29929_, _29928_, _06921_);
  or (_29930_, _29929_, _29925_);
  and (_29931_, _29930_, _13030_);
  nor (_29932_, _29674_, _13030_);
  or (_29934_, _29932_, _29931_);
  nand (_29935_, _29934_, _06926_);
  nor (_29936_, _12403_, _06926_);
  nor (_29937_, _29936_, _13038_);
  nand (_29938_, _29937_, _29935_);
  nor (_29939_, _29689_, _13037_);
  nor (_29940_, _29939_, _06361_);
  nand (_29941_, _29940_, _29938_);
  and (_29942_, _06361_, _06317_);
  nor (_29943_, _29942_, _05940_);
  nand (_29945_, _29943_, _29941_);
  and (_29946_, _12403_, _05940_);
  nor (_29947_, _29946_, _05927_);
  nand (_29948_, _29947_, _29945_);
  nor (_29949_, _29928_, _05928_);
  nor (_29950_, _29949_, _13053_);
  nand (_29951_, _29950_, _29948_);
  nor (_29952_, _29689_, _13052_);
  nor (_29953_, _29952_, _06278_);
  nand (_29954_, _29953_, _29951_);
  nor (_29956_, _12403_, _06279_);
  nor (_29957_, _29956_, _13059_);
  nand (_29958_, _29957_, _29954_);
  nor (_29959_, _29689_, _12141_);
  nor (_29960_, _29959_, _06379_);
  and (_29961_, _29960_, _29958_);
  and (_29962_, _06379_, _06317_);
  or (_29963_, _29962_, _29961_);
  nand (_29964_, _29963_, _29058_);
  nor (_29965_, _12403_, _29058_);
  nor (_29967_, _29965_, _13068_);
  and (_29968_, _29967_, _29964_);
  and (_29969_, _29674_, _13068_);
  or (_29970_, _29969_, _29968_);
  or (_29971_, _29970_, _01351_);
  or (_29972_, _01347_, \oc8051_golden_model_1.PC [14]);
  and (_29973_, _29972_, _42618_);
  and (_43261_, _29973_, _29971_);
  nand (_29974_, _11263_, _07904_);
  and (_29975_, _13077_, \oc8051_golden_model_1.P2 [0]);
  nor (_29977_, _29975_, _07234_);
  nand (_29978_, _29977_, _29974_);
  and (_29979_, _07904_, _07133_);
  or (_29980_, _29979_, _29975_);
  or (_29981_, _29980_, _07215_);
  nor (_29982_, _08390_, _13077_);
  or (_29983_, _29982_, _29975_);
  or (_29984_, _29983_, _07151_);
  and (_29985_, _07904_, \oc8051_golden_model_1.ACC [0]);
  or (_29986_, _29985_, _29975_);
  and (_29988_, _29986_, _07141_);
  and (_29989_, _07142_, \oc8051_golden_model_1.P2 [0]);
  or (_29990_, _29989_, _06341_);
  or (_29991_, _29990_, _29988_);
  and (_29992_, _29991_, _06273_);
  and (_29993_, _29992_, _29984_);
  and (_29994_, _13085_, \oc8051_golden_model_1.P2 [0]);
  and (_29995_, _14382_, _08624_);
  or (_29996_, _29995_, _29994_);
  and (_29997_, _29996_, _06272_);
  or (_29999_, _29997_, _29993_);
  and (_30000_, _29999_, _07166_);
  and (_30001_, _29980_, _06461_);
  or (_30002_, _30001_, _06464_);
  or (_30003_, _30002_, _30000_);
  or (_30004_, _29986_, _06465_);
  and (_30005_, _30004_, _06269_);
  and (_30006_, _30005_, _30003_);
  and (_30007_, _29975_, _06268_);
  or (_30008_, _30007_, _06261_);
  or (_30010_, _30008_, _30006_);
  or (_30011_, _29983_, _06262_);
  and (_30012_, _30011_, _06258_);
  and (_30013_, _30012_, _30010_);
  and (_30014_, _14413_, _08624_);
  or (_30015_, _30014_, _29994_);
  and (_30016_, _30015_, _06257_);
  or (_30017_, _30016_, _10080_);
  or (_30018_, _30017_, _30013_);
  and (_30019_, _30018_, _29981_);
  or (_30021_, _30019_, _07460_);
  and (_30022_, _09392_, _07904_);
  or (_30023_, _29975_, _07208_);
  or (_30024_, _30023_, _30022_);
  and (_30025_, _30024_, _30021_);
  or (_30026_, _30025_, _10094_);
  and (_30027_, _14467_, _07904_);
  or (_30028_, _29975_, _05982_);
  or (_30029_, _30028_, _30027_);
  and (_30030_, _30029_, _06219_);
  and (_30032_, _30030_, _30026_);
  and (_30033_, _07904_, _08954_);
  or (_30034_, _30033_, _29975_);
  and (_30035_, _30034_, _06218_);
  or (_30036_, _30035_, _06369_);
  or (_30037_, _30036_, _30032_);
  and (_30038_, _14366_, _07904_);
  or (_30039_, _30038_, _29975_);
  or (_30040_, _30039_, _07237_);
  and (_30041_, _30040_, _07240_);
  and (_30043_, _30041_, _30037_);
  nor (_30044_, _12580_, _13077_);
  or (_30045_, _30044_, _29975_);
  and (_30046_, _29974_, _06536_);
  and (_30047_, _30046_, _30045_);
  or (_30048_, _30047_, _30043_);
  and (_30049_, _30048_, _07242_);
  nand (_30050_, _30034_, _06375_);
  nor (_30051_, _30050_, _29982_);
  or (_30052_, _30051_, _06545_);
  or (_30054_, _30052_, _30049_);
  and (_30055_, _30054_, _29978_);
  or (_30056_, _30055_, _06366_);
  and (_30057_, _14363_, _07904_);
  or (_30058_, _29975_, _09056_);
  or (_30059_, _30058_, _30057_);
  and (_30060_, _30059_, _09061_);
  and (_30061_, _30060_, _30056_);
  and (_30062_, _30045_, _06528_);
  or (_30063_, _30062_, _06568_);
  or (_30065_, _30063_, _30061_);
  or (_30066_, _29983_, _06926_);
  and (_30067_, _30066_, _30065_);
  or (_30068_, _30067_, _05927_);
  or (_30069_, _29975_, _05928_);
  and (_30070_, _30069_, _30068_);
  or (_30071_, _30070_, _06278_);
  or (_30072_, _29983_, _06279_);
  and (_30073_, _30072_, _01347_);
  and (_30074_, _30073_, _30071_);
  nor (_30076_, \oc8051_golden_model_1.P2 [0], rst);
  nor (_30077_, _30076_, _01354_);
  or (_43262_, _30077_, _30074_);
  nor (_30078_, \oc8051_golden_model_1.P2 [1], rst);
  nor (_30079_, _30078_, _01354_);
  and (_30080_, _13077_, \oc8051_golden_model_1.P2 [1]);
  nor (_30081_, _11261_, _13077_);
  or (_30082_, _30081_, _30080_);
  or (_30083_, _30082_, _09061_);
  nand (_30084_, _07904_, _07038_);
  or (_30086_, _07904_, \oc8051_golden_model_1.P2 [1]);
  and (_30087_, _30086_, _06218_);
  and (_30088_, _30087_, _30084_);
  nor (_30089_, _13077_, _07357_);
  or (_30090_, _30089_, _30080_);
  and (_30091_, _30090_, _06461_);
  and (_30092_, _13085_, \oc8051_golden_model_1.P2 [1]);
  and (_30093_, _14557_, _08624_);
  or (_30094_, _30093_, _30092_);
  or (_30095_, _30094_, _06273_);
  and (_30097_, _14562_, _07904_);
  not (_30098_, _30097_);
  and (_30099_, _30098_, _30086_);
  and (_30100_, _30099_, _06341_);
  and (_30101_, _07142_, \oc8051_golden_model_1.P2 [1]);
  and (_30102_, _07904_, \oc8051_golden_model_1.ACC [1]);
  or (_30103_, _30102_, _30080_);
  and (_30104_, _30103_, _07141_);
  or (_30105_, _30104_, _30101_);
  and (_30106_, _30105_, _07151_);
  or (_30108_, _30106_, _06272_);
  or (_30109_, _30108_, _30100_);
  and (_30110_, _30109_, _30095_);
  and (_30111_, _30110_, _07166_);
  or (_30112_, _30111_, _30091_);
  or (_30113_, _30112_, _06464_);
  or (_30114_, _30103_, _06465_);
  and (_30115_, _30114_, _06269_);
  and (_30116_, _30115_, _30113_);
  and (_30117_, _14560_, _08624_);
  or (_30119_, _30117_, _30092_);
  and (_30120_, _30119_, _06268_);
  or (_30121_, _30120_, _06261_);
  or (_30122_, _30121_, _30116_);
  or (_30123_, _30092_, _14556_);
  and (_30124_, _30123_, _30094_);
  or (_30125_, _30124_, _06262_);
  and (_30126_, _30125_, _06258_);
  and (_30127_, _30126_, _30122_);
  or (_30128_, _30092_, _14597_);
  and (_30130_, _30128_, _06257_);
  and (_30131_, _30130_, _30094_);
  or (_30132_, _30131_, _10080_);
  or (_30133_, _30132_, _30127_);
  or (_30134_, _30090_, _07215_);
  and (_30135_, _30134_, _30133_);
  or (_30136_, _30135_, _07460_);
  and (_30137_, _09451_, _07904_);
  or (_30138_, _30080_, _07208_);
  or (_30139_, _30138_, _30137_);
  and (_30141_, _30139_, _05982_);
  and (_30142_, _30141_, _30136_);
  and (_30143_, _14653_, _07904_);
  or (_30144_, _30143_, _30080_);
  and (_30145_, _30144_, _10094_);
  or (_30146_, _30145_, _30142_);
  and (_30147_, _30146_, _06219_);
  or (_30148_, _30147_, _30088_);
  and (_30149_, _30148_, _07237_);
  or (_30150_, _14668_, _13077_);
  and (_30152_, _30086_, _06369_);
  and (_30153_, _30152_, _30150_);
  or (_30154_, _30153_, _06536_);
  or (_30155_, _30154_, _30149_);
  nand (_30156_, _11260_, _07904_);
  and (_30157_, _30156_, _30082_);
  or (_30158_, _30157_, _07240_);
  and (_30159_, _30158_, _07242_);
  and (_30160_, _30159_, _30155_);
  or (_30161_, _14666_, _13077_);
  and (_30163_, _30086_, _06375_);
  and (_30164_, _30163_, _30161_);
  or (_30165_, _30164_, _06545_);
  or (_30166_, _30165_, _30160_);
  nor (_30167_, _30080_, _07234_);
  nand (_30168_, _30167_, _30156_);
  and (_30169_, _30168_, _09056_);
  and (_30170_, _30169_, _30166_);
  or (_30171_, _30084_, _08341_);
  and (_30172_, _30086_, _06366_);
  and (_30174_, _30172_, _30171_);
  or (_30175_, _30174_, _06528_);
  or (_30176_, _30175_, _30170_);
  and (_30177_, _30176_, _30083_);
  or (_30178_, _30177_, _06568_);
  or (_30179_, _30099_, _06926_);
  and (_30180_, _30179_, _05928_);
  and (_30181_, _30180_, _30178_);
  and (_30182_, _30119_, _05927_);
  or (_30183_, _30182_, _06278_);
  or (_30185_, _30183_, _30181_);
  or (_30186_, _30080_, _06279_);
  or (_30187_, _30186_, _30097_);
  and (_30188_, _30187_, _01347_);
  and (_30189_, _30188_, _30185_);
  or (_43264_, _30189_, _30079_);
  and (_30190_, _13077_, \oc8051_golden_model_1.P2 [2]);
  nor (_30191_, _13077_, _07776_);
  or (_30192_, _30191_, _30190_);
  or (_30193_, _30192_, _07215_);
  or (_30195_, _30192_, _07166_);
  and (_30196_, _14770_, _07904_);
  or (_30197_, _30196_, _30190_);
  or (_30198_, _30197_, _07151_);
  and (_30199_, _07904_, \oc8051_golden_model_1.ACC [2]);
  or (_30200_, _30199_, _30190_);
  and (_30201_, _30200_, _07141_);
  and (_30202_, _07142_, \oc8051_golden_model_1.P2 [2]);
  or (_30203_, _30202_, _06341_);
  or (_30204_, _30203_, _30201_);
  and (_30206_, _30204_, _06273_);
  and (_30207_, _30206_, _30198_);
  and (_30208_, _13085_, \oc8051_golden_model_1.P2 [2]);
  and (_30209_, _14774_, _08624_);
  or (_30210_, _30209_, _30208_);
  and (_30211_, _30210_, _06272_);
  or (_30212_, _30211_, _06461_);
  or (_30213_, _30212_, _30207_);
  and (_30214_, _30213_, _30195_);
  or (_30215_, _30214_, _06464_);
  or (_30217_, _30200_, _06465_);
  and (_30218_, _30217_, _06269_);
  and (_30219_, _30218_, _30215_);
  and (_30220_, _14756_, _08624_);
  or (_30221_, _30220_, _30208_);
  and (_30222_, _30221_, _06268_);
  or (_30223_, _30222_, _06261_);
  or (_30224_, _30223_, _30219_);
  and (_30225_, _30209_, _14789_);
  or (_30226_, _30208_, _06262_);
  or (_30228_, _30226_, _30225_);
  and (_30229_, _30228_, _06258_);
  and (_30230_, _30229_, _30224_);
  and (_30231_, _14804_, _08624_);
  or (_30232_, _30231_, _30208_);
  and (_30233_, _30232_, _06257_);
  or (_30234_, _30233_, _10080_);
  or (_30235_, _30234_, _30230_);
  and (_30236_, _30235_, _30193_);
  or (_30237_, _30236_, _07460_);
  and (_30239_, _09450_, _07904_);
  or (_30240_, _30190_, _07208_);
  or (_30241_, _30240_, _30239_);
  and (_30242_, _30241_, _05982_);
  and (_30243_, _30242_, _30237_);
  and (_30244_, _14859_, _07904_);
  or (_30245_, _30244_, _30190_);
  and (_30246_, _30245_, _10094_);
  or (_30247_, _30246_, _06218_);
  or (_30248_, _30247_, _30243_);
  and (_30250_, _07904_, _08973_);
  or (_30251_, _30250_, _30190_);
  or (_30252_, _30251_, _06219_);
  and (_30253_, _30252_, _30248_);
  or (_30254_, _30253_, _06369_);
  and (_30255_, _14751_, _07904_);
  or (_30256_, _30255_, _30190_);
  or (_30257_, _30256_, _07237_);
  and (_30258_, _30257_, _07240_);
  and (_30259_, _30258_, _30254_);
  and (_30261_, _11259_, _07904_);
  or (_30262_, _30261_, _30190_);
  and (_30263_, _30262_, _06536_);
  or (_30264_, _30263_, _30259_);
  and (_30265_, _30264_, _07242_);
  or (_30266_, _30190_, _08440_);
  and (_30267_, _30251_, _06375_);
  and (_30268_, _30267_, _30266_);
  or (_30269_, _30268_, _30265_);
  and (_30270_, _30269_, _07234_);
  and (_30272_, _30200_, _06545_);
  and (_30273_, _30272_, _30266_);
  or (_30274_, _30273_, _06366_);
  or (_30275_, _30274_, _30270_);
  and (_30276_, _14748_, _07904_);
  or (_30277_, _30190_, _09056_);
  or (_30278_, _30277_, _30276_);
  and (_30279_, _30278_, _09061_);
  and (_30280_, _30279_, _30275_);
  nor (_30281_, _11258_, _13077_);
  or (_30283_, _30281_, _30190_);
  and (_30284_, _30283_, _06528_);
  or (_30285_, _30284_, _06568_);
  or (_30286_, _30285_, _30280_);
  or (_30287_, _30197_, _06926_);
  and (_30288_, _30287_, _05928_);
  and (_30289_, _30288_, _30286_);
  and (_30290_, _30221_, _05927_);
  or (_30291_, _30290_, _06278_);
  or (_30292_, _30291_, _30289_);
  and (_30294_, _14926_, _07904_);
  or (_30295_, _30190_, _06279_);
  or (_30296_, _30295_, _30294_);
  and (_30297_, _30296_, _01347_);
  and (_30298_, _30297_, _30292_);
  nor (_30299_, \oc8051_golden_model_1.P2 [2], rst);
  nor (_30300_, _30299_, _01354_);
  or (_43265_, _30300_, _30298_);
  and (_30301_, _13077_, \oc8051_golden_model_1.P2 [3]);
  nor (_30302_, _13077_, _07594_);
  or (_30304_, _30302_, _30301_);
  or (_30305_, _30304_, _07215_);
  and (_30306_, _14953_, _07904_);
  or (_30307_, _30306_, _30301_);
  or (_30308_, _30307_, _07151_);
  and (_30309_, _07904_, \oc8051_golden_model_1.ACC [3]);
  or (_30310_, _30309_, _30301_);
  and (_30311_, _30310_, _07141_);
  and (_30312_, _07142_, \oc8051_golden_model_1.P2 [3]);
  or (_30313_, _30312_, _06341_);
  or (_30315_, _30313_, _30311_);
  and (_30316_, _30315_, _06273_);
  and (_30317_, _30316_, _30308_);
  and (_30318_, _13085_, \oc8051_golden_model_1.P2 [3]);
  and (_30319_, _14950_, _08624_);
  or (_30320_, _30319_, _30318_);
  and (_30321_, _30320_, _06272_);
  or (_30322_, _30321_, _06461_);
  or (_30323_, _30322_, _30317_);
  or (_30324_, _30304_, _07166_);
  and (_30325_, _30324_, _30323_);
  or (_30326_, _30325_, _06464_);
  or (_30327_, _30310_, _06465_);
  and (_30328_, _30327_, _06269_);
  and (_30329_, _30328_, _30326_);
  and (_30330_, _14948_, _08624_);
  or (_30331_, _30330_, _30318_);
  and (_30332_, _30331_, _06268_);
  or (_30333_, _30332_, _06261_);
  or (_30334_, _30333_, _30329_);
  or (_30337_, _30318_, _14979_);
  and (_30338_, _30337_, _30320_);
  or (_30339_, _30338_, _06262_);
  and (_30340_, _30339_, _06258_);
  and (_30341_, _30340_, _30334_);
  or (_30342_, _30318_, _14992_);
  and (_30343_, _30342_, _06257_);
  and (_30344_, _30343_, _30320_);
  or (_30345_, _30344_, _10080_);
  or (_30346_, _30345_, _30341_);
  and (_30348_, _30346_, _30305_);
  or (_30349_, _30348_, _07460_);
  and (_30350_, _09449_, _07904_);
  or (_30351_, _30301_, _07208_);
  or (_30352_, _30351_, _30350_);
  and (_30353_, _30352_, _05982_);
  and (_30354_, _30353_, _30349_);
  and (_30355_, _15048_, _07904_);
  or (_30356_, _30355_, _30301_);
  and (_30357_, _30356_, _10094_);
  or (_30359_, _30357_, _06218_);
  or (_30360_, _30359_, _30354_);
  and (_30361_, _07904_, _08930_);
  or (_30362_, _30361_, _30301_);
  or (_30363_, _30362_, _06219_);
  and (_30364_, _30363_, _30360_);
  or (_30365_, _30364_, _06369_);
  and (_30366_, _14943_, _07904_);
  or (_30367_, _30366_, _30301_);
  or (_30368_, _30367_, _07237_);
  and (_30370_, _30368_, _07240_);
  and (_30371_, _30370_, _30365_);
  and (_30372_, _12577_, _07904_);
  or (_30373_, _30372_, _30301_);
  and (_30374_, _30373_, _06536_);
  or (_30375_, _30374_, _30371_);
  and (_30376_, _30375_, _07242_);
  or (_30377_, _30301_, _08292_);
  and (_30378_, _30362_, _06375_);
  and (_30379_, _30378_, _30377_);
  or (_30381_, _30379_, _30376_);
  and (_30382_, _30381_, _07234_);
  and (_30383_, _30310_, _06545_);
  and (_30384_, _30383_, _30377_);
  or (_30385_, _30384_, _06366_);
  or (_30386_, _30385_, _30382_);
  and (_30387_, _14940_, _07904_);
  or (_30388_, _30301_, _09056_);
  or (_30389_, _30388_, _30387_);
  and (_30390_, _30389_, _09061_);
  and (_30392_, _30390_, _30386_);
  nor (_30393_, _11256_, _13077_);
  or (_30394_, _30393_, _30301_);
  and (_30395_, _30394_, _06528_);
  or (_30396_, _30395_, _06568_);
  or (_30397_, _30396_, _30392_);
  or (_30398_, _30307_, _06926_);
  and (_30399_, _30398_, _05928_);
  and (_30400_, _30399_, _30397_);
  and (_30401_, _30331_, _05927_);
  or (_30403_, _30401_, _06278_);
  or (_30404_, _30403_, _30400_);
  and (_30405_, _15128_, _07904_);
  or (_30406_, _30301_, _06279_);
  or (_30407_, _30406_, _30405_);
  and (_30408_, _30407_, _01347_);
  and (_30409_, _30408_, _30404_);
  nor (_30410_, \oc8051_golden_model_1.P2 [3], rst);
  nor (_30411_, _30410_, _01354_);
  or (_43266_, _30411_, _30409_);
  nor (_30413_, \oc8051_golden_model_1.P2 [4], rst);
  nor (_30414_, _30413_, _01354_);
  and (_30415_, _13077_, \oc8051_golden_model_1.P2 [4]);
  nor (_30416_, _08541_, _13077_);
  or (_30417_, _30416_, _30415_);
  or (_30418_, _30417_, _07215_);
  and (_30419_, _13085_, \oc8051_golden_model_1.P2 [4]);
  and (_30420_, _15176_, _08624_);
  or (_30421_, _30420_, _30419_);
  and (_30422_, _30421_, _06268_);
  and (_30424_, _15162_, _07904_);
  or (_30425_, _30424_, _30415_);
  or (_30426_, _30425_, _07151_);
  and (_30427_, _07904_, \oc8051_golden_model_1.ACC [4]);
  or (_30428_, _30427_, _30415_);
  and (_30429_, _30428_, _07141_);
  and (_30430_, _07142_, \oc8051_golden_model_1.P2 [4]);
  or (_30431_, _30430_, _06341_);
  or (_30432_, _30431_, _30429_);
  and (_30433_, _30432_, _06273_);
  and (_30435_, _30433_, _30426_);
  and (_30436_, _15166_, _08624_);
  or (_30437_, _30436_, _30419_);
  and (_30438_, _30437_, _06272_);
  or (_30439_, _30438_, _06461_);
  or (_30440_, _30439_, _30435_);
  or (_30441_, _30417_, _07166_);
  and (_30442_, _30441_, _30440_);
  or (_30443_, _30442_, _06464_);
  or (_30444_, _30428_, _06465_);
  and (_30446_, _30444_, _06269_);
  and (_30447_, _30446_, _30443_);
  or (_30448_, _30447_, _30422_);
  and (_30449_, _30448_, _06262_);
  and (_30450_, _15184_, _08624_);
  or (_30451_, _30450_, _30419_);
  and (_30452_, _30451_, _06261_);
  or (_30453_, _30452_, _30449_);
  and (_30454_, _30453_, _06258_);
  and (_30455_, _15200_, _08624_);
  or (_30457_, _30455_, _30419_);
  and (_30458_, _30457_, _06257_);
  or (_30459_, _30458_, _10080_);
  or (_30460_, _30459_, _30454_);
  and (_30461_, _30460_, _30418_);
  or (_30462_, _30461_, _07460_);
  and (_30463_, _09448_, _07904_);
  or (_30464_, _30415_, _07208_);
  or (_30465_, _30464_, _30463_);
  and (_30466_, _30465_, _05982_);
  and (_30468_, _30466_, _30462_);
  and (_30469_, _15254_, _07904_);
  or (_30470_, _30469_, _30415_);
  and (_30471_, _30470_, _10094_);
  or (_30472_, _30471_, _06218_);
  or (_30473_, _30472_, _30468_);
  and (_30474_, _08959_, _07904_);
  or (_30475_, _30474_, _30415_);
  or (_30476_, _30475_, _06219_);
  and (_30477_, _30476_, _30473_);
  or (_30479_, _30477_, _06369_);
  and (_30480_, _15269_, _07904_);
  or (_30481_, _30480_, _30415_);
  or (_30482_, _30481_, _07237_);
  and (_30483_, _30482_, _07240_);
  and (_30484_, _30483_, _30479_);
  and (_30485_, _11254_, _07904_);
  or (_30486_, _30485_, _30415_);
  and (_30487_, _30486_, _06536_);
  or (_30488_, _30487_, _30484_);
  and (_30490_, _30488_, _07242_);
  or (_30491_, _30415_, _08544_);
  and (_30492_, _30475_, _06375_);
  and (_30493_, _30492_, _30491_);
  or (_30494_, _30493_, _30490_);
  and (_30495_, _30494_, _07234_);
  and (_30496_, _30428_, _06545_);
  and (_30497_, _30496_, _30491_);
  or (_30498_, _30497_, _06366_);
  or (_30499_, _30498_, _30495_);
  and (_30501_, _15266_, _07904_);
  or (_30502_, _30415_, _09056_);
  or (_30503_, _30502_, _30501_);
  and (_30504_, _30503_, _09061_);
  and (_30505_, _30504_, _30499_);
  nor (_30506_, _11253_, _13077_);
  or (_30507_, _30506_, _30415_);
  and (_30508_, _30507_, _06528_);
  or (_30509_, _30508_, _06568_);
  or (_30510_, _30509_, _30505_);
  or (_30512_, _30425_, _06926_);
  and (_30513_, _30512_, _05928_);
  and (_30514_, _30513_, _30510_);
  and (_30515_, _30421_, _05927_);
  or (_30516_, _30515_, _06278_);
  or (_30517_, _30516_, _30514_);
  and (_30518_, _15329_, _07904_);
  or (_30519_, _30415_, _06279_);
  or (_30520_, _30519_, _30518_);
  and (_30521_, _30520_, _01347_);
  and (_30523_, _30521_, _30517_);
  or (_43267_, _30523_, _30414_);
  and (_30524_, _13077_, \oc8051_golden_model_1.P2 [5]);
  and (_30525_, _15358_, _07904_);
  or (_30526_, _30525_, _30524_);
  or (_30527_, _30526_, _07151_);
  and (_30528_, _07904_, \oc8051_golden_model_1.ACC [5]);
  or (_30529_, _30528_, _30524_);
  and (_30530_, _30529_, _07141_);
  and (_30531_, _07142_, \oc8051_golden_model_1.P2 [5]);
  or (_30533_, _30531_, _06341_);
  or (_30534_, _30533_, _30530_);
  and (_30535_, _30534_, _06273_);
  and (_30536_, _30535_, _30527_);
  and (_30537_, _13085_, \oc8051_golden_model_1.P2 [5]);
  and (_30538_, _15372_, _08624_);
  or (_30539_, _30538_, _30537_);
  and (_30540_, _30539_, _06272_);
  or (_30541_, _30540_, _06461_);
  or (_30542_, _30541_, _30536_);
  nor (_30544_, _08244_, _13077_);
  or (_30545_, _30544_, _30524_);
  or (_30546_, _30545_, _07166_);
  and (_30547_, _30546_, _30542_);
  or (_30548_, _30547_, _06464_);
  or (_30549_, _30529_, _06465_);
  and (_30550_, _30549_, _06269_);
  and (_30551_, _30550_, _30548_);
  and (_30552_, _15355_, _08624_);
  or (_30553_, _30552_, _30537_);
  and (_30555_, _30553_, _06268_);
  or (_30556_, _30555_, _06261_);
  or (_30557_, _30556_, _30551_);
  or (_30558_, _30537_, _15387_);
  and (_30559_, _30558_, _30539_);
  or (_30560_, _30559_, _06262_);
  and (_30561_, _30560_, _06258_);
  and (_30562_, _30561_, _30557_);
  or (_30563_, _30537_, _15403_);
  and (_30564_, _30563_, _06257_);
  and (_30566_, _30564_, _30539_);
  or (_30567_, _30566_, _10080_);
  or (_30568_, _30567_, _30562_);
  or (_30569_, _30545_, _07215_);
  and (_30570_, _30569_, _30568_);
  or (_30571_, _30570_, _07460_);
  and (_30572_, _09447_, _07904_);
  or (_30573_, _30524_, _07208_);
  or (_30574_, _30573_, _30572_);
  and (_30575_, _30574_, _05982_);
  and (_30577_, _30575_, _30571_);
  and (_30578_, _15459_, _07904_);
  or (_30579_, _30578_, _30524_);
  and (_30580_, _30579_, _10094_);
  or (_30581_, _30580_, _06218_);
  or (_30582_, _30581_, _30577_);
  and (_30583_, _08946_, _07904_);
  or (_30584_, _30583_, _30524_);
  or (_30585_, _30584_, _06219_);
  and (_30586_, _30585_, _30582_);
  or (_30588_, _30586_, _06369_);
  and (_30589_, _15353_, _07904_);
  or (_30590_, _30589_, _30524_);
  or (_30591_, _30590_, _07237_);
  and (_30592_, _30591_, _07240_);
  and (_30593_, _30592_, _30588_);
  and (_30594_, _11250_, _07904_);
  or (_30595_, _30594_, _30524_);
  and (_30596_, _30595_, _06536_);
  or (_30597_, _30596_, _30593_);
  and (_30599_, _30597_, _07242_);
  or (_30600_, _30524_, _08247_);
  and (_30601_, _30584_, _06375_);
  and (_30602_, _30601_, _30600_);
  or (_30603_, _30602_, _30599_);
  and (_30604_, _30603_, _07234_);
  and (_30605_, _30529_, _06545_);
  and (_30606_, _30605_, _30600_);
  or (_30607_, _30606_, _06366_);
  or (_30608_, _30607_, _30604_);
  and (_30610_, _15350_, _07904_);
  or (_30611_, _30524_, _09056_);
  or (_30612_, _30611_, _30610_);
  and (_30613_, _30612_, _09061_);
  and (_30614_, _30613_, _30608_);
  nor (_30615_, _11249_, _13077_);
  or (_30616_, _30615_, _30524_);
  and (_30617_, _30616_, _06528_);
  or (_30618_, _30617_, _06568_);
  or (_30619_, _30618_, _30614_);
  or (_30621_, _30526_, _06926_);
  and (_30622_, _30621_, _05928_);
  and (_30623_, _30622_, _30619_);
  and (_30624_, _30553_, _05927_);
  or (_30625_, _30624_, _06278_);
  or (_30626_, _30625_, _30623_);
  and (_30627_, _15532_, _07904_);
  or (_30628_, _30524_, _06279_);
  or (_30629_, _30628_, _30627_);
  and (_30630_, _30629_, _01347_);
  and (_30632_, _30630_, _30626_);
  nor (_30633_, \oc8051_golden_model_1.P2 [5], rst);
  nor (_30634_, _30633_, _01354_);
  or (_43268_, _30634_, _30632_);
  nor (_30635_, \oc8051_golden_model_1.P2 [6], rst);
  nor (_30636_, _30635_, _01354_);
  and (_30637_, _13077_, \oc8051_golden_model_1.P2 [6]);
  and (_30638_, _15554_, _07904_);
  or (_30639_, _30638_, _30637_);
  or (_30640_, _30639_, _07151_);
  and (_30642_, _07904_, \oc8051_golden_model_1.ACC [6]);
  or (_30643_, _30642_, _30637_);
  and (_30644_, _30643_, _07141_);
  and (_30645_, _07142_, \oc8051_golden_model_1.P2 [6]);
  or (_30646_, _30645_, _06341_);
  or (_30647_, _30646_, _30644_);
  and (_30648_, _30647_, _06273_);
  and (_30649_, _30648_, _30640_);
  and (_30650_, _13085_, \oc8051_golden_model_1.P2 [6]);
  and (_30651_, _15570_, _08624_);
  or (_30653_, _30651_, _30650_);
  and (_30654_, _30653_, _06272_);
  or (_30655_, _30654_, _06461_);
  or (_30656_, _30655_, _30649_);
  nor (_30657_, _08142_, _13077_);
  or (_30658_, _30657_, _30637_);
  or (_30659_, _30658_, _07166_);
  and (_30660_, _30659_, _30656_);
  or (_30661_, _30660_, _06464_);
  or (_30662_, _30643_, _06465_);
  and (_30664_, _30662_, _06269_);
  and (_30665_, _30664_, _30661_);
  and (_30666_, _15551_, _08624_);
  or (_30667_, _30666_, _30650_);
  and (_30668_, _30667_, _06268_);
  or (_30669_, _30668_, _06261_);
  or (_30670_, _30669_, _30665_);
  or (_30671_, _30650_, _15585_);
  and (_30672_, _30671_, _30653_);
  or (_30673_, _30672_, _06262_);
  and (_30675_, _30673_, _06258_);
  and (_30676_, _30675_, _30670_);
  and (_30677_, _15602_, _08624_);
  or (_30678_, _30677_, _30650_);
  and (_30679_, _30678_, _06257_);
  or (_30680_, _30679_, _10080_);
  or (_30681_, _30680_, _30676_);
  or (_30682_, _30658_, _07215_);
  and (_30683_, _30682_, _30681_);
  or (_30684_, _30683_, _07460_);
  and (_30686_, _09446_, _07904_);
  or (_30687_, _30637_, _07208_);
  or (_30688_, _30687_, _30686_);
  and (_30689_, _30688_, _05982_);
  and (_30690_, _30689_, _30684_);
  and (_30691_, _15657_, _07904_);
  or (_30692_, _30691_, _30637_);
  and (_30693_, _30692_, _10094_);
  or (_30694_, _30693_, _06218_);
  or (_30695_, _30694_, _30690_);
  and (_30697_, _15664_, _07904_);
  or (_30698_, _30697_, _30637_);
  or (_30699_, _30698_, _06219_);
  and (_30700_, _30699_, _30695_);
  or (_30701_, _30700_, _06369_);
  and (_30702_, _15549_, _07904_);
  or (_30703_, _30702_, _30637_);
  or (_30704_, _30703_, _07237_);
  and (_30705_, _30704_, _07240_);
  and (_30706_, _30705_, _30701_);
  and (_30708_, _11247_, _07904_);
  or (_30709_, _30708_, _30637_);
  and (_30710_, _30709_, _06536_);
  or (_30711_, _30710_, _30706_);
  and (_30712_, _30711_, _07242_);
  or (_30713_, _30637_, _08145_);
  and (_30714_, _30698_, _06375_);
  and (_30715_, _30714_, _30713_);
  or (_30716_, _30715_, _30712_);
  and (_30717_, _30716_, _07234_);
  and (_30719_, _30643_, _06545_);
  and (_30720_, _30719_, _30713_);
  or (_30721_, _30720_, _06366_);
  or (_30722_, _30721_, _30717_);
  and (_30723_, _15546_, _07904_);
  or (_30724_, _30637_, _09056_);
  or (_30725_, _30724_, _30723_);
  and (_30726_, _30725_, _09061_);
  and (_30727_, _30726_, _30722_);
  nor (_30728_, _11246_, _13077_);
  or (_30730_, _30728_, _30637_);
  and (_30731_, _30730_, _06528_);
  or (_30732_, _30731_, _06568_);
  or (_30733_, _30732_, _30727_);
  or (_30734_, _30639_, _06926_);
  and (_30735_, _30734_, _05928_);
  and (_30736_, _30735_, _30733_);
  and (_30737_, _30667_, _05927_);
  or (_30738_, _30737_, _06278_);
  or (_30739_, _30738_, _30736_);
  and (_30741_, _15734_, _07904_);
  or (_30742_, _30637_, _06279_);
  or (_30743_, _30742_, _30741_);
  and (_30744_, _30743_, _01347_);
  and (_30745_, _30744_, _30739_);
  or (_43269_, _30745_, _30636_);
  and (_30746_, _07894_, \oc8051_golden_model_1.ACC [0]);
  and (_30747_, _30746_, _08390_);
  and (_30748_, _13180_, \oc8051_golden_model_1.P3 [0]);
  or (_30749_, _30748_, _07234_);
  or (_30751_, _30749_, _30747_);
  and (_30752_, _07894_, _07133_);
  or (_30753_, _30752_, _30748_);
  or (_30754_, _30753_, _07215_);
  nor (_30755_, _08390_, _13180_);
  or (_30756_, _30755_, _30748_);
  and (_30757_, _30756_, _06341_);
  and (_30758_, _07142_, \oc8051_golden_model_1.P3 [0]);
  or (_30759_, _30746_, _30748_);
  and (_30760_, _30759_, _07141_);
  or (_30762_, _30760_, _30758_);
  and (_30763_, _30762_, _07151_);
  or (_30764_, _30763_, _06272_);
  or (_30765_, _30764_, _30757_);
  and (_30766_, _14382_, _08628_);
  and (_30767_, _13188_, \oc8051_golden_model_1.P3 [0]);
  or (_30768_, _30767_, _06273_);
  or (_30769_, _30768_, _30766_);
  and (_30770_, _30769_, _07166_);
  and (_30771_, _30770_, _30765_);
  and (_30773_, _30753_, _06461_);
  or (_30774_, _30773_, _06464_);
  or (_30775_, _30774_, _30771_);
  or (_30776_, _30759_, _06465_);
  and (_30777_, _30776_, _06269_);
  and (_30778_, _30777_, _30775_);
  and (_30779_, _30748_, _06268_);
  or (_30780_, _30779_, _06261_);
  or (_30781_, _30780_, _30778_);
  or (_30782_, _30756_, _06262_);
  and (_30784_, _30782_, _06258_);
  and (_30785_, _30784_, _30781_);
  and (_30786_, _14413_, _08628_);
  or (_30787_, _30786_, _30767_);
  and (_30788_, _30787_, _06257_);
  or (_30789_, _30788_, _10080_);
  or (_30790_, _30789_, _30785_);
  and (_30791_, _30790_, _30754_);
  or (_30792_, _30791_, _07460_);
  and (_30793_, _09392_, _07894_);
  or (_30795_, _30748_, _07208_);
  or (_30796_, _30795_, _30793_);
  and (_30797_, _30796_, _30792_);
  or (_30798_, _30797_, _10094_);
  and (_30799_, _14467_, _07894_);
  or (_30800_, _30748_, _05982_);
  or (_30801_, _30800_, _30799_);
  and (_30802_, _30801_, _06219_);
  and (_30803_, _30802_, _30798_);
  and (_30804_, _07894_, _08954_);
  or (_30806_, _30804_, _30748_);
  and (_30807_, _30806_, _06218_);
  or (_30808_, _30807_, _06369_);
  or (_30809_, _30808_, _30803_);
  and (_30810_, _14366_, _07894_);
  or (_30811_, _30810_, _30748_);
  or (_30812_, _30811_, _07237_);
  and (_30813_, _30812_, _07240_);
  and (_30814_, _30813_, _30809_);
  nor (_30815_, _12580_, _13180_);
  or (_30817_, _30815_, _30748_);
  nor (_30818_, _30747_, _07240_);
  and (_30819_, _30818_, _30817_);
  or (_30820_, _30819_, _30814_);
  and (_30821_, _30820_, _07242_);
  nand (_30822_, _30806_, _06375_);
  nor (_30823_, _30822_, _30755_);
  or (_30824_, _30823_, _06545_);
  or (_30825_, _30824_, _30821_);
  and (_30826_, _30825_, _30751_);
  or (_30828_, _30826_, _06366_);
  and (_30829_, _14363_, _07894_);
  or (_30830_, _30748_, _09056_);
  or (_30831_, _30830_, _30829_);
  and (_30832_, _30831_, _09061_);
  and (_30833_, _30832_, _30828_);
  and (_30834_, _30817_, _06528_);
  or (_30835_, _30834_, _06568_);
  or (_30836_, _30835_, _30833_);
  or (_30837_, _30756_, _06926_);
  and (_30839_, _30837_, _30836_);
  or (_30840_, _30839_, _05927_);
  or (_30841_, _30748_, _05928_);
  and (_30842_, _30841_, _30840_);
  or (_30843_, _30842_, _06278_);
  or (_30844_, _30756_, _06279_);
  and (_30845_, _30844_, _01347_);
  and (_30846_, _30845_, _30843_);
  nor (_30847_, \oc8051_golden_model_1.P3 [0], rst);
  nor (_30848_, _30847_, _01354_);
  or (_43271_, _30848_, _30846_);
  and (_30850_, _13180_, \oc8051_golden_model_1.P3 [1]);
  nor (_30851_, _11261_, _13180_);
  or (_30852_, _30851_, _30850_);
  or (_30853_, _30852_, _09061_);
  nand (_30854_, _07894_, _07038_);
  or (_30855_, _07894_, \oc8051_golden_model_1.P3 [1]);
  and (_30856_, _30855_, _06218_);
  and (_30857_, _30856_, _30854_);
  nor (_30858_, _13180_, _07357_);
  or (_30860_, _30858_, _30850_);
  or (_30861_, _30860_, _07166_);
  and (_30862_, _14562_, _07894_);
  not (_30863_, _30862_);
  and (_30864_, _30863_, _30855_);
  or (_30865_, _30864_, _07151_);
  and (_30866_, _07894_, \oc8051_golden_model_1.ACC [1]);
  or (_30867_, _30866_, _30850_);
  and (_30868_, _30867_, _07141_);
  and (_30869_, _07142_, \oc8051_golden_model_1.P3 [1]);
  or (_30871_, _30869_, _06341_);
  or (_30872_, _30871_, _30868_);
  and (_30873_, _30872_, _06273_);
  and (_30874_, _30873_, _30865_);
  and (_30875_, _13188_, \oc8051_golden_model_1.P3 [1]);
  and (_30876_, _14557_, _08628_);
  or (_30877_, _30876_, _30875_);
  and (_30878_, _30877_, _06272_);
  or (_30879_, _30878_, _06461_);
  or (_30880_, _30879_, _30874_);
  and (_30882_, _30880_, _30861_);
  or (_30883_, _30882_, _06464_);
  or (_30884_, _30867_, _06465_);
  and (_30885_, _30884_, _06269_);
  and (_30886_, _30885_, _30883_);
  and (_30887_, _14560_, _08628_);
  or (_30888_, _30887_, _30875_);
  and (_30889_, _30888_, _06268_);
  or (_30890_, _30889_, _06261_);
  or (_30891_, _30890_, _30886_);
  and (_30893_, _30876_, _14556_);
  or (_30894_, _30875_, _06262_);
  or (_30895_, _30894_, _30893_);
  and (_30896_, _30895_, _06258_);
  and (_30897_, _30896_, _30891_);
  or (_30898_, _30875_, _14597_);
  and (_30899_, _30898_, _06257_);
  and (_30900_, _30899_, _30877_);
  or (_30901_, _30900_, _10080_);
  or (_30902_, _30901_, _30897_);
  or (_30904_, _30860_, _07215_);
  and (_30905_, _30904_, _30902_);
  or (_30906_, _30905_, _07460_);
  and (_30907_, _09451_, _07894_);
  or (_30908_, _30850_, _07208_);
  or (_30909_, _30908_, _30907_);
  and (_30910_, _30909_, _05982_);
  and (_30911_, _30910_, _30906_);
  and (_30912_, _14653_, _07894_);
  or (_30913_, _30912_, _30850_);
  and (_30915_, _30913_, _10094_);
  or (_30916_, _30915_, _30911_);
  and (_30917_, _30916_, _06219_);
  or (_30918_, _30917_, _30857_);
  and (_30919_, _30918_, _07237_);
  or (_30920_, _14668_, _13180_);
  and (_30921_, _30855_, _06369_);
  and (_30922_, _30921_, _30920_);
  or (_30923_, _30922_, _06536_);
  or (_30924_, _30923_, _30919_);
  and (_30926_, _11262_, _07894_);
  or (_30927_, _30926_, _30850_);
  or (_30928_, _30927_, _07240_);
  and (_30929_, _30928_, _07242_);
  and (_30930_, _30929_, _30924_);
  or (_30931_, _14666_, _13180_);
  and (_30932_, _30855_, _06375_);
  and (_30933_, _30932_, _30931_);
  or (_30934_, _30933_, _06545_);
  or (_30935_, _30934_, _30930_);
  and (_30937_, _30866_, _08341_);
  or (_30938_, _30850_, _07234_);
  or (_30939_, _30938_, _30937_);
  and (_30940_, _30939_, _09056_);
  and (_30941_, _30940_, _30935_);
  or (_30942_, _30854_, _08341_);
  and (_30943_, _30855_, _06366_);
  and (_30944_, _30943_, _30942_);
  or (_30945_, _30944_, _06528_);
  or (_30946_, _30945_, _30941_);
  and (_30948_, _30946_, _30853_);
  or (_30949_, _30948_, _06568_);
  or (_30950_, _30864_, _06926_);
  and (_30951_, _30950_, _05928_);
  and (_30952_, _30951_, _30949_);
  and (_30953_, _30888_, _05927_);
  or (_30954_, _30953_, _06278_);
  or (_30955_, _30954_, _30952_);
  or (_30956_, _30850_, _06279_);
  or (_30957_, _30956_, _30862_);
  and (_30959_, _30957_, _01347_);
  and (_30960_, _30959_, _30955_);
  nor (_30961_, \oc8051_golden_model_1.P3 [1], rst);
  nor (_30962_, _30961_, _01354_);
  or (_43272_, _30962_, _30960_);
  and (_30963_, _13180_, \oc8051_golden_model_1.P3 [2]);
  nor (_30964_, _13180_, _07776_);
  or (_30965_, _30964_, _30963_);
  or (_30966_, _30965_, _07215_);
  or (_30967_, _30965_, _07166_);
  and (_30969_, _14770_, _07894_);
  or (_30970_, _30969_, _30963_);
  or (_30971_, _30970_, _07151_);
  and (_30972_, _07894_, \oc8051_golden_model_1.ACC [2]);
  or (_30973_, _30972_, _30963_);
  and (_30974_, _30973_, _07141_);
  and (_30975_, _07142_, \oc8051_golden_model_1.P3 [2]);
  or (_30976_, _30975_, _06341_);
  or (_30977_, _30976_, _30974_);
  and (_30978_, _30977_, _06273_);
  and (_30980_, _30978_, _30971_);
  and (_30981_, _13188_, \oc8051_golden_model_1.P3 [2]);
  and (_30982_, _14774_, _08628_);
  or (_30983_, _30982_, _30981_);
  and (_30984_, _30983_, _06272_);
  or (_30985_, _30984_, _06461_);
  or (_30986_, _30985_, _30980_);
  and (_30987_, _30986_, _30967_);
  or (_30988_, _30987_, _06464_);
  or (_30989_, _30973_, _06465_);
  and (_30991_, _30989_, _06269_);
  and (_30992_, _30991_, _30988_);
  and (_30993_, _14756_, _08628_);
  or (_30994_, _30993_, _30981_);
  and (_30995_, _30994_, _06268_);
  or (_30996_, _30995_, _06261_);
  or (_30997_, _30996_, _30992_);
  and (_30998_, _30982_, _14789_);
  or (_30999_, _30981_, _06262_);
  or (_31000_, _30999_, _30998_);
  and (_31002_, _31000_, _06258_);
  and (_31003_, _31002_, _30997_);
  and (_31004_, _14804_, _08628_);
  or (_31005_, _31004_, _30981_);
  and (_31006_, _31005_, _06257_);
  or (_31007_, _31006_, _10080_);
  or (_31008_, _31007_, _31003_);
  and (_31009_, _31008_, _30966_);
  or (_31010_, _31009_, _07460_);
  and (_31011_, _09450_, _07894_);
  or (_31013_, _30963_, _07208_);
  or (_31014_, _31013_, _31011_);
  and (_31015_, _31014_, _05982_);
  and (_31016_, _31015_, _31010_);
  and (_31017_, _14859_, _07894_);
  or (_31018_, _31017_, _30963_);
  and (_31019_, _31018_, _10094_);
  or (_31020_, _31019_, _06218_);
  or (_31021_, _31020_, _31016_);
  and (_31022_, _07894_, _08973_);
  or (_31024_, _31022_, _30963_);
  or (_31025_, _31024_, _06219_);
  and (_31026_, _31025_, _31021_);
  or (_31027_, _31026_, _06369_);
  and (_31028_, _14751_, _07894_);
  or (_31029_, _31028_, _30963_);
  or (_31030_, _31029_, _07237_);
  and (_31031_, _31030_, _07240_);
  and (_31032_, _31031_, _31027_);
  and (_31033_, _11259_, _07894_);
  or (_31035_, _31033_, _30963_);
  and (_31036_, _31035_, _06536_);
  or (_31037_, _31036_, _31032_);
  and (_31038_, _31037_, _07242_);
  or (_31039_, _30963_, _08440_);
  and (_31040_, _31024_, _06375_);
  and (_31041_, _31040_, _31039_);
  or (_31042_, _31041_, _31038_);
  and (_31043_, _31042_, _07234_);
  and (_31044_, _30973_, _06545_);
  and (_31047_, _31044_, _31039_);
  or (_31048_, _31047_, _06366_);
  or (_31049_, _31048_, _31043_);
  and (_31050_, _14748_, _07894_);
  or (_31051_, _30963_, _09056_);
  or (_31052_, _31051_, _31050_);
  and (_31053_, _31052_, _09061_);
  and (_31054_, _31053_, _31049_);
  nor (_31055_, _11258_, _13180_);
  or (_31056_, _31055_, _30963_);
  and (_31058_, _31056_, _06528_);
  or (_31059_, _31058_, _06568_);
  or (_31060_, _31059_, _31054_);
  or (_31061_, _30970_, _06926_);
  and (_31062_, _31061_, _05928_);
  and (_31063_, _31062_, _31060_);
  and (_31064_, _30994_, _05927_);
  or (_31065_, _31064_, _06278_);
  or (_31066_, _31065_, _31063_);
  and (_31067_, _14926_, _07894_);
  or (_31070_, _30963_, _06279_);
  or (_31071_, _31070_, _31067_);
  and (_31072_, _31071_, _01347_);
  and (_31073_, _31072_, _31066_);
  nor (_31074_, \oc8051_golden_model_1.P3 [2], rst);
  nor (_31075_, _31074_, _01354_);
  or (_43273_, _31075_, _31073_);
  nor (_31076_, \oc8051_golden_model_1.P3 [3], rst);
  nor (_31077_, _31076_, _01354_);
  and (_31078_, _13180_, \oc8051_golden_model_1.P3 [3]);
  nor (_31080_, _13180_, _07594_);
  or (_31081_, _31080_, _31078_);
  or (_31082_, _31081_, _07215_);
  and (_31083_, _14953_, _07894_);
  or (_31084_, _31083_, _31078_);
  or (_31085_, _31084_, _07151_);
  and (_31086_, _07894_, \oc8051_golden_model_1.ACC [3]);
  or (_31087_, _31086_, _31078_);
  and (_31088_, _31087_, _07141_);
  and (_31089_, _07142_, \oc8051_golden_model_1.P3 [3]);
  or (_31092_, _31089_, _06341_);
  or (_31093_, _31092_, _31088_);
  and (_31094_, _31093_, _06273_);
  and (_31095_, _31094_, _31085_);
  and (_31096_, _13188_, \oc8051_golden_model_1.P3 [3]);
  and (_31097_, _14950_, _08628_);
  or (_31098_, _31097_, _31096_);
  and (_31099_, _31098_, _06272_);
  or (_31100_, _31099_, _06461_);
  or (_31101_, _31100_, _31095_);
  or (_31103_, _31081_, _07166_);
  and (_31104_, _31103_, _31101_);
  or (_31105_, _31104_, _06464_);
  or (_31106_, _31087_, _06465_);
  and (_31107_, _31106_, _06269_);
  and (_31108_, _31107_, _31105_);
  and (_31109_, _14948_, _08628_);
  or (_31110_, _31109_, _31096_);
  and (_31111_, _31110_, _06268_);
  or (_31112_, _31111_, _06261_);
  or (_31115_, _31112_, _31108_);
  or (_31116_, _31096_, _14979_);
  and (_31117_, _31116_, _31098_);
  or (_31118_, _31117_, _06262_);
  and (_31119_, _31118_, _06258_);
  and (_31120_, _31119_, _31115_);
  or (_31121_, _31096_, _14992_);
  and (_31122_, _31121_, _06257_);
  and (_31123_, _31122_, _31098_);
  or (_31124_, _31123_, _10080_);
  or (_31126_, _31124_, _31120_);
  and (_31127_, _31126_, _31082_);
  or (_31128_, _31127_, _07460_);
  and (_31129_, _09449_, _07894_);
  or (_31130_, _31078_, _07208_);
  or (_31131_, _31130_, _31129_);
  and (_31132_, _31131_, _05982_);
  and (_31133_, _31132_, _31128_);
  and (_31134_, _15048_, _07894_);
  or (_31135_, _31134_, _31078_);
  and (_31137_, _31135_, _10094_);
  or (_31138_, _31137_, _06218_);
  or (_31139_, _31138_, _31133_);
  and (_31140_, _07894_, _08930_);
  or (_31141_, _31140_, _31078_);
  or (_31142_, _31141_, _06219_);
  and (_31143_, _31142_, _31139_);
  or (_31144_, _31143_, _06369_);
  and (_31145_, _14943_, _07894_);
  or (_31146_, _31145_, _31078_);
  or (_31148_, _31146_, _07237_);
  and (_31149_, _31148_, _07240_);
  and (_31150_, _31149_, _31144_);
  and (_31151_, _12577_, _07894_);
  or (_31152_, _31151_, _31078_);
  and (_31153_, _31152_, _06536_);
  or (_31154_, _31153_, _31150_);
  and (_31155_, _31154_, _07242_);
  or (_31156_, _31078_, _08292_);
  and (_31157_, _31141_, _06375_);
  and (_31158_, _31157_, _31156_);
  or (_31159_, _31158_, _31155_);
  and (_31160_, _31159_, _07234_);
  and (_31161_, _31087_, _06545_);
  and (_31162_, _31161_, _31156_);
  or (_31163_, _31162_, _06366_);
  or (_31164_, _31163_, _31160_);
  and (_31165_, _14940_, _07894_);
  or (_31166_, _31078_, _09056_);
  or (_31167_, _31166_, _31165_);
  and (_31170_, _31167_, _09061_);
  and (_31171_, _31170_, _31164_);
  nor (_31172_, _11256_, _13180_);
  or (_31173_, _31172_, _31078_);
  and (_31174_, _31173_, _06528_);
  or (_31175_, _31174_, _06568_);
  or (_31176_, _31175_, _31171_);
  or (_31177_, _31084_, _06926_);
  and (_31178_, _31177_, _05928_);
  and (_31179_, _31178_, _31176_);
  and (_31180_, _31110_, _05927_);
  or (_31181_, _31180_, _06278_);
  or (_31182_, _31181_, _31179_);
  and (_31183_, _15128_, _07894_);
  or (_31184_, _31078_, _06279_);
  or (_31185_, _31184_, _31183_);
  and (_31186_, _31185_, _01347_);
  and (_31187_, _31186_, _31182_);
  or (_43274_, _31187_, _31077_);
  and (_31188_, _13180_, \oc8051_golden_model_1.P3 [4]);
  nor (_31191_, _08541_, _13180_);
  or (_31192_, _31191_, _31188_);
  or (_31193_, _31192_, _07215_);
  and (_31194_, _13188_, \oc8051_golden_model_1.P3 [4]);
  and (_31195_, _15176_, _08628_);
  or (_31196_, _31195_, _31194_);
  and (_31197_, _31196_, _06268_);
  and (_31198_, _15162_, _07894_);
  or (_31199_, _31198_, _31188_);
  or (_31200_, _31199_, _07151_);
  and (_31201_, _07894_, \oc8051_golden_model_1.ACC [4]);
  or (_31202_, _31201_, _31188_);
  and (_31203_, _31202_, _07141_);
  and (_31204_, _07142_, \oc8051_golden_model_1.P3 [4]);
  or (_31205_, _31204_, _06341_);
  or (_31206_, _31205_, _31203_);
  and (_31207_, _31206_, _06273_);
  and (_31208_, _31207_, _31200_);
  and (_31209_, _15166_, _08628_);
  or (_31210_, _31209_, _31194_);
  and (_31213_, _31210_, _06272_);
  or (_31214_, _31213_, _06461_);
  or (_31215_, _31214_, _31208_);
  or (_31216_, _31192_, _07166_);
  and (_31217_, _31216_, _31215_);
  or (_31218_, _31217_, _06464_);
  or (_31219_, _31202_, _06465_);
  and (_31220_, _31219_, _06269_);
  and (_31221_, _31220_, _31218_);
  or (_31222_, _31221_, _31197_);
  and (_31223_, _31222_, _06262_);
  and (_31224_, _15184_, _08628_);
  or (_31225_, _31224_, _31194_);
  and (_31226_, _31225_, _06261_);
  or (_31227_, _31226_, _31223_);
  and (_31228_, _31227_, _06258_);
  and (_31229_, _15200_, _08628_);
  or (_31230_, _31229_, _31194_);
  and (_31231_, _31230_, _06257_);
  or (_31232_, _31231_, _10080_);
  or (_31235_, _31232_, _31228_);
  and (_31236_, _31235_, _31193_);
  or (_31237_, _31236_, _07460_);
  and (_31238_, _09448_, _07894_);
  or (_31239_, _31188_, _07208_);
  or (_31240_, _31239_, _31238_);
  and (_31241_, _31240_, _05982_);
  and (_31242_, _31241_, _31237_);
  and (_31243_, _15254_, _07894_);
  or (_31244_, _31243_, _31188_);
  and (_31245_, _31244_, _10094_);
  or (_31246_, _31245_, _06218_);
  or (_31247_, _31246_, _31242_);
  and (_31248_, _08959_, _07894_);
  or (_31249_, _31248_, _31188_);
  or (_31250_, _31249_, _06219_);
  and (_31251_, _31250_, _31247_);
  or (_31252_, _31251_, _06369_);
  and (_31253_, _15269_, _07894_);
  or (_31254_, _31253_, _31188_);
  or (_31257_, _31254_, _07237_);
  and (_31258_, _31257_, _07240_);
  and (_31259_, _31258_, _31252_);
  and (_31260_, _11254_, _07894_);
  or (_31261_, _31260_, _31188_);
  and (_31262_, _31261_, _06536_);
  or (_31263_, _31262_, _31259_);
  and (_31264_, _31263_, _07242_);
  or (_31265_, _31188_, _08544_);
  and (_31266_, _31249_, _06375_);
  and (_31267_, _31266_, _31265_);
  or (_31268_, _31267_, _31264_);
  and (_31269_, _31268_, _07234_);
  and (_31270_, _31202_, _06545_);
  and (_31271_, _31270_, _31265_);
  or (_31272_, _31271_, _06366_);
  or (_31273_, _31272_, _31269_);
  and (_31274_, _15266_, _07894_);
  or (_31275_, _31188_, _09056_);
  or (_31276_, _31275_, _31274_);
  and (_31279_, _31276_, _09061_);
  and (_31280_, _31279_, _31273_);
  nor (_31281_, _11253_, _13180_);
  or (_31282_, _31281_, _31188_);
  and (_31283_, _31282_, _06528_);
  or (_31284_, _31283_, _06568_);
  or (_31285_, _31284_, _31280_);
  or (_31286_, _31199_, _06926_);
  and (_31287_, _31286_, _05928_);
  and (_31288_, _31287_, _31285_);
  and (_31289_, _31196_, _05927_);
  or (_31290_, _31289_, _06278_);
  or (_31291_, _31290_, _31288_);
  and (_31292_, _15329_, _07894_);
  or (_31293_, _31188_, _06279_);
  or (_31294_, _31293_, _31292_);
  and (_31295_, _31294_, _01347_);
  and (_31296_, _31295_, _31291_);
  nor (_31297_, \oc8051_golden_model_1.P3 [4], rst);
  nor (_31298_, _31297_, _01354_);
  or (_43275_, _31298_, _31296_);
  nor (_31301_, \oc8051_golden_model_1.P3 [5], rst);
  nor (_31302_, _31301_, _01354_);
  and (_31303_, _13180_, \oc8051_golden_model_1.P3 [5]);
  and (_31304_, _15358_, _07894_);
  or (_31305_, _31304_, _31303_);
  or (_31306_, _31305_, _07151_);
  and (_31307_, _07894_, \oc8051_golden_model_1.ACC [5]);
  or (_31308_, _31307_, _31303_);
  and (_31309_, _31308_, _07141_);
  and (_31310_, _07142_, \oc8051_golden_model_1.P3 [5]);
  or (_31311_, _31310_, _06341_);
  or (_31312_, _31311_, _31309_);
  and (_31313_, _31312_, _06273_);
  and (_31314_, _31313_, _31306_);
  and (_31315_, _13188_, \oc8051_golden_model_1.P3 [5]);
  and (_31316_, _15372_, _08628_);
  or (_31317_, _31316_, _31315_);
  and (_31318_, _31317_, _06272_);
  or (_31319_, _31318_, _06461_);
  or (_31322_, _31319_, _31314_);
  nor (_31323_, _08244_, _13180_);
  or (_31324_, _31323_, _31303_);
  or (_31325_, _31324_, _07166_);
  and (_31326_, _31325_, _31322_);
  or (_31327_, _31326_, _06464_);
  or (_31328_, _31308_, _06465_);
  and (_31329_, _31328_, _06269_);
  and (_31330_, _31329_, _31327_);
  and (_31331_, _15355_, _08628_);
  or (_31332_, _31331_, _31315_);
  and (_31333_, _31332_, _06268_);
  or (_31334_, _31333_, _06261_);
  or (_31335_, _31334_, _31330_);
  or (_31336_, _31315_, _15387_);
  and (_31337_, _31336_, _31317_);
  or (_31338_, _31337_, _06262_);
  and (_31339_, _31338_, _06258_);
  and (_31340_, _31339_, _31335_);
  or (_31341_, _31315_, _15403_);
  and (_31344_, _31341_, _06257_);
  and (_31345_, _31344_, _31317_);
  or (_31346_, _31345_, _10080_);
  or (_31347_, _31346_, _31340_);
  or (_31348_, _31324_, _07215_);
  and (_31349_, _31348_, _31347_);
  or (_31350_, _31349_, _07460_);
  and (_31351_, _09447_, _07894_);
  or (_31352_, _31303_, _07208_);
  or (_31353_, _31352_, _31351_);
  and (_31354_, _31353_, _05982_);
  and (_31355_, _31354_, _31350_);
  and (_31356_, _15459_, _07894_);
  or (_31357_, _31356_, _31303_);
  and (_31358_, _31357_, _10094_);
  or (_31359_, _31358_, _06218_);
  or (_31360_, _31359_, _31355_);
  and (_31361_, _08946_, _07894_);
  or (_31362_, _31361_, _31303_);
  or (_31363_, _31362_, _06219_);
  and (_31366_, _31363_, _31360_);
  or (_31367_, _31366_, _06369_);
  and (_31368_, _15353_, _07894_);
  or (_31369_, _31368_, _31303_);
  or (_31370_, _31369_, _07237_);
  and (_31371_, _31370_, _07240_);
  and (_31372_, _31371_, _31367_);
  and (_31373_, _11250_, _07894_);
  or (_31374_, _31373_, _31303_);
  and (_31375_, _31374_, _06536_);
  or (_31376_, _31375_, _31372_);
  and (_31377_, _31376_, _07242_);
  or (_31378_, _31303_, _08247_);
  and (_31379_, _31362_, _06375_);
  and (_31380_, _31379_, _31378_);
  or (_31381_, _31380_, _31377_);
  and (_31382_, _31381_, _07234_);
  and (_31383_, _31308_, _06545_);
  and (_31384_, _31383_, _31378_);
  or (_31385_, _31384_, _06366_);
  or (_31388_, _31385_, _31382_);
  and (_31389_, _15350_, _07894_);
  or (_31390_, _31303_, _09056_);
  or (_31391_, _31390_, _31389_);
  and (_31392_, _31391_, _09061_);
  and (_31393_, _31392_, _31388_);
  nor (_31394_, _11249_, _13180_);
  or (_31395_, _31394_, _31303_);
  and (_31396_, _31395_, _06528_);
  or (_31397_, _31396_, _06568_);
  or (_31398_, _31397_, _31393_);
  or (_31399_, _31305_, _06926_);
  and (_31400_, _31399_, _05928_);
  and (_31401_, _31400_, _31398_);
  and (_31402_, _31332_, _05927_);
  or (_31403_, _31402_, _06278_);
  or (_31404_, _31403_, _31401_);
  and (_31405_, _15532_, _07894_);
  or (_31406_, _31303_, _06279_);
  or (_31407_, _31406_, _31405_);
  and (_31410_, _31407_, _01347_);
  and (_31411_, _31410_, _31404_);
  or (_43276_, _31411_, _31302_);
  and (_31412_, _13180_, \oc8051_golden_model_1.P3 [6]);
  and (_31413_, _15554_, _07894_);
  or (_31414_, _31413_, _31412_);
  or (_31415_, _31414_, _07151_);
  and (_31416_, _07894_, \oc8051_golden_model_1.ACC [6]);
  or (_31417_, _31416_, _31412_);
  and (_31418_, _31417_, _07141_);
  and (_31419_, _07142_, \oc8051_golden_model_1.P3 [6]);
  or (_31420_, _31419_, _06341_);
  or (_31421_, _31420_, _31418_);
  and (_31422_, _31421_, _06273_);
  and (_31423_, _31422_, _31415_);
  and (_31424_, _13188_, \oc8051_golden_model_1.P3 [6]);
  and (_31425_, _15570_, _08628_);
  or (_31426_, _31425_, _31424_);
  and (_31427_, _31426_, _06272_);
  or (_31428_, _31427_, _06461_);
  or (_31431_, _31428_, _31423_);
  nor (_31432_, _08142_, _13180_);
  or (_31433_, _31432_, _31412_);
  or (_31434_, _31433_, _07166_);
  and (_31435_, _31434_, _31431_);
  or (_31436_, _31435_, _06464_);
  or (_31437_, _31417_, _06465_);
  and (_31438_, _31437_, _06269_);
  and (_31439_, _31438_, _31436_);
  and (_31440_, _15551_, _08628_);
  or (_31441_, _31440_, _31424_);
  and (_31442_, _31441_, _06268_);
  or (_31443_, _31442_, _06261_);
  or (_31444_, _31443_, _31439_);
  or (_31445_, _31424_, _15585_);
  and (_31446_, _31445_, _31426_);
  or (_31447_, _31446_, _06262_);
  and (_31448_, _31447_, _06258_);
  and (_31449_, _31448_, _31444_);
  and (_31450_, _15602_, _08628_);
  or (_31453_, _31450_, _31424_);
  and (_31454_, _31453_, _06257_);
  or (_31455_, _31454_, _10080_);
  or (_31456_, _31455_, _31449_);
  or (_31457_, _31433_, _07215_);
  and (_31458_, _31457_, _31456_);
  or (_31459_, _31458_, _07460_);
  and (_31460_, _09446_, _07894_);
  or (_31461_, _31412_, _07208_);
  or (_31462_, _31461_, _31460_);
  and (_31463_, _31462_, _05982_);
  and (_31464_, _31463_, _31459_);
  and (_31465_, _15657_, _07894_);
  or (_31466_, _31465_, _31412_);
  and (_31467_, _31466_, _10094_);
  or (_31468_, _31467_, _06218_);
  or (_31469_, _31468_, _31464_);
  and (_31470_, _15664_, _07894_);
  or (_31471_, _31470_, _31412_);
  or (_31472_, _31471_, _06219_);
  and (_31475_, _31472_, _31469_);
  or (_31476_, _31475_, _06369_);
  and (_31477_, _15549_, _07894_);
  or (_31478_, _31477_, _31412_);
  or (_31479_, _31478_, _07237_);
  and (_31480_, _31479_, _07240_);
  and (_31481_, _31480_, _31476_);
  and (_31482_, _11247_, _07894_);
  or (_31483_, _31482_, _31412_);
  and (_31484_, _31483_, _06536_);
  or (_31485_, _31484_, _31481_);
  and (_31486_, _31485_, _07242_);
  or (_31487_, _31412_, _08145_);
  and (_31488_, _31471_, _06375_);
  and (_31489_, _31488_, _31487_);
  or (_31490_, _31489_, _31486_);
  and (_31491_, _31490_, _07234_);
  and (_31492_, _31417_, _06545_);
  and (_31493_, _31492_, _31487_);
  or (_31494_, _31493_, _06366_);
  or (_31497_, _31494_, _31491_);
  and (_31498_, _15546_, _07894_);
  or (_31499_, _31412_, _09056_);
  or (_31500_, _31499_, _31498_);
  and (_31501_, _31500_, _09061_);
  and (_31502_, _31501_, _31497_);
  nor (_31503_, _11246_, _13180_);
  or (_31504_, _31503_, _31412_);
  and (_31505_, _31504_, _06528_);
  or (_31506_, _31505_, _06568_);
  or (_31507_, _31506_, _31502_);
  or (_31508_, _31414_, _06926_);
  and (_31509_, _31508_, _05928_);
  and (_31510_, _31509_, _31507_);
  and (_31511_, _31441_, _05927_);
  or (_31512_, _31511_, _06278_);
  or (_31513_, _31512_, _31510_);
  and (_31514_, _15734_, _07894_);
  or (_31515_, _31412_, _06279_);
  or (_31516_, _31515_, _31514_);
  and (_31519_, _31516_, _01347_);
  and (_31520_, _31519_, _31513_);
  nor (_31521_, \oc8051_golden_model_1.P3 [6], rst);
  nor (_31522_, _31521_, _01354_);
  or (_43277_, _31522_, _31520_);
  nand (_31523_, _11263_, _07926_);
  not (_31524_, \oc8051_golden_model_1.P0 [0]);
  nor (_31525_, _07926_, _31524_);
  nor (_31526_, _31525_, _07234_);
  nand (_31527_, _31526_, _31523_);
  and (_31528_, _07926_, _07133_);
  or (_31529_, _31528_, _31525_);
  or (_31530_, _31529_, _07215_);
  nor (_31531_, _08390_, _13283_);
  or (_31532_, _31531_, _31525_);
  or (_31533_, _31532_, _07151_);
  and (_31534_, _07926_, \oc8051_golden_model_1.ACC [0]);
  or (_31535_, _31534_, _31525_);
  and (_31536_, _31535_, _07141_);
  nor (_31537_, _07141_, _31524_);
  or (_31540_, _31537_, _06341_);
  or (_31541_, _31540_, _31536_);
  and (_31542_, _31541_, _06273_);
  and (_31543_, _31542_, _31533_);
  nor (_31544_, _07948_, _31524_);
  and (_31545_, _14382_, _07948_);
  or (_31546_, _31545_, _31544_);
  and (_31547_, _31546_, _06272_);
  or (_31548_, _31547_, _31543_);
  and (_31549_, _31548_, _07166_);
  and (_31550_, _31529_, _06461_);
  or (_31551_, _31550_, _06464_);
  or (_31552_, _31551_, _31549_);
  or (_31553_, _31535_, _06465_);
  and (_31554_, _31553_, _06269_);
  and (_31555_, _31554_, _31552_);
  and (_31556_, _31525_, _06268_);
  or (_31557_, _31556_, _06261_);
  or (_31558_, _31557_, _31555_);
  or (_31559_, _31532_, _06262_);
  and (_31562_, _31559_, _06258_);
  and (_31563_, _31562_, _31558_);
  and (_31564_, _14413_, _07948_);
  or (_31565_, _31564_, _31544_);
  and (_31566_, _31565_, _06257_);
  or (_31567_, _31566_, _10080_);
  or (_31568_, _31567_, _31563_);
  and (_31569_, _31568_, _31530_);
  or (_31570_, _31569_, _07460_);
  and (_31571_, _09392_, _07926_);
  or (_31572_, _31525_, _07208_);
  or (_31573_, _31572_, _31571_);
  and (_31574_, _31573_, _31570_);
  or (_31575_, _31574_, _10094_);
  and (_31576_, _14467_, _07926_);
  or (_31577_, _31525_, _05982_);
  or (_31578_, _31577_, _31576_);
  and (_31579_, _31578_, _06219_);
  and (_31580_, _31579_, _31575_);
  and (_31581_, _07926_, _08954_);
  or (_31584_, _31581_, _31525_);
  and (_31585_, _31584_, _06218_);
  or (_31586_, _31585_, _06369_);
  or (_31587_, _31586_, _31580_);
  and (_31588_, _14366_, _07926_);
  or (_31589_, _31588_, _31525_);
  or (_31590_, _31589_, _07237_);
  and (_31591_, _31590_, _07240_);
  and (_31592_, _31591_, _31587_);
  nor (_31593_, _12580_, _13283_);
  or (_31594_, _31593_, _31525_);
  and (_31595_, _31523_, _06536_);
  and (_31596_, _31595_, _31594_);
  or (_31597_, _31596_, _31592_);
  and (_31598_, _31597_, _07242_);
  nand (_31599_, _31584_, _06375_);
  nor (_31600_, _31599_, _31531_);
  or (_31601_, _31600_, _06545_);
  or (_31602_, _31601_, _31598_);
  and (_31603_, _31602_, _31527_);
  or (_31606_, _31603_, _06366_);
  and (_31607_, _14363_, _07926_);
  or (_31608_, _31607_, _31525_);
  or (_31609_, _31608_, _09056_);
  and (_31610_, _31609_, _09061_);
  and (_31611_, _31610_, _31606_);
  and (_31612_, _31594_, _06528_);
  or (_31613_, _31612_, _06568_);
  or (_31614_, _31613_, _31611_);
  or (_31615_, _31532_, _06926_);
  and (_31616_, _31615_, _31614_);
  or (_31617_, _31616_, _05927_);
  or (_31618_, _31525_, _05928_);
  and (_31619_, _31618_, _31617_);
  or (_31620_, _31619_, _06278_);
  or (_31621_, _31532_, _06279_);
  and (_31622_, _31621_, _01347_);
  and (_31623_, _31622_, _31620_);
  nor (_31624_, \oc8051_golden_model_1.P0 [0], rst);
  nor (_31625_, _31624_, _01354_);
  or (_43279_, _31625_, _31623_);
  nor (_31628_, \oc8051_golden_model_1.P0 [1], rst);
  nor (_31629_, _31628_, _01354_);
  not (_31630_, \oc8051_golden_model_1.P0 [1]);
  nor (_31631_, _07926_, _31630_);
  nor (_31632_, _11261_, _13283_);
  or (_31633_, _31632_, _31631_);
  or (_31634_, _31633_, _09061_);
  nor (_31635_, _13283_, _07357_);
  or (_31636_, _31635_, _31631_);
  or (_31637_, _31636_, _07166_);
  or (_31638_, _07926_, \oc8051_golden_model_1.P0 [1]);
  and (_31639_, _14562_, _07926_);
  not (_31640_, _31639_);
  and (_31641_, _31640_, _31638_);
  or (_31642_, _31641_, _07151_);
  and (_31643_, _07926_, \oc8051_golden_model_1.ACC [1]);
  or (_31644_, _31643_, _31631_);
  and (_31645_, _31644_, _07141_);
  nor (_31646_, _07141_, _31630_);
  or (_31649_, _31646_, _06341_);
  or (_31650_, _31649_, _31645_);
  and (_31651_, _31650_, _06273_);
  and (_31652_, _31651_, _31642_);
  nor (_31653_, _07948_, _31630_);
  and (_31654_, _14557_, _07948_);
  or (_31655_, _31654_, _31653_);
  and (_31656_, _31655_, _06272_);
  or (_31657_, _31656_, _06461_);
  or (_31658_, _31657_, _31652_);
  and (_31659_, _31658_, _31637_);
  or (_31660_, _31659_, _06464_);
  or (_31661_, _31644_, _06465_);
  and (_31662_, _31661_, _06269_);
  and (_31663_, _31662_, _31660_);
  and (_31664_, _14560_, _07948_);
  or (_31665_, _31664_, _31653_);
  and (_31666_, _31665_, _06268_);
  or (_31667_, _31666_, _06261_);
  or (_31668_, _31667_, _31663_);
  and (_31671_, _31654_, _14556_);
  or (_31672_, _31653_, _06262_);
  or (_31673_, _31672_, _31671_);
  and (_31674_, _31673_, _06258_);
  and (_31675_, _31674_, _31668_);
  or (_31676_, _31653_, _14597_);
  and (_31677_, _31676_, _06257_);
  and (_31678_, _31677_, _31655_);
  or (_31679_, _31678_, _10080_);
  or (_31680_, _31679_, _31675_);
  or (_31681_, _31636_, _07215_);
  and (_31682_, _31681_, _31680_);
  or (_31683_, _31682_, _07460_);
  and (_31684_, _09451_, _07926_);
  or (_31685_, _31631_, _07208_);
  or (_31686_, _31685_, _31684_);
  and (_31687_, _31686_, _05982_);
  and (_31688_, _31687_, _31683_);
  and (_31689_, _14653_, _07926_);
  or (_31690_, _31689_, _31631_);
  and (_31693_, _31690_, _10094_);
  or (_31694_, _31693_, _31688_);
  and (_31695_, _31694_, _06219_);
  nand (_31696_, _07926_, _07038_);
  and (_31697_, _31638_, _06218_);
  and (_31698_, _31697_, _31696_);
  or (_31699_, _31698_, _31695_);
  and (_31700_, _31699_, _07237_);
  or (_31701_, _14668_, _13283_);
  and (_31702_, _31638_, _06369_);
  and (_31703_, _31702_, _31701_);
  or (_31704_, _31703_, _06536_);
  or (_31705_, _31704_, _31700_);
  nand (_31706_, _11260_, _07926_);
  and (_31707_, _31706_, _31633_);
  or (_31708_, _31707_, _07240_);
  and (_31709_, _31708_, _07242_);
  and (_31710_, _31709_, _31705_);
  or (_31711_, _14666_, _13283_);
  and (_31712_, _31638_, _06375_);
  and (_31715_, _31712_, _31711_);
  or (_31716_, _31715_, _06545_);
  or (_31717_, _31716_, _31710_);
  nor (_31718_, _31631_, _07234_);
  nand (_31719_, _31718_, _31706_);
  and (_31720_, _31719_, _09056_);
  and (_31721_, _31720_, _31717_);
  or (_31722_, _31696_, _08341_);
  and (_31723_, _31638_, _06366_);
  and (_31724_, _31723_, _31722_);
  or (_31725_, _31724_, _06528_);
  or (_31726_, _31725_, _31721_);
  and (_31727_, _31726_, _31634_);
  or (_31728_, _31727_, _06568_);
  or (_31729_, _31641_, _06926_);
  and (_31730_, _31729_, _05928_);
  and (_31731_, _31730_, _31728_);
  and (_31732_, _31665_, _05927_);
  or (_31733_, _31732_, _06278_);
  or (_31734_, _31733_, _31731_);
  or (_31737_, _31631_, _06279_);
  or (_31738_, _31737_, _31639_);
  and (_31739_, _31738_, _01347_);
  and (_31740_, _31739_, _31734_);
  or (_43280_, _31740_, _31629_);
  and (_31741_, _13283_, \oc8051_golden_model_1.P0 [2]);
  nor (_31742_, _13283_, _07776_);
  or (_31743_, _31742_, _31741_);
  or (_31744_, _31743_, _07215_);
  or (_31745_, _31743_, _07166_);
  and (_31746_, _14770_, _07926_);
  or (_31747_, _31746_, _31741_);
  or (_31748_, _31747_, _07151_);
  and (_31749_, _07926_, \oc8051_golden_model_1.ACC [2]);
  or (_31750_, _31749_, _31741_);
  and (_31751_, _31750_, _07141_);
  and (_31752_, _07142_, \oc8051_golden_model_1.P0 [2]);
  or (_31753_, _31752_, _06341_);
  or (_31754_, _31753_, _31751_);
  and (_31755_, _31754_, _06273_);
  and (_31758_, _31755_, _31748_);
  and (_31759_, _13291_, \oc8051_golden_model_1.P0 [2]);
  and (_31760_, _14774_, _07948_);
  or (_31761_, _31760_, _31759_);
  and (_31762_, _31761_, _06272_);
  or (_31763_, _31762_, _06461_);
  or (_31764_, _31763_, _31758_);
  and (_31765_, _31764_, _31745_);
  or (_31766_, _31765_, _06464_);
  or (_31767_, _31750_, _06465_);
  and (_31769_, _31767_, _06269_);
  and (_31770_, _31769_, _31766_);
  and (_31771_, _14756_, _07948_);
  or (_31772_, _31771_, _31759_);
  and (_31773_, _31772_, _06268_);
  or (_31774_, _31773_, _06261_);
  or (_31775_, _31774_, _31770_);
  and (_31776_, _31760_, _14789_);
  or (_31777_, _31759_, _06262_);
  or (_31778_, _31777_, _31776_);
  and (_31780_, _31778_, _06258_);
  and (_31781_, _31780_, _31775_);
  and (_31782_, _14804_, _07948_);
  or (_31783_, _31782_, _31759_);
  and (_31784_, _31783_, _06257_);
  or (_31785_, _31784_, _10080_);
  or (_31786_, _31785_, _31781_);
  and (_31787_, _31786_, _31744_);
  or (_31788_, _31787_, _07460_);
  and (_31789_, _09450_, _07926_);
  or (_31791_, _31741_, _07208_);
  or (_31792_, _31791_, _31789_);
  and (_31793_, _31792_, _05982_);
  and (_31794_, _31793_, _31788_);
  and (_31795_, _14859_, _07926_);
  or (_31796_, _31795_, _31741_);
  and (_31797_, _31796_, _10094_);
  or (_31798_, _31797_, _06218_);
  or (_31799_, _31798_, _31794_);
  and (_31800_, _07926_, _08973_);
  or (_31802_, _31800_, _31741_);
  or (_31803_, _31802_, _06219_);
  and (_31804_, _31803_, _31799_);
  or (_31805_, _31804_, _06369_);
  and (_31806_, _14751_, _07926_);
  or (_31807_, _31806_, _31741_);
  or (_31808_, _31807_, _07237_);
  and (_31809_, _31808_, _07240_);
  and (_31810_, _31809_, _31805_);
  and (_31811_, _11259_, _07926_);
  or (_31813_, _31811_, _31741_);
  and (_31814_, _31813_, _06536_);
  or (_31815_, _31814_, _31810_);
  and (_31816_, _31815_, _07242_);
  or (_31817_, _31741_, _08440_);
  and (_31818_, _31802_, _06375_);
  and (_31819_, _31818_, _31817_);
  or (_31820_, _31819_, _31816_);
  and (_31821_, _31820_, _07234_);
  and (_31822_, _31750_, _06545_);
  and (_31824_, _31822_, _31817_);
  or (_31825_, _31824_, _06366_);
  or (_31826_, _31825_, _31821_);
  and (_31827_, _14748_, _07926_);
  or (_31828_, _31741_, _09056_);
  or (_31829_, _31828_, _31827_);
  and (_31830_, _31829_, _09061_);
  and (_31831_, _31830_, _31826_);
  nor (_31832_, _11258_, _13283_);
  or (_31833_, _31832_, _31741_);
  and (_31835_, _31833_, _06528_);
  or (_31836_, _31835_, _06568_);
  or (_31837_, _31836_, _31831_);
  or (_31838_, _31747_, _06926_);
  and (_31839_, _31838_, _05928_);
  and (_31840_, _31839_, _31837_);
  and (_31841_, _31772_, _05927_);
  or (_31842_, _31841_, _06278_);
  or (_31843_, _31842_, _31840_);
  and (_31844_, _14926_, _07926_);
  or (_31846_, _31741_, _06279_);
  or (_31847_, _31846_, _31844_);
  and (_31848_, _31847_, _01347_);
  and (_31849_, _31848_, _31843_);
  nor (_31850_, \oc8051_golden_model_1.P0 [2], rst);
  nor (_31851_, _31850_, _01354_);
  or (_43281_, _31851_, _31849_);
  and (_31852_, _13283_, \oc8051_golden_model_1.P0 [3]);
  nor (_31853_, _13283_, _07594_);
  or (_31854_, _31853_, _31852_);
  or (_31856_, _31854_, _07215_);
  and (_31857_, _14953_, _07926_);
  or (_31858_, _31857_, _31852_);
  or (_31859_, _31858_, _07151_);
  and (_31860_, _07926_, \oc8051_golden_model_1.ACC [3]);
  or (_31861_, _31860_, _31852_);
  and (_31862_, _31861_, _07141_);
  and (_31863_, _07142_, \oc8051_golden_model_1.P0 [3]);
  or (_31864_, _31863_, _06341_);
  or (_31865_, _31864_, _31862_);
  and (_31867_, _31865_, _06273_);
  and (_31868_, _31867_, _31859_);
  and (_31869_, _13291_, \oc8051_golden_model_1.P0 [3]);
  and (_31870_, _14950_, _07948_);
  or (_31871_, _31870_, _31869_);
  and (_31872_, _31871_, _06272_);
  or (_31873_, _31872_, _06461_);
  or (_31874_, _31873_, _31868_);
  or (_31875_, _31854_, _07166_);
  and (_31876_, _31875_, _31874_);
  or (_31878_, _31876_, _06464_);
  or (_31879_, _31861_, _06465_);
  and (_31880_, _31879_, _06269_);
  and (_31881_, _31880_, _31878_);
  and (_31882_, _14948_, _07948_);
  or (_31883_, _31882_, _31869_);
  and (_31884_, _31883_, _06268_);
  or (_31885_, _31884_, _06261_);
  or (_31886_, _31885_, _31881_);
  or (_31887_, _31869_, _14979_);
  and (_31889_, _31887_, _31871_);
  or (_31890_, _31889_, _06262_);
  and (_31891_, _31890_, _06258_);
  and (_31892_, _31891_, _31886_);
  or (_31893_, _31869_, _14992_);
  and (_31894_, _31893_, _06257_);
  and (_31895_, _31894_, _31871_);
  or (_31896_, _31895_, _10080_);
  or (_31897_, _31896_, _31892_);
  and (_31898_, _31897_, _31856_);
  or (_31900_, _31898_, _07460_);
  and (_31901_, _09449_, _07926_);
  or (_31902_, _31852_, _07208_);
  or (_31903_, _31902_, _31901_);
  and (_31904_, _31903_, _05982_);
  and (_31905_, _31904_, _31900_);
  and (_31906_, _15048_, _07926_);
  or (_31907_, _31906_, _31852_);
  and (_31908_, _31907_, _10094_);
  or (_31909_, _31908_, _06218_);
  or (_31911_, _31909_, _31905_);
  and (_31912_, _07926_, _08930_);
  or (_31913_, _31912_, _31852_);
  or (_31914_, _31913_, _06219_);
  and (_31915_, _31914_, _31911_);
  or (_31916_, _31915_, _06369_);
  and (_31917_, _14943_, _07926_);
  or (_31918_, _31917_, _31852_);
  or (_31919_, _31918_, _07237_);
  and (_31920_, _31919_, _07240_);
  and (_31922_, _31920_, _31916_);
  and (_31923_, _12577_, _07926_);
  or (_31924_, _31923_, _31852_);
  and (_31925_, _31924_, _06536_);
  or (_31926_, _31925_, _31922_);
  and (_31927_, _31926_, _07242_);
  or (_31928_, _31852_, _08292_);
  and (_31929_, _31913_, _06375_);
  and (_31930_, _31929_, _31928_);
  or (_31931_, _31930_, _31927_);
  and (_31933_, _31931_, _07234_);
  and (_31934_, _31861_, _06545_);
  and (_31935_, _31934_, _31928_);
  or (_31936_, _31935_, _06366_);
  or (_31937_, _31936_, _31933_);
  and (_31938_, _14940_, _07926_);
  or (_31939_, _31852_, _09056_);
  or (_31940_, _31939_, _31938_);
  and (_31941_, _31940_, _09061_);
  and (_31942_, _31941_, _31937_);
  nor (_31944_, _11256_, _13283_);
  or (_31945_, _31944_, _31852_);
  and (_31946_, _31945_, _06528_);
  or (_31947_, _31946_, _06568_);
  or (_31948_, _31947_, _31942_);
  or (_31949_, _31858_, _06926_);
  and (_31950_, _31949_, _05928_);
  and (_31951_, _31950_, _31948_);
  and (_31952_, _31883_, _05927_);
  or (_31953_, _31952_, _06278_);
  or (_31954_, _31953_, _31951_);
  and (_31955_, _15128_, _07926_);
  or (_31956_, _31852_, _06279_);
  or (_31957_, _31956_, _31955_);
  and (_31958_, _31957_, _01347_);
  and (_31959_, _31958_, _31954_);
  nor (_31960_, \oc8051_golden_model_1.P0 [3], rst);
  nor (_31961_, _31960_, _01354_);
  or (_43283_, _31961_, _31959_);
  nor (_31962_, \oc8051_golden_model_1.P0 [4], rst);
  nor (_31964_, _31962_, _01354_);
  and (_31965_, _13283_, \oc8051_golden_model_1.P0 [4]);
  nor (_31966_, _08541_, _13283_);
  or (_31967_, _31966_, _31965_);
  or (_31968_, _31967_, _07215_);
  and (_31969_, _13291_, \oc8051_golden_model_1.P0 [4]);
  and (_31970_, _15176_, _07948_);
  or (_31971_, _31970_, _31969_);
  and (_31972_, _31971_, _06268_);
  and (_31973_, _15162_, _07926_);
  or (_31975_, _31973_, _31965_);
  or (_31976_, _31975_, _07151_);
  and (_31977_, _07926_, \oc8051_golden_model_1.ACC [4]);
  or (_31978_, _31977_, _31965_);
  and (_31979_, _31978_, _07141_);
  and (_31980_, _07142_, \oc8051_golden_model_1.P0 [4]);
  or (_31981_, _31980_, _06341_);
  or (_31982_, _31981_, _31979_);
  and (_31983_, _31982_, _06273_);
  and (_31984_, _31983_, _31976_);
  and (_31986_, _15166_, _07948_);
  or (_31987_, _31986_, _31969_);
  and (_31988_, _31987_, _06272_);
  or (_31989_, _31988_, _06461_);
  or (_31990_, _31989_, _31984_);
  or (_31991_, _31967_, _07166_);
  and (_31992_, _31991_, _31990_);
  or (_31993_, _31992_, _06464_);
  or (_31994_, _31978_, _06465_);
  and (_31995_, _31994_, _06269_);
  and (_31997_, _31995_, _31993_);
  or (_31998_, _31997_, _31972_);
  and (_31999_, _31998_, _06262_);
  and (_32000_, _15184_, _07948_);
  or (_32001_, _32000_, _31969_);
  and (_32002_, _32001_, _06261_);
  or (_32003_, _32002_, _31999_);
  and (_32004_, _32003_, _06258_);
  and (_32005_, _15200_, _07948_);
  or (_32006_, _32005_, _31969_);
  and (_32008_, _32006_, _06257_);
  or (_32009_, _32008_, _10080_);
  or (_32010_, _32009_, _32004_);
  and (_32011_, _32010_, _31968_);
  or (_32012_, _32011_, _07460_);
  and (_32013_, _09448_, _07926_);
  or (_32014_, _31965_, _07208_);
  or (_32015_, _32014_, _32013_);
  and (_32016_, _32015_, _05982_);
  and (_32017_, _32016_, _32012_);
  and (_32019_, _15254_, _07926_);
  or (_32020_, _32019_, _31965_);
  and (_32021_, _32020_, _10094_);
  or (_32022_, _32021_, _06218_);
  or (_32023_, _32022_, _32017_);
  and (_32024_, _08959_, _07926_);
  or (_32025_, _32024_, _31965_);
  or (_32026_, _32025_, _06219_);
  and (_32027_, _32026_, _32023_);
  or (_32028_, _32027_, _06369_);
  and (_32030_, _15269_, _07926_);
  or (_32031_, _32030_, _31965_);
  or (_32032_, _32031_, _07237_);
  and (_32033_, _32032_, _07240_);
  and (_32034_, _32033_, _32028_);
  and (_32035_, _11254_, _07926_);
  or (_32036_, _32035_, _31965_);
  and (_32037_, _32036_, _06536_);
  or (_32038_, _32037_, _32034_);
  and (_32039_, _32038_, _07242_);
  or (_32041_, _31965_, _08544_);
  and (_32042_, _32025_, _06375_);
  and (_32043_, _32042_, _32041_);
  or (_32044_, _32043_, _32039_);
  and (_32045_, _32044_, _07234_);
  and (_32046_, _31978_, _06545_);
  and (_32047_, _32046_, _32041_);
  or (_32048_, _32047_, _06366_);
  or (_32049_, _32048_, _32045_);
  and (_32050_, _15266_, _07926_);
  or (_32052_, _31965_, _09056_);
  or (_32053_, _32052_, _32050_);
  and (_32054_, _32053_, _09061_);
  and (_32055_, _32054_, _32049_);
  nor (_32056_, _11253_, _13283_);
  or (_32057_, _32056_, _31965_);
  and (_32058_, _32057_, _06528_);
  or (_32059_, _32058_, _06568_);
  or (_32060_, _32059_, _32055_);
  or (_32061_, _31975_, _06926_);
  and (_32063_, _32061_, _05928_);
  and (_32064_, _32063_, _32060_);
  and (_32065_, _31971_, _05927_);
  or (_32066_, _32065_, _06278_);
  or (_32067_, _32066_, _32064_);
  and (_32068_, _15329_, _07926_);
  or (_32069_, _31965_, _06279_);
  or (_32070_, _32069_, _32068_);
  and (_32071_, _32070_, _01347_);
  and (_32072_, _32071_, _32067_);
  or (_43284_, _32072_, _31964_);
  and (_32074_, _13283_, \oc8051_golden_model_1.P0 [5]);
  and (_32075_, _15358_, _07926_);
  or (_32076_, _32075_, _32074_);
  or (_32077_, _32076_, _07151_);
  and (_32078_, _07926_, \oc8051_golden_model_1.ACC [5]);
  or (_32079_, _32078_, _32074_);
  and (_32080_, _32079_, _07141_);
  and (_32081_, _07142_, \oc8051_golden_model_1.P0 [5]);
  or (_32082_, _32081_, _06341_);
  or (_32084_, _32082_, _32080_);
  and (_32085_, _32084_, _06273_);
  and (_32086_, _32085_, _32077_);
  and (_32087_, _13291_, \oc8051_golden_model_1.P0 [5]);
  and (_32088_, _15372_, _07948_);
  or (_32089_, _32088_, _32087_);
  and (_32090_, _32089_, _06272_);
  or (_32091_, _32090_, _06461_);
  or (_32092_, _32091_, _32086_);
  nor (_32093_, _08244_, _13283_);
  or (_32095_, _32093_, _32074_);
  or (_32096_, _32095_, _07166_);
  and (_32097_, _32096_, _32092_);
  or (_32098_, _32097_, _06464_);
  or (_32099_, _32079_, _06465_);
  and (_32100_, _32099_, _06269_);
  and (_32101_, _32100_, _32098_);
  and (_32102_, _15355_, _07948_);
  or (_32103_, _32102_, _32087_);
  and (_32104_, _32103_, _06268_);
  or (_32106_, _32104_, _06261_);
  or (_32107_, _32106_, _32101_);
  or (_32108_, _32087_, _15387_);
  and (_32109_, _32108_, _32089_);
  or (_32110_, _32109_, _06262_);
  and (_32111_, _32110_, _06258_);
  and (_32112_, _32111_, _32107_);
  or (_32113_, _32087_, _15403_);
  and (_32114_, _32113_, _06257_);
  and (_32115_, _32114_, _32089_);
  or (_32117_, _32115_, _10080_);
  or (_32118_, _32117_, _32112_);
  or (_32119_, _32095_, _07215_);
  and (_32120_, _32119_, _32118_);
  or (_32121_, _32120_, _07460_);
  and (_32122_, _09447_, _07926_);
  or (_32123_, _32074_, _07208_);
  or (_32124_, _32123_, _32122_);
  and (_32125_, _32124_, _05982_);
  and (_32126_, _32125_, _32121_);
  and (_32128_, _15459_, _07926_);
  or (_32129_, _32128_, _32074_);
  and (_32130_, _32129_, _10094_);
  or (_32131_, _32130_, _06218_);
  or (_32132_, _32131_, _32126_);
  and (_32133_, _08946_, _07926_);
  or (_32134_, _32133_, _32074_);
  or (_32135_, _32134_, _06219_);
  and (_32136_, _32135_, _32132_);
  or (_32137_, _32136_, _06369_);
  and (_32139_, _15353_, _07926_);
  or (_32140_, _32139_, _32074_);
  or (_32141_, _32140_, _07237_);
  and (_32142_, _32141_, _07240_);
  and (_32143_, _32142_, _32137_);
  and (_32144_, _11250_, _07926_);
  or (_32145_, _32144_, _32074_);
  and (_32146_, _32145_, _06536_);
  or (_32147_, _32146_, _32143_);
  and (_32148_, _32147_, _07242_);
  or (_32150_, _32074_, _08247_);
  and (_32151_, _32134_, _06375_);
  and (_32152_, _32151_, _32150_);
  or (_32153_, _32152_, _32148_);
  and (_32154_, _32153_, _07234_);
  and (_32155_, _32079_, _06545_);
  and (_32156_, _32155_, _32150_);
  or (_32157_, _32156_, _06366_);
  or (_32158_, _32157_, _32154_);
  and (_32159_, _15350_, _07926_);
  or (_32161_, _32074_, _09056_);
  or (_32162_, _32161_, _32159_);
  and (_32163_, _32162_, _09061_);
  and (_32164_, _32163_, _32158_);
  nor (_32165_, _11249_, _13283_);
  or (_32166_, _32165_, _32074_);
  and (_32167_, _32166_, _06528_);
  or (_32168_, _32167_, _06568_);
  or (_32169_, _32168_, _32164_);
  or (_32170_, _32076_, _06926_);
  and (_32172_, _32170_, _05928_);
  and (_32173_, _32172_, _32169_);
  and (_32174_, _32103_, _05927_);
  or (_32175_, _32174_, _06278_);
  or (_32176_, _32175_, _32173_);
  and (_32177_, _15532_, _07926_);
  or (_32178_, _32074_, _06279_);
  or (_32179_, _32178_, _32177_);
  and (_32180_, _32179_, _01347_);
  and (_32181_, _32180_, _32176_);
  nor (_32183_, \oc8051_golden_model_1.P0 [5], rst);
  nor (_32184_, _32183_, _01354_);
  or (_43285_, _32184_, _32181_);
  and (_32185_, _13283_, \oc8051_golden_model_1.P0 [6]);
  and (_32186_, _15554_, _07926_);
  or (_32187_, _32186_, _32185_);
  or (_32188_, _32187_, _07151_);
  and (_32189_, _07926_, \oc8051_golden_model_1.ACC [6]);
  or (_32190_, _32189_, _32185_);
  and (_32191_, _32190_, _07141_);
  and (_32193_, _07142_, \oc8051_golden_model_1.P0 [6]);
  or (_32194_, _32193_, _06341_);
  or (_32195_, _32194_, _32191_);
  and (_32196_, _32195_, _06273_);
  and (_32197_, _32196_, _32188_);
  and (_32198_, _13291_, \oc8051_golden_model_1.P0 [6]);
  and (_32199_, _15570_, _07948_);
  or (_32200_, _32199_, _32198_);
  and (_32201_, _32200_, _06272_);
  or (_32202_, _32201_, _06461_);
  or (_32204_, _32202_, _32197_);
  nor (_32205_, _08142_, _13283_);
  or (_32206_, _32205_, _32185_);
  or (_32207_, _32206_, _07166_);
  and (_32208_, _32207_, _32204_);
  or (_32209_, _32208_, _06464_);
  or (_32210_, _32190_, _06465_);
  and (_32211_, _32210_, _06269_);
  and (_32212_, _32211_, _32209_);
  and (_32213_, _15551_, _07948_);
  or (_32215_, _32213_, _32198_);
  and (_32216_, _32215_, _06268_);
  or (_32217_, _32216_, _06261_);
  or (_32218_, _32217_, _32212_);
  or (_32219_, _32198_, _15585_);
  and (_32220_, _32219_, _32200_);
  or (_32221_, _32220_, _06262_);
  and (_32222_, _32221_, _06258_);
  and (_32223_, _32222_, _32218_);
  and (_32224_, _15602_, _07948_);
  or (_32226_, _32224_, _32198_);
  and (_32227_, _32226_, _06257_);
  or (_32228_, _32227_, _10080_);
  or (_32229_, _32228_, _32223_);
  or (_32230_, _32206_, _07215_);
  and (_32231_, _32230_, _32229_);
  or (_32232_, _32231_, _07460_);
  and (_32233_, _09446_, _07926_);
  or (_32234_, _32185_, _07208_);
  or (_32235_, _32234_, _32233_);
  and (_32237_, _32235_, _05982_);
  and (_32238_, _32237_, _32232_);
  and (_32239_, _15657_, _07926_);
  or (_32240_, _32239_, _32185_);
  and (_32241_, _32240_, _10094_);
  or (_32242_, _32241_, _06218_);
  or (_32243_, _32242_, _32238_);
  and (_32244_, _15664_, _07926_);
  or (_32245_, _32244_, _32185_);
  or (_32246_, _32245_, _06219_);
  and (_32248_, _32246_, _32243_);
  or (_32249_, _32248_, _06369_);
  and (_32250_, _15549_, _07926_);
  or (_32251_, _32250_, _32185_);
  or (_32252_, _32251_, _07237_);
  and (_32253_, _32252_, _07240_);
  and (_32254_, _32253_, _32249_);
  and (_32255_, _11247_, _07926_);
  or (_32256_, _32255_, _32185_);
  and (_32257_, _32256_, _06536_);
  or (_32259_, _32257_, _32254_);
  and (_32260_, _32259_, _07242_);
  or (_32261_, _32185_, _08145_);
  and (_32262_, _32245_, _06375_);
  and (_32263_, _32262_, _32261_);
  or (_32264_, _32263_, _32260_);
  and (_32265_, _32264_, _07234_);
  and (_32266_, _32190_, _06545_);
  and (_32267_, _32266_, _32261_);
  or (_32268_, _32267_, _06366_);
  or (_32270_, _32268_, _32265_);
  and (_32271_, _15546_, _07926_);
  or (_32272_, _32185_, _09056_);
  or (_32273_, _32272_, _32271_);
  and (_32274_, _32273_, _09061_);
  and (_32275_, _32274_, _32270_);
  nor (_32276_, _11246_, _13283_);
  or (_32277_, _32276_, _32185_);
  and (_32278_, _32277_, _06528_);
  or (_32279_, _32278_, _06568_);
  or (_32281_, _32279_, _32275_);
  or (_32282_, _32187_, _06926_);
  and (_32283_, _32282_, _05928_);
  and (_32284_, _32283_, _32281_);
  and (_32285_, _32215_, _05927_);
  or (_32286_, _32285_, _06278_);
  or (_32287_, _32286_, _32284_);
  and (_32288_, _15734_, _07926_);
  or (_32289_, _32185_, _06279_);
  or (_32290_, _32289_, _32288_);
  and (_32292_, _32290_, _01347_);
  and (_32293_, _32292_, _32287_);
  nor (_32294_, \oc8051_golden_model_1.P0 [6], rst);
  nor (_32295_, _32294_, _01354_);
  or (_43286_, _32295_, _32293_);
  nor (_32296_, \oc8051_golden_model_1.P1 [0], rst);
  nor (_32297_, _32296_, _01354_);
  nand (_32298_, _11263_, _07971_);
  and (_32299_, _13388_, \oc8051_golden_model_1.P1 [0]);
  nor (_32300_, _32299_, _07234_);
  nand (_32302_, _32300_, _32298_);
  and (_32303_, _07971_, _07133_);
  or (_32304_, _32303_, _32299_);
  or (_32305_, _32304_, _07215_);
  nor (_32306_, _08390_, _13388_);
  or (_32307_, _32306_, _32299_);
  and (_32308_, _32307_, _06341_);
  and (_32309_, _07142_, \oc8051_golden_model_1.P1 [0]);
  and (_32310_, _07971_, \oc8051_golden_model_1.ACC [0]);
  or (_32311_, _32310_, _32299_);
  and (_32313_, _32311_, _07141_);
  or (_32314_, _32313_, _32309_);
  and (_32315_, _32314_, _07151_);
  or (_32316_, _32315_, _06272_);
  or (_32317_, _32316_, _32308_);
  and (_32318_, _14382_, _08620_);
  and (_32319_, _13396_, \oc8051_golden_model_1.P1 [0]);
  or (_32320_, _32319_, _06273_);
  or (_32321_, _32320_, _32318_);
  and (_32322_, _32321_, _07166_);
  and (_32324_, _32322_, _32317_);
  and (_32325_, _32304_, _06461_);
  or (_32326_, _32325_, _06464_);
  or (_32327_, _32326_, _32324_);
  or (_32328_, _32311_, _06465_);
  and (_32329_, _32328_, _06269_);
  and (_32330_, _32329_, _32327_);
  and (_32331_, _32299_, _06268_);
  or (_32332_, _32331_, _06261_);
  or (_32333_, _32332_, _32330_);
  or (_32335_, _32307_, _06262_);
  and (_32336_, _32335_, _06258_);
  and (_32337_, _32336_, _32333_);
  and (_32338_, _14413_, _08620_);
  or (_32339_, _32338_, _32319_);
  and (_32340_, _32339_, _06257_);
  or (_32341_, _32340_, _10080_);
  or (_32342_, _32341_, _32337_);
  and (_32343_, _32342_, _32305_);
  or (_32344_, _32343_, _07460_);
  and (_32346_, _09392_, _07971_);
  or (_32347_, _32299_, _07208_);
  or (_32348_, _32347_, _32346_);
  and (_32349_, _32348_, _32344_);
  or (_32350_, _32349_, _10094_);
  and (_32351_, _14467_, _07971_);
  or (_32352_, _32299_, _05982_);
  or (_32353_, _32352_, _32351_);
  and (_32354_, _32353_, _06219_);
  and (_32355_, _32354_, _32350_);
  and (_32357_, _07971_, _08954_);
  or (_32358_, _32357_, _32299_);
  and (_32359_, _32358_, _06218_);
  or (_32360_, _32359_, _06369_);
  or (_32361_, _32360_, _32355_);
  and (_32362_, _14366_, _07971_);
  or (_32363_, _32362_, _32299_);
  or (_32364_, _32363_, _07237_);
  and (_32365_, _32364_, _07240_);
  and (_32366_, _32365_, _32361_);
  nor (_32368_, _12580_, _13388_);
  or (_32369_, _32368_, _32299_);
  and (_32370_, _32298_, _06536_);
  and (_32371_, _32370_, _32369_);
  or (_32372_, _32371_, _32366_);
  and (_32373_, _32372_, _07242_);
  nand (_32374_, _32358_, _06375_);
  nor (_32375_, _32374_, _32306_);
  or (_32376_, _32375_, _06545_);
  or (_32377_, _32376_, _32373_);
  and (_32379_, _32377_, _32302_);
  or (_32380_, _32379_, _06366_);
  and (_32381_, _14363_, _07971_);
  or (_32382_, _32299_, _09056_);
  or (_32383_, _32382_, _32381_);
  and (_32384_, _32383_, _09061_);
  and (_32385_, _32384_, _32380_);
  and (_32386_, _32369_, _06528_);
  or (_32387_, _32386_, _06568_);
  or (_32388_, _32387_, _32385_);
  or (_32390_, _32307_, _06926_);
  and (_32391_, _32390_, _32388_);
  or (_32392_, _32391_, _05927_);
  or (_32393_, _32299_, _05928_);
  and (_32394_, _32393_, _32392_);
  or (_32395_, _32394_, _06278_);
  or (_32396_, _32307_, _06279_);
  and (_32397_, _32396_, _01347_);
  and (_32398_, _32397_, _32395_);
  or (_43288_, _32398_, _32297_);
  and (_32400_, _13388_, \oc8051_golden_model_1.P1 [1]);
  nor (_32401_, _11261_, _13388_);
  or (_32402_, _32401_, _32400_);
  or (_32403_, _32402_, _09061_);
  nand (_32404_, _07971_, _07038_);
  or (_32405_, _07971_, \oc8051_golden_model_1.P1 [1]);
  and (_32406_, _32405_, _06218_);
  and (_32407_, _32406_, _32404_);
  nor (_32408_, _13388_, _07357_);
  or (_32409_, _32408_, _32400_);
  or (_32411_, _32409_, _07166_);
  and (_32412_, _14562_, _07971_);
  not (_32413_, _32412_);
  and (_32414_, _32413_, _32405_);
  or (_32415_, _32414_, _07151_);
  and (_32416_, _07971_, \oc8051_golden_model_1.ACC [1]);
  or (_32417_, _32416_, _32400_);
  and (_32418_, _32417_, _07141_);
  and (_32419_, _07142_, \oc8051_golden_model_1.P1 [1]);
  or (_32420_, _32419_, _06341_);
  or (_32422_, _32420_, _32418_);
  and (_32423_, _32422_, _06273_);
  and (_32424_, _32423_, _32415_);
  and (_32425_, _13396_, \oc8051_golden_model_1.P1 [1]);
  and (_32426_, _14557_, _08620_);
  or (_32427_, _32426_, _32425_);
  and (_32428_, _32427_, _06272_);
  or (_32429_, _32428_, _06461_);
  or (_32430_, _32429_, _32424_);
  and (_32431_, _32430_, _32411_);
  or (_32433_, _32431_, _06464_);
  or (_32434_, _32417_, _06465_);
  and (_32435_, _32434_, _06269_);
  and (_32436_, _32435_, _32433_);
  and (_32437_, _14560_, _08620_);
  or (_32438_, _32437_, _32425_);
  and (_32439_, _32438_, _06268_);
  or (_32440_, _32439_, _06261_);
  or (_32441_, _32440_, _32436_);
  and (_32442_, _32426_, _14556_);
  or (_32444_, _32425_, _06262_);
  or (_32445_, _32444_, _32442_);
  and (_32446_, _32445_, _06258_);
  and (_32447_, _32446_, _32441_);
  or (_32448_, _32425_, _14597_);
  and (_32449_, _32448_, _06257_);
  and (_32450_, _32449_, _32427_);
  or (_32451_, _32450_, _10080_);
  or (_32452_, _32451_, _32447_);
  or (_32453_, _32409_, _07215_);
  and (_32455_, _32453_, _32452_);
  or (_32456_, _32455_, _07460_);
  and (_32457_, _09451_, _07971_);
  or (_32458_, _32400_, _07208_);
  or (_32459_, _32458_, _32457_);
  and (_32460_, _32459_, _05982_);
  and (_32461_, _32460_, _32456_);
  and (_32462_, _14653_, _07971_);
  or (_32463_, _32462_, _32400_);
  and (_32464_, _32463_, _10094_);
  or (_32466_, _32464_, _32461_);
  and (_32467_, _32466_, _06219_);
  or (_32468_, _32467_, _32407_);
  and (_32469_, _32468_, _07237_);
  or (_32470_, _14668_, _13388_);
  and (_32471_, _32405_, _06369_);
  and (_32472_, _32471_, _32470_);
  or (_32473_, _32472_, _06536_);
  or (_32474_, _32473_, _32469_);
  and (_32475_, _11262_, _07971_);
  or (_32476_, _32475_, _32400_);
  or (_32477_, _32476_, _07240_);
  and (_32478_, _32477_, _07242_);
  and (_32479_, _32478_, _32474_);
  or (_32480_, _14666_, _13388_);
  and (_32481_, _32405_, _06375_);
  and (_32482_, _32481_, _32480_);
  or (_32483_, _32482_, _06545_);
  or (_32484_, _32483_, _32479_);
  and (_32485_, _32416_, _08341_);
  or (_32487_, _32400_, _07234_);
  or (_32488_, _32487_, _32485_);
  and (_32489_, _32488_, _09056_);
  and (_32490_, _32489_, _32484_);
  or (_32491_, _32404_, _08341_);
  and (_32492_, _32405_, _06366_);
  and (_32493_, _32492_, _32491_);
  or (_32494_, _32493_, _06528_);
  or (_32495_, _32494_, _32490_);
  and (_32496_, _32495_, _32403_);
  or (_32498_, _32496_, _06568_);
  or (_32499_, _32414_, _06926_);
  and (_32500_, _32499_, _05928_);
  and (_32501_, _32500_, _32498_);
  and (_32502_, _32438_, _05927_);
  or (_32503_, _32502_, _06278_);
  or (_32504_, _32503_, _32501_);
  or (_32505_, _32400_, _06279_);
  or (_32506_, _32505_, _32412_);
  and (_32507_, _32506_, _01347_);
  and (_32509_, _32507_, _32504_);
  nor (_32510_, \oc8051_golden_model_1.P1 [1], rst);
  nor (_32511_, _32510_, _01354_);
  or (_43289_, _32511_, _32509_);
  nor (_32512_, \oc8051_golden_model_1.P1 [2], rst);
  nor (_32513_, _32512_, _01354_);
  and (_32514_, _13388_, \oc8051_golden_model_1.P1 [2]);
  nor (_32515_, _13388_, _07776_);
  or (_32516_, _32515_, _32514_);
  or (_32517_, _32516_, _07215_);
  or (_32519_, _32516_, _07166_);
  and (_32520_, _14770_, _07971_);
  or (_32521_, _32520_, _32514_);
  or (_32522_, _32521_, _07151_);
  and (_32523_, _07971_, \oc8051_golden_model_1.ACC [2]);
  or (_32524_, _32523_, _32514_);
  and (_32525_, _32524_, _07141_);
  and (_32526_, _07142_, \oc8051_golden_model_1.P1 [2]);
  or (_32527_, _32526_, _06341_);
  or (_32528_, _32527_, _32525_);
  and (_32530_, _32528_, _06273_);
  and (_32531_, _32530_, _32522_);
  and (_32532_, _13396_, \oc8051_golden_model_1.P1 [2]);
  and (_32533_, _14774_, _08620_);
  or (_32534_, _32533_, _32532_);
  and (_32535_, _32534_, _06272_);
  or (_32536_, _32535_, _06461_);
  or (_32537_, _32536_, _32531_);
  and (_32538_, _32537_, _32519_);
  or (_32539_, _32538_, _06464_);
  or (_32541_, _32524_, _06465_);
  and (_32542_, _32541_, _06269_);
  and (_32543_, _32542_, _32539_);
  and (_32544_, _14756_, _08620_);
  or (_32545_, _32544_, _32532_);
  and (_32546_, _32545_, _06268_);
  or (_32547_, _32546_, _06261_);
  or (_32548_, _32547_, _32543_);
  and (_32549_, _32533_, _14789_);
  or (_32550_, _32532_, _06262_);
  or (_32552_, _32550_, _32549_);
  and (_32553_, _32552_, _06258_);
  and (_32554_, _32553_, _32548_);
  and (_32555_, _14804_, _08620_);
  or (_32556_, _32555_, _32532_);
  and (_32557_, _32556_, _06257_);
  or (_32558_, _32557_, _10080_);
  or (_32559_, _32558_, _32554_);
  and (_32560_, _32559_, _32517_);
  or (_32561_, _32560_, _07460_);
  and (_32563_, _09450_, _07971_);
  or (_32564_, _32514_, _07208_);
  or (_32565_, _32564_, _32563_);
  and (_32566_, _32565_, _05982_);
  and (_32567_, _32566_, _32561_);
  and (_32568_, _14859_, _07971_);
  or (_32569_, _32568_, _32514_);
  and (_32570_, _32569_, _10094_);
  or (_32571_, _32570_, _06218_);
  or (_32572_, _32571_, _32567_);
  and (_32574_, _07971_, _08973_);
  or (_32575_, _32574_, _32514_);
  or (_32576_, _32575_, _06219_);
  and (_32577_, _32576_, _32572_);
  or (_32578_, _32577_, _06369_);
  and (_32579_, _14751_, _07971_);
  or (_32580_, _32579_, _32514_);
  or (_32581_, _32580_, _07237_);
  and (_32582_, _32581_, _07240_);
  and (_32583_, _32582_, _32578_);
  and (_32585_, _11259_, _07971_);
  or (_32586_, _32585_, _32514_);
  and (_32587_, _32586_, _06536_);
  or (_32588_, _32587_, _32583_);
  and (_32589_, _32588_, _07242_);
  or (_32590_, _32514_, _08440_);
  and (_32591_, _32575_, _06375_);
  and (_32592_, _32591_, _32590_);
  or (_32593_, _32592_, _32589_);
  and (_32594_, _32593_, _07234_);
  and (_32596_, _32524_, _06545_);
  and (_32597_, _32596_, _32590_);
  or (_32598_, _32597_, _06366_);
  or (_32599_, _32598_, _32594_);
  and (_32600_, _14748_, _07971_);
  or (_32601_, _32514_, _09056_);
  or (_32602_, _32601_, _32600_);
  and (_32603_, _32602_, _09061_);
  and (_32604_, _32603_, _32599_);
  nor (_32605_, _11258_, _13388_);
  or (_32607_, _32605_, _32514_);
  and (_32608_, _32607_, _06528_);
  or (_32609_, _32608_, _06568_);
  or (_32610_, _32609_, _32604_);
  or (_32611_, _32521_, _06926_);
  and (_32612_, _32611_, _05928_);
  and (_32613_, _32612_, _32610_);
  and (_32614_, _32545_, _05927_);
  or (_32615_, _32614_, _06278_);
  or (_32616_, _32615_, _32613_);
  and (_32618_, _14926_, _07971_);
  or (_32619_, _32514_, _06279_);
  or (_32620_, _32619_, _32618_);
  and (_32621_, _32620_, _01347_);
  and (_32622_, _32621_, _32616_);
  or (_43290_, _32622_, _32513_);
  and (_32623_, _13388_, \oc8051_golden_model_1.P1 [3]);
  nor (_32624_, _13388_, _07594_);
  or (_32625_, _32624_, _32623_);
  or (_32626_, _32625_, _07215_);
  and (_32628_, _14953_, _07971_);
  or (_32629_, _32628_, _32623_);
  or (_32630_, _32629_, _07151_);
  and (_32631_, _07971_, \oc8051_golden_model_1.ACC [3]);
  or (_32632_, _32631_, _32623_);
  and (_32633_, _32632_, _07141_);
  and (_32634_, _07142_, \oc8051_golden_model_1.P1 [3]);
  or (_32635_, _32634_, _06341_);
  or (_32636_, _32635_, _32633_);
  and (_32637_, _32636_, _06273_);
  and (_32639_, _32637_, _32630_);
  and (_32640_, _13396_, \oc8051_golden_model_1.P1 [3]);
  and (_32641_, _14950_, _08620_);
  or (_32642_, _32641_, _32640_);
  and (_32643_, _32642_, _06272_);
  or (_32644_, _32643_, _06461_);
  or (_32645_, _32644_, _32639_);
  or (_32646_, _32625_, _07166_);
  and (_32647_, _32646_, _32645_);
  or (_32648_, _32647_, _06464_);
  or (_32650_, _32632_, _06465_);
  and (_32651_, _32650_, _06269_);
  and (_32652_, _32651_, _32648_);
  and (_32653_, _14948_, _08620_);
  or (_32654_, _32653_, _32640_);
  and (_32655_, _32654_, _06268_);
  or (_32656_, _32655_, _06261_);
  or (_32657_, _32656_, _32652_);
  or (_32658_, _32640_, _14979_);
  and (_32659_, _32658_, _32642_);
  or (_32661_, _32659_, _06262_);
  and (_32662_, _32661_, _06258_);
  and (_32663_, _32662_, _32657_);
  or (_32664_, _32640_, _14992_);
  and (_32665_, _32664_, _06257_);
  and (_32666_, _32665_, _32642_);
  or (_32667_, _32666_, _10080_);
  or (_32668_, _32667_, _32663_);
  and (_32669_, _32668_, _32626_);
  or (_32670_, _32669_, _07460_);
  and (_32672_, _09449_, _07971_);
  or (_32673_, _32623_, _07208_);
  or (_32674_, _32673_, _32672_);
  and (_32675_, _32674_, _05982_);
  and (_32676_, _32675_, _32670_);
  and (_32677_, _15048_, _07971_);
  or (_32678_, _32677_, _32623_);
  and (_32679_, _32678_, _10094_);
  or (_32680_, _32679_, _06218_);
  or (_32681_, _32680_, _32676_);
  and (_32683_, _07971_, _08930_);
  or (_32684_, _32683_, _32623_);
  or (_32685_, _32684_, _06219_);
  and (_32686_, _32685_, _32681_);
  or (_32687_, _32686_, _06369_);
  and (_32688_, _14943_, _07971_);
  or (_32689_, _32688_, _32623_);
  or (_32690_, _32689_, _07237_);
  and (_32691_, _32690_, _07240_);
  and (_32692_, _32691_, _32687_);
  and (_32694_, _12577_, _07971_);
  or (_32695_, _32694_, _32623_);
  and (_32696_, _32695_, _06536_);
  or (_32697_, _32696_, _32692_);
  and (_32698_, _32697_, _07242_);
  or (_32699_, _32623_, _08292_);
  and (_32700_, _32684_, _06375_);
  and (_32701_, _32700_, _32699_);
  or (_32702_, _32701_, _32698_);
  and (_32703_, _32702_, _07234_);
  and (_32705_, _32632_, _06545_);
  and (_32706_, _32705_, _32699_);
  or (_32707_, _32706_, _06366_);
  or (_32708_, _32707_, _32703_);
  and (_32709_, _14940_, _07971_);
  or (_32710_, _32623_, _09056_);
  or (_32711_, _32710_, _32709_);
  and (_32712_, _32711_, _09061_);
  and (_32713_, _32712_, _32708_);
  nor (_32714_, _11256_, _13388_);
  or (_32716_, _32714_, _32623_);
  and (_32717_, _32716_, _06528_);
  or (_32718_, _32717_, _06568_);
  or (_32719_, _32718_, _32713_);
  or (_32720_, _32629_, _06926_);
  and (_32721_, _32720_, _05928_);
  and (_32722_, _32721_, _32719_);
  and (_32723_, _32654_, _05927_);
  or (_32724_, _32723_, _06278_);
  or (_32725_, _32724_, _32722_);
  and (_32727_, _15128_, _07971_);
  or (_32728_, _32623_, _06279_);
  or (_32729_, _32728_, _32727_);
  and (_32730_, _32729_, _01347_);
  and (_32731_, _32730_, _32725_);
  nor (_32732_, \oc8051_golden_model_1.P1 [3], rst);
  nor (_32733_, _32732_, _01354_);
  or (_43291_, _32733_, _32731_);
  nor (_32734_, \oc8051_golden_model_1.P1 [4], rst);
  nor (_32735_, _32734_, _01354_);
  and (_32737_, _13388_, \oc8051_golden_model_1.P1 [4]);
  nor (_32738_, _08541_, _13388_);
  or (_32739_, _32738_, _32737_);
  or (_32740_, _32739_, _07215_);
  and (_32741_, _13396_, \oc8051_golden_model_1.P1 [4]);
  and (_32742_, _15176_, _08620_);
  or (_32743_, _32742_, _32741_);
  and (_32744_, _32743_, _06268_);
  and (_32745_, _15162_, _07971_);
  or (_32746_, _32745_, _32737_);
  or (_32748_, _32746_, _07151_);
  and (_32749_, _07971_, \oc8051_golden_model_1.ACC [4]);
  or (_32750_, _32749_, _32737_);
  and (_32751_, _32750_, _07141_);
  and (_32752_, _07142_, \oc8051_golden_model_1.P1 [4]);
  or (_32753_, _32752_, _06341_);
  or (_32754_, _32753_, _32751_);
  and (_32755_, _32754_, _06273_);
  and (_32756_, _32755_, _32748_);
  and (_32757_, _15166_, _08620_);
  or (_32759_, _32757_, _32741_);
  and (_32760_, _32759_, _06272_);
  or (_32761_, _32760_, _06461_);
  or (_32762_, _32761_, _32756_);
  or (_32763_, _32739_, _07166_);
  and (_32764_, _32763_, _32762_);
  or (_32765_, _32764_, _06464_);
  or (_32766_, _32750_, _06465_);
  and (_32767_, _32766_, _06269_);
  and (_32768_, _32767_, _32765_);
  or (_32770_, _32768_, _32744_);
  and (_32771_, _32770_, _06262_);
  and (_32772_, _15184_, _08620_);
  or (_32773_, _32772_, _32741_);
  and (_32774_, _32773_, _06261_);
  or (_32775_, _32774_, _32771_);
  and (_32776_, _32775_, _06258_);
  and (_32777_, _15200_, _08620_);
  or (_32778_, _32777_, _32741_);
  and (_32779_, _32778_, _06257_);
  or (_32781_, _32779_, _10080_);
  or (_32782_, _32781_, _32776_);
  and (_32783_, _32782_, _32740_);
  or (_32784_, _32783_, _07460_);
  and (_32785_, _09448_, _07971_);
  or (_32786_, _32737_, _07208_);
  or (_32787_, _32786_, _32785_);
  and (_32788_, _32787_, _05982_);
  and (_32789_, _32788_, _32784_);
  and (_32790_, _15254_, _07971_);
  or (_32792_, _32790_, _32737_);
  and (_32793_, _32792_, _10094_);
  or (_32794_, _32793_, _06218_);
  or (_32795_, _32794_, _32789_);
  and (_32796_, _08959_, _07971_);
  or (_32797_, _32796_, _32737_);
  or (_32798_, _32797_, _06219_);
  and (_32799_, _32798_, _32795_);
  or (_32800_, _32799_, _06369_);
  and (_32801_, _15269_, _07971_);
  or (_32803_, _32801_, _32737_);
  or (_32804_, _32803_, _07237_);
  and (_32805_, _32804_, _07240_);
  and (_32806_, _32805_, _32800_);
  and (_32807_, _11254_, _07971_);
  or (_32808_, _32807_, _32737_);
  and (_32809_, _32808_, _06536_);
  or (_32810_, _32809_, _32806_);
  and (_32811_, _32810_, _07242_);
  or (_32812_, _32737_, _08544_);
  and (_32814_, _32797_, _06375_);
  and (_32815_, _32814_, _32812_);
  or (_32816_, _32815_, _32811_);
  and (_32817_, _32816_, _07234_);
  and (_32818_, _32750_, _06545_);
  and (_32819_, _32818_, _32812_);
  or (_32820_, _32819_, _06366_);
  or (_32821_, _32820_, _32817_);
  and (_32822_, _15266_, _07971_);
  or (_32823_, _32737_, _09056_);
  or (_32825_, _32823_, _32822_);
  and (_32826_, _32825_, _09061_);
  and (_32827_, _32826_, _32821_);
  nor (_32828_, _11253_, _13388_);
  or (_32829_, _32828_, _32737_);
  and (_32830_, _32829_, _06528_);
  or (_32831_, _32830_, _06568_);
  or (_32832_, _32831_, _32827_);
  or (_32833_, _32746_, _06926_);
  and (_32834_, _32833_, _05928_);
  and (_32836_, _32834_, _32832_);
  and (_32837_, _32743_, _05927_);
  or (_32838_, _32837_, _06278_);
  or (_32839_, _32838_, _32836_);
  and (_32840_, _15329_, _07971_);
  or (_32841_, _32737_, _06279_);
  or (_32842_, _32841_, _32840_);
  and (_32843_, _32842_, _01347_);
  and (_32844_, _32843_, _32839_);
  or (_43292_, _32844_, _32735_);
  and (_32846_, _13388_, \oc8051_golden_model_1.P1 [5]);
  and (_32847_, _15358_, _07971_);
  or (_32848_, _32847_, _32846_);
  or (_32849_, _32848_, _07151_);
  and (_32850_, _07971_, \oc8051_golden_model_1.ACC [5]);
  or (_32851_, _32850_, _32846_);
  and (_32852_, _32851_, _07141_);
  and (_32853_, _07142_, \oc8051_golden_model_1.P1 [5]);
  or (_32854_, _32853_, _06341_);
  or (_32855_, _32854_, _32852_);
  and (_32857_, _32855_, _06273_);
  and (_32858_, _32857_, _32849_);
  and (_32859_, _13396_, \oc8051_golden_model_1.P1 [5]);
  and (_32860_, _15372_, _08620_);
  or (_32861_, _32860_, _32859_);
  and (_32862_, _32861_, _06272_);
  or (_32863_, _32862_, _06461_);
  or (_32864_, _32863_, _32858_);
  nor (_32865_, _08244_, _13388_);
  or (_32866_, _32865_, _32846_);
  or (_32868_, _32866_, _07166_);
  and (_32869_, _32868_, _32864_);
  or (_32870_, _32869_, _06464_);
  or (_32871_, _32851_, _06465_);
  and (_32872_, _32871_, _06269_);
  and (_32873_, _32872_, _32870_);
  and (_32874_, _15355_, _08620_);
  or (_32875_, _32874_, _32859_);
  and (_32876_, _32875_, _06268_);
  or (_32877_, _32876_, _06261_);
  or (_32879_, _32877_, _32873_);
  or (_32880_, _32859_, _15387_);
  and (_32881_, _32880_, _32861_);
  or (_32882_, _32881_, _06262_);
  and (_32883_, _32882_, _06258_);
  and (_32884_, _32883_, _32879_);
  or (_32885_, _32859_, _15403_);
  and (_32886_, _32885_, _06257_);
  and (_32887_, _32886_, _32861_);
  or (_32888_, _32887_, _10080_);
  or (_32890_, _32888_, _32884_);
  or (_32891_, _32866_, _07215_);
  and (_32892_, _32891_, _32890_);
  or (_32893_, _32892_, _07460_);
  and (_32894_, _09447_, _07971_);
  or (_32895_, _32846_, _07208_);
  or (_32896_, _32895_, _32894_);
  and (_32897_, _32896_, _05982_);
  and (_32898_, _32897_, _32893_);
  and (_32899_, _15459_, _07971_);
  or (_32901_, _32899_, _32846_);
  and (_32902_, _32901_, _10094_);
  or (_32903_, _32902_, _06218_);
  or (_32904_, _32903_, _32898_);
  and (_32905_, _08946_, _07971_);
  or (_32906_, _32905_, _32846_);
  or (_32907_, _32906_, _06219_);
  and (_32908_, _32907_, _32904_);
  or (_32909_, _32908_, _06369_);
  and (_32910_, _15353_, _07971_);
  or (_32912_, _32910_, _32846_);
  or (_32913_, _32912_, _07237_);
  and (_32914_, _32913_, _07240_);
  and (_32915_, _32914_, _32909_);
  and (_32916_, _11250_, _07971_);
  or (_32917_, _32916_, _32846_);
  and (_32918_, _32917_, _06536_);
  or (_32919_, _32918_, _32915_);
  and (_32920_, _32919_, _07242_);
  or (_32921_, _32846_, _08247_);
  and (_32923_, _32906_, _06375_);
  and (_32924_, _32923_, _32921_);
  or (_32925_, _32924_, _32920_);
  and (_32926_, _32925_, _07234_);
  and (_32927_, _32851_, _06545_);
  and (_32928_, _32927_, _32921_);
  or (_32929_, _32928_, _06366_);
  or (_32930_, _32929_, _32926_);
  and (_32931_, _15350_, _07971_);
  or (_32932_, _32846_, _09056_);
  or (_32934_, _32932_, _32931_);
  and (_32935_, _32934_, _09061_);
  and (_32936_, _32935_, _32930_);
  nor (_32937_, _11249_, _13388_);
  or (_32938_, _32937_, _32846_);
  and (_32939_, _32938_, _06528_);
  or (_32940_, _32939_, _06568_);
  or (_32941_, _32940_, _32936_);
  or (_32942_, _32848_, _06926_);
  and (_32943_, _32942_, _05928_);
  and (_32945_, _32943_, _32941_);
  and (_32946_, _32875_, _05927_);
  or (_32947_, _32946_, _06278_);
  or (_32948_, _32947_, _32945_);
  and (_32949_, _15532_, _07971_);
  or (_32950_, _32846_, _06279_);
  or (_32951_, _32950_, _32949_);
  and (_32952_, _32951_, _01347_);
  and (_32953_, _32952_, _32948_);
  nor (_32954_, \oc8051_golden_model_1.P1 [5], rst);
  nor (_32956_, _32954_, _01354_);
  or (_43293_, _32956_, _32953_);
  and (_32957_, _13388_, \oc8051_golden_model_1.P1 [6]);
  and (_32958_, _15554_, _07971_);
  or (_32959_, _32958_, _32957_);
  or (_32960_, _32959_, _07151_);
  and (_32961_, _07971_, \oc8051_golden_model_1.ACC [6]);
  or (_32962_, _32961_, _32957_);
  and (_32963_, _32962_, _07141_);
  and (_32964_, _07142_, \oc8051_golden_model_1.P1 [6]);
  or (_32966_, _32964_, _06341_);
  or (_32967_, _32966_, _32963_);
  and (_32968_, _32967_, _06273_);
  and (_32969_, _32968_, _32960_);
  and (_32970_, _13396_, \oc8051_golden_model_1.P1 [6]);
  and (_32971_, _15570_, _08620_);
  or (_32972_, _32971_, _32970_);
  and (_32973_, _32972_, _06272_);
  or (_32974_, _32973_, _06461_);
  or (_32975_, _32974_, _32969_);
  nor (_32977_, _08142_, _13388_);
  or (_32978_, _32977_, _32957_);
  or (_32979_, _32978_, _07166_);
  and (_32980_, _32979_, _32975_);
  or (_32981_, _32980_, _06464_);
  or (_32982_, _32962_, _06465_);
  and (_32983_, _32982_, _06269_);
  and (_32984_, _32983_, _32981_);
  and (_32985_, _15551_, _08620_);
  or (_32986_, _32985_, _32970_);
  and (_32988_, _32986_, _06268_);
  or (_32989_, _32988_, _06261_);
  or (_32990_, _32989_, _32984_);
  or (_32991_, _32970_, _15585_);
  and (_32992_, _32991_, _32972_);
  or (_32993_, _32992_, _06262_);
  and (_32994_, _32993_, _06258_);
  and (_32995_, _32994_, _32990_);
  and (_32996_, _15602_, _08620_);
  or (_32997_, _32996_, _32970_);
  and (_32999_, _32997_, _06257_);
  or (_33000_, _32999_, _10080_);
  or (_33001_, _33000_, _32995_);
  or (_33002_, _32978_, _07215_);
  and (_33003_, _33002_, _33001_);
  or (_33004_, _33003_, _07460_);
  and (_33005_, _09446_, _07971_);
  or (_33006_, _32957_, _07208_);
  or (_33007_, _33006_, _33005_);
  and (_33008_, _33007_, _05982_);
  and (_33010_, _33008_, _33004_);
  and (_33011_, _15657_, _07971_);
  or (_33012_, _33011_, _32957_);
  and (_33013_, _33012_, _10094_);
  or (_33014_, _33013_, _06218_);
  or (_33015_, _33014_, _33010_);
  and (_33016_, _15664_, _07971_);
  or (_33017_, _33016_, _32957_);
  or (_33018_, _33017_, _06219_);
  and (_33019_, _33018_, _33015_);
  or (_33021_, _33019_, _06369_);
  and (_33022_, _15549_, _07971_);
  or (_33023_, _33022_, _32957_);
  or (_33024_, _33023_, _07237_);
  and (_33025_, _33024_, _07240_);
  and (_33026_, _33025_, _33021_);
  and (_33027_, _11247_, _07971_);
  or (_33028_, _33027_, _32957_);
  and (_33029_, _33028_, _06536_);
  or (_33030_, _33029_, _33026_);
  and (_33032_, _33030_, _07242_);
  or (_33033_, _32957_, _08145_);
  and (_33034_, _33017_, _06375_);
  and (_33035_, _33034_, _33033_);
  or (_33036_, _33035_, _33032_);
  and (_33037_, _33036_, _07234_);
  and (_33038_, _32962_, _06545_);
  and (_33039_, _33038_, _33033_);
  or (_33040_, _33039_, _06366_);
  or (_33041_, _33040_, _33037_);
  and (_33043_, _15546_, _07971_);
  or (_33044_, _32957_, _09056_);
  or (_33045_, _33044_, _33043_);
  and (_33046_, _33045_, _09061_);
  and (_33047_, _33046_, _33041_);
  nor (_33048_, _11246_, _13388_);
  or (_33049_, _33048_, _32957_);
  and (_33050_, _33049_, _06528_);
  or (_33051_, _33050_, _06568_);
  or (_33052_, _33051_, _33047_);
  or (_33054_, _32959_, _06926_);
  and (_33055_, _33054_, _05928_);
  and (_33056_, _33055_, _33052_);
  and (_33057_, _32986_, _05927_);
  or (_33058_, _33057_, _06278_);
  or (_33059_, _33058_, _33056_);
  and (_33060_, _15734_, _07971_);
  or (_33061_, _32957_, _06279_);
  or (_33062_, _33061_, _33060_);
  and (_33063_, _33062_, _01347_);
  and (_33065_, _33063_, _33059_);
  nor (_33066_, \oc8051_golden_model_1.P1 [6], rst);
  nor (_33067_, _33066_, _01354_);
  or (_43294_, _33067_, _33065_);
  and (_33068_, _01351_, \oc8051_golden_model_1.IP [0]);
  and (_33069_, _07946_, \oc8051_golden_model_1.ACC [0]);
  and (_33070_, _33069_, _08390_);
  and (_33071_, _13490_, \oc8051_golden_model_1.IP [0]);
  or (_33072_, _33071_, _07234_);
  or (_33073_, _33072_, _33070_);
  and (_33075_, _07946_, _07133_);
  or (_33076_, _33075_, _33071_);
  or (_33077_, _33076_, _07215_);
  nor (_33078_, _08390_, _13490_);
  or (_33079_, _33078_, _33071_);
  and (_33080_, _33079_, _06341_);
  and (_33081_, _07142_, \oc8051_golden_model_1.IP [0]);
  or (_33082_, _33069_, _33071_);
  and (_33083_, _33082_, _07141_);
  or (_33084_, _33083_, _33081_);
  and (_33086_, _33084_, _07151_);
  or (_33087_, _33086_, _06272_);
  or (_33088_, _33087_, _33080_);
  and (_33089_, _14382_, _08632_);
  and (_33090_, _13498_, \oc8051_golden_model_1.IP [0]);
  or (_33091_, _33090_, _06273_);
  or (_33092_, _33091_, _33089_);
  and (_33093_, _33092_, _07166_);
  and (_33094_, _33093_, _33088_);
  and (_33095_, _33076_, _06461_);
  or (_33097_, _33095_, _06464_);
  or (_33098_, _33097_, _33094_);
  or (_33099_, _33082_, _06465_);
  and (_33100_, _33099_, _06269_);
  and (_33101_, _33100_, _33098_);
  and (_33102_, _33071_, _06268_);
  or (_33103_, _33102_, _06261_);
  or (_33104_, _33103_, _33101_);
  or (_33105_, _33079_, _06262_);
  and (_33106_, _33105_, _06258_);
  and (_33108_, _33106_, _33104_);
  and (_33109_, _14413_, _08632_);
  or (_33110_, _33109_, _33090_);
  and (_33111_, _33110_, _06257_);
  or (_33112_, _33111_, _10080_);
  or (_33113_, _33112_, _33108_);
  and (_33114_, _33113_, _33077_);
  or (_33115_, _33114_, _07460_);
  and (_33116_, _09392_, _07946_);
  or (_33117_, _33071_, _07208_);
  or (_33119_, _33117_, _33116_);
  and (_33120_, _33119_, _33115_);
  or (_33121_, _33120_, _10094_);
  and (_33122_, _14467_, _07946_);
  or (_33123_, _33071_, _05982_);
  or (_33124_, _33123_, _33122_);
  and (_33125_, _33124_, _06219_);
  and (_33126_, _33125_, _33121_);
  and (_33127_, _07946_, _08954_);
  or (_33128_, _33127_, _33071_);
  and (_33130_, _33128_, _06218_);
  or (_33131_, _33130_, _06369_);
  or (_33132_, _33131_, _33126_);
  and (_33133_, _14366_, _07946_);
  or (_33134_, _33133_, _33071_);
  or (_33135_, _33134_, _07237_);
  and (_33136_, _33135_, _07240_);
  and (_33137_, _33136_, _33132_);
  nor (_33138_, _12580_, _13490_);
  or (_33139_, _33138_, _33071_);
  nor (_33141_, _33070_, _07240_);
  and (_33142_, _33141_, _33139_);
  or (_33143_, _33142_, _33137_);
  and (_33144_, _33143_, _07242_);
  nand (_33145_, _33128_, _06375_);
  nor (_33146_, _33145_, _33078_);
  or (_33147_, _33146_, _06545_);
  or (_33148_, _33147_, _33144_);
  and (_33149_, _33148_, _33073_);
  or (_33150_, _33149_, _06366_);
  and (_33152_, _14363_, _07946_);
  or (_33153_, _33071_, _09056_);
  or (_33154_, _33153_, _33152_);
  and (_33155_, _33154_, _09061_);
  and (_33156_, _33155_, _33150_);
  and (_33157_, _33139_, _06528_);
  or (_33158_, _33157_, _06568_);
  or (_33159_, _33158_, _33156_);
  or (_33160_, _33079_, _06926_);
  and (_33161_, _33160_, _33159_);
  or (_33163_, _33161_, _05927_);
  or (_33164_, _33071_, _05928_);
  and (_33165_, _33164_, _33163_);
  or (_33166_, _33165_, _06278_);
  or (_33167_, _33079_, _06279_);
  and (_33168_, _33167_, _01347_);
  and (_33169_, _33168_, _33166_);
  or (_33170_, _33169_, _33068_);
  and (_43296_, _33170_, _42618_);
  not (_33171_, \oc8051_golden_model_1.IP [1]);
  nor (_33173_, _01347_, _33171_);
  nor (_33174_, _07946_, _33171_);
  nor (_33175_, _11261_, _13490_);
  or (_33176_, _33175_, _33174_);
  or (_33177_, _33176_, _09061_);
  nand (_33178_, _07946_, _07038_);
  or (_33179_, _07946_, \oc8051_golden_model_1.IP [1]);
  and (_33180_, _33179_, _06218_);
  and (_33181_, _33180_, _33178_);
  nor (_33182_, _13490_, _07357_);
  or (_33184_, _33182_, _33174_);
  or (_33185_, _33184_, _07166_);
  and (_33186_, _14562_, _07946_);
  not (_33187_, _33186_);
  and (_33188_, _33187_, _33179_);
  or (_33189_, _33188_, _07151_);
  and (_33190_, _07946_, \oc8051_golden_model_1.ACC [1]);
  or (_33191_, _33190_, _33174_);
  and (_33192_, _33191_, _07141_);
  nor (_33193_, _07141_, _33171_);
  or (_33195_, _33193_, _06341_);
  or (_33196_, _33195_, _33192_);
  and (_33197_, _33196_, _06273_);
  and (_33198_, _33197_, _33189_);
  nor (_33199_, _08632_, _33171_);
  and (_33200_, _14557_, _08632_);
  or (_33201_, _33200_, _33199_);
  and (_33202_, _33201_, _06272_);
  or (_33203_, _33202_, _06461_);
  or (_33204_, _33203_, _33198_);
  and (_33206_, _33204_, _33185_);
  or (_33207_, _33206_, _06464_);
  or (_33208_, _33191_, _06465_);
  and (_33209_, _33208_, _06269_);
  and (_33210_, _33209_, _33207_);
  and (_33211_, _14560_, _08632_);
  or (_33212_, _33211_, _33199_);
  and (_33213_, _33212_, _06268_);
  or (_33214_, _33213_, _06261_);
  or (_33215_, _33214_, _33210_);
  and (_33216_, _33200_, _14556_);
  or (_33217_, _33199_, _06262_);
  or (_33218_, _33217_, _33216_);
  and (_33219_, _33218_, _06258_);
  and (_33220_, _33219_, _33215_);
  or (_33221_, _33199_, _14597_);
  and (_33222_, _33221_, _06257_);
  and (_33223_, _33222_, _33201_);
  or (_33224_, _33223_, _10080_);
  or (_33225_, _33224_, _33220_);
  or (_33227_, _33184_, _07215_);
  and (_33228_, _33227_, _33225_);
  or (_33229_, _33228_, _07460_);
  and (_33230_, _09451_, _07946_);
  or (_33231_, _33174_, _07208_);
  or (_33232_, _33231_, _33230_);
  and (_33233_, _33232_, _05982_);
  and (_33234_, _33233_, _33229_);
  and (_33235_, _14653_, _07946_);
  or (_33236_, _33235_, _33174_);
  and (_33238_, _33236_, _10094_);
  or (_33239_, _33238_, _33234_);
  and (_33240_, _33239_, _06219_);
  or (_33241_, _33240_, _33181_);
  and (_33242_, _33241_, _07237_);
  or (_33243_, _14668_, _13490_);
  and (_33244_, _33179_, _06369_);
  and (_33245_, _33244_, _33243_);
  or (_33246_, _33245_, _06536_);
  or (_33247_, _33246_, _33242_);
  nand (_33249_, _11260_, _07946_);
  and (_33250_, _33249_, _33176_);
  or (_33251_, _33250_, _07240_);
  and (_33252_, _33251_, _07242_);
  and (_33253_, _33252_, _33247_);
  or (_33254_, _14666_, _13490_);
  and (_33255_, _33179_, _06375_);
  and (_33256_, _33255_, _33254_);
  or (_33257_, _33256_, _06545_);
  or (_33258_, _33257_, _33253_);
  nor (_33260_, _33174_, _07234_);
  nand (_33261_, _33260_, _33249_);
  and (_33262_, _33261_, _09056_);
  and (_33263_, _33262_, _33258_);
  or (_33264_, _33178_, _08341_);
  and (_33265_, _33179_, _06366_);
  and (_33266_, _33265_, _33264_);
  or (_33267_, _33266_, _06528_);
  or (_33268_, _33267_, _33263_);
  and (_33269_, _33268_, _33177_);
  or (_33271_, _33269_, _06568_);
  or (_33272_, _33188_, _06926_);
  and (_33273_, _33272_, _05928_);
  and (_33274_, _33273_, _33271_);
  and (_33275_, _33212_, _05927_);
  or (_33276_, _33275_, _06278_);
  or (_33277_, _33276_, _33274_);
  or (_33278_, _33174_, _06279_);
  or (_33279_, _33278_, _33186_);
  and (_33280_, _33279_, _01347_);
  and (_33282_, _33280_, _33277_);
  or (_33283_, _33282_, _33173_);
  and (_43297_, _33283_, _42618_);
  and (_33284_, _01351_, \oc8051_golden_model_1.IP [2]);
  and (_33285_, _13490_, \oc8051_golden_model_1.IP [2]);
  nor (_33286_, _13490_, _07776_);
  or (_33287_, _33286_, _33285_);
  or (_33288_, _33287_, _07215_);
  or (_33289_, _33287_, _07166_);
  and (_33290_, _14770_, _07946_);
  or (_33292_, _33290_, _33285_);
  or (_33293_, _33292_, _07151_);
  and (_33294_, _07946_, \oc8051_golden_model_1.ACC [2]);
  or (_33295_, _33294_, _33285_);
  and (_33296_, _33295_, _07141_);
  and (_33297_, _07142_, \oc8051_golden_model_1.IP [2]);
  or (_33298_, _33297_, _06341_);
  or (_33299_, _33298_, _33296_);
  and (_33300_, _33299_, _06273_);
  and (_33301_, _33300_, _33293_);
  and (_33303_, _13498_, \oc8051_golden_model_1.IP [2]);
  and (_33304_, _14774_, _08632_);
  or (_33305_, _33304_, _33303_);
  and (_33306_, _33305_, _06272_);
  or (_33307_, _33306_, _06461_);
  or (_33308_, _33307_, _33301_);
  and (_33309_, _33308_, _33289_);
  or (_33310_, _33309_, _06464_);
  or (_33311_, _33295_, _06465_);
  and (_33312_, _33311_, _06269_);
  and (_33314_, _33312_, _33310_);
  and (_33315_, _14756_, _08632_);
  or (_33316_, _33315_, _33303_);
  and (_33317_, _33316_, _06268_);
  or (_33318_, _33317_, _06261_);
  or (_33319_, _33318_, _33314_);
  and (_33320_, _33304_, _14789_);
  or (_33321_, _33303_, _06262_);
  or (_33322_, _33321_, _33320_);
  and (_33323_, _33322_, _06258_);
  and (_33325_, _33323_, _33319_);
  and (_33326_, _14804_, _08632_);
  or (_33327_, _33326_, _33303_);
  and (_33328_, _33327_, _06257_);
  or (_33329_, _33328_, _10080_);
  or (_33330_, _33329_, _33325_);
  and (_33331_, _33330_, _33288_);
  or (_33332_, _33331_, _07460_);
  and (_33333_, _09450_, _07946_);
  or (_33334_, _33285_, _07208_);
  or (_33336_, _33334_, _33333_);
  and (_33337_, _33336_, _05982_);
  and (_33338_, _33337_, _33332_);
  and (_33339_, _14859_, _07946_);
  or (_33340_, _33339_, _33285_);
  and (_33341_, _33340_, _10094_);
  or (_33342_, _33341_, _06218_);
  or (_33343_, _33342_, _33338_);
  and (_33344_, _07946_, _08973_);
  or (_33345_, _33344_, _33285_);
  or (_33347_, _33345_, _06219_);
  and (_33348_, _33347_, _33343_);
  or (_33349_, _33348_, _06369_);
  and (_33350_, _14751_, _07946_);
  or (_33351_, _33350_, _33285_);
  or (_33352_, _33351_, _07237_);
  and (_33353_, _33352_, _07240_);
  and (_33354_, _33353_, _33349_);
  and (_33355_, _11259_, _07946_);
  or (_33356_, _33355_, _33285_);
  and (_33358_, _33356_, _06536_);
  or (_33359_, _33358_, _33354_);
  and (_33360_, _33359_, _07242_);
  or (_33361_, _33285_, _08440_);
  and (_33362_, _33345_, _06375_);
  and (_33363_, _33362_, _33361_);
  or (_33364_, _33363_, _33360_);
  and (_33365_, _33364_, _07234_);
  and (_33366_, _33295_, _06545_);
  and (_33367_, _33366_, _33361_);
  or (_33369_, _33367_, _06366_);
  or (_33370_, _33369_, _33365_);
  and (_33371_, _14748_, _07946_);
  or (_33372_, _33285_, _09056_);
  or (_33373_, _33372_, _33371_);
  and (_33374_, _33373_, _09061_);
  and (_33375_, _33374_, _33370_);
  nor (_33376_, _11258_, _13490_);
  or (_33377_, _33376_, _33285_);
  and (_33378_, _33377_, _06528_);
  or (_33380_, _33378_, _06568_);
  or (_33381_, _33380_, _33375_);
  or (_33382_, _33292_, _06926_);
  and (_33383_, _33382_, _05928_);
  and (_33384_, _33383_, _33381_);
  and (_33385_, _33316_, _05927_);
  or (_33386_, _33385_, _06278_);
  or (_33387_, _33386_, _33384_);
  and (_33388_, _14926_, _07946_);
  or (_33389_, _33285_, _06279_);
  or (_33391_, _33389_, _33388_);
  and (_33392_, _33391_, _01347_);
  and (_33393_, _33392_, _33387_);
  or (_33394_, _33393_, _33284_);
  and (_43298_, _33394_, _42618_);
  and (_33395_, _01351_, \oc8051_golden_model_1.IP [3]);
  and (_33396_, _13490_, \oc8051_golden_model_1.IP [3]);
  nor (_33397_, _13490_, _07594_);
  or (_33398_, _33397_, _33396_);
  or (_33399_, _33398_, _07215_);
  and (_33401_, _14953_, _07946_);
  or (_33402_, _33401_, _33396_);
  or (_33403_, _33402_, _07151_);
  and (_33404_, _07946_, \oc8051_golden_model_1.ACC [3]);
  or (_33405_, _33404_, _33396_);
  and (_33406_, _33405_, _07141_);
  and (_33407_, _07142_, \oc8051_golden_model_1.IP [3]);
  or (_33408_, _33407_, _06341_);
  or (_33409_, _33408_, _33406_);
  and (_33410_, _33409_, _06273_);
  and (_33412_, _33410_, _33403_);
  and (_33413_, _13498_, \oc8051_golden_model_1.IP [3]);
  and (_33414_, _14950_, _08632_);
  or (_33415_, _33414_, _33413_);
  and (_33416_, _33415_, _06272_);
  or (_33417_, _33416_, _06461_);
  or (_33418_, _33417_, _33412_);
  or (_33419_, _33398_, _07166_);
  and (_33420_, _33419_, _33418_);
  or (_33421_, _33420_, _06464_);
  or (_33423_, _33405_, _06465_);
  and (_33424_, _33423_, _06269_);
  and (_33425_, _33424_, _33421_);
  and (_33426_, _14948_, _08632_);
  or (_33427_, _33426_, _33413_);
  and (_33428_, _33427_, _06268_);
  or (_33429_, _33428_, _06261_);
  or (_33430_, _33429_, _33425_);
  or (_33431_, _33413_, _14979_);
  and (_33432_, _33431_, _33415_);
  or (_33434_, _33432_, _06262_);
  and (_33435_, _33434_, _06258_);
  and (_33436_, _33435_, _33430_);
  or (_33437_, _33413_, _14992_);
  and (_33438_, _33437_, _06257_);
  and (_33439_, _33438_, _33415_);
  or (_33440_, _33439_, _10080_);
  or (_33441_, _33440_, _33436_);
  and (_33442_, _33441_, _33399_);
  or (_33443_, _33442_, _07460_);
  and (_33445_, _09449_, _07946_);
  or (_33446_, _33396_, _07208_);
  or (_33447_, _33446_, _33445_);
  and (_33448_, _33447_, _05982_);
  and (_33449_, _33448_, _33443_);
  and (_33450_, _15048_, _07946_);
  or (_33451_, _33450_, _33396_);
  and (_33452_, _33451_, _10094_);
  or (_33453_, _33452_, _06218_);
  or (_33454_, _33453_, _33449_);
  and (_33456_, _07946_, _08930_);
  or (_33457_, _33456_, _33396_);
  or (_33458_, _33457_, _06219_);
  and (_33459_, _33458_, _33454_);
  or (_33460_, _33459_, _06369_);
  and (_33461_, _14943_, _07946_);
  or (_33462_, _33461_, _33396_);
  or (_33463_, _33462_, _07237_);
  and (_33464_, _33463_, _07240_);
  and (_33465_, _33464_, _33460_);
  and (_33467_, _12577_, _07946_);
  or (_33468_, _33467_, _33396_);
  and (_33469_, _33468_, _06536_);
  or (_33470_, _33469_, _33465_);
  and (_33471_, _33470_, _07242_);
  or (_33472_, _33396_, _08292_);
  and (_33473_, _33457_, _06375_);
  and (_33474_, _33473_, _33472_);
  or (_33475_, _33474_, _33471_);
  and (_33476_, _33475_, _07234_);
  and (_33478_, _33405_, _06545_);
  and (_33479_, _33478_, _33472_);
  or (_33480_, _33479_, _06366_);
  or (_33481_, _33480_, _33476_);
  and (_33482_, _14940_, _07946_);
  or (_33483_, _33396_, _09056_);
  or (_33484_, _33483_, _33482_);
  and (_33485_, _33484_, _09061_);
  and (_33486_, _33485_, _33481_);
  nor (_33487_, _11256_, _13490_);
  or (_33489_, _33487_, _33396_);
  and (_33490_, _33489_, _06528_);
  or (_33491_, _33490_, _06568_);
  or (_33492_, _33491_, _33486_);
  or (_33493_, _33402_, _06926_);
  and (_33494_, _33493_, _05928_);
  and (_33495_, _33494_, _33492_);
  and (_33496_, _33427_, _05927_);
  or (_33497_, _33496_, _06278_);
  or (_33498_, _33497_, _33495_);
  and (_33500_, _15128_, _07946_);
  or (_33501_, _33396_, _06279_);
  or (_33502_, _33501_, _33500_);
  and (_33503_, _33502_, _01347_);
  and (_33504_, _33503_, _33498_);
  or (_33505_, _33504_, _33395_);
  and (_43299_, _33505_, _42618_);
  and (_33506_, _01351_, \oc8051_golden_model_1.IP [4]);
  and (_33507_, _13490_, \oc8051_golden_model_1.IP [4]);
  nor (_33508_, _08541_, _13490_);
  or (_33510_, _33508_, _33507_);
  or (_33511_, _33510_, _07215_);
  and (_33512_, _13498_, \oc8051_golden_model_1.IP [4]);
  and (_33513_, _15176_, _08632_);
  or (_33514_, _33513_, _33512_);
  and (_33515_, _33514_, _06268_);
  and (_33516_, _15162_, _07946_);
  or (_33517_, _33516_, _33507_);
  or (_33518_, _33517_, _07151_);
  and (_33519_, _07946_, \oc8051_golden_model_1.ACC [4]);
  or (_33521_, _33519_, _33507_);
  and (_33522_, _33521_, _07141_);
  and (_33523_, _07142_, \oc8051_golden_model_1.IP [4]);
  or (_33524_, _33523_, _06341_);
  or (_33525_, _33524_, _33522_);
  and (_33526_, _33525_, _06273_);
  and (_33527_, _33526_, _33518_);
  and (_33528_, _15166_, _08632_);
  or (_33529_, _33528_, _33512_);
  and (_33530_, _33529_, _06272_);
  or (_33532_, _33530_, _06461_);
  or (_33533_, _33532_, _33527_);
  or (_33534_, _33510_, _07166_);
  and (_33535_, _33534_, _33533_);
  or (_33536_, _33535_, _06464_);
  or (_33537_, _33521_, _06465_);
  and (_33538_, _33537_, _06269_);
  and (_33539_, _33538_, _33536_);
  or (_33540_, _33539_, _33515_);
  and (_33541_, _33540_, _06262_);
  or (_33543_, _33512_, _15183_);
  and (_33544_, _33543_, _06261_);
  and (_33545_, _33544_, _33529_);
  or (_33546_, _33545_, _33541_);
  and (_33547_, _33546_, _06258_);
  and (_33548_, _15200_, _08632_);
  or (_33549_, _33548_, _33512_);
  and (_33550_, _33549_, _06257_);
  or (_33551_, _33550_, _10080_);
  or (_33552_, _33551_, _33547_);
  and (_33554_, _33552_, _33511_);
  or (_33555_, _33554_, _07460_);
  and (_33556_, _09448_, _07946_);
  or (_33557_, _33507_, _07208_);
  or (_33558_, _33557_, _33556_);
  and (_33559_, _33558_, _05982_);
  and (_33560_, _33559_, _33555_);
  and (_33561_, _15254_, _07946_);
  or (_33562_, _33561_, _33507_);
  and (_33563_, _33562_, _10094_);
  or (_33565_, _33563_, _06218_);
  or (_33566_, _33565_, _33560_);
  and (_33567_, _08959_, _07946_);
  or (_33568_, _33567_, _33507_);
  or (_33569_, _33568_, _06219_);
  and (_33570_, _33569_, _33566_);
  or (_33571_, _33570_, _06369_);
  and (_33572_, _15269_, _07946_);
  or (_33573_, _33572_, _33507_);
  or (_33574_, _33573_, _07237_);
  and (_33576_, _33574_, _07240_);
  and (_33577_, _33576_, _33571_);
  and (_33578_, _11254_, _07946_);
  or (_33579_, _33578_, _33507_);
  and (_33580_, _33579_, _06536_);
  or (_33581_, _33580_, _33577_);
  and (_33582_, _33581_, _07242_);
  or (_33583_, _33507_, _08544_);
  and (_33584_, _33568_, _06375_);
  and (_33585_, _33584_, _33583_);
  or (_33587_, _33585_, _33582_);
  and (_33588_, _33587_, _07234_);
  and (_33589_, _33521_, _06545_);
  and (_33590_, _33589_, _33583_);
  or (_33591_, _33590_, _06366_);
  or (_33592_, _33591_, _33588_);
  and (_33593_, _15266_, _07946_);
  or (_33594_, _33507_, _09056_);
  or (_33595_, _33594_, _33593_);
  and (_33596_, _33595_, _09061_);
  and (_33598_, _33596_, _33592_);
  nor (_33599_, _11253_, _13490_);
  or (_33600_, _33599_, _33507_);
  and (_33601_, _33600_, _06528_);
  or (_33602_, _33601_, _06568_);
  or (_33603_, _33602_, _33598_);
  or (_33604_, _33517_, _06926_);
  and (_33605_, _33604_, _05928_);
  and (_33606_, _33605_, _33603_);
  and (_33607_, _33514_, _05927_);
  or (_33609_, _33607_, _06278_);
  or (_33610_, _33609_, _33606_);
  and (_33611_, _15329_, _07946_);
  or (_33612_, _33507_, _06279_);
  or (_33613_, _33612_, _33611_);
  and (_33614_, _33613_, _01347_);
  and (_33615_, _33614_, _33610_);
  or (_33616_, _33615_, _33506_);
  and (_43300_, _33616_, _42618_);
  and (_33617_, _01351_, \oc8051_golden_model_1.IP [5]);
  and (_33619_, _13490_, \oc8051_golden_model_1.IP [5]);
  and (_33620_, _15358_, _07946_);
  or (_33621_, _33620_, _33619_);
  or (_33622_, _33621_, _07151_);
  and (_33623_, _07946_, \oc8051_golden_model_1.ACC [5]);
  or (_33624_, _33623_, _33619_);
  and (_33625_, _33624_, _07141_);
  and (_33626_, _07142_, \oc8051_golden_model_1.IP [5]);
  or (_33627_, _33626_, _06341_);
  or (_33628_, _33627_, _33625_);
  and (_33630_, _33628_, _06273_);
  and (_33631_, _33630_, _33622_);
  and (_33632_, _13498_, \oc8051_golden_model_1.IP [5]);
  and (_33633_, _15372_, _08632_);
  or (_33634_, _33633_, _33632_);
  and (_33635_, _33634_, _06272_);
  or (_33636_, _33635_, _06461_);
  or (_33637_, _33636_, _33631_);
  nor (_33638_, _08244_, _13490_);
  or (_33639_, _33638_, _33619_);
  or (_33641_, _33639_, _07166_);
  and (_33642_, _33641_, _33637_);
  or (_33643_, _33642_, _06464_);
  or (_33644_, _33624_, _06465_);
  and (_33645_, _33644_, _06269_);
  and (_33646_, _33645_, _33643_);
  and (_33647_, _15355_, _08632_);
  or (_33648_, _33647_, _33632_);
  and (_33649_, _33648_, _06268_);
  or (_33650_, _33649_, _06261_);
  or (_33652_, _33650_, _33646_);
  or (_33653_, _33632_, _15387_);
  and (_33654_, _33653_, _33634_);
  or (_33655_, _33654_, _06262_);
  and (_33656_, _33655_, _06258_);
  and (_33657_, _33656_, _33652_);
  or (_33658_, _33632_, _15403_);
  and (_33659_, _33658_, _06257_);
  and (_33660_, _33659_, _33634_);
  or (_33661_, _33660_, _10080_);
  or (_33663_, _33661_, _33657_);
  or (_33664_, _33639_, _07215_);
  and (_33665_, _33664_, _33663_);
  or (_33666_, _33665_, _07460_);
  and (_33667_, _09447_, _07946_);
  or (_33668_, _33619_, _07208_);
  or (_33669_, _33668_, _33667_);
  and (_33670_, _33669_, _05982_);
  and (_33671_, _33670_, _33666_);
  and (_33672_, _15459_, _07946_);
  or (_33674_, _33672_, _33619_);
  and (_33675_, _33674_, _10094_);
  or (_33676_, _33675_, _06218_);
  or (_33677_, _33676_, _33671_);
  and (_33678_, _08946_, _07946_);
  or (_33679_, _33678_, _33619_);
  or (_33680_, _33679_, _06219_);
  and (_33681_, _33680_, _33677_);
  or (_33682_, _33681_, _06369_);
  and (_33683_, _15353_, _07946_);
  or (_33685_, _33683_, _33619_);
  or (_33686_, _33685_, _07237_);
  and (_33687_, _33686_, _07240_);
  and (_33688_, _33687_, _33682_);
  and (_33689_, _11250_, _07946_);
  or (_33690_, _33689_, _33619_);
  and (_33691_, _33690_, _06536_);
  or (_33692_, _33691_, _33688_);
  and (_33693_, _33692_, _07242_);
  or (_33694_, _33619_, _08247_);
  and (_33696_, _33679_, _06375_);
  and (_33697_, _33696_, _33694_);
  or (_33698_, _33697_, _33693_);
  and (_33699_, _33698_, _07234_);
  and (_33700_, _33624_, _06545_);
  and (_33701_, _33700_, _33694_);
  or (_33702_, _33701_, _06366_);
  or (_33703_, _33702_, _33699_);
  and (_33704_, _15350_, _07946_);
  or (_33705_, _33619_, _09056_);
  or (_33707_, _33705_, _33704_);
  and (_33708_, _33707_, _09061_);
  and (_33709_, _33708_, _33703_);
  nor (_33710_, _11249_, _13490_);
  or (_33711_, _33710_, _33619_);
  and (_33712_, _33711_, _06528_);
  or (_33713_, _33712_, _06568_);
  or (_33714_, _33713_, _33709_);
  or (_33715_, _33621_, _06926_);
  and (_33716_, _33715_, _05928_);
  and (_33718_, _33716_, _33714_);
  and (_33719_, _33648_, _05927_);
  or (_33720_, _33719_, _06278_);
  or (_33721_, _33720_, _33718_);
  and (_33722_, _15532_, _07946_);
  or (_33723_, _33619_, _06279_);
  or (_33724_, _33723_, _33722_);
  and (_33725_, _33724_, _01347_);
  and (_33726_, _33725_, _33721_);
  or (_33727_, _33726_, _33617_);
  and (_43302_, _33727_, _42618_);
  and (_33729_, _01351_, \oc8051_golden_model_1.IP [6]);
  and (_33730_, _13490_, \oc8051_golden_model_1.IP [6]);
  and (_33731_, _15554_, _07946_);
  or (_33732_, _33731_, _33730_);
  or (_33733_, _33732_, _07151_);
  and (_33734_, _07946_, \oc8051_golden_model_1.ACC [6]);
  or (_33735_, _33734_, _33730_);
  and (_33736_, _33735_, _07141_);
  and (_33737_, _07142_, \oc8051_golden_model_1.IP [6]);
  or (_33739_, _33737_, _06341_);
  or (_33740_, _33739_, _33736_);
  and (_33741_, _33740_, _06273_);
  and (_33742_, _33741_, _33733_);
  and (_33743_, _13498_, \oc8051_golden_model_1.IP [6]);
  and (_33744_, _15570_, _08632_);
  or (_33745_, _33744_, _33743_);
  and (_33746_, _33745_, _06272_);
  or (_33747_, _33746_, _06461_);
  or (_33748_, _33747_, _33742_);
  nor (_33750_, _08142_, _13490_);
  or (_33751_, _33750_, _33730_);
  or (_33752_, _33751_, _07166_);
  and (_33753_, _33752_, _33748_);
  or (_33754_, _33753_, _06464_);
  or (_33755_, _33735_, _06465_);
  and (_33756_, _33755_, _06269_);
  and (_33757_, _33756_, _33754_);
  and (_33758_, _15551_, _08632_);
  or (_33759_, _33758_, _33743_);
  and (_33761_, _33759_, _06268_);
  or (_33762_, _33761_, _06261_);
  or (_33763_, _33762_, _33757_);
  or (_33764_, _33743_, _15585_);
  and (_33765_, _33764_, _33745_);
  or (_33766_, _33765_, _06262_);
  and (_33767_, _33766_, _06258_);
  and (_33768_, _33767_, _33763_);
  and (_33769_, _15602_, _08632_);
  or (_33770_, _33769_, _33743_);
  and (_33772_, _33770_, _06257_);
  or (_33773_, _33772_, _10080_);
  or (_33774_, _33773_, _33768_);
  or (_33775_, _33751_, _07215_);
  and (_33776_, _33775_, _33774_);
  or (_33777_, _33776_, _07460_);
  and (_33778_, _09446_, _07946_);
  or (_33779_, _33730_, _07208_);
  or (_33780_, _33779_, _33778_);
  and (_33781_, _33780_, _05982_);
  and (_33783_, _33781_, _33777_);
  and (_33784_, _15657_, _07946_);
  or (_33785_, _33784_, _33730_);
  and (_33786_, _33785_, _10094_);
  or (_33787_, _33786_, _06218_);
  or (_33788_, _33787_, _33783_);
  and (_33789_, _15664_, _07946_);
  or (_33790_, _33789_, _33730_);
  or (_33791_, _33790_, _06219_);
  and (_33792_, _33791_, _33788_);
  or (_33794_, _33792_, _06369_);
  and (_33795_, _15549_, _07946_);
  or (_33796_, _33795_, _33730_);
  or (_33797_, _33796_, _07237_);
  and (_33798_, _33797_, _07240_);
  and (_33799_, _33798_, _33794_);
  and (_33800_, _11247_, _07946_);
  or (_33801_, _33800_, _33730_);
  and (_33802_, _33801_, _06536_);
  or (_33803_, _33802_, _33799_);
  and (_33805_, _33803_, _07242_);
  or (_33806_, _33730_, _08145_);
  and (_33807_, _33790_, _06375_);
  and (_33808_, _33807_, _33806_);
  or (_33809_, _33808_, _33805_);
  and (_33810_, _33809_, _07234_);
  and (_33811_, _33735_, _06545_);
  and (_33812_, _33811_, _33806_);
  or (_33813_, _33812_, _06366_);
  or (_33814_, _33813_, _33810_);
  and (_33816_, _15546_, _07946_);
  or (_33817_, _33730_, _09056_);
  or (_33818_, _33817_, _33816_);
  and (_33819_, _33818_, _09061_);
  and (_33820_, _33819_, _33814_);
  nor (_33821_, _11246_, _13490_);
  or (_33822_, _33821_, _33730_);
  and (_33823_, _33822_, _06528_);
  or (_33824_, _33823_, _06568_);
  or (_33825_, _33824_, _33820_);
  or (_33827_, _33732_, _06926_);
  and (_33828_, _33827_, _05928_);
  and (_33829_, _33828_, _33825_);
  and (_33830_, _33759_, _05927_);
  or (_33831_, _33830_, _06278_);
  or (_33832_, _33831_, _33829_);
  and (_33833_, _15734_, _07946_);
  or (_33834_, _33730_, _06279_);
  or (_33835_, _33834_, _33833_);
  and (_33836_, _33835_, _01347_);
  and (_33838_, _33836_, _33832_);
  or (_33839_, _33838_, _33729_);
  and (_43303_, _33839_, _42618_);
  and (_33840_, _01351_, \oc8051_golden_model_1.IE [0]);
  and (_33841_, _07900_, \oc8051_golden_model_1.ACC [0]);
  and (_33842_, _33841_, _08390_);
  and (_33843_, _13593_, \oc8051_golden_model_1.IE [0]);
  or (_33844_, _33843_, _07234_);
  or (_33845_, _33844_, _33842_);
  and (_33846_, _07900_, _07133_);
  or (_33848_, _33846_, _33843_);
  or (_33849_, _33848_, _07215_);
  nor (_33850_, _08390_, _13593_);
  or (_33851_, _33850_, _33843_);
  and (_33852_, _33851_, _06341_);
  and (_33853_, _07142_, \oc8051_golden_model_1.IE [0]);
  or (_33854_, _33841_, _33843_);
  and (_33855_, _33854_, _07141_);
  or (_33856_, _33855_, _33853_);
  and (_33857_, _33856_, _07151_);
  or (_33859_, _33857_, _06272_);
  or (_33860_, _33859_, _33852_);
  and (_33861_, _14382_, _08626_);
  and (_33862_, _13601_, \oc8051_golden_model_1.IE [0]);
  or (_33863_, _33862_, _06273_);
  or (_33864_, _33863_, _33861_);
  and (_33865_, _33864_, _07166_);
  and (_33866_, _33865_, _33860_);
  and (_33867_, _33848_, _06461_);
  or (_33868_, _33867_, _06464_);
  or (_33870_, _33868_, _33866_);
  or (_33871_, _33854_, _06465_);
  and (_33872_, _33871_, _06269_);
  and (_33873_, _33872_, _33870_);
  and (_33874_, _33843_, _06268_);
  or (_33875_, _33874_, _06261_);
  or (_33876_, _33875_, _33873_);
  or (_33877_, _33851_, _06262_);
  and (_33878_, _33877_, _06258_);
  and (_33879_, _33878_, _33876_);
  and (_33881_, _14413_, _08626_);
  or (_33882_, _33881_, _33862_);
  and (_33883_, _33882_, _06257_);
  or (_33884_, _33883_, _10080_);
  or (_33885_, _33884_, _33879_);
  and (_33886_, _33885_, _33849_);
  or (_33887_, _33886_, _07460_);
  and (_33888_, _09392_, _07900_);
  or (_33889_, _33843_, _07208_);
  or (_33890_, _33889_, _33888_);
  and (_33892_, _33890_, _33887_);
  or (_33893_, _33892_, _10094_);
  and (_33894_, _14467_, _07900_);
  or (_33895_, _33843_, _05982_);
  or (_33896_, _33895_, _33894_);
  and (_33897_, _33896_, _06219_);
  and (_33898_, _33897_, _33893_);
  and (_33899_, _07900_, _08954_);
  or (_33900_, _33899_, _33843_);
  and (_33901_, _33900_, _06218_);
  or (_33903_, _33901_, _06369_);
  or (_33904_, _33903_, _33898_);
  and (_33905_, _14366_, _07900_);
  or (_33906_, _33905_, _33843_);
  or (_33907_, _33906_, _07237_);
  and (_33908_, _33907_, _07240_);
  and (_33909_, _33908_, _33904_);
  nor (_33910_, _12580_, _13593_);
  or (_33911_, _33910_, _33843_);
  nor (_33912_, _33842_, _07240_);
  and (_33914_, _33912_, _33911_);
  or (_33915_, _33914_, _33909_);
  and (_33916_, _33915_, _07242_);
  nand (_33917_, _33900_, _06375_);
  nor (_33918_, _33917_, _33850_);
  or (_33919_, _33918_, _06545_);
  or (_33920_, _33919_, _33916_);
  and (_33921_, _33920_, _33845_);
  or (_33922_, _33921_, _06366_);
  and (_33923_, _14363_, _07900_);
  or (_33925_, _33843_, _09056_);
  or (_33926_, _33925_, _33923_);
  and (_33927_, _33926_, _09061_);
  and (_33928_, _33927_, _33922_);
  and (_33929_, _33911_, _06528_);
  or (_33930_, _33929_, _06568_);
  or (_33931_, _33930_, _33928_);
  or (_33932_, _33851_, _06926_);
  and (_33933_, _33932_, _33931_);
  or (_33934_, _33933_, _05927_);
  or (_33936_, _33843_, _05928_);
  and (_33937_, _33936_, _33934_);
  or (_33938_, _33937_, _06278_);
  or (_33939_, _33851_, _06279_);
  and (_33940_, _33939_, _01347_);
  and (_33941_, _33940_, _33938_);
  or (_33942_, _33941_, _33840_);
  and (_43304_, _33942_, _42618_);
  not (_33943_, \oc8051_golden_model_1.IE [1]);
  nor (_33944_, _01347_, _33943_);
  nor (_33946_, _07900_, _33943_);
  nor (_33947_, _11261_, _13593_);
  or (_33948_, _33947_, _33946_);
  or (_33949_, _33948_, _09061_);
  nand (_33950_, _07900_, _07038_);
  or (_33951_, _07900_, \oc8051_golden_model_1.IE [1]);
  and (_33952_, _33951_, _06218_);
  and (_33953_, _33952_, _33950_);
  nor (_33954_, _13593_, _07357_);
  or (_33955_, _33954_, _33946_);
  or (_33957_, _33955_, _07166_);
  and (_33958_, _14562_, _07900_);
  not (_33959_, _33958_);
  and (_33960_, _33959_, _33951_);
  or (_33961_, _33960_, _07151_);
  and (_33962_, _07900_, \oc8051_golden_model_1.ACC [1]);
  or (_33963_, _33962_, _33946_);
  and (_33964_, _33963_, _07141_);
  nor (_33965_, _07141_, _33943_);
  or (_33966_, _33965_, _06341_);
  or (_33967_, _33966_, _33964_);
  and (_33968_, _33967_, _06273_);
  and (_33969_, _33968_, _33961_);
  nor (_33970_, _08626_, _33943_);
  and (_33971_, _14557_, _08626_);
  or (_33972_, _33971_, _33970_);
  and (_33973_, _33972_, _06272_);
  or (_33974_, _33973_, _06461_);
  or (_33975_, _33974_, _33969_);
  and (_33976_, _33975_, _33957_);
  or (_33978_, _33976_, _06464_);
  or (_33979_, _33963_, _06465_);
  and (_33980_, _33979_, _06269_);
  and (_33981_, _33980_, _33978_);
  and (_33982_, _14560_, _08626_);
  or (_33983_, _33982_, _33970_);
  and (_33984_, _33983_, _06268_);
  or (_33985_, _33984_, _06261_);
  or (_33986_, _33985_, _33981_);
  and (_33987_, _33971_, _14556_);
  or (_33989_, _33970_, _06262_);
  or (_33990_, _33989_, _33987_);
  and (_33991_, _33990_, _06258_);
  and (_33992_, _33991_, _33986_);
  or (_33993_, _33970_, _14597_);
  and (_33994_, _33993_, _06257_);
  and (_33995_, _33994_, _33972_);
  or (_33996_, _33995_, _10080_);
  or (_33997_, _33996_, _33992_);
  or (_33998_, _33955_, _07215_);
  and (_34000_, _33998_, _33997_);
  or (_34001_, _34000_, _07460_);
  and (_34002_, _09451_, _07900_);
  or (_34003_, _33946_, _07208_);
  or (_34004_, _34003_, _34002_);
  and (_34005_, _34004_, _05982_);
  and (_34006_, _34005_, _34001_);
  and (_34007_, _14653_, _07900_);
  or (_34008_, _34007_, _33946_);
  and (_34009_, _34008_, _10094_);
  or (_34011_, _34009_, _34006_);
  and (_34012_, _34011_, _06219_);
  or (_34013_, _34012_, _33953_);
  and (_34014_, _34013_, _07237_);
  or (_34015_, _14668_, _13593_);
  and (_34016_, _33951_, _06369_);
  and (_34017_, _34016_, _34015_);
  or (_34018_, _34017_, _06536_);
  or (_34019_, _34018_, _34014_);
  nand (_34020_, _11260_, _07900_);
  and (_34022_, _34020_, _33948_);
  or (_34023_, _34022_, _07240_);
  and (_34024_, _34023_, _07242_);
  and (_34025_, _34024_, _34019_);
  or (_34026_, _14666_, _13593_);
  and (_34027_, _33951_, _06375_);
  and (_34028_, _34027_, _34026_);
  or (_34029_, _34028_, _06545_);
  or (_34030_, _34029_, _34025_);
  nor (_34031_, _33946_, _07234_);
  nand (_34033_, _34031_, _34020_);
  and (_34034_, _34033_, _09056_);
  and (_34035_, _34034_, _34030_);
  or (_34036_, _33950_, _08341_);
  and (_34037_, _33951_, _06366_);
  and (_34038_, _34037_, _34036_);
  or (_34039_, _34038_, _06528_);
  or (_34040_, _34039_, _34035_);
  and (_34041_, _34040_, _33949_);
  or (_34042_, _34041_, _06568_);
  or (_34044_, _33960_, _06926_);
  and (_34045_, _34044_, _05928_);
  and (_34046_, _34045_, _34042_);
  and (_34047_, _33983_, _05927_);
  or (_34048_, _34047_, _06278_);
  or (_34049_, _34048_, _34046_);
  or (_34050_, _33946_, _06279_);
  or (_34051_, _34050_, _33958_);
  and (_34052_, _34051_, _01347_);
  and (_34053_, _34052_, _34049_);
  or (_34055_, _34053_, _33944_);
  and (_43306_, _34055_, _42618_);
  and (_34056_, _01351_, \oc8051_golden_model_1.IE [2]);
  and (_34057_, _13593_, \oc8051_golden_model_1.IE [2]);
  nor (_34058_, _13593_, _07776_);
  or (_34059_, _34058_, _34057_);
  or (_34060_, _34059_, _07215_);
  or (_34061_, _34059_, _07166_);
  and (_34062_, _14770_, _07900_);
  or (_34063_, _34062_, _34057_);
  or (_34065_, _34063_, _07151_);
  and (_34066_, _07900_, \oc8051_golden_model_1.ACC [2]);
  or (_34067_, _34066_, _34057_);
  and (_34068_, _34067_, _07141_);
  and (_34069_, _07142_, \oc8051_golden_model_1.IE [2]);
  or (_34070_, _34069_, _06341_);
  or (_34071_, _34070_, _34068_);
  and (_34072_, _34071_, _06273_);
  and (_34073_, _34072_, _34065_);
  and (_34074_, _13601_, \oc8051_golden_model_1.IE [2]);
  and (_34076_, _14774_, _08626_);
  or (_34077_, _34076_, _34074_);
  and (_34078_, _34077_, _06272_);
  or (_34079_, _34078_, _06461_);
  or (_34080_, _34079_, _34073_);
  and (_34081_, _34080_, _34061_);
  or (_34082_, _34081_, _06464_);
  or (_34083_, _34067_, _06465_);
  and (_34084_, _34083_, _06269_);
  and (_34085_, _34084_, _34082_);
  and (_34087_, _14756_, _08626_);
  or (_34088_, _34087_, _34074_);
  and (_34089_, _34088_, _06268_);
  or (_34090_, _34089_, _06261_);
  or (_34091_, _34090_, _34085_);
  and (_34092_, _34076_, _14789_);
  or (_34093_, _34074_, _06262_);
  or (_34094_, _34093_, _34092_);
  and (_34095_, _34094_, _06258_);
  and (_34096_, _34095_, _34091_);
  and (_34098_, _14804_, _08626_);
  or (_34099_, _34098_, _34074_);
  and (_34100_, _34099_, _06257_);
  or (_34101_, _34100_, _10080_);
  or (_34102_, _34101_, _34096_);
  and (_34103_, _34102_, _34060_);
  or (_34104_, _34103_, _07460_);
  and (_34105_, _09450_, _07900_);
  or (_34106_, _34057_, _07208_);
  or (_34107_, _34106_, _34105_);
  and (_34109_, _34107_, _05982_);
  and (_34110_, _34109_, _34104_);
  and (_34111_, _14859_, _07900_);
  or (_34112_, _34111_, _34057_);
  and (_34113_, _34112_, _10094_);
  or (_34114_, _34113_, _06218_);
  or (_34115_, _34114_, _34110_);
  and (_34116_, _07900_, _08973_);
  or (_34117_, _34116_, _34057_);
  or (_34118_, _34117_, _06219_);
  and (_34120_, _34118_, _34115_);
  or (_34121_, _34120_, _06369_);
  and (_34122_, _14751_, _07900_);
  or (_34123_, _34122_, _34057_);
  or (_34124_, _34123_, _07237_);
  and (_34125_, _34124_, _07240_);
  and (_34126_, _34125_, _34121_);
  and (_34127_, _11259_, _07900_);
  or (_34128_, _34127_, _34057_);
  and (_34129_, _34128_, _06536_);
  or (_34131_, _34129_, _34126_);
  and (_34132_, _34131_, _07242_);
  or (_34133_, _34057_, _08440_);
  and (_34134_, _34117_, _06375_);
  and (_34135_, _34134_, _34133_);
  or (_34136_, _34135_, _34132_);
  and (_34137_, _34136_, _07234_);
  and (_34138_, _34067_, _06545_);
  and (_34139_, _34138_, _34133_);
  or (_34140_, _34139_, _06366_);
  or (_34142_, _34140_, _34137_);
  and (_34143_, _14748_, _07900_);
  or (_34144_, _34057_, _09056_);
  or (_34145_, _34144_, _34143_);
  and (_34146_, _34145_, _09061_);
  and (_34147_, _34146_, _34142_);
  nor (_34148_, _11258_, _13593_);
  or (_34149_, _34148_, _34057_);
  and (_34150_, _34149_, _06528_);
  or (_34151_, _34150_, _06568_);
  or (_34153_, _34151_, _34147_);
  or (_34154_, _34063_, _06926_);
  and (_34155_, _34154_, _05928_);
  and (_34156_, _34155_, _34153_);
  and (_34157_, _34088_, _05927_);
  or (_34158_, _34157_, _06278_);
  or (_34159_, _34158_, _34156_);
  and (_34160_, _14926_, _07900_);
  or (_34161_, _34057_, _06279_);
  or (_34162_, _34161_, _34160_);
  and (_34164_, _34162_, _01347_);
  and (_34165_, _34164_, _34159_);
  or (_34166_, _34165_, _34056_);
  and (_43307_, _34166_, _42618_);
  and (_34167_, _01351_, \oc8051_golden_model_1.IE [3]);
  and (_34168_, _13593_, \oc8051_golden_model_1.IE [3]);
  nor (_34169_, _13593_, _07594_);
  or (_34170_, _34169_, _34168_);
  or (_34171_, _34170_, _07215_);
  and (_34172_, _14953_, _07900_);
  or (_34174_, _34172_, _34168_);
  or (_34175_, _34174_, _07151_);
  and (_34176_, _07900_, \oc8051_golden_model_1.ACC [3]);
  or (_34177_, _34176_, _34168_);
  and (_34178_, _34177_, _07141_);
  and (_34179_, _07142_, \oc8051_golden_model_1.IE [3]);
  or (_34180_, _34179_, _06341_);
  or (_34181_, _34180_, _34178_);
  and (_34183_, _34181_, _06273_);
  and (_34185_, _34183_, _34175_);
  and (_34188_, _13601_, \oc8051_golden_model_1.IE [3]);
  and (_34190_, _14950_, _08626_);
  or (_34192_, _34190_, _34188_);
  and (_34194_, _34192_, _06272_);
  or (_34196_, _34194_, _06461_);
  or (_34198_, _34196_, _34185_);
  or (_34200_, _34170_, _07166_);
  and (_34202_, _34200_, _34198_);
  or (_34203_, _34202_, _06464_);
  or (_34204_, _34177_, _06465_);
  and (_34206_, _34204_, _06269_);
  and (_34207_, _34206_, _34203_);
  and (_34208_, _14948_, _08626_);
  or (_34209_, _34208_, _34188_);
  and (_34210_, _34209_, _06268_);
  or (_34211_, _34210_, _06261_);
  or (_34212_, _34211_, _34207_);
  or (_34213_, _34188_, _14979_);
  and (_34214_, _34213_, _34192_);
  or (_34215_, _34214_, _06262_);
  and (_34217_, _34215_, _06258_);
  and (_34218_, _34217_, _34212_);
  or (_34219_, _34188_, _14992_);
  and (_34220_, _34219_, _06257_);
  and (_34221_, _34220_, _34192_);
  or (_34222_, _34221_, _10080_);
  or (_34223_, _34222_, _34218_);
  and (_34224_, _34223_, _34171_);
  or (_34225_, _34224_, _07460_);
  and (_34226_, _09449_, _07900_);
  or (_34228_, _34168_, _07208_);
  or (_34229_, _34228_, _34226_);
  and (_34230_, _34229_, _05982_);
  and (_34231_, _34230_, _34225_);
  and (_34232_, _15048_, _07900_);
  or (_34233_, _34232_, _34168_);
  and (_34234_, _34233_, _10094_);
  or (_34235_, _34234_, _06218_);
  or (_34236_, _34235_, _34231_);
  and (_34237_, _07900_, _08930_);
  or (_34239_, _34237_, _34168_);
  or (_34240_, _34239_, _06219_);
  and (_34241_, _34240_, _34236_);
  or (_34242_, _34241_, _06369_);
  and (_34243_, _14943_, _07900_);
  or (_34244_, _34243_, _34168_);
  or (_34245_, _34244_, _07237_);
  and (_34246_, _34245_, _07240_);
  and (_34247_, _34246_, _34242_);
  and (_34248_, _12577_, _07900_);
  or (_34250_, _34248_, _34168_);
  and (_34251_, _34250_, _06536_);
  or (_34252_, _34251_, _34247_);
  and (_34253_, _34252_, _07242_);
  or (_34254_, _34168_, _08292_);
  and (_34255_, _34239_, _06375_);
  and (_34256_, _34255_, _34254_);
  or (_34257_, _34256_, _34253_);
  and (_34258_, _34257_, _07234_);
  and (_34259_, _34177_, _06545_);
  and (_34261_, _34259_, _34254_);
  or (_34262_, _34261_, _06366_);
  or (_34263_, _34262_, _34258_);
  and (_34264_, _14940_, _07900_);
  or (_34265_, _34168_, _09056_);
  or (_34266_, _34265_, _34264_);
  and (_34267_, _34266_, _09061_);
  and (_34268_, _34267_, _34263_);
  nor (_34269_, _11256_, _13593_);
  or (_34270_, _34269_, _34168_);
  and (_34272_, _34270_, _06528_);
  or (_34273_, _34272_, _06568_);
  or (_34274_, _34273_, _34268_);
  or (_34275_, _34174_, _06926_);
  and (_34276_, _34275_, _05928_);
  and (_34277_, _34276_, _34274_);
  and (_34278_, _34209_, _05927_);
  or (_34279_, _34278_, _06278_);
  or (_34280_, _34279_, _34277_);
  and (_34281_, _15128_, _07900_);
  or (_34283_, _34168_, _06279_);
  or (_34284_, _34283_, _34281_);
  and (_34285_, _34284_, _01347_);
  and (_34286_, _34285_, _34280_);
  or (_34287_, _34286_, _34167_);
  and (_43308_, _34287_, _42618_);
  and (_34288_, _01351_, \oc8051_golden_model_1.IE [4]);
  and (_34289_, _13593_, \oc8051_golden_model_1.IE [4]);
  nor (_34290_, _08541_, _13593_);
  or (_34291_, _34290_, _34289_);
  or (_34293_, _34291_, _07215_);
  and (_34294_, _13601_, \oc8051_golden_model_1.IE [4]);
  and (_34295_, _15176_, _08626_);
  or (_34296_, _34295_, _34294_);
  and (_34297_, _34296_, _06268_);
  and (_34298_, _15162_, _07900_);
  or (_34299_, _34298_, _34289_);
  or (_34300_, _34299_, _07151_);
  and (_34301_, _07900_, \oc8051_golden_model_1.ACC [4]);
  or (_34302_, _34301_, _34289_);
  and (_34304_, _34302_, _07141_);
  and (_34305_, _07142_, \oc8051_golden_model_1.IE [4]);
  or (_34306_, _34305_, _06341_);
  or (_34307_, _34306_, _34304_);
  and (_34308_, _34307_, _06273_);
  and (_34309_, _34308_, _34300_);
  and (_34310_, _15166_, _08626_);
  or (_34311_, _34310_, _34294_);
  and (_34312_, _34311_, _06272_);
  or (_34313_, _34312_, _06461_);
  or (_34315_, _34313_, _34309_);
  or (_34316_, _34291_, _07166_);
  and (_34317_, _34316_, _34315_);
  or (_34318_, _34317_, _06464_);
  or (_34319_, _34302_, _06465_);
  and (_34320_, _34319_, _06269_);
  and (_34321_, _34320_, _34318_);
  or (_34322_, _34321_, _34297_);
  and (_34323_, _34322_, _06262_);
  and (_34324_, _15184_, _08626_);
  or (_34326_, _34324_, _34294_);
  and (_34327_, _34326_, _06261_);
  or (_34328_, _34327_, _34323_);
  and (_34329_, _34328_, _06258_);
  and (_34330_, _15200_, _08626_);
  or (_34331_, _34330_, _34294_);
  and (_34332_, _34331_, _06257_);
  or (_34333_, _34332_, _10080_);
  or (_34334_, _34333_, _34329_);
  and (_34335_, _34334_, _34293_);
  or (_34337_, _34335_, _07460_);
  and (_34338_, _09448_, _07900_);
  or (_34339_, _34289_, _07208_);
  or (_34340_, _34339_, _34338_);
  and (_34341_, _34340_, _05982_);
  and (_34342_, _34341_, _34337_);
  and (_34343_, _15254_, _07900_);
  or (_34344_, _34343_, _34289_);
  and (_34345_, _34344_, _10094_);
  or (_34346_, _34345_, _06218_);
  or (_34348_, _34346_, _34342_);
  and (_34349_, _08959_, _07900_);
  or (_34350_, _34349_, _34289_);
  or (_34351_, _34350_, _06219_);
  and (_34352_, _34351_, _34348_);
  or (_34353_, _34352_, _06369_);
  and (_34354_, _15269_, _07900_);
  or (_34355_, _34354_, _34289_);
  or (_34356_, _34355_, _07237_);
  and (_34357_, _34356_, _07240_);
  and (_34359_, _34357_, _34353_);
  and (_34360_, _11254_, _07900_);
  or (_34361_, _34360_, _34289_);
  and (_34362_, _34361_, _06536_);
  or (_34363_, _34362_, _34359_);
  and (_34364_, _34363_, _07242_);
  or (_34365_, _34289_, _08544_);
  and (_34366_, _34350_, _06375_);
  and (_34367_, _34366_, _34365_);
  or (_34368_, _34367_, _34364_);
  and (_34370_, _34368_, _07234_);
  and (_34371_, _34302_, _06545_);
  and (_34372_, _34371_, _34365_);
  or (_34373_, _34372_, _06366_);
  or (_34374_, _34373_, _34370_);
  and (_34375_, _15266_, _07900_);
  or (_34376_, _34289_, _09056_);
  or (_34377_, _34376_, _34375_);
  and (_34378_, _34377_, _09061_);
  and (_34379_, _34378_, _34374_);
  nor (_34381_, _11253_, _13593_);
  or (_34382_, _34381_, _34289_);
  and (_34383_, _34382_, _06528_);
  or (_34384_, _34383_, _06568_);
  or (_34385_, _34384_, _34379_);
  or (_34386_, _34299_, _06926_);
  and (_34387_, _34386_, _05928_);
  and (_34388_, _34387_, _34385_);
  and (_34389_, _34296_, _05927_);
  or (_34390_, _34389_, _06278_);
  or (_34392_, _34390_, _34388_);
  and (_34393_, _15329_, _07900_);
  or (_34394_, _34289_, _06279_);
  or (_34395_, _34394_, _34393_);
  and (_34396_, _34395_, _01347_);
  and (_34397_, _34396_, _34392_);
  or (_34398_, _34397_, _34288_);
  and (_43309_, _34398_, _42618_);
  and (_34399_, _01351_, \oc8051_golden_model_1.IE [5]);
  and (_34400_, _13593_, \oc8051_golden_model_1.IE [5]);
  and (_34402_, _15358_, _07900_);
  or (_34403_, _34402_, _34400_);
  or (_34404_, _34403_, _07151_);
  and (_34405_, _07900_, \oc8051_golden_model_1.ACC [5]);
  or (_34406_, _34405_, _34400_);
  and (_34407_, _34406_, _07141_);
  and (_34408_, _07142_, \oc8051_golden_model_1.IE [5]);
  or (_34409_, _34408_, _06341_);
  or (_34410_, _34409_, _34407_);
  and (_34411_, _34410_, _06273_);
  and (_34413_, _34411_, _34404_);
  and (_34414_, _13601_, \oc8051_golden_model_1.IE [5]);
  and (_34415_, _15372_, _08626_);
  or (_34416_, _34415_, _34414_);
  and (_34417_, _34416_, _06272_);
  or (_34418_, _34417_, _06461_);
  or (_34419_, _34418_, _34413_);
  nor (_34420_, _08244_, _13593_);
  or (_34421_, _34420_, _34400_);
  or (_34422_, _34421_, _07166_);
  and (_34424_, _34422_, _34419_);
  or (_34425_, _34424_, _06464_);
  or (_34426_, _34406_, _06465_);
  and (_34427_, _34426_, _06269_);
  and (_34428_, _34427_, _34425_);
  and (_34429_, _15355_, _08626_);
  or (_34430_, _34429_, _34414_);
  and (_34431_, _34430_, _06268_);
  or (_34432_, _34431_, _06261_);
  or (_34433_, _34432_, _34428_);
  or (_34435_, _34414_, _15387_);
  and (_34436_, _34435_, _34416_);
  or (_34437_, _34436_, _06262_);
  and (_34438_, _34437_, _06258_);
  and (_34439_, _34438_, _34433_);
  or (_34440_, _34414_, _15403_);
  and (_34441_, _34440_, _06257_);
  and (_34442_, _34441_, _34416_);
  or (_34443_, _34442_, _10080_);
  or (_34444_, _34443_, _34439_);
  or (_34446_, _34421_, _07215_);
  and (_34447_, _34446_, _34444_);
  or (_34448_, _34447_, _07460_);
  and (_34449_, _09447_, _07900_);
  or (_34450_, _34400_, _07208_);
  or (_34451_, _34450_, _34449_);
  and (_34452_, _34451_, _05982_);
  and (_34453_, _34452_, _34448_);
  and (_34454_, _15459_, _07900_);
  or (_34455_, _34454_, _34400_);
  and (_34457_, _34455_, _10094_);
  or (_34458_, _34457_, _06218_);
  or (_34459_, _34458_, _34453_);
  and (_34460_, _08946_, _07900_);
  or (_34461_, _34460_, _34400_);
  or (_34462_, _34461_, _06219_);
  and (_34463_, _34462_, _34459_);
  or (_34464_, _34463_, _06369_);
  and (_34465_, _15353_, _07900_);
  or (_34466_, _34465_, _34400_);
  or (_34468_, _34466_, _07237_);
  and (_34469_, _34468_, _07240_);
  and (_34470_, _34469_, _34464_);
  and (_34471_, _11250_, _07900_);
  or (_34472_, _34471_, _34400_);
  and (_34473_, _34472_, _06536_);
  or (_34474_, _34473_, _34470_);
  and (_34475_, _34474_, _07242_);
  or (_34476_, _34400_, _08247_);
  and (_34477_, _34461_, _06375_);
  and (_34479_, _34477_, _34476_);
  or (_34480_, _34479_, _34475_);
  and (_34481_, _34480_, _07234_);
  and (_34482_, _34406_, _06545_);
  and (_34483_, _34482_, _34476_);
  or (_34484_, _34483_, _06366_);
  or (_34485_, _34484_, _34481_);
  and (_34486_, _15350_, _07900_);
  or (_34487_, _34400_, _09056_);
  or (_34488_, _34487_, _34486_);
  and (_34490_, _34488_, _09061_);
  and (_34491_, _34490_, _34485_);
  nor (_34492_, _11249_, _13593_);
  or (_34493_, _34492_, _34400_);
  and (_34494_, _34493_, _06528_);
  or (_34495_, _34494_, _06568_);
  or (_34496_, _34495_, _34491_);
  or (_34497_, _34403_, _06926_);
  and (_34498_, _34497_, _05928_);
  and (_34499_, _34498_, _34496_);
  and (_34501_, _34430_, _05927_);
  or (_34502_, _34501_, _06278_);
  or (_34503_, _34502_, _34499_);
  and (_34504_, _15532_, _07900_);
  or (_34505_, _34400_, _06279_);
  or (_34506_, _34505_, _34504_);
  and (_34507_, _34506_, _01347_);
  and (_34508_, _34507_, _34503_);
  or (_34509_, _34508_, _34399_);
  and (_43310_, _34509_, _42618_);
  and (_34511_, _01351_, \oc8051_golden_model_1.IE [6]);
  and (_34512_, _13593_, \oc8051_golden_model_1.IE [6]);
  and (_34513_, _15554_, _07900_);
  or (_34514_, _34513_, _34512_);
  or (_34515_, _34514_, _07151_);
  and (_34516_, _07900_, \oc8051_golden_model_1.ACC [6]);
  or (_34517_, _34516_, _34512_);
  and (_34518_, _34517_, _07141_);
  and (_34519_, _07142_, \oc8051_golden_model_1.IE [6]);
  or (_34520_, _34519_, _06341_);
  or (_34522_, _34520_, _34518_);
  and (_34523_, _34522_, _06273_);
  and (_34524_, _34523_, _34515_);
  and (_34525_, _13601_, \oc8051_golden_model_1.IE [6]);
  and (_34526_, _15570_, _08626_);
  or (_34527_, _34526_, _34525_);
  and (_34528_, _34527_, _06272_);
  or (_34529_, _34528_, _06461_);
  or (_34530_, _34529_, _34524_);
  nor (_34531_, _08142_, _13593_);
  or (_34533_, _34531_, _34512_);
  or (_34534_, _34533_, _07166_);
  and (_34535_, _34534_, _34530_);
  or (_34536_, _34535_, _06464_);
  or (_34537_, _34517_, _06465_);
  and (_34538_, _34537_, _06269_);
  and (_34539_, _34538_, _34536_);
  and (_34540_, _15551_, _08626_);
  or (_34541_, _34540_, _34525_);
  and (_34542_, _34541_, _06268_);
  or (_34544_, _34542_, _06261_);
  or (_34545_, _34544_, _34539_);
  or (_34546_, _34525_, _15585_);
  and (_34547_, _34546_, _34527_);
  or (_34548_, _34547_, _06262_);
  and (_34549_, _34548_, _06258_);
  and (_34550_, _34549_, _34545_);
  and (_34551_, _15602_, _08626_);
  or (_34552_, _34551_, _34525_);
  and (_34553_, _34552_, _06257_);
  or (_34555_, _34553_, _10080_);
  or (_34556_, _34555_, _34550_);
  or (_34557_, _34533_, _07215_);
  and (_34558_, _34557_, _34556_);
  or (_34559_, _34558_, _07460_);
  and (_34560_, _09446_, _07900_);
  or (_34561_, _34512_, _07208_);
  or (_34562_, _34561_, _34560_);
  and (_34563_, _34562_, _05982_);
  and (_34564_, _34563_, _34559_);
  and (_34566_, _15657_, _07900_);
  or (_34567_, _34566_, _34512_);
  and (_34568_, _34567_, _10094_);
  or (_34569_, _34568_, _06218_);
  or (_34570_, _34569_, _34564_);
  and (_34571_, _15664_, _07900_);
  or (_34572_, _34571_, _34512_);
  or (_34573_, _34572_, _06219_);
  and (_34574_, _34573_, _34570_);
  or (_34575_, _34574_, _06369_);
  and (_34577_, _15549_, _07900_);
  or (_34578_, _34577_, _34512_);
  or (_34579_, _34578_, _07237_);
  and (_34580_, _34579_, _07240_);
  and (_34581_, _34580_, _34575_);
  and (_34582_, _11247_, _07900_);
  or (_34583_, _34582_, _34512_);
  and (_34584_, _34583_, _06536_);
  or (_34585_, _34584_, _34581_);
  and (_34586_, _34585_, _07242_);
  or (_34588_, _34512_, _08145_);
  and (_34589_, _34572_, _06375_);
  and (_34590_, _34589_, _34588_);
  or (_34591_, _34590_, _34586_);
  and (_34592_, _34591_, _07234_);
  and (_34593_, _34517_, _06545_);
  and (_34594_, _34593_, _34588_);
  or (_34595_, _34594_, _06366_);
  or (_34596_, _34595_, _34592_);
  and (_34597_, _15546_, _07900_);
  or (_34599_, _34512_, _09056_);
  or (_34600_, _34599_, _34597_);
  and (_34601_, _34600_, _09061_);
  and (_34602_, _34601_, _34596_);
  nor (_34603_, _11246_, _13593_);
  or (_34604_, _34603_, _34512_);
  and (_34605_, _34604_, _06528_);
  or (_34606_, _34605_, _06568_);
  or (_34607_, _34606_, _34602_);
  or (_34608_, _34514_, _06926_);
  and (_34610_, _34608_, _05928_);
  and (_34611_, _34610_, _34607_);
  and (_34612_, _34541_, _05927_);
  or (_34613_, _34612_, _06278_);
  or (_34614_, _34613_, _34611_);
  and (_34615_, _15734_, _07900_);
  or (_34616_, _34512_, _06279_);
  or (_34617_, _34616_, _34615_);
  and (_34618_, _34617_, _01347_);
  and (_34619_, _34618_, _34614_);
  or (_34621_, _34619_, _34511_);
  and (_43311_, _34621_, _42618_);
  not (_34622_, \oc8051_golden_model_1.SCON [0]);
  nor (_34623_, _01347_, _34622_);
  nand (_34624_, _11263_, _07973_);
  nor (_34625_, _07973_, _34622_);
  nor (_34626_, _34625_, _07234_);
  nand (_34627_, _34626_, _34624_);
  and (_34628_, _07973_, _07133_);
  or (_34629_, _34628_, _34625_);
  or (_34631_, _34629_, _07215_);
  nor (_34632_, _08390_, _13705_);
  or (_34633_, _34632_, _34625_);
  or (_34634_, _34633_, _07151_);
  and (_34635_, _07973_, \oc8051_golden_model_1.ACC [0]);
  or (_34636_, _34635_, _34625_);
  and (_34637_, _34636_, _07141_);
  nor (_34638_, _07141_, _34622_);
  or (_34639_, _34638_, _06341_);
  or (_34640_, _34639_, _34637_);
  and (_34642_, _34640_, _06273_);
  and (_34643_, _34642_, _34634_);
  nor (_34644_, _08622_, _34622_);
  and (_34645_, _14382_, _08622_);
  or (_34646_, _34645_, _34644_);
  and (_34647_, _34646_, _06272_);
  or (_34648_, _34647_, _34643_);
  and (_34649_, _34648_, _07166_);
  and (_34650_, _34629_, _06461_);
  or (_34651_, _34650_, _06464_);
  or (_34653_, _34651_, _34649_);
  or (_34654_, _34636_, _06465_);
  and (_34655_, _34654_, _06269_);
  and (_34656_, _34655_, _34653_);
  and (_34657_, _34625_, _06268_);
  or (_34658_, _34657_, _06261_);
  or (_34659_, _34658_, _34656_);
  or (_34660_, _34633_, _06262_);
  and (_34661_, _34660_, _06258_);
  and (_34662_, _34661_, _34659_);
  and (_34664_, _14413_, _08622_);
  or (_34665_, _34664_, _34644_);
  and (_34666_, _34665_, _06257_);
  or (_34667_, _34666_, _10080_);
  or (_34668_, _34667_, _34662_);
  and (_34669_, _34668_, _34631_);
  or (_34670_, _34669_, _07460_);
  and (_34671_, _09392_, _07973_);
  or (_34672_, _34625_, _07208_);
  or (_34673_, _34672_, _34671_);
  and (_34675_, _34673_, _34670_);
  or (_34676_, _34675_, _10094_);
  and (_34677_, _14467_, _07973_);
  or (_34678_, _34625_, _05982_);
  or (_34679_, _34678_, _34677_);
  and (_34680_, _34679_, _06219_);
  and (_34681_, _34680_, _34676_);
  and (_34682_, _07973_, _08954_);
  or (_34683_, _34682_, _34625_);
  and (_34684_, _34683_, _06218_);
  or (_34686_, _34684_, _06369_);
  or (_34687_, _34686_, _34681_);
  and (_34688_, _14366_, _07973_);
  or (_34689_, _34688_, _34625_);
  or (_34690_, _34689_, _07237_);
  and (_34691_, _34690_, _07240_);
  and (_34692_, _34691_, _34687_);
  nor (_34693_, _12580_, _13705_);
  or (_34694_, _34693_, _34625_);
  and (_34695_, _34624_, _06536_);
  and (_34696_, _34695_, _34694_);
  or (_34697_, _34696_, _34692_);
  and (_34698_, _34697_, _07242_);
  nand (_34699_, _34683_, _06375_);
  nor (_34700_, _34699_, _34632_);
  or (_34701_, _34700_, _06545_);
  or (_34702_, _34701_, _34698_);
  and (_34703_, _34702_, _34627_);
  or (_34704_, _34703_, _06366_);
  and (_34705_, _14363_, _07973_);
  or (_34707_, _34625_, _09056_);
  or (_34708_, _34707_, _34705_);
  and (_34709_, _34708_, _09061_);
  and (_34710_, _34709_, _34704_);
  and (_34711_, _34694_, _06528_);
  or (_34712_, _34711_, _06568_);
  or (_34713_, _34712_, _34710_);
  or (_34714_, _34633_, _06926_);
  and (_34715_, _34714_, _34713_);
  or (_34716_, _34715_, _05927_);
  or (_34718_, _34625_, _05928_);
  and (_34719_, _34718_, _34716_);
  or (_34720_, _34719_, _06278_);
  or (_34721_, _34633_, _06279_);
  and (_34722_, _34721_, _01347_);
  and (_34723_, _34722_, _34720_);
  or (_34724_, _34723_, _34623_);
  and (_43313_, _34724_, _42618_);
  not (_34725_, \oc8051_golden_model_1.SCON [1]);
  nor (_34726_, _01347_, _34725_);
  nor (_34728_, _07973_, _34725_);
  nor (_34729_, _11261_, _13705_);
  or (_34730_, _34729_, _34728_);
  or (_34731_, _34730_, _09061_);
  nand (_34732_, _07973_, _07038_);
  or (_34733_, _07973_, \oc8051_golden_model_1.SCON [1]);
  and (_34734_, _34733_, _06218_);
  and (_34735_, _34734_, _34732_);
  nor (_34736_, _13705_, _07357_);
  or (_34737_, _34736_, _34728_);
  or (_34739_, _34737_, _07166_);
  and (_34740_, _14562_, _07973_);
  not (_34741_, _34740_);
  and (_34742_, _34741_, _34733_);
  or (_34743_, _34742_, _07151_);
  and (_34744_, _07973_, \oc8051_golden_model_1.ACC [1]);
  or (_34745_, _34744_, _34728_);
  and (_34746_, _34745_, _07141_);
  nor (_34747_, _07141_, _34725_);
  or (_34748_, _34747_, _06341_);
  or (_34750_, _34748_, _34746_);
  and (_34751_, _34750_, _06273_);
  and (_34752_, _34751_, _34743_);
  nor (_34753_, _08622_, _34725_);
  and (_34754_, _14557_, _08622_);
  or (_34755_, _34754_, _34753_);
  and (_34756_, _34755_, _06272_);
  or (_34757_, _34756_, _06461_);
  or (_34758_, _34757_, _34752_);
  and (_34759_, _34758_, _34739_);
  or (_34761_, _34759_, _06464_);
  or (_34762_, _34745_, _06465_);
  and (_34763_, _34762_, _06269_);
  and (_34764_, _34763_, _34761_);
  and (_34765_, _14560_, _08622_);
  or (_34766_, _34765_, _34753_);
  and (_34767_, _34766_, _06268_);
  or (_34768_, _34767_, _06261_);
  or (_34769_, _34768_, _34764_);
  and (_34770_, _34754_, _14556_);
  or (_34772_, _34753_, _06262_);
  or (_34773_, _34772_, _34770_);
  and (_34774_, _34773_, _06258_);
  and (_34775_, _34774_, _34769_);
  or (_34776_, _34753_, _14597_);
  and (_34777_, _34776_, _06257_);
  and (_34778_, _34777_, _34755_);
  or (_34779_, _34778_, _10080_);
  or (_34780_, _34779_, _34775_);
  or (_34781_, _34737_, _07215_);
  and (_34783_, _34781_, _34780_);
  or (_34784_, _34783_, _07460_);
  and (_34785_, _09451_, _07973_);
  or (_34786_, _34728_, _07208_);
  or (_34787_, _34786_, _34785_);
  and (_34788_, _34787_, _05982_);
  and (_34789_, _34788_, _34784_);
  and (_34790_, _14653_, _07973_);
  or (_34791_, _34790_, _34728_);
  and (_34792_, _34791_, _10094_);
  or (_34794_, _34792_, _34789_);
  and (_34795_, _34794_, _06219_);
  or (_34796_, _34795_, _34735_);
  and (_34797_, _34796_, _07237_);
  or (_34798_, _14668_, _13705_);
  and (_34799_, _34733_, _06369_);
  and (_34800_, _34799_, _34798_);
  or (_34801_, _34800_, _06536_);
  or (_34802_, _34801_, _34797_);
  nand (_34803_, _11260_, _07973_);
  and (_34805_, _34803_, _34730_);
  or (_34806_, _34805_, _07240_);
  and (_34807_, _34806_, _07242_);
  and (_34808_, _34807_, _34802_);
  or (_34809_, _14666_, _13705_);
  and (_34810_, _34733_, _06375_);
  and (_34811_, _34810_, _34809_);
  or (_34812_, _34811_, _06545_);
  or (_34813_, _34812_, _34808_);
  nor (_34814_, _34728_, _07234_);
  nand (_34816_, _34814_, _34803_);
  and (_34817_, _34816_, _09056_);
  and (_34818_, _34817_, _34813_);
  or (_34819_, _34732_, _08341_);
  and (_34820_, _34733_, _06366_);
  and (_34821_, _34820_, _34819_);
  or (_34822_, _34821_, _06528_);
  or (_34823_, _34822_, _34818_);
  and (_34824_, _34823_, _34731_);
  or (_34825_, _34824_, _06568_);
  or (_34827_, _34742_, _06926_);
  and (_34828_, _34827_, _05928_);
  and (_34829_, _34828_, _34825_);
  and (_34830_, _34766_, _05927_);
  or (_34831_, _34830_, _06278_);
  or (_34832_, _34831_, _34829_);
  or (_34833_, _34728_, _06279_);
  or (_34834_, _34833_, _34740_);
  and (_34835_, _34834_, _01347_);
  and (_34836_, _34835_, _34832_);
  or (_34838_, _34836_, _34726_);
  and (_43314_, _34838_, _42618_);
  and (_34839_, _01351_, \oc8051_golden_model_1.SCON [2]);
  and (_34840_, _13705_, \oc8051_golden_model_1.SCON [2]);
  nor (_34841_, _13705_, _07776_);
  or (_34842_, _34841_, _34840_);
  or (_34843_, _34842_, _07215_);
  and (_34844_, _34842_, _06461_);
  and (_34845_, _13714_, \oc8051_golden_model_1.SCON [2]);
  and (_34846_, _14774_, _08622_);
  or (_34848_, _34846_, _34845_);
  or (_34849_, _34848_, _06273_);
  and (_34850_, _14770_, _07973_);
  or (_34851_, _34850_, _34840_);
  and (_34852_, _34851_, _06341_);
  and (_34853_, _07142_, \oc8051_golden_model_1.SCON [2]);
  and (_34854_, _07973_, \oc8051_golden_model_1.ACC [2]);
  or (_34855_, _34854_, _34840_);
  and (_34856_, _34855_, _07141_);
  or (_34857_, _34856_, _34853_);
  and (_34859_, _34857_, _07151_);
  or (_34860_, _34859_, _06272_);
  or (_34861_, _34860_, _34852_);
  and (_34862_, _34861_, _34849_);
  and (_34863_, _34862_, _07166_);
  or (_34864_, _34863_, _34844_);
  or (_34865_, _34864_, _06464_);
  or (_34866_, _34855_, _06465_);
  and (_34867_, _34866_, _06269_);
  and (_34868_, _34867_, _34865_);
  and (_34870_, _14756_, _08622_);
  or (_34871_, _34870_, _34845_);
  and (_34872_, _34871_, _06268_);
  or (_34873_, _34872_, _06261_);
  or (_34874_, _34873_, _34868_);
  or (_34875_, _34845_, _14789_);
  and (_34876_, _34875_, _34848_);
  or (_34877_, _34876_, _06262_);
  and (_34878_, _34877_, _06258_);
  and (_34879_, _34878_, _34874_);
  and (_34881_, _14804_, _08622_);
  or (_34882_, _34881_, _34845_);
  and (_34883_, _34882_, _06257_);
  or (_34884_, _34883_, _10080_);
  or (_34885_, _34884_, _34879_);
  and (_34886_, _34885_, _34843_);
  or (_34887_, _34886_, _07460_);
  and (_34888_, _09450_, _07973_);
  or (_34889_, _34840_, _07208_);
  or (_34890_, _34889_, _34888_);
  and (_34892_, _34890_, _05982_);
  and (_34893_, _34892_, _34887_);
  and (_34894_, _14859_, _07973_);
  or (_34895_, _34894_, _34840_);
  and (_34896_, _34895_, _10094_);
  or (_34897_, _34896_, _06218_);
  or (_34898_, _34897_, _34893_);
  and (_34899_, _07973_, _08973_);
  or (_34900_, _34899_, _34840_);
  or (_34901_, _34900_, _06219_);
  and (_34903_, _34901_, _34898_);
  or (_34904_, _34903_, _06369_);
  and (_34905_, _14751_, _07973_);
  or (_34906_, _34905_, _34840_);
  or (_34907_, _34906_, _07237_);
  and (_34908_, _34907_, _07240_);
  and (_34909_, _34908_, _34904_);
  and (_34910_, _11259_, _07973_);
  or (_34911_, _34910_, _34840_);
  and (_34912_, _34911_, _06536_);
  or (_34914_, _34912_, _34909_);
  and (_34915_, _34914_, _07242_);
  or (_34916_, _34840_, _08440_);
  and (_34917_, _34900_, _06375_);
  and (_34918_, _34917_, _34916_);
  or (_34919_, _34918_, _34915_);
  and (_34920_, _34919_, _07234_);
  and (_34921_, _34855_, _06545_);
  and (_34922_, _34921_, _34916_);
  or (_34923_, _34922_, _06366_);
  or (_34925_, _34923_, _34920_);
  and (_34926_, _14748_, _07973_);
  or (_34927_, _34840_, _09056_);
  or (_34928_, _34927_, _34926_);
  and (_34929_, _34928_, _09061_);
  and (_34930_, _34929_, _34925_);
  nor (_34931_, _11258_, _13705_);
  or (_34932_, _34931_, _34840_);
  and (_34933_, _34932_, _06528_);
  or (_34934_, _34933_, _06568_);
  or (_34936_, _34934_, _34930_);
  or (_34937_, _34851_, _06926_);
  and (_34938_, _34937_, _05928_);
  and (_34939_, _34938_, _34936_);
  and (_34940_, _34871_, _05927_);
  or (_34941_, _34940_, _06278_);
  or (_34942_, _34941_, _34939_);
  and (_34943_, _14926_, _07973_);
  or (_34944_, _34840_, _06279_);
  or (_34945_, _34944_, _34943_);
  and (_34947_, _34945_, _01347_);
  and (_34948_, _34947_, _34942_);
  or (_34949_, _34948_, _34839_);
  and (_43315_, _34949_, _42618_);
  and (_34950_, _01351_, \oc8051_golden_model_1.SCON [3]);
  and (_34951_, _13705_, \oc8051_golden_model_1.SCON [3]);
  nor (_34952_, _13705_, _07594_);
  or (_34953_, _34952_, _34951_);
  or (_34954_, _34953_, _07215_);
  and (_34955_, _14953_, _07973_);
  or (_34957_, _34955_, _34951_);
  or (_34958_, _34957_, _07151_);
  and (_34959_, _07973_, \oc8051_golden_model_1.ACC [3]);
  or (_34960_, _34959_, _34951_);
  and (_34961_, _34960_, _07141_);
  and (_34962_, _07142_, \oc8051_golden_model_1.SCON [3]);
  or (_34963_, _34962_, _06341_);
  or (_34964_, _34963_, _34961_);
  and (_34965_, _34964_, _06273_);
  and (_34966_, _34965_, _34958_);
  and (_34968_, _13714_, \oc8051_golden_model_1.SCON [3]);
  and (_34969_, _14950_, _08622_);
  or (_34970_, _34969_, _34968_);
  and (_34971_, _34970_, _06272_);
  or (_34972_, _34971_, _06461_);
  or (_34973_, _34972_, _34966_);
  or (_34974_, _34953_, _07166_);
  and (_34975_, _34974_, _34973_);
  or (_34976_, _34975_, _06464_);
  or (_34977_, _34960_, _06465_);
  and (_34979_, _34977_, _06269_);
  and (_34980_, _34979_, _34976_);
  and (_34981_, _14948_, _08622_);
  or (_34982_, _34981_, _34968_);
  and (_34983_, _34982_, _06268_);
  or (_34984_, _34983_, _06261_);
  or (_34985_, _34984_, _34980_);
  or (_34986_, _34968_, _14979_);
  and (_34987_, _34986_, _34970_);
  or (_34988_, _34987_, _06262_);
  and (_34990_, _34988_, _06258_);
  and (_34991_, _34990_, _34985_);
  or (_34992_, _34968_, _14992_);
  and (_34993_, _34992_, _06257_);
  and (_34994_, _34993_, _34970_);
  or (_34995_, _34994_, _10080_);
  or (_34996_, _34995_, _34991_);
  and (_34997_, _34996_, _34954_);
  or (_34998_, _34997_, _07460_);
  and (_34999_, _09449_, _07973_);
  or (_35001_, _34951_, _07208_);
  or (_35002_, _35001_, _34999_);
  and (_35003_, _35002_, _05982_);
  and (_35004_, _35003_, _34998_);
  and (_35005_, _15048_, _07973_);
  or (_35006_, _35005_, _34951_);
  and (_35007_, _35006_, _10094_);
  or (_35008_, _35007_, _06218_);
  or (_35009_, _35008_, _35004_);
  and (_35010_, _07973_, _08930_);
  or (_35012_, _35010_, _34951_);
  or (_35013_, _35012_, _06219_);
  and (_35014_, _35013_, _35009_);
  or (_35015_, _35014_, _06369_);
  and (_35016_, _14943_, _07973_);
  or (_35017_, _35016_, _34951_);
  or (_35018_, _35017_, _07237_);
  and (_35019_, _35018_, _07240_);
  and (_35020_, _35019_, _35015_);
  and (_35021_, _12577_, _07973_);
  or (_35023_, _35021_, _34951_);
  and (_35024_, _35023_, _06536_);
  or (_35025_, _35024_, _35020_);
  and (_35026_, _35025_, _07242_);
  or (_35027_, _34951_, _08292_);
  and (_35028_, _35012_, _06375_);
  and (_35029_, _35028_, _35027_);
  or (_35030_, _35029_, _35026_);
  and (_35031_, _35030_, _07234_);
  and (_35032_, _34960_, _06545_);
  and (_35034_, _35032_, _35027_);
  or (_35035_, _35034_, _06366_);
  or (_35036_, _35035_, _35031_);
  and (_35037_, _14940_, _07973_);
  or (_35038_, _34951_, _09056_);
  or (_35039_, _35038_, _35037_);
  and (_35040_, _35039_, _09061_);
  and (_35041_, _35040_, _35036_);
  nor (_35042_, _11256_, _13705_);
  or (_35043_, _35042_, _34951_);
  and (_35045_, _35043_, _06528_);
  or (_35046_, _35045_, _06568_);
  or (_35047_, _35046_, _35041_);
  or (_35048_, _34957_, _06926_);
  and (_35049_, _35048_, _05928_);
  and (_35050_, _35049_, _35047_);
  and (_35051_, _34982_, _05927_);
  or (_35052_, _35051_, _06278_);
  or (_35053_, _35052_, _35050_);
  and (_35054_, _15128_, _07973_);
  or (_35056_, _34951_, _06279_);
  or (_35057_, _35056_, _35054_);
  and (_35058_, _35057_, _01347_);
  and (_35059_, _35058_, _35053_);
  or (_35060_, _35059_, _34950_);
  and (_43316_, _35060_, _42618_);
  and (_35061_, _01351_, \oc8051_golden_model_1.SCON [4]);
  and (_35062_, _13705_, \oc8051_golden_model_1.SCON [4]);
  nor (_35063_, _08541_, _13705_);
  or (_35064_, _35063_, _35062_);
  or (_35066_, _35064_, _07215_);
  and (_35067_, _13714_, \oc8051_golden_model_1.SCON [4]);
  and (_35068_, _15176_, _08622_);
  or (_35069_, _35068_, _35067_);
  and (_35070_, _35069_, _06268_);
  and (_35071_, _15162_, _07973_);
  or (_35072_, _35071_, _35062_);
  or (_35073_, _35072_, _07151_);
  and (_35074_, _07973_, \oc8051_golden_model_1.ACC [4]);
  or (_35075_, _35074_, _35062_);
  and (_35077_, _35075_, _07141_);
  and (_35078_, _07142_, \oc8051_golden_model_1.SCON [4]);
  or (_35079_, _35078_, _06341_);
  or (_35080_, _35079_, _35077_);
  and (_35081_, _35080_, _06273_);
  and (_35082_, _35081_, _35073_);
  and (_35083_, _15166_, _08622_);
  or (_35084_, _35083_, _35067_);
  and (_35085_, _35084_, _06272_);
  or (_35086_, _35085_, _06461_);
  or (_35088_, _35086_, _35082_);
  or (_35089_, _35064_, _07166_);
  and (_35090_, _35089_, _35088_);
  or (_35091_, _35090_, _06464_);
  or (_35092_, _35075_, _06465_);
  and (_35093_, _35092_, _06269_);
  and (_35094_, _35093_, _35091_);
  or (_35095_, _35094_, _35070_);
  and (_35096_, _35095_, _06262_);
  or (_35097_, _35067_, _15183_);
  and (_35099_, _35097_, _06261_);
  and (_35100_, _35099_, _35084_);
  or (_35101_, _35100_, _35096_);
  and (_35102_, _35101_, _06258_);
  and (_35103_, _15200_, _08622_);
  or (_35104_, _35103_, _35067_);
  and (_35105_, _35104_, _06257_);
  or (_35106_, _35105_, _10080_);
  or (_35107_, _35106_, _35102_);
  and (_35108_, _35107_, _35066_);
  or (_35110_, _35108_, _07460_);
  and (_35111_, _09448_, _07973_);
  or (_35112_, _35062_, _07208_);
  or (_35113_, _35112_, _35111_);
  and (_35114_, _35113_, _05982_);
  and (_35115_, _35114_, _35110_);
  and (_35116_, _15254_, _07973_);
  or (_35117_, _35116_, _35062_);
  and (_35118_, _35117_, _10094_);
  or (_35119_, _35118_, _06218_);
  or (_35121_, _35119_, _35115_);
  and (_35122_, _08959_, _07973_);
  or (_35123_, _35122_, _35062_);
  or (_35124_, _35123_, _06219_);
  and (_35125_, _35124_, _35121_);
  or (_35126_, _35125_, _06369_);
  and (_35127_, _15269_, _07973_);
  or (_35128_, _35127_, _35062_);
  or (_35129_, _35128_, _07237_);
  and (_35130_, _35129_, _07240_);
  and (_35132_, _35130_, _35126_);
  and (_35133_, _11254_, _07973_);
  or (_35134_, _35133_, _35062_);
  and (_35135_, _35134_, _06536_);
  or (_35136_, _35135_, _35132_);
  and (_35137_, _35136_, _07242_);
  or (_35138_, _35062_, _08544_);
  and (_35139_, _35123_, _06375_);
  and (_35140_, _35139_, _35138_);
  or (_35141_, _35140_, _35137_);
  and (_35143_, _35141_, _07234_);
  and (_35144_, _35075_, _06545_);
  and (_35145_, _35144_, _35138_);
  or (_35146_, _35145_, _06366_);
  or (_35147_, _35146_, _35143_);
  and (_35148_, _15266_, _07973_);
  or (_35149_, _35062_, _09056_);
  or (_35150_, _35149_, _35148_);
  and (_35151_, _35150_, _09061_);
  and (_35152_, _35151_, _35147_);
  nor (_35154_, _11253_, _13705_);
  or (_35155_, _35154_, _35062_);
  and (_35156_, _35155_, _06528_);
  or (_35157_, _35156_, _06568_);
  or (_35158_, _35157_, _35152_);
  or (_35159_, _35072_, _06926_);
  and (_35160_, _35159_, _05928_);
  and (_35161_, _35160_, _35158_);
  and (_35162_, _35069_, _05927_);
  or (_35163_, _35162_, _06278_);
  or (_35165_, _35163_, _35161_);
  and (_35166_, _15329_, _07973_);
  or (_35167_, _35062_, _06279_);
  or (_35168_, _35167_, _35166_);
  and (_35169_, _35168_, _01347_);
  and (_35170_, _35169_, _35165_);
  or (_35171_, _35170_, _35061_);
  and (_43317_, _35171_, _42618_);
  and (_35172_, _01351_, \oc8051_golden_model_1.SCON [5]);
  and (_35173_, _13705_, \oc8051_golden_model_1.SCON [5]);
  and (_35175_, _15358_, _07973_);
  or (_35176_, _35175_, _35173_);
  or (_35177_, _35176_, _07151_);
  and (_35178_, _07973_, \oc8051_golden_model_1.ACC [5]);
  or (_35179_, _35178_, _35173_);
  and (_35180_, _35179_, _07141_);
  and (_35181_, _07142_, \oc8051_golden_model_1.SCON [5]);
  or (_35182_, _35181_, _06341_);
  or (_35183_, _35182_, _35180_);
  and (_35184_, _35183_, _06273_);
  and (_35186_, _35184_, _35177_);
  and (_35187_, _13714_, \oc8051_golden_model_1.SCON [5]);
  and (_35188_, _15372_, _08622_);
  or (_35189_, _35188_, _35187_);
  and (_35190_, _35189_, _06272_);
  or (_35191_, _35190_, _06461_);
  or (_35192_, _35191_, _35186_);
  nor (_35193_, _08244_, _13705_);
  or (_35194_, _35193_, _35173_);
  or (_35195_, _35194_, _07166_);
  and (_35197_, _35195_, _35192_);
  or (_35198_, _35197_, _06464_);
  or (_35199_, _35179_, _06465_);
  and (_35200_, _35199_, _06269_);
  and (_35201_, _35200_, _35198_);
  and (_35202_, _15355_, _08622_);
  or (_35203_, _35202_, _35187_);
  and (_35204_, _35203_, _06268_);
  or (_35205_, _35204_, _06261_);
  or (_35206_, _35205_, _35201_);
  or (_35208_, _35187_, _15387_);
  and (_35209_, _35208_, _35189_);
  or (_35210_, _35209_, _06262_);
  and (_35211_, _35210_, _06258_);
  and (_35212_, _35211_, _35206_);
  or (_35213_, _35187_, _15403_);
  and (_35214_, _35213_, _06257_);
  and (_35215_, _35214_, _35189_);
  or (_35216_, _35215_, _10080_);
  or (_35217_, _35216_, _35212_);
  or (_35219_, _35194_, _07215_);
  and (_35220_, _35219_, _35217_);
  or (_35221_, _35220_, _07460_);
  and (_35222_, _09447_, _07973_);
  or (_35223_, _35173_, _07208_);
  or (_35224_, _35223_, _35222_);
  and (_35225_, _35224_, _05982_);
  and (_35226_, _35225_, _35221_);
  and (_35227_, _15459_, _07973_);
  or (_35228_, _35227_, _35173_);
  and (_35230_, _35228_, _10094_);
  or (_35231_, _35230_, _06218_);
  or (_35232_, _35231_, _35226_);
  and (_35233_, _08946_, _07973_);
  or (_35234_, _35233_, _35173_);
  or (_35235_, _35234_, _06219_);
  and (_35236_, _35235_, _35232_);
  or (_35237_, _35236_, _06369_);
  and (_35238_, _15353_, _07973_);
  or (_35239_, _35238_, _35173_);
  or (_35241_, _35239_, _07237_);
  and (_35242_, _35241_, _07240_);
  and (_35243_, _35242_, _35237_);
  and (_35244_, _11250_, _07973_);
  or (_35245_, _35244_, _35173_);
  and (_35246_, _35245_, _06536_);
  or (_35247_, _35246_, _35243_);
  and (_35248_, _35247_, _07242_);
  or (_35249_, _35173_, _08247_);
  and (_35250_, _35234_, _06375_);
  and (_35252_, _35250_, _35249_);
  or (_35253_, _35252_, _35248_);
  and (_35254_, _35253_, _07234_);
  and (_35255_, _35179_, _06545_);
  and (_35256_, _35255_, _35249_);
  or (_35257_, _35256_, _06366_);
  or (_35258_, _35257_, _35254_);
  and (_35259_, _15350_, _07973_);
  or (_35260_, _35173_, _09056_);
  or (_35261_, _35260_, _35259_);
  and (_35263_, _35261_, _09061_);
  and (_35264_, _35263_, _35258_);
  nor (_35265_, _11249_, _13705_);
  or (_35266_, _35265_, _35173_);
  and (_35267_, _35266_, _06528_);
  or (_35268_, _35267_, _06568_);
  or (_35269_, _35268_, _35264_);
  or (_35270_, _35176_, _06926_);
  and (_35271_, _35270_, _05928_);
  and (_35272_, _35271_, _35269_);
  and (_35274_, _35203_, _05927_);
  or (_35275_, _35274_, _06278_);
  or (_35276_, _35275_, _35272_);
  and (_35277_, _15532_, _07973_);
  or (_35278_, _35173_, _06279_);
  or (_35279_, _35278_, _35277_);
  and (_35280_, _35279_, _01347_);
  and (_35281_, _35280_, _35276_);
  or (_35282_, _35281_, _35172_);
  and (_43318_, _35282_, _42618_);
  and (_35284_, _01351_, \oc8051_golden_model_1.SCON [6]);
  and (_35285_, _13705_, \oc8051_golden_model_1.SCON [6]);
  and (_35286_, _15554_, _07973_);
  or (_35287_, _35286_, _35285_);
  or (_35288_, _35287_, _07151_);
  and (_35289_, _07973_, \oc8051_golden_model_1.ACC [6]);
  or (_35290_, _35289_, _35285_);
  and (_35291_, _35290_, _07141_);
  and (_35292_, _07142_, \oc8051_golden_model_1.SCON [6]);
  or (_35293_, _35292_, _06341_);
  or (_35295_, _35293_, _35291_);
  and (_35296_, _35295_, _06273_);
  and (_35297_, _35296_, _35288_);
  and (_35298_, _13714_, \oc8051_golden_model_1.SCON [6]);
  and (_35299_, _15570_, _08622_);
  or (_35300_, _35299_, _35298_);
  and (_35301_, _35300_, _06272_);
  or (_35302_, _35301_, _06461_);
  or (_35303_, _35302_, _35297_);
  nor (_35304_, _08142_, _13705_);
  or (_35306_, _35304_, _35285_);
  or (_35307_, _35306_, _07166_);
  and (_35308_, _35307_, _35303_);
  or (_35309_, _35308_, _06464_);
  or (_35310_, _35290_, _06465_);
  and (_35311_, _35310_, _06269_);
  and (_35312_, _35311_, _35309_);
  and (_35313_, _15551_, _08622_);
  or (_35314_, _35313_, _35298_);
  and (_35315_, _35314_, _06268_);
  or (_35317_, _35315_, _06261_);
  or (_35318_, _35317_, _35312_);
  or (_35319_, _35298_, _15585_);
  and (_35320_, _35319_, _35300_);
  or (_35321_, _35320_, _06262_);
  and (_35322_, _35321_, _06258_);
  and (_35323_, _35322_, _35318_);
  and (_35324_, _15602_, _08622_);
  or (_35325_, _35324_, _35298_);
  and (_35326_, _35325_, _06257_);
  or (_35328_, _35326_, _10080_);
  or (_35329_, _35328_, _35323_);
  or (_35330_, _35306_, _07215_);
  and (_35331_, _35330_, _35329_);
  or (_35332_, _35331_, _07460_);
  and (_35333_, _09446_, _07973_);
  or (_35334_, _35285_, _07208_);
  or (_35335_, _35334_, _35333_);
  and (_35336_, _35335_, _05982_);
  and (_35337_, _35336_, _35332_);
  and (_35339_, _15657_, _07973_);
  or (_35340_, _35339_, _35285_);
  and (_35341_, _35340_, _10094_);
  or (_35342_, _35341_, _06218_);
  or (_35343_, _35342_, _35337_);
  and (_35344_, _15664_, _07973_);
  or (_35345_, _35344_, _35285_);
  or (_35346_, _35345_, _06219_);
  and (_35347_, _35346_, _35343_);
  or (_35348_, _35347_, _06369_);
  and (_35350_, _15549_, _07973_);
  or (_35351_, _35350_, _35285_);
  or (_35352_, _35351_, _07237_);
  and (_35353_, _35352_, _07240_);
  and (_35354_, _35353_, _35348_);
  and (_35355_, _11247_, _07973_);
  or (_35356_, _35355_, _35285_);
  and (_35357_, _35356_, _06536_);
  or (_35358_, _35357_, _35354_);
  and (_35359_, _35358_, _07242_);
  or (_35361_, _35285_, _08145_);
  and (_35362_, _35345_, _06375_);
  and (_35363_, _35362_, _35361_);
  or (_35364_, _35363_, _35359_);
  and (_35365_, _35364_, _07234_);
  and (_35366_, _35290_, _06545_);
  and (_35367_, _35366_, _35361_);
  or (_35368_, _35367_, _06366_);
  or (_35369_, _35368_, _35365_);
  and (_35370_, _15546_, _07973_);
  or (_35372_, _35285_, _09056_);
  or (_35373_, _35372_, _35370_);
  and (_35374_, _35373_, _09061_);
  and (_35375_, _35374_, _35369_);
  nor (_35376_, _11246_, _13705_);
  or (_35377_, _35376_, _35285_);
  and (_35378_, _35377_, _06528_);
  or (_35379_, _35378_, _06568_);
  or (_35380_, _35379_, _35375_);
  or (_35381_, _35287_, _06926_);
  and (_35383_, _35381_, _05928_);
  and (_35384_, _35383_, _35380_);
  and (_35385_, _35314_, _05927_);
  or (_35386_, _35385_, _06278_);
  or (_35387_, _35386_, _35384_);
  and (_35388_, _15734_, _07973_);
  or (_35389_, _35285_, _06279_);
  or (_35390_, _35389_, _35388_);
  and (_35391_, _35390_, _01347_);
  and (_35392_, _35391_, _35387_);
  or (_35394_, _35392_, _35284_);
  and (_43319_, _35394_, _42618_);
  nor (_35395_, _01347_, _06800_);
  nor (_35396_, _07956_, _06800_);
  and (_35397_, _07956_, \oc8051_golden_model_1.ACC [0]);
  and (_35398_, _35397_, _08390_);
  or (_35399_, _35398_, _35396_);
  or (_35400_, _35399_, _07234_);
  nor (_35401_, _08390_, _13872_);
  or (_35402_, _35401_, _35396_);
  or (_35404_, _35402_, _07151_);
  or (_35405_, _35397_, _35396_);
  and (_35406_, _35405_, _07141_);
  nor (_35407_, _07141_, _06800_);
  or (_35408_, _35407_, _06341_);
  or (_35409_, _35408_, _35406_);
  and (_35410_, _35409_, _07166_);
  nand (_35411_, _35410_, _35404_);
  nand (_35412_, _35411_, _06802_);
  or (_35413_, _35405_, _06465_);
  and (_35415_, _35413_, _07303_);
  and (_35416_, _35415_, _35412_);
  nand (_35417_, _07215_, _07186_);
  or (_35418_, _35417_, _35416_);
  and (_35419_, _08173_, _07133_);
  or (_35420_, _35396_, _07215_);
  or (_35421_, _35420_, _35419_);
  and (_35422_, _35421_, _35418_);
  or (_35423_, _35422_, _07460_);
  or (_35424_, _35396_, _07208_);
  and (_35426_, _09392_, _07956_);
  or (_35427_, _35426_, _35424_);
  and (_35428_, _35427_, _35423_);
  or (_35429_, _35428_, _10094_);
  and (_35430_, _14467_, _08173_);
  or (_35431_, _35396_, _05982_);
  or (_35432_, _35431_, _35430_);
  and (_35433_, _35432_, _06219_);
  and (_35434_, _35433_, _35429_);
  and (_35435_, _07956_, _08954_);
  or (_35437_, _35435_, _35396_);
  and (_35438_, _35437_, _06218_);
  or (_35439_, _35438_, _06369_);
  or (_35440_, _35439_, _35434_);
  and (_35441_, _14366_, _07956_);
  or (_35442_, _35441_, _35396_);
  or (_35443_, _35442_, _07237_);
  and (_35444_, _35443_, _07240_);
  and (_35445_, _35444_, _35440_);
  nor (_35446_, _12580_, _13872_);
  or (_35448_, _35446_, _35396_);
  nor (_35449_, _35398_, _07240_);
  and (_35450_, _35449_, _35448_);
  or (_35451_, _35450_, _35445_);
  and (_35452_, _35451_, _07242_);
  nand (_35453_, _35437_, _06375_);
  nor (_35454_, _35453_, _35401_);
  or (_35455_, _35454_, _06545_);
  or (_35456_, _35455_, _35452_);
  and (_35457_, _35456_, _35400_);
  or (_35459_, _35457_, _06366_);
  and (_35460_, _14363_, _07956_);
  or (_35461_, _35460_, _35396_);
  or (_35462_, _35461_, _09056_);
  and (_35463_, _35462_, _09061_);
  and (_35464_, _35463_, _35459_);
  and (_35465_, _35448_, _06528_);
  or (_35466_, _35465_, _19502_);
  or (_35467_, _35466_, _35464_);
  or (_35468_, _35402_, _06661_);
  and (_35470_, _35468_, _01347_);
  and (_35471_, _35470_, _35467_);
  or (_35472_, _35471_, _35395_);
  and (_43321_, _35472_, _42618_);
  nand (_35473_, _08173_, _07038_);
  or (_35474_, _35473_, _08341_);
  or (_35475_, _07956_, \oc8051_golden_model_1.SP [1]);
  and (_35476_, _35475_, _06366_);
  and (_35477_, _35476_, _35474_);
  and (_35478_, _11260_, _08173_);
  nor (_35479_, _07956_, _07067_);
  or (_35480_, _35479_, _07234_);
  or (_35481_, _35480_, _35478_);
  and (_35482_, _14562_, _08173_);
  not (_35483_, _35482_);
  and (_35484_, _35483_, _35475_);
  or (_35485_, _35484_, _07151_);
  nand (_35486_, _06758_, \oc8051_golden_model_1.SP [1]);
  and (_35487_, _07956_, \oc8051_golden_model_1.ACC [1]);
  or (_35488_, _35487_, _35479_);
  and (_35490_, _35488_, _07141_);
  nor (_35491_, _07141_, _07067_);
  or (_35492_, _35491_, _06758_);
  or (_35493_, _35492_, _35490_);
  and (_35494_, _35493_, _35486_);
  or (_35495_, _35494_, _06341_);
  and (_35496_, _35495_, _06010_);
  and (_35497_, _35496_, _35485_);
  nor (_35498_, _06010_, \oc8051_golden_model_1.SP [1]);
  or (_35499_, _35498_, _06461_);
  or (_35501_, _35499_, _35497_);
  nand (_35502_, _07301_, _06461_);
  and (_35503_, _35502_, _35501_);
  or (_35504_, _35503_, _06464_);
  or (_35505_, _35488_, _06465_);
  and (_35506_, _35505_, _07303_);
  and (_35507_, _35506_, _35504_);
  not (_35508_, _07494_);
  or (_35509_, _35508_, _07302_);
  or (_35510_, _35509_, _35507_);
  or (_35512_, _07494_, _07067_);
  and (_35513_, _35512_, _07215_);
  and (_35514_, _35513_, _35510_);
  nand (_35515_, _08173_, _07357_);
  and (_35516_, _35475_, _10080_);
  and (_35517_, _35516_, _35515_);
  or (_35518_, _35517_, _07460_);
  or (_35519_, _35518_, _35514_);
  or (_35520_, _35479_, _07208_);
  and (_35521_, _09451_, _07956_);
  or (_35523_, _35521_, _35520_);
  and (_35524_, _35523_, _05982_);
  and (_35525_, _35524_, _35519_);
  and (_35526_, _35475_, _10094_);
  or (_35527_, _14653_, _13872_);
  and (_35528_, _35527_, _35526_);
  or (_35529_, _35528_, _35525_);
  and (_35530_, _35529_, _06219_);
  and (_35531_, _35475_, _06218_);
  and (_35532_, _35531_, _35473_);
  or (_35534_, _35532_, _06217_);
  or (_35535_, _35534_, _35530_);
  nor (_35536_, _05952_, _07067_);
  nor (_35537_, _35536_, _06369_);
  and (_35538_, _35537_, _35535_);
  or (_35539_, _14668_, _13872_);
  and (_35540_, _35475_, _06369_);
  and (_35541_, _35540_, _35539_);
  or (_35542_, _35541_, _06536_);
  or (_35543_, _35542_, _35538_);
  and (_35545_, _11262_, _07956_);
  or (_35546_, _35545_, _35479_);
  or (_35547_, _35546_, _07240_);
  and (_35548_, _35547_, _07242_);
  and (_35549_, _35548_, _35543_);
  or (_35550_, _14666_, _13872_);
  and (_35551_, _35475_, _06375_);
  and (_35552_, _35551_, _35550_);
  or (_35553_, _35552_, _06545_);
  or (_35554_, _35553_, _35549_);
  and (_35556_, _35554_, _35481_);
  or (_35557_, _35556_, _07233_);
  nor (_35558_, _05961_, _07067_);
  nor (_35559_, _35558_, _06366_);
  and (_35560_, _35559_, _35557_);
  or (_35561_, _35560_, _35477_);
  and (_35562_, _35561_, _09061_);
  nor (_35563_, _11261_, _13872_);
  or (_35564_, _35563_, _35479_);
  and (_35565_, _35564_, _06528_);
  or (_35567_, _35565_, _06551_);
  nor (_35568_, _35567_, _35562_);
  or (_35569_, _35568_, _07044_);
  nor (_35570_, _06281_, _07253_);
  nand (_35571_, _35570_, _35569_);
  or (_35572_, _35570_, _07067_);
  and (_35573_, _35572_, _06926_);
  and (_35574_, _35573_, _35571_);
  and (_35575_, _35484_, _06568_);
  or (_35576_, _35575_, _07695_);
  or (_35578_, _35576_, _35574_);
  or (_35579_, _07271_, _07067_);
  and (_35580_, _35579_, _06279_);
  and (_35581_, _35580_, _35578_);
  or (_35582_, _35482_, _35479_);
  and (_35583_, _35582_, _06278_);
  or (_35584_, _35583_, _01351_);
  or (_35585_, _35584_, _35581_);
  or (_35586_, _01347_, \oc8051_golden_model_1.SP [1]);
  and (_35587_, _35586_, _42618_);
  and (_43322_, _35587_, _35585_);
  nor (_35589_, _01347_, _06715_);
  or (_35590_, _07866_, _05952_);
  nor (_35591_, _13872_, _07776_);
  nor (_35592_, _07956_, _06715_);
  or (_35593_, _35592_, _07215_);
  or (_35594_, _35593_, _35591_);
  or (_35595_, _07866_, _06007_);
  and (_35596_, _35595_, _05978_);
  and (_35597_, _14770_, _08173_);
  or (_35599_, _35597_, _35592_);
  and (_35600_, _35599_, _06341_);
  and (_35601_, _07956_, \oc8051_golden_model_1.ACC [2]);
  or (_35602_, _35601_, _35592_);
  and (_35603_, _35602_, _07141_);
  nor (_35604_, _07141_, _06715_);
  or (_35605_, _35604_, _06758_);
  or (_35606_, _35605_, _35603_);
  nand (_35607_, _16081_, _06758_);
  and (_35608_, _35607_, _07151_);
  and (_35610_, _35608_, _35606_);
  or (_35611_, _35610_, _27826_);
  or (_35612_, _35611_, _35600_);
  or (_35613_, _07866_, _06010_);
  nand (_35614_, _08684_, _06461_);
  and (_35615_, _35614_, _35613_);
  and (_35616_, _35615_, _35612_);
  or (_35617_, _35616_, _06464_);
  or (_35618_, _35602_, _06465_);
  and (_35619_, _35618_, _07303_);
  and (_35621_, _35619_, _35617_);
  or (_35622_, _07720_, _12613_);
  or (_35623_, _35622_, _35621_);
  and (_35624_, _35623_, _35596_);
  or (_35625_, _16081_, _05978_);
  nand (_35626_, _35625_, _07215_);
  or (_35627_, _35626_, _35624_);
  and (_35628_, _35627_, _35594_);
  or (_35629_, _35628_, _07460_);
  or (_35630_, _35592_, _07208_);
  and (_35632_, _09450_, _07956_);
  or (_35633_, _35632_, _35630_);
  and (_35634_, _35633_, _05982_);
  and (_35635_, _35634_, _35629_);
  and (_35636_, _14859_, _07956_);
  or (_35637_, _35636_, _35592_);
  and (_35638_, _35637_, _10094_);
  or (_35639_, _35638_, _06218_);
  or (_35640_, _35639_, _35635_);
  and (_35641_, _07956_, _08973_);
  or (_35643_, _35641_, _35592_);
  or (_35644_, _35643_, _06219_);
  and (_35645_, _35644_, _35640_);
  or (_35646_, _35645_, _06217_);
  and (_35647_, _35646_, _35590_);
  or (_35648_, _35647_, _06369_);
  and (_35649_, _14751_, _07956_);
  or (_35650_, _35649_, _35592_);
  or (_35651_, _35650_, _07237_);
  and (_35652_, _35651_, _07240_);
  and (_35654_, _35652_, _35648_);
  and (_35655_, _11259_, _07956_);
  or (_35656_, _35655_, _35592_);
  and (_35657_, _35656_, _06536_);
  or (_35658_, _35657_, _35654_);
  and (_35659_, _35658_, _07242_);
  or (_35660_, _35592_, _08440_);
  and (_35661_, _35643_, _06375_);
  and (_35662_, _35661_, _35660_);
  or (_35663_, _35662_, _35659_);
  and (_35665_, _35663_, _12772_);
  and (_35666_, _35602_, _06545_);
  and (_35667_, _35666_, _35660_);
  nor (_35668_, _16081_, _05961_);
  or (_35669_, _35668_, _06366_);
  or (_35670_, _35669_, _35667_);
  or (_35671_, _35670_, _35665_);
  and (_35672_, _14748_, _07956_);
  or (_35673_, _35672_, _35592_);
  or (_35674_, _35673_, _09056_);
  and (_35676_, _35674_, _35671_);
  or (_35677_, _35676_, _06528_);
  nor (_35678_, _11258_, _13872_);
  or (_35679_, _35678_, _35592_);
  or (_35680_, _35679_, _09061_);
  and (_35681_, _35680_, _06716_);
  and (_35682_, _35681_, _35677_);
  and (_35683_, _16081_, _06551_);
  or (_35684_, _35683_, _07253_);
  or (_35685_, _35684_, _35682_);
  nor (_35687_, _07866_, _05959_);
  nor (_35688_, _35687_, _06281_);
  and (_35689_, _35688_, _35685_);
  and (_35690_, _16081_, _06281_);
  or (_35691_, _35690_, _06568_);
  or (_35692_, _35691_, _35689_);
  or (_35693_, _35599_, _06926_);
  and (_35694_, _35693_, _07271_);
  and (_35695_, _35694_, _35692_);
  nor (_35696_, _16081_, _07271_);
  or (_35698_, _35696_, _06278_);
  or (_35699_, _35698_, _35695_);
  and (_35700_, _14926_, _08173_);
  or (_35701_, _35592_, _06279_);
  or (_35702_, _35701_, _35700_);
  and (_35703_, _35702_, _01347_);
  and (_35704_, _35703_, _35699_);
  or (_35705_, _35704_, _35589_);
  and (_43323_, _35705_, _42618_);
  nor (_35706_, _01347_, _06460_);
  or (_35708_, _07869_, _07271_);
  or (_35709_, _07869_, _05959_);
  or (_35710_, _07869_, _05952_);
  nor (_35711_, _13872_, _07594_);
  nor (_35712_, _07956_, _06460_);
  or (_35713_, _35712_, _07460_);
  or (_35714_, _35713_, _35711_);
  and (_35715_, _35714_, _12659_);
  and (_35716_, _14953_, _08173_);
  or (_35717_, _35716_, _35712_);
  or (_35719_, _35717_, _07151_);
  and (_35720_, _07956_, \oc8051_golden_model_1.ACC [3]);
  or (_35721_, _35720_, _35712_);
  or (_35722_, _35721_, _07142_);
  or (_35723_, _07141_, \oc8051_golden_model_1.SP [3]);
  and (_35724_, _35723_, _07504_);
  and (_35725_, _35724_, _35722_);
  and (_35726_, _07869_, _06758_);
  or (_35727_, _35726_, _06341_);
  or (_35728_, _35727_, _35725_);
  and (_35730_, _35728_, _06010_);
  and (_35731_, _35730_, _35719_);
  nor (_35732_, _15897_, _06010_);
  or (_35733_, _35732_, _06461_);
  or (_35734_, _35733_, _35731_);
  nand (_35735_, _08674_, _06461_);
  and (_35736_, _35735_, _35734_);
  or (_35737_, _35736_, _06464_);
  or (_35738_, _35721_, _06465_);
  and (_35739_, _35738_, _07303_);
  and (_35741_, _35739_, _35737_);
  or (_35742_, _07652_, _35508_);
  or (_35743_, _35742_, _35741_);
  or (_35744_, _07869_, _07494_);
  and (_35745_, _35744_, _07215_);
  and (_35746_, _35745_, _35743_);
  or (_35747_, _35746_, _35715_);
  or (_35748_, _35712_, _07208_);
  and (_35749_, _09449_, _07956_);
  or (_35750_, _35749_, _35748_);
  and (_35752_, _35750_, _05982_);
  and (_35753_, _35752_, _35747_);
  and (_35754_, _15048_, _07956_);
  or (_35755_, _35754_, _35712_);
  and (_35756_, _35755_, _10094_);
  or (_35757_, _35756_, _06218_);
  or (_35758_, _35757_, _35753_);
  and (_35759_, _07956_, _08930_);
  or (_35760_, _35759_, _35712_);
  or (_35761_, _35760_, _06219_);
  and (_35763_, _35761_, _35758_);
  or (_35764_, _35763_, _06217_);
  and (_35765_, _35764_, _35710_);
  or (_35766_, _35765_, _06369_);
  and (_35767_, _14943_, _07956_);
  or (_35768_, _35767_, _35712_);
  or (_35769_, _35768_, _07237_);
  and (_35770_, _35769_, _07240_);
  and (_35771_, _35770_, _35766_);
  and (_35772_, _12577_, _07956_);
  or (_35774_, _35772_, _35712_);
  and (_35775_, _35774_, _06536_);
  or (_35776_, _35775_, _35771_);
  and (_35777_, _35776_, _07242_);
  or (_35778_, _35712_, _08292_);
  and (_35779_, _35760_, _06375_);
  and (_35780_, _35779_, _35778_);
  or (_35781_, _35780_, _35777_);
  and (_35782_, _35781_, _12772_);
  and (_35783_, _35721_, _06545_);
  and (_35785_, _35783_, _35778_);
  nor (_35786_, _15897_, _05961_);
  or (_35787_, _35786_, _06366_);
  or (_35788_, _35787_, _35785_);
  or (_35789_, _35788_, _35782_);
  and (_35790_, _14940_, _08173_);
  or (_35791_, _35712_, _09056_);
  or (_35792_, _35791_, _35790_);
  and (_35793_, _35792_, _35789_);
  or (_35794_, _35793_, _06528_);
  nor (_35796_, _11256_, _13872_);
  or (_35797_, _35796_, _35712_);
  or (_35798_, _35797_, _09061_);
  and (_35799_, _35798_, _06716_);
  and (_35800_, _35799_, _35794_);
  nor (_35801_, _08671_, _06460_);
  or (_35802_, _35801_, _08672_);
  and (_35803_, _35802_, _06551_);
  or (_35804_, _35803_, _07253_);
  or (_35805_, _35804_, _35800_);
  and (_35807_, _35805_, _35709_);
  or (_35808_, _35807_, _06281_);
  or (_35809_, _35802_, _06282_);
  and (_35810_, _35809_, _06926_);
  and (_35811_, _35810_, _35808_);
  and (_35812_, _35717_, _06568_);
  or (_35813_, _35812_, _07695_);
  or (_35814_, _35813_, _35811_);
  and (_35815_, _35814_, _35708_);
  or (_35816_, _35815_, _06278_);
  and (_35818_, _15128_, _08173_);
  or (_35819_, _35712_, _06279_);
  or (_35820_, _35819_, _35818_);
  and (_35821_, _35820_, _01347_);
  and (_35822_, _35821_, _35816_);
  or (_35823_, _35822_, _35706_);
  and (_43325_, _35823_, _42618_);
  nor (_35824_, _01347_, _13845_);
  nor (_35825_, _07602_, \oc8051_golden_model_1.SP [4]);
  nor (_35826_, _35825_, _13814_);
  or (_35828_, _35826_, _07271_);
  nor (_35829_, _08541_, _13872_);
  nor (_35830_, _07956_, _13845_);
  or (_35831_, _35830_, _07460_);
  or (_35832_, _35831_, _35829_);
  and (_35833_, _35832_, _12659_);
  and (_35834_, _15162_, _08173_);
  or (_35835_, _35834_, _35830_);
  or (_35836_, _35835_, _07151_);
  and (_35837_, _07956_, \oc8051_golden_model_1.ACC [4]);
  or (_35839_, _35837_, _35830_);
  or (_35840_, _35839_, _07142_);
  or (_35841_, _07141_, \oc8051_golden_model_1.SP [4]);
  and (_35842_, _35841_, _07504_);
  and (_35843_, _35842_, _35840_);
  and (_35844_, _35826_, _06758_);
  or (_35845_, _35844_, _06341_);
  or (_35846_, _35845_, _35843_);
  and (_35847_, _35846_, _06010_);
  and (_35848_, _35847_, _35836_);
  and (_35850_, _35826_, _07611_);
  or (_35851_, _35850_, _06461_);
  or (_35852_, _35851_, _35848_);
  and (_35853_, _13846_, _06800_);
  nor (_35854_, _08673_, _13845_);
  nor (_35855_, _35854_, _35853_);
  nand (_35856_, _35855_, _06461_);
  and (_35857_, _35856_, _35852_);
  or (_35858_, _35857_, _06464_);
  or (_35859_, _35839_, _06465_);
  and (_35861_, _35859_, _07303_);
  and (_35862_, _35861_, _35858_);
  and (_35863_, _07603_, \oc8051_golden_model_1.SP [4]);
  nor (_35864_, _07603_, \oc8051_golden_model_1.SP [4]);
  nor (_35865_, _35864_, _35863_);
  nand (_35866_, _35865_, _06267_);
  nand (_35867_, _35866_, _07494_);
  or (_35868_, _35867_, _35862_);
  or (_35869_, _35826_, _07494_);
  and (_35870_, _35869_, _07215_);
  and (_35872_, _35870_, _35868_);
  or (_35873_, _35872_, _35833_);
  or (_35874_, _35830_, _07208_);
  and (_35875_, _09448_, _07956_);
  or (_35876_, _35875_, _35874_);
  and (_35877_, _35876_, _05982_);
  and (_35878_, _35877_, _35873_);
  and (_35879_, _15254_, _07956_);
  or (_35880_, _35879_, _35830_);
  and (_35881_, _35880_, _10094_);
  or (_35883_, _35881_, _06218_);
  or (_35884_, _35883_, _35878_);
  and (_35885_, _08959_, _07956_);
  or (_35886_, _35885_, _35830_);
  or (_35887_, _35886_, _06219_);
  and (_35888_, _35887_, _35884_);
  or (_35889_, _35888_, _06217_);
  or (_35890_, _35826_, _05952_);
  and (_35891_, _35890_, _35889_);
  or (_35892_, _35891_, _06369_);
  and (_35894_, _15269_, _07956_);
  or (_35895_, _35894_, _35830_);
  or (_35896_, _35895_, _07237_);
  and (_35897_, _35896_, _07240_);
  and (_35898_, _35897_, _35892_);
  and (_35899_, _11254_, _07956_);
  or (_35900_, _35899_, _35830_);
  and (_35901_, _35900_, _06536_);
  or (_35902_, _35901_, _35898_);
  and (_35903_, _35902_, _07242_);
  or (_35905_, _35830_, _08544_);
  and (_35906_, _35886_, _06375_);
  and (_35907_, _35906_, _35905_);
  or (_35908_, _35907_, _35903_);
  and (_35909_, _35908_, _12772_);
  and (_35910_, _35839_, _06545_);
  and (_35911_, _35910_, _35905_);
  and (_35912_, _35826_, _07233_);
  or (_35913_, _35912_, _06366_);
  or (_35914_, _35913_, _35911_);
  or (_35916_, _35914_, _35909_);
  and (_35917_, _15266_, _07956_);
  or (_35918_, _35917_, _35830_);
  or (_35919_, _35918_, _09056_);
  and (_35920_, _35919_, _35916_);
  or (_35921_, _35920_, _06528_);
  nor (_35922_, _11253_, _13872_);
  or (_35923_, _35922_, _35830_);
  or (_35924_, _35923_, _09061_);
  and (_35925_, _35924_, _06716_);
  and (_35927_, _35925_, _35921_);
  nor (_35928_, _08672_, _13845_);
  or (_35929_, _35928_, _13846_);
  and (_35930_, _35929_, _06551_);
  or (_35931_, _35930_, _07253_);
  or (_35932_, _35931_, _35927_);
  or (_35933_, _35826_, _05959_);
  and (_35934_, _35933_, _35932_);
  or (_35935_, _35934_, _06281_);
  or (_35936_, _35929_, _06282_);
  and (_35938_, _35936_, _06926_);
  and (_35939_, _35938_, _35935_);
  and (_35940_, _35835_, _06568_);
  or (_35941_, _35940_, _07695_);
  or (_35942_, _35941_, _35939_);
  and (_35943_, _35942_, _35828_);
  or (_35944_, _35943_, _06278_);
  and (_35945_, _15329_, _08173_);
  or (_35946_, _35830_, _06279_);
  or (_35947_, _35946_, _35945_);
  and (_35949_, _35947_, _01347_);
  and (_35950_, _35949_, _35944_);
  or (_35951_, _35950_, _35824_);
  and (_43326_, _35951_, _42618_);
  nor (_35952_, _01347_, _13844_);
  nor (_35953_, _13814_, \oc8051_golden_model_1.SP [5]);
  nor (_35954_, _35953_, _13815_);
  or (_35955_, _35954_, _07271_);
  nor (_35956_, _08244_, _13872_);
  nor (_35957_, _07956_, _13844_);
  or (_35959_, _35957_, _07460_);
  or (_35960_, _35959_, _35956_);
  and (_35961_, _35960_, _12659_);
  and (_35962_, _15358_, _08173_);
  or (_35963_, _35962_, _35957_);
  or (_35964_, _35963_, _07151_);
  and (_35965_, _07956_, \oc8051_golden_model_1.ACC [5]);
  or (_35966_, _35965_, _35957_);
  and (_35967_, _35966_, _07141_);
  nor (_35968_, _07141_, _13844_);
  or (_35970_, _35968_, _06758_);
  or (_35971_, _35970_, _35967_);
  or (_35972_, _35954_, _07504_);
  and (_35973_, _35972_, _35971_);
  or (_35974_, _35973_, _06341_);
  and (_35975_, _35974_, _06010_);
  and (_35976_, _35975_, _35964_);
  and (_35977_, _35954_, _07611_);
  or (_35978_, _35977_, _06461_);
  or (_35979_, _35978_, _35976_);
  and (_35981_, _13847_, _06800_);
  nor (_35982_, _35853_, _13844_);
  nor (_35983_, _35982_, _35981_);
  nand (_35984_, _35983_, _06461_);
  and (_35985_, _35984_, _35979_);
  or (_35986_, _35985_, _06464_);
  or (_35987_, _35966_, _06465_);
  and (_35988_, _35987_, _07303_);
  and (_35989_, _35988_, _35986_);
  nor (_35990_, _35863_, \oc8051_golden_model_1.SP [5]);
  nor (_35992_, _35990_, _13859_);
  nand (_35993_, _35992_, _06267_);
  nand (_35994_, _35993_, _07494_);
  or (_35995_, _35994_, _35989_);
  or (_35996_, _35954_, _07494_);
  and (_35997_, _35996_, _07215_);
  and (_35998_, _35997_, _35995_);
  or (_35999_, _35998_, _35961_);
  or (_36000_, _35957_, _07208_);
  and (_36001_, _09447_, _07956_);
  or (_36003_, _36001_, _36000_);
  and (_36004_, _36003_, _05982_);
  and (_36005_, _36004_, _35999_);
  and (_36006_, _15459_, _07956_);
  or (_36007_, _36006_, _35957_);
  and (_36008_, _36007_, _10094_);
  or (_36009_, _36008_, _06218_);
  or (_36010_, _36009_, _36005_);
  and (_36011_, _08946_, _07956_);
  or (_36012_, _36011_, _35957_);
  or (_36014_, _36012_, _06219_);
  and (_36015_, _36014_, _36010_);
  or (_36016_, _36015_, _06217_);
  or (_36017_, _35954_, _05952_);
  and (_36018_, _36017_, _36016_);
  or (_36019_, _36018_, _06369_);
  and (_36020_, _15353_, _07956_);
  or (_36021_, _36020_, _35957_);
  or (_36022_, _36021_, _07237_);
  and (_36023_, _36022_, _07240_);
  and (_36025_, _36023_, _36019_);
  and (_36026_, _11250_, _07956_);
  or (_36027_, _36026_, _35957_);
  and (_36028_, _36027_, _06536_);
  or (_36029_, _36028_, _36025_);
  and (_36030_, _36029_, _07242_);
  or (_36031_, _35957_, _08247_);
  and (_36032_, _36012_, _06375_);
  and (_36033_, _36032_, _36031_);
  or (_36034_, _36033_, _36030_);
  and (_36036_, _36034_, _12772_);
  and (_36037_, _35966_, _06545_);
  and (_36038_, _36037_, _36031_);
  and (_36039_, _35954_, _07233_);
  or (_36040_, _36039_, _06366_);
  or (_36041_, _36040_, _36038_);
  or (_36042_, _36041_, _36036_);
  and (_36043_, _15350_, _07956_);
  or (_36044_, _36043_, _35957_);
  or (_36045_, _36044_, _09056_);
  and (_36047_, _36045_, _36042_);
  or (_36048_, _36047_, _06528_);
  nor (_36049_, _11249_, _13872_);
  or (_36050_, _36049_, _35957_);
  or (_36051_, _36050_, _09061_);
  and (_36052_, _36051_, _06716_);
  and (_36053_, _36052_, _36048_);
  nor (_36054_, _13846_, _13844_);
  or (_36055_, _36054_, _13847_);
  and (_36056_, _36055_, _06551_);
  or (_36058_, _36056_, _07253_);
  or (_36059_, _36058_, _36053_);
  or (_36060_, _35954_, _05959_);
  and (_36061_, _36060_, _36059_);
  or (_36062_, _36061_, _06281_);
  or (_36063_, _36055_, _06282_);
  and (_36064_, _36063_, _06926_);
  and (_36065_, _36064_, _36062_);
  and (_36066_, _35963_, _06568_);
  or (_36067_, _36066_, _07695_);
  or (_36069_, _36067_, _36065_);
  and (_36070_, _36069_, _35955_);
  or (_36071_, _36070_, _06278_);
  and (_36072_, _15532_, _08173_);
  or (_36073_, _35957_, _06279_);
  or (_36074_, _36073_, _36072_);
  and (_36075_, _36074_, _01347_);
  and (_36076_, _36075_, _36071_);
  or (_36077_, _36076_, _35952_);
  and (_43327_, _36077_, _42618_);
  nor (_36079_, _01347_, _13843_);
  nor (_36080_, _07956_, _13843_);
  and (_36081_, _15554_, _08173_);
  or (_36082_, _36081_, _36080_);
  or (_36083_, _36082_, _07151_);
  and (_36084_, _07956_, \oc8051_golden_model_1.ACC [6]);
  or (_36085_, _36084_, _36080_);
  and (_36086_, _36085_, _07141_);
  nor (_36087_, _07141_, _13843_);
  or (_36088_, _36087_, _06758_);
  or (_36090_, _36088_, _36086_);
  nor (_36091_, _13815_, \oc8051_golden_model_1.SP [6]);
  nor (_36092_, _36091_, _13816_);
  or (_36093_, _36092_, _07504_);
  and (_36094_, _36093_, _36090_);
  or (_36095_, _36094_, _06341_);
  and (_36096_, _36095_, _06010_);
  and (_36097_, _36096_, _36083_);
  and (_36098_, _36092_, _07611_);
  or (_36099_, _36098_, _06461_);
  or (_36101_, _36099_, _36097_);
  nor (_36102_, _35981_, _13843_);
  nor (_36103_, _36102_, _13849_);
  nand (_36104_, _36103_, _06461_);
  and (_36105_, _36104_, _36101_);
  or (_36106_, _36105_, _06464_);
  or (_36107_, _36085_, _06465_);
  and (_36108_, _36107_, _07303_);
  and (_36109_, _36108_, _36106_);
  nor (_36110_, _13859_, \oc8051_golden_model_1.SP [6]);
  nor (_36112_, _36110_, _13860_);
  and (_36113_, _36112_, _06267_);
  or (_36114_, _36113_, _36109_);
  and (_36115_, _36114_, _07494_);
  nand (_36116_, _36092_, _35508_);
  nand (_36117_, _36116_, _07215_);
  or (_36118_, _36117_, _36115_);
  nor (_36119_, _08142_, _13872_);
  or (_36120_, _36080_, _07215_);
  or (_36121_, _36120_, _36119_);
  and (_36123_, _36121_, _36118_);
  or (_36124_, _36123_, _07460_);
  and (_36125_, _09446_, _07956_);
  or (_36126_, _36080_, _07208_);
  or (_36127_, _36126_, _36125_);
  and (_36128_, _36127_, _05982_);
  and (_36129_, _36128_, _36124_);
  and (_36130_, _15657_, _08173_);
  or (_36131_, _36130_, _36080_);
  and (_36132_, _36131_, _10094_);
  or (_36134_, _36132_, _06218_);
  or (_36135_, _36134_, _36129_);
  and (_36136_, _15664_, _07956_);
  or (_36137_, _36136_, _36080_);
  or (_36138_, _36137_, _06219_);
  and (_36139_, _36138_, _36135_);
  or (_36140_, _36139_, _06217_);
  or (_36141_, _36092_, _05952_);
  and (_36142_, _36141_, _36140_);
  or (_36143_, _36142_, _06369_);
  and (_36145_, _15549_, _07956_);
  or (_36146_, _36145_, _36080_);
  or (_36147_, _36146_, _07237_);
  and (_36148_, _36147_, _07240_);
  and (_36149_, _36148_, _36143_);
  and (_36150_, _11247_, _07956_);
  or (_36151_, _36150_, _36080_);
  and (_36152_, _36151_, _06536_);
  or (_36153_, _36152_, _36149_);
  and (_36154_, _36153_, _07242_);
  or (_36156_, _36080_, _08145_);
  and (_36157_, _36137_, _06375_);
  and (_36158_, _36157_, _36156_);
  or (_36159_, _36158_, _36154_);
  and (_36160_, _36159_, _12772_);
  and (_36161_, _36085_, _06545_);
  and (_36162_, _36161_, _36156_);
  and (_36163_, _36092_, _07233_);
  or (_36164_, _36163_, _06366_);
  or (_36165_, _36164_, _36162_);
  or (_36167_, _36165_, _36160_);
  and (_36168_, _15546_, _07956_);
  or (_36169_, _36168_, _36080_);
  or (_36170_, _36169_, _09056_);
  and (_36171_, _36170_, _36167_);
  or (_36172_, _36171_, _06528_);
  nor (_36173_, _11246_, _13872_);
  or (_36174_, _36173_, _36080_);
  or (_36175_, _36174_, _09061_);
  and (_36176_, _36175_, _06716_);
  and (_36178_, _36176_, _36172_);
  nor (_36179_, _13847_, _13843_);
  or (_36180_, _36179_, _13848_);
  and (_36181_, _36180_, _06551_);
  or (_36182_, _36181_, _07253_);
  or (_36183_, _36182_, _36178_);
  nor (_36184_, _36092_, _05959_);
  nor (_36185_, _36184_, _06281_);
  and (_36186_, _36185_, _36183_);
  and (_36187_, _36180_, _06281_);
  or (_36189_, _36187_, _06568_);
  or (_36190_, _36189_, _36186_);
  or (_36191_, _36082_, _06926_);
  and (_36192_, _36191_, _07271_);
  and (_36193_, _36192_, _36190_);
  and (_36194_, _36092_, _07695_);
  or (_36195_, _36194_, _06278_);
  or (_36196_, _36195_, _36193_);
  and (_36197_, _15734_, _08173_);
  or (_36198_, _36080_, _06279_);
  or (_36200_, _36198_, _36197_);
  and (_36201_, _36200_, _01347_);
  and (_36202_, _36201_, _36196_);
  or (_36203_, _36202_, _36079_);
  and (_43328_, _36203_, _42618_);
  not (_36204_, \oc8051_golden_model_1.SBUF [0]);
  nor (_36205_, _01347_, _36204_);
  nand (_36206_, _11263_, _07886_);
  nor (_36207_, _07886_, _36204_);
  nor (_36208_, _36207_, _07234_);
  nand (_36210_, _36208_, _36206_);
  and (_36211_, _07886_, \oc8051_golden_model_1.ACC [0]);
  or (_36212_, _36211_, _36207_);
  and (_36213_, _36212_, _06464_);
  or (_36214_, _36213_, _10080_);
  nor (_36215_, _08390_, _13951_);
  or (_36216_, _36215_, _36207_);
  and (_36217_, _36216_, _06341_);
  nor (_36218_, _07141_, _36204_);
  and (_36219_, _36212_, _07141_);
  or (_36220_, _36219_, _36218_);
  and (_36221_, _36220_, _07151_);
  or (_36222_, _36221_, _06461_);
  or (_36223_, _36222_, _36217_);
  and (_36224_, _36223_, _06465_);
  or (_36225_, _36224_, _36214_);
  and (_36226_, _07886_, _07133_);
  or (_36227_, _36207_, _22611_);
  or (_36228_, _36227_, _36226_);
  and (_36229_, _36228_, _36225_);
  or (_36231_, _36229_, _07460_);
  and (_36232_, _09392_, _07886_);
  or (_36233_, _36207_, _07208_);
  or (_36234_, _36233_, _36232_);
  and (_36235_, _36234_, _36231_);
  or (_36236_, _36235_, _10094_);
  and (_36237_, _14467_, _07886_);
  or (_36238_, _36207_, _05982_);
  or (_36239_, _36238_, _36237_);
  and (_36240_, _36239_, _06219_);
  and (_36242_, _36240_, _36236_);
  and (_36243_, _07886_, _08954_);
  or (_36244_, _36243_, _36207_);
  and (_36245_, _36244_, _06218_);
  or (_36246_, _36245_, _06369_);
  or (_36247_, _36246_, _36242_);
  and (_36248_, _14366_, _07886_);
  or (_36249_, _36248_, _36207_);
  or (_36250_, _36249_, _07237_);
  and (_36251_, _36250_, _07240_);
  and (_36253_, _36251_, _36247_);
  nor (_36254_, _12580_, _13951_);
  or (_36255_, _36254_, _36207_);
  and (_36256_, _36206_, _06536_);
  and (_36257_, _36256_, _36255_);
  or (_36258_, _36257_, _36253_);
  and (_36259_, _36258_, _07242_);
  nand (_36260_, _36244_, _06375_);
  nor (_36261_, _36260_, _36215_);
  or (_36262_, _36261_, _06545_);
  or (_36264_, _36262_, _36259_);
  and (_36265_, _36264_, _36210_);
  or (_36266_, _36265_, _06366_);
  and (_36267_, _14363_, _07886_);
  or (_36268_, _36207_, _09056_);
  or (_36269_, _36268_, _36267_);
  and (_36270_, _36269_, _09061_);
  and (_36271_, _36270_, _36266_);
  and (_36272_, _36255_, _06528_);
  or (_36273_, _36272_, _19502_);
  or (_36275_, _36273_, _36271_);
  or (_36276_, _36216_, _06661_);
  and (_36277_, _36276_, _01347_);
  and (_36278_, _36277_, _36275_);
  or (_36279_, _36278_, _36205_);
  and (_43330_, _36279_, _42618_);
  not (_36280_, \oc8051_golden_model_1.SBUF [1]);
  nor (_36281_, _01347_, _36280_);
  nand (_36282_, _07886_, _07038_);
  or (_36283_, _07886_, \oc8051_golden_model_1.SBUF [1]);
  and (_36285_, _36283_, _06218_);
  and (_36286_, _36285_, _36282_);
  nor (_36287_, _07886_, _36280_);
  nor (_36288_, _13951_, _07357_);
  or (_36289_, _36288_, _36287_);
  or (_36290_, _36289_, _07215_);
  and (_36291_, _14562_, _07886_);
  not (_36292_, _36291_);
  and (_36293_, _36292_, _36283_);
  or (_36294_, _36293_, _07151_);
  and (_36296_, _07886_, \oc8051_golden_model_1.ACC [1]);
  or (_36297_, _36296_, _36287_);
  and (_36298_, _36297_, _07141_);
  nor (_36299_, _07141_, _36280_);
  or (_36300_, _36299_, _06341_);
  or (_36301_, _36300_, _36298_);
  and (_36302_, _36301_, _07166_);
  and (_36303_, _36302_, _36294_);
  and (_36304_, _36289_, _06461_);
  or (_36305_, _36304_, _36303_);
  and (_36307_, _36305_, _06465_);
  and (_36308_, _36297_, _06464_);
  or (_36309_, _36308_, _10080_);
  or (_36310_, _36309_, _36307_);
  and (_36311_, _36310_, _36290_);
  or (_36312_, _36311_, _07460_);
  and (_36313_, _09451_, _07886_);
  or (_36314_, _36287_, _07208_);
  or (_36315_, _36314_, _36313_);
  and (_36316_, _36315_, _05982_);
  and (_36318_, _36316_, _36312_);
  or (_36319_, _14653_, _13951_);
  and (_36320_, _36283_, _10094_);
  and (_36321_, _36320_, _36319_);
  or (_36322_, _36321_, _36318_);
  and (_36323_, _36322_, _06219_);
  or (_36324_, _36323_, _36286_);
  and (_36325_, _36324_, _07237_);
  or (_36326_, _14668_, _13951_);
  and (_36327_, _36283_, _06369_);
  and (_36329_, _36327_, _36326_);
  or (_36330_, _36329_, _06536_);
  or (_36331_, _36330_, _36325_);
  nor (_36332_, _11261_, _13951_);
  or (_36333_, _36332_, _36287_);
  nand (_36334_, _11260_, _07886_);
  and (_36335_, _36334_, _36333_);
  or (_36336_, _36335_, _07240_);
  and (_36337_, _36336_, _07242_);
  and (_36338_, _36337_, _36331_);
  or (_36340_, _14666_, _13951_);
  and (_36341_, _36283_, _06375_);
  and (_36342_, _36341_, _36340_);
  or (_36343_, _36342_, _06545_);
  or (_36344_, _36343_, _36338_);
  nor (_36345_, _36287_, _07234_);
  nand (_36346_, _36345_, _36334_);
  and (_36347_, _36346_, _09056_);
  and (_36348_, _36347_, _36344_);
  or (_36349_, _36282_, _08341_);
  and (_36351_, _36283_, _06366_);
  and (_36352_, _36351_, _36349_);
  or (_36353_, _36352_, _06528_);
  or (_36354_, _36353_, _36348_);
  or (_36355_, _36333_, _09061_);
  and (_36356_, _36355_, _06926_);
  and (_36357_, _36356_, _36354_);
  and (_36358_, _36293_, _06568_);
  or (_36359_, _36358_, _06278_);
  or (_36360_, _36359_, _36357_);
  or (_36362_, _36287_, _06279_);
  or (_36363_, _36362_, _36291_);
  and (_36364_, _36363_, _01347_);
  and (_36365_, _36364_, _36360_);
  or (_36366_, _36365_, _36281_);
  and (_43331_, _36366_, _42618_);
  and (_36367_, _01351_, \oc8051_golden_model_1.SBUF [2]);
  and (_36368_, _13951_, \oc8051_golden_model_1.SBUF [2]);
  and (_36369_, _09450_, _07886_);
  or (_36370_, _36369_, _36368_);
  and (_36372_, _36370_, _07460_);
  and (_36373_, _14770_, _07886_);
  or (_36374_, _36373_, _36368_);
  or (_36375_, _36374_, _07151_);
  and (_36376_, _07886_, \oc8051_golden_model_1.ACC [2]);
  or (_36377_, _36376_, _36368_);
  and (_36378_, _36377_, _07141_);
  and (_36379_, _07142_, \oc8051_golden_model_1.SBUF [2]);
  or (_36380_, _36379_, _06341_);
  or (_36381_, _36380_, _36378_);
  and (_36383_, _36381_, _07166_);
  and (_36384_, _36383_, _36375_);
  nor (_36385_, _13951_, _07776_);
  or (_36386_, _36385_, _36368_);
  and (_36387_, _36386_, _06461_);
  or (_36388_, _36387_, _36384_);
  and (_36389_, _36388_, _06465_);
  and (_36390_, _36377_, _06464_);
  or (_36391_, _36390_, _10080_);
  or (_36392_, _36391_, _36389_);
  or (_36394_, _36386_, _07215_);
  and (_36395_, _36394_, _07208_);
  and (_36396_, _36395_, _36392_);
  or (_36397_, _36396_, _10094_);
  or (_36398_, _36397_, _36372_);
  and (_36399_, _14859_, _07886_);
  or (_36400_, _36368_, _05982_);
  or (_36401_, _36400_, _36399_);
  and (_36402_, _36401_, _06219_);
  and (_36403_, _36402_, _36398_);
  and (_36405_, _07886_, _08973_);
  or (_36406_, _36405_, _36368_);
  and (_36407_, _36406_, _06218_);
  or (_36408_, _36407_, _06369_);
  or (_36409_, _36408_, _36403_);
  and (_36410_, _14751_, _07886_);
  or (_36411_, _36410_, _36368_);
  or (_36412_, _36411_, _07237_);
  and (_36413_, _36412_, _07240_);
  and (_36414_, _36413_, _36409_);
  and (_36416_, _11259_, _07886_);
  or (_36417_, _36416_, _36368_);
  and (_36418_, _36417_, _06536_);
  or (_36419_, _36418_, _36414_);
  and (_36420_, _36419_, _07242_);
  or (_36421_, _36368_, _08440_);
  and (_36422_, _36406_, _06375_);
  and (_36423_, _36422_, _36421_);
  or (_36424_, _36423_, _36420_);
  and (_36425_, _36424_, _07234_);
  and (_36427_, _36377_, _06545_);
  and (_36428_, _36427_, _36421_);
  or (_36429_, _36428_, _06366_);
  or (_36430_, _36429_, _36425_);
  and (_36431_, _14748_, _07886_);
  or (_36432_, _36368_, _09056_);
  or (_36433_, _36432_, _36431_);
  and (_36434_, _36433_, _09061_);
  and (_36435_, _36434_, _36430_);
  nor (_36436_, _11258_, _13951_);
  or (_36438_, _36436_, _36368_);
  and (_36439_, _36438_, _06528_);
  or (_36440_, _36439_, _36435_);
  and (_36441_, _36440_, _06926_);
  and (_36442_, _36374_, _06568_);
  or (_36443_, _36442_, _06278_);
  or (_36444_, _36443_, _36441_);
  and (_36445_, _14926_, _07886_);
  or (_36446_, _36368_, _06279_);
  or (_36447_, _36446_, _36445_);
  and (_36449_, _36447_, _01347_);
  and (_36450_, _36449_, _36444_);
  or (_36451_, _36450_, _36367_);
  and (_43332_, _36451_, _42618_);
  and (_36452_, _01351_, \oc8051_golden_model_1.SBUF [3]);
  and (_36453_, _13951_, \oc8051_golden_model_1.SBUF [3]);
  and (_36454_, _14953_, _07886_);
  or (_36455_, _36454_, _36453_);
  or (_36456_, _36455_, _07151_);
  and (_36457_, _07886_, \oc8051_golden_model_1.ACC [3]);
  or (_36459_, _36457_, _36453_);
  and (_36460_, _36459_, _07141_);
  and (_36461_, _07142_, \oc8051_golden_model_1.SBUF [3]);
  or (_36462_, _36461_, _06341_);
  or (_36463_, _36462_, _36460_);
  and (_36464_, _36463_, _07166_);
  and (_36465_, _36464_, _36456_);
  nor (_36466_, _13951_, _07594_);
  or (_36467_, _36466_, _36453_);
  and (_36468_, _36467_, _06461_);
  or (_36470_, _36468_, _36465_);
  and (_36471_, _36470_, _06465_);
  and (_36472_, _36459_, _06464_);
  or (_36473_, _36472_, _10080_);
  or (_36474_, _36473_, _36471_);
  or (_36475_, _36467_, _07215_);
  and (_36476_, _36475_, _36474_);
  or (_36477_, _36476_, _07460_);
  and (_36478_, _09449_, _07886_);
  or (_36479_, _36453_, _07208_);
  or (_36481_, _36479_, _36478_);
  and (_36482_, _36481_, _05982_);
  and (_36483_, _36482_, _36477_);
  and (_36484_, _15048_, _07886_);
  or (_36485_, _36484_, _36453_);
  and (_36486_, _36485_, _10094_);
  or (_36487_, _36486_, _06218_);
  or (_36488_, _36487_, _36483_);
  and (_36489_, _07886_, _08930_);
  or (_36490_, _36489_, _36453_);
  or (_36492_, _36490_, _06219_);
  and (_36493_, _36492_, _36488_);
  or (_36494_, _36493_, _06369_);
  and (_36495_, _14943_, _07886_);
  or (_36496_, _36495_, _36453_);
  or (_36497_, _36496_, _07237_);
  and (_36498_, _36497_, _07240_);
  and (_36499_, _36498_, _36494_);
  and (_36500_, _12577_, _07886_);
  or (_36501_, _36500_, _36453_);
  and (_36503_, _36501_, _06536_);
  or (_36504_, _36503_, _36499_);
  and (_36505_, _36504_, _07242_);
  or (_36506_, _36453_, _08292_);
  and (_36507_, _36490_, _06375_);
  and (_36508_, _36507_, _36506_);
  or (_36509_, _36508_, _36505_);
  and (_36510_, _36509_, _07234_);
  and (_36511_, _36459_, _06545_);
  and (_36512_, _36511_, _36506_);
  or (_36514_, _36512_, _06366_);
  or (_36515_, _36514_, _36510_);
  and (_36516_, _14940_, _07886_);
  or (_36517_, _36453_, _09056_);
  or (_36518_, _36517_, _36516_);
  and (_36519_, _36518_, _09061_);
  and (_36520_, _36519_, _36515_);
  nor (_36521_, _11256_, _13951_);
  or (_36522_, _36521_, _36453_);
  and (_36523_, _36522_, _06528_);
  or (_36525_, _36523_, _36520_);
  and (_36526_, _36525_, _06926_);
  and (_36527_, _36455_, _06568_);
  or (_36528_, _36527_, _06278_);
  or (_36529_, _36528_, _36526_);
  and (_36530_, _15128_, _07886_);
  or (_36531_, _36453_, _06279_);
  or (_36532_, _36531_, _36530_);
  and (_36533_, _36532_, _01347_);
  and (_36534_, _36533_, _36529_);
  or (_36536_, _36534_, _36452_);
  and (_43333_, _36536_, _42618_);
  and (_36537_, _01351_, \oc8051_golden_model_1.SBUF [4]);
  and (_36538_, _13951_, \oc8051_golden_model_1.SBUF [4]);
  nor (_36539_, _08541_, _13951_);
  or (_36540_, _36539_, _36538_);
  or (_36541_, _36540_, _07215_);
  and (_36542_, _15162_, _07886_);
  or (_36543_, _36542_, _36538_);
  or (_36544_, _36543_, _07151_);
  and (_36546_, _07886_, \oc8051_golden_model_1.ACC [4]);
  or (_36547_, _36546_, _36538_);
  and (_36548_, _36547_, _07141_);
  and (_36549_, _07142_, \oc8051_golden_model_1.SBUF [4]);
  or (_36550_, _36549_, _06341_);
  or (_36551_, _36550_, _36548_);
  and (_36552_, _36551_, _07166_);
  and (_36553_, _36552_, _36544_);
  and (_36554_, _36540_, _06461_);
  or (_36555_, _36554_, _36553_);
  and (_36557_, _36555_, _06465_);
  and (_36558_, _36547_, _06464_);
  or (_36559_, _36558_, _10080_);
  or (_36560_, _36559_, _36557_);
  and (_36561_, _36560_, _07208_);
  and (_36562_, _36561_, _36541_);
  and (_36563_, _09448_, _07886_);
  or (_36564_, _36563_, _36538_);
  and (_36565_, _36564_, _07460_);
  or (_36566_, _36565_, _10094_);
  or (_36568_, _36566_, _36562_);
  and (_36569_, _15254_, _07886_);
  or (_36570_, _36538_, _05982_);
  or (_36571_, _36570_, _36569_);
  and (_36572_, _36571_, _06219_);
  and (_36573_, _36572_, _36568_);
  and (_36574_, _08959_, _07886_);
  or (_36575_, _36574_, _36538_);
  and (_36576_, _36575_, _06218_);
  or (_36577_, _36576_, _06369_);
  or (_36579_, _36577_, _36573_);
  and (_36580_, _15269_, _07886_);
  or (_36581_, _36580_, _36538_);
  or (_36582_, _36581_, _07237_);
  and (_36583_, _36582_, _07240_);
  and (_36584_, _36583_, _36579_);
  and (_36585_, _11254_, _07886_);
  or (_36586_, _36585_, _36538_);
  and (_36587_, _36586_, _06536_);
  or (_36588_, _36587_, _36584_);
  and (_36590_, _36588_, _07242_);
  or (_36591_, _36538_, _08544_);
  and (_36592_, _36575_, _06375_);
  and (_36593_, _36592_, _36591_);
  or (_36594_, _36593_, _36590_);
  and (_36595_, _36594_, _07234_);
  and (_36596_, _36547_, _06545_);
  and (_36597_, _36596_, _36591_);
  or (_36598_, _36597_, _06366_);
  or (_36599_, _36598_, _36595_);
  and (_36601_, _15266_, _07886_);
  or (_36602_, _36538_, _09056_);
  or (_36603_, _36602_, _36601_);
  and (_36604_, _36603_, _09061_);
  and (_36605_, _36604_, _36599_);
  nor (_36606_, _11253_, _13951_);
  or (_36607_, _36606_, _36538_);
  and (_36608_, _36607_, _06528_);
  or (_36609_, _36608_, _36605_);
  and (_36610_, _36609_, _06926_);
  and (_36612_, _36543_, _06568_);
  or (_36613_, _36612_, _06278_);
  or (_36614_, _36613_, _36610_);
  and (_36615_, _15329_, _07886_);
  or (_36616_, _36538_, _06279_);
  or (_36617_, _36616_, _36615_);
  and (_36618_, _36617_, _01347_);
  and (_36619_, _36618_, _36614_);
  or (_36620_, _36619_, _36537_);
  and (_43334_, _36620_, _42618_);
  and (_36622_, _01351_, \oc8051_golden_model_1.SBUF [5]);
  and (_36623_, _13951_, \oc8051_golden_model_1.SBUF [5]);
  nor (_36624_, _08244_, _13951_);
  or (_36625_, _36624_, _36623_);
  or (_36626_, _36625_, _07215_);
  and (_36627_, _15358_, _07886_);
  or (_36628_, _36627_, _36623_);
  or (_36629_, _36628_, _07151_);
  and (_36630_, _07886_, \oc8051_golden_model_1.ACC [5]);
  or (_36631_, _36630_, _36623_);
  and (_36633_, _36631_, _07141_);
  and (_36634_, _07142_, \oc8051_golden_model_1.SBUF [5]);
  or (_36635_, _36634_, _06341_);
  or (_36636_, _36635_, _36633_);
  and (_36637_, _36636_, _07166_);
  and (_36638_, _36637_, _36629_);
  and (_36639_, _36625_, _06461_);
  or (_36640_, _36639_, _36638_);
  and (_36641_, _36640_, _06465_);
  and (_36642_, _36631_, _06464_);
  or (_36644_, _36642_, _10080_);
  or (_36645_, _36644_, _36641_);
  and (_36646_, _36645_, _36626_);
  or (_36647_, _36646_, _07460_);
  and (_36648_, _09447_, _07886_);
  or (_36649_, _36623_, _07208_);
  or (_36650_, _36649_, _36648_);
  and (_36651_, _36650_, _05982_);
  and (_36652_, _36651_, _36647_);
  and (_36653_, _15459_, _07886_);
  or (_36655_, _36653_, _36623_);
  and (_36656_, _36655_, _10094_);
  or (_36657_, _36656_, _06218_);
  or (_36658_, _36657_, _36652_);
  and (_36659_, _08946_, _07886_);
  or (_36660_, _36659_, _36623_);
  or (_36661_, _36660_, _06219_);
  and (_36662_, _36661_, _36658_);
  or (_36663_, _36662_, _06369_);
  and (_36664_, _15353_, _07886_);
  or (_36666_, _36664_, _36623_);
  or (_36667_, _36666_, _07237_);
  and (_36668_, _36667_, _07240_);
  and (_36669_, _36668_, _36663_);
  and (_36670_, _11250_, _07886_);
  or (_36671_, _36670_, _36623_);
  and (_36672_, _36671_, _06536_);
  or (_36673_, _36672_, _36669_);
  and (_36674_, _36673_, _07242_);
  or (_36675_, _36623_, _08247_);
  and (_36677_, _36660_, _06375_);
  and (_36678_, _36677_, _36675_);
  or (_36679_, _36678_, _36674_);
  and (_36680_, _36679_, _07234_);
  and (_36681_, _36631_, _06545_);
  and (_36682_, _36681_, _36675_);
  or (_36683_, _36682_, _06366_);
  or (_36684_, _36683_, _36680_);
  and (_36685_, _15350_, _07886_);
  or (_36686_, _36623_, _09056_);
  or (_36688_, _36686_, _36685_);
  and (_36689_, _36688_, _09061_);
  and (_36690_, _36689_, _36684_);
  nor (_36691_, _11249_, _13951_);
  or (_36692_, _36691_, _36623_);
  and (_36693_, _36692_, _06528_);
  or (_36694_, _36693_, _36690_);
  and (_36695_, _36694_, _06926_);
  and (_36696_, _36628_, _06568_);
  or (_36697_, _36696_, _06278_);
  or (_36699_, _36697_, _36695_);
  and (_36700_, _15532_, _07886_);
  or (_36701_, _36623_, _06279_);
  or (_36702_, _36701_, _36700_);
  and (_36703_, _36702_, _01347_);
  and (_36704_, _36703_, _36699_);
  or (_36705_, _36704_, _36622_);
  and (_43335_, _36705_, _42618_);
  and (_36706_, _01351_, \oc8051_golden_model_1.SBUF [6]);
  and (_36707_, _13951_, \oc8051_golden_model_1.SBUF [6]);
  and (_36709_, _15554_, _07886_);
  or (_36710_, _36709_, _36707_);
  or (_36711_, _36710_, _07151_);
  and (_36712_, _07886_, \oc8051_golden_model_1.ACC [6]);
  or (_36713_, _36712_, _36707_);
  and (_36714_, _36713_, _07141_);
  and (_36715_, _07142_, \oc8051_golden_model_1.SBUF [6]);
  or (_36716_, _36715_, _06341_);
  or (_36717_, _36716_, _36714_);
  and (_36718_, _36717_, _07166_);
  and (_36720_, _36718_, _36711_);
  nor (_36721_, _08142_, _13951_);
  or (_36722_, _36721_, _36707_);
  and (_36723_, _36722_, _06461_);
  or (_36724_, _36723_, _36720_);
  and (_36725_, _36724_, _06465_);
  and (_36726_, _36713_, _06464_);
  or (_36727_, _36726_, _10080_);
  or (_36728_, _36727_, _36725_);
  or (_36729_, _36722_, _07215_);
  and (_36731_, _36729_, _36728_);
  or (_36732_, _36731_, _07460_);
  and (_36733_, _09446_, _07886_);
  or (_36734_, _36707_, _07208_);
  or (_36735_, _36734_, _36733_);
  and (_36736_, _36735_, _05982_);
  and (_36737_, _36736_, _36732_);
  and (_36738_, _15657_, _07886_);
  or (_36739_, _36738_, _36707_);
  and (_36740_, _36739_, _10094_);
  or (_36742_, _36740_, _06218_);
  or (_36743_, _36742_, _36737_);
  and (_36744_, _15664_, _07886_);
  or (_36745_, _36744_, _36707_);
  or (_36746_, _36745_, _06219_);
  and (_36747_, _36746_, _36743_);
  or (_36748_, _36747_, _06369_);
  and (_36749_, _15549_, _07886_);
  or (_36750_, _36749_, _36707_);
  or (_36751_, _36750_, _07237_);
  and (_36753_, _36751_, _07240_);
  and (_36754_, _36753_, _36748_);
  and (_36755_, _11247_, _07886_);
  or (_36756_, _36755_, _36707_);
  and (_36757_, _36756_, _06536_);
  or (_36758_, _36757_, _36754_);
  and (_36759_, _36758_, _07242_);
  or (_36760_, _36707_, _08145_);
  and (_36761_, _36745_, _06375_);
  and (_36762_, _36761_, _36760_);
  or (_36764_, _36762_, _36759_);
  and (_36765_, _36764_, _07234_);
  and (_36766_, _36713_, _06545_);
  and (_36767_, _36766_, _36760_);
  or (_36768_, _36767_, _06366_);
  or (_36769_, _36768_, _36765_);
  and (_36770_, _15546_, _07886_);
  or (_36771_, _36707_, _09056_);
  or (_36772_, _36771_, _36770_);
  and (_36773_, _36772_, _09061_);
  and (_36775_, _36773_, _36769_);
  nor (_36776_, _11246_, _13951_);
  or (_36777_, _36776_, _36707_);
  and (_36778_, _36777_, _06528_);
  or (_36779_, _36778_, _36775_);
  and (_36780_, _36779_, _06926_);
  and (_36781_, _36710_, _06568_);
  or (_36782_, _36781_, _06278_);
  or (_36783_, _36782_, _36780_);
  and (_36784_, _15734_, _07886_);
  or (_36786_, _36707_, _06279_);
  or (_36787_, _36786_, _36784_);
  and (_36788_, _36787_, _01347_);
  and (_36789_, _36788_, _36783_);
  or (_36790_, _36789_, _36706_);
  and (_43336_, _36790_, _42618_);
  not (_36791_, \oc8051_golden_model_1.PSW [0]);
  nor (_36792_, _01347_, _36791_);
  nand (_36793_, _11263_, _07935_);
  nor (_36794_, _07935_, _36791_);
  nor (_36796_, _36794_, _07234_);
  nand (_36797_, _36796_, _36793_);
  and (_36798_, _07935_, _07133_);
  or (_36799_, _36798_, _36794_);
  or (_36800_, _36799_, _07215_);
  nor (_36801_, _08390_, _14045_);
  or (_36802_, _36801_, _36794_);
  or (_36803_, _36802_, _07151_);
  and (_36804_, _07935_, \oc8051_golden_model_1.ACC [0]);
  or (_36805_, _36804_, _36794_);
  and (_36807_, _36805_, _07141_);
  nor (_36808_, _07141_, _36791_);
  or (_36809_, _36808_, _06341_);
  or (_36810_, _36809_, _36807_);
  and (_36811_, _36810_, _06273_);
  and (_36812_, _36811_, _36803_);
  nor (_36813_, _08630_, _36791_);
  and (_36814_, _14382_, _08630_);
  or (_36815_, _36814_, _36813_);
  and (_36816_, _36815_, _06272_);
  or (_36818_, _36816_, _36812_);
  and (_36819_, _36818_, _07166_);
  and (_36820_, _36799_, _06461_);
  or (_36821_, _36820_, _06464_);
  or (_36822_, _36821_, _36819_);
  or (_36823_, _36805_, _06465_);
  and (_36824_, _36823_, _06269_);
  and (_36825_, _36824_, _36822_);
  and (_36826_, _36794_, _06268_);
  or (_36827_, _36826_, _06261_);
  or (_36829_, _36827_, _36825_);
  or (_36830_, _36802_, _06262_);
  and (_36831_, _36830_, _06258_);
  and (_36832_, _36831_, _36829_);
  and (_36833_, _14413_, _08630_);
  or (_36834_, _36833_, _36813_);
  and (_36835_, _36834_, _06257_);
  or (_36836_, _36835_, _10080_);
  or (_36837_, _36836_, _36832_);
  and (_36838_, _36837_, _36800_);
  or (_36840_, _36838_, _07460_);
  and (_36841_, _09392_, _07935_);
  or (_36842_, _36794_, _07208_);
  or (_36843_, _36842_, _36841_);
  and (_36844_, _36843_, _36840_);
  or (_36845_, _36844_, _10094_);
  and (_36846_, _14467_, _07935_);
  or (_36847_, _36794_, _05982_);
  or (_36848_, _36847_, _36846_);
  and (_36849_, _36848_, _06219_);
  and (_36851_, _36849_, _36845_);
  and (_36852_, _07935_, _08954_);
  or (_36853_, _36852_, _36794_);
  and (_36854_, _36853_, _06218_);
  or (_36855_, _36854_, _06369_);
  or (_36856_, _36855_, _36851_);
  and (_36857_, _14366_, _07935_);
  or (_36858_, _36857_, _36794_);
  or (_36859_, _36858_, _07237_);
  and (_36860_, _36859_, _07240_);
  and (_36862_, _36860_, _36856_);
  nor (_36863_, _12580_, _14045_);
  or (_36864_, _36863_, _36794_);
  and (_36865_, _36793_, _06536_);
  and (_36866_, _36865_, _36864_);
  or (_36867_, _36866_, _36862_);
  and (_36868_, _36867_, _07242_);
  nand (_36869_, _36853_, _06375_);
  nor (_36870_, _36869_, _36801_);
  or (_36871_, _36870_, _06545_);
  or (_36872_, _36871_, _36868_);
  and (_36873_, _36872_, _36797_);
  or (_36874_, _36873_, _06366_);
  and (_36875_, _14363_, _07935_);
  or (_36876_, _36794_, _09056_);
  or (_36877_, _36876_, _36875_);
  and (_36878_, _36877_, _09061_);
  and (_36879_, _36878_, _36874_);
  and (_36880_, _36864_, _06528_);
  or (_36881_, _36880_, _06568_);
  or (_36883_, _36881_, _36879_);
  or (_36884_, _36802_, _06926_);
  and (_36885_, _36884_, _36883_);
  or (_36886_, _36885_, _05927_);
  or (_36887_, _36794_, _05928_);
  and (_36888_, _36887_, _36886_);
  or (_36889_, _36888_, _06278_);
  or (_36890_, _36802_, _06279_);
  and (_36891_, _36890_, _01347_);
  and (_36892_, _36891_, _36889_);
  or (_36894_, _36892_, _36792_);
  and (_43338_, _36894_, _42618_);
  not (_36895_, \oc8051_golden_model_1.PSW [1]);
  nor (_36896_, _01347_, _36895_);
  nor (_36897_, _07935_, _36895_);
  nor (_36898_, _11261_, _14045_);
  or (_36899_, _36898_, _36897_);
  or (_36900_, _36899_, _09061_);
  nor (_36901_, _14045_, _07357_);
  or (_36902_, _36901_, _36897_);
  or (_36904_, _36902_, _07215_);
  and (_36905_, _36902_, _06461_);
  nor (_36906_, _08630_, _36895_);
  and (_36907_, _14557_, _08630_);
  or (_36908_, _36907_, _36906_);
  or (_36909_, _36908_, _06273_);
  or (_36910_, _07935_, \oc8051_golden_model_1.PSW [1]);
  and (_36911_, _14562_, _07935_);
  not (_36912_, _36911_);
  and (_36913_, _36912_, _36910_);
  and (_36915_, _36913_, _06341_);
  nor (_36916_, _07141_, _36895_);
  and (_36917_, _07935_, \oc8051_golden_model_1.ACC [1]);
  or (_36918_, _36917_, _36897_);
  and (_36919_, _36918_, _07141_);
  or (_36920_, _36919_, _36916_);
  and (_36921_, _36920_, _07151_);
  or (_36922_, _36921_, _06272_);
  or (_36923_, _36922_, _36915_);
  and (_36924_, _36923_, _36909_);
  and (_36926_, _36924_, _07166_);
  or (_36927_, _36926_, _36905_);
  or (_36928_, _36927_, _06464_);
  or (_36929_, _36918_, _06465_);
  and (_36930_, _36929_, _06269_);
  and (_36931_, _36930_, _36928_);
  and (_36932_, _14560_, _08630_);
  or (_36933_, _36932_, _36906_);
  and (_36934_, _36933_, _06268_);
  or (_36935_, _36934_, _06261_);
  or (_36937_, _36935_, _36931_);
  or (_36938_, _36906_, _14556_);
  and (_36939_, _36938_, _36908_);
  or (_36940_, _36939_, _06262_);
  and (_36941_, _36940_, _06258_);
  and (_36942_, _36941_, _36937_);
  or (_36943_, _36906_, _14597_);
  and (_36944_, _36943_, _06257_);
  and (_36945_, _36944_, _36908_);
  or (_36946_, _36945_, _10080_);
  or (_36948_, _36946_, _36942_);
  and (_36949_, _36948_, _36904_);
  or (_36950_, _36949_, _07460_);
  and (_36951_, _09451_, _07935_);
  or (_36952_, _36897_, _07208_);
  or (_36953_, _36952_, _36951_);
  and (_36954_, _36953_, _05982_);
  and (_36955_, _36954_, _36950_);
  or (_36956_, _14653_, _14045_);
  and (_36957_, _36910_, _10094_);
  and (_36959_, _36957_, _36956_);
  or (_36960_, _36959_, _36955_);
  and (_36961_, _36960_, _06219_);
  nand (_36962_, _07935_, _07038_);
  and (_36963_, _36910_, _06218_);
  and (_36964_, _36963_, _36962_);
  or (_36965_, _36964_, _36961_);
  and (_36966_, _36965_, _07237_);
  or (_36967_, _14668_, _14045_);
  and (_36968_, _36910_, _06369_);
  and (_36970_, _36968_, _36967_);
  or (_36971_, _36970_, _06536_);
  or (_36972_, _36971_, _36966_);
  nand (_36973_, _11260_, _07935_);
  and (_36974_, _36973_, _36899_);
  or (_36975_, _36974_, _07240_);
  and (_36976_, _36975_, _07242_);
  and (_36977_, _36976_, _36972_);
  or (_36978_, _14666_, _14045_);
  and (_36979_, _36910_, _06375_);
  and (_36981_, _36979_, _36978_);
  or (_36982_, _36981_, _06545_);
  or (_36983_, _36982_, _36977_);
  nor (_36984_, _36897_, _07234_);
  nand (_36985_, _36984_, _36973_);
  and (_36986_, _36985_, _09056_);
  and (_36987_, _36986_, _36983_);
  or (_36988_, _36962_, _08341_);
  and (_36989_, _36910_, _06366_);
  and (_36990_, _36989_, _36988_);
  or (_36992_, _36990_, _06528_);
  or (_36993_, _36992_, _36987_);
  and (_36994_, _36993_, _36900_);
  or (_36995_, _36994_, _06568_);
  or (_36996_, _36913_, _06926_);
  and (_36997_, _36996_, _05928_);
  and (_36998_, _36997_, _36995_);
  and (_36999_, _36933_, _05927_);
  or (_37000_, _36999_, _06278_);
  or (_37001_, _37000_, _36998_);
  or (_37003_, _36897_, _06279_);
  or (_37004_, _37003_, _36911_);
  and (_37005_, _37004_, _01347_);
  and (_37006_, _37005_, _37001_);
  or (_37007_, _37006_, _36896_);
  and (_43339_, _37007_, _42618_);
  and (_37008_, _01351_, \oc8051_golden_model_1.PSW [2]);
  not (_37009_, _10960_);
  and (_37010_, _11319_, _37009_);
  or (_37011_, _37010_, _14336_);
  nand (_37013_, _37011_, _06926_);
  not (_37014_, _10499_);
  nand (_37015_, _11236_, _37014_);
  or (_37016_, _11236_, _10498_);
  and (_37017_, _37016_, _37015_);
  or (_37018_, _37017_, _17800_);
  not (_37019_, _11035_);
  nand (_37020_, _11062_, \oc8051_golden_model_1.ACC [7]);
  nand (_37021_, _37020_, _10666_);
  not (_37022_, _10669_);
  and (_37024_, _11062_, _37022_);
  nor (_37025_, _37024_, _11064_);
  or (_37026_, _37025_, _10666_);
  and (_37027_, _37026_, _37021_);
  or (_37028_, _37027_, _37019_);
  and (_37029_, _14045_, \oc8051_golden_model_1.PSW [2]);
  nor (_37030_, _14045_, _07776_);
  or (_37031_, _37030_, _37029_);
  or (_37032_, _37031_, _07215_);
  and (_37033_, _14234_, _10522_);
  nor (_37035_, _14234_, _10522_);
  or (_37036_, _37035_, _37033_);
  or (_37037_, _37036_, _10581_);
  nand (_37038_, _37036_, _10581_);
  and (_37039_, _37038_, _37037_);
  and (_37040_, _37039_, _10516_);
  nor (_37041_, _10596_, \oc8051_golden_model_1.ACC [7]);
  nor (_37042_, _10595_, _37014_);
  nor (_37043_, _37042_, _37041_);
  not (_37044_, _37043_);
  or (_37046_, _37044_, _14053_);
  nand (_37047_, _37044_, _14053_);
  and (_37048_, _37047_, _37046_);
  and (_37049_, _37048_, _10654_);
  nor (_37050_, _37048_, _10654_);
  or (_37051_, _37050_, _37049_);
  or (_37052_, _37051_, _10588_);
  and (_37053_, _14209_, _10665_);
  nor (_37054_, _14209_, _10665_);
  or (_37055_, _37054_, _37053_);
  or (_37057_, _37055_, _10724_);
  nand (_37058_, _37055_, _10724_);
  and (_37059_, _37058_, _10737_);
  and (_37060_, _37059_, _37057_);
  or (_37061_, _37031_, _07166_);
  and (_37062_, _14770_, _07935_);
  or (_37063_, _37062_, _37029_);
  or (_37064_, _37063_, _07151_);
  and (_37065_, _07935_, \oc8051_golden_model_1.ACC [2]);
  or (_37066_, _37065_, _37029_);
  and (_37068_, _37066_, _07141_);
  and (_37069_, _07142_, \oc8051_golden_model_1.PSW [2]);
  or (_37070_, _37069_, _06341_);
  or (_37071_, _37070_, _37068_);
  and (_37072_, _37071_, _06273_);
  and (_37073_, _37072_, _37064_);
  not (_37074_, _08630_);
  and (_37075_, _37074_, \oc8051_golden_model_1.PSW [2]);
  and (_37076_, _14774_, _08630_);
  or (_37077_, _37076_, _37075_);
  and (_37079_, _37077_, _06272_);
  or (_37080_, _37079_, _06461_);
  or (_37081_, _37080_, _37073_);
  and (_37082_, _37081_, _37061_);
  or (_37083_, _37082_, _06464_);
  or (_37084_, _37066_, _06465_);
  and (_37085_, _37084_, _06269_);
  and (_37086_, _37085_, _37083_);
  and (_37087_, _14756_, _08630_);
  or (_37088_, _37087_, _37075_);
  and (_37090_, _37088_, _06268_);
  or (_37091_, _37090_, _06261_);
  or (_37092_, _37091_, _37086_);
  and (_37093_, _37076_, _14789_);
  or (_37094_, _37075_, _06262_);
  or (_37095_, _37094_, _37093_);
  and (_37096_, _37095_, _37092_);
  or (_37097_, _37096_, _09531_);
  or (_37098_, _16582_, _16472_);
  or (_37099_, _37098_, _16694_);
  or (_37101_, _37099_, _16814_);
  or (_37102_, _37101_, _16931_);
  or (_37103_, _37102_, _17045_);
  or (_37104_, _37103_, _17165_);
  or (_37105_, _37104_, _10076_);
  and (_37106_, _37105_, _10735_);
  and (_37107_, _37106_, _37097_);
  or (_37108_, _37107_, _10656_);
  or (_37109_, _37108_, _37060_);
  and (_37110_, _37109_, _06517_);
  and (_37112_, _37110_, _37052_);
  nor (_37113_, _10840_, _14329_);
  nor (_37114_, _10841_, \oc8051_golden_model_1.ACC [7]);
  nor (_37115_, _37114_, _37113_);
  not (_37116_, _37115_);
  or (_37117_, _37116_, _14223_);
  nand (_37118_, _37116_, _14223_);
  and (_37119_, _37118_, _37117_);
  and (_37120_, _37119_, _10898_);
  nor (_37121_, _37119_, _10898_);
  or (_37123_, _37121_, _37120_);
  and (_37124_, _37123_, _06512_);
  or (_37125_, _37124_, _37112_);
  and (_37126_, _37125_, _10517_);
  or (_37127_, _37126_, _37040_);
  and (_37128_, _37127_, _06258_);
  and (_37129_, _14804_, _08630_);
  or (_37130_, _37129_, _37075_);
  and (_37131_, _37130_, _06257_);
  or (_37132_, _37131_, _10080_);
  or (_37134_, _37132_, _37128_);
  and (_37135_, _37134_, _37032_);
  or (_37136_, _37135_, _07460_);
  and (_37137_, _09450_, _07935_);
  or (_37138_, _37029_, _07208_);
  or (_37139_, _37138_, _37137_);
  and (_37140_, _37139_, _05982_);
  and (_37141_, _37140_, _37136_);
  and (_37142_, _14859_, _07935_);
  or (_37143_, _37142_, _37029_);
  and (_37145_, _37143_, _10094_);
  or (_37146_, _37145_, _10093_);
  or (_37147_, _37146_, _37141_);
  nand (_37148_, _10113_, _10106_);
  nand (_37149_, _37148_, _10093_);
  and (_37150_, _37149_, _37147_);
  and (_37151_, _37150_, _06219_);
  and (_37152_, _07935_, _08973_);
  or (_37153_, _37152_, _37029_);
  and (_37154_, _37153_, _06218_);
  or (_37156_, _37154_, _06369_);
  or (_37157_, _37156_, _37151_);
  and (_37158_, _14751_, _07935_);
  or (_37159_, _37158_, _37029_);
  or (_37160_, _37159_, _07237_);
  and (_37161_, _37160_, _07240_);
  and (_37162_, _37161_, _37157_);
  and (_37163_, _11259_, _07935_);
  or (_37164_, _37163_, _37029_);
  and (_37165_, _37164_, _06536_);
  or (_37167_, _37165_, _37162_);
  and (_37168_, _37167_, _07242_);
  or (_37169_, _37029_, _08440_);
  and (_37170_, _37153_, _06375_);
  and (_37171_, _37170_, _37169_);
  or (_37172_, _37171_, _37168_);
  and (_37173_, _37172_, _07234_);
  and (_37174_, _37066_, _06545_);
  and (_37175_, _37174_, _37169_);
  or (_37176_, _37175_, _06366_);
  or (_37178_, _37176_, _37173_);
  and (_37179_, _14748_, _07935_);
  or (_37180_, _37179_, _37029_);
  or (_37181_, _37180_, _09056_);
  and (_37182_, _37181_, _09061_);
  and (_37183_, _37182_, _37178_);
  nor (_37184_, _11258_, _14045_);
  or (_37185_, _37184_, _37029_);
  and (_37186_, _37185_, _06528_);
  or (_37187_, _37186_, _11035_);
  or (_37189_, _37187_, _37183_);
  and (_37190_, _37189_, _37028_);
  or (_37191_, _37190_, _11036_);
  not (_37192_, _11036_);
  or (_37193_, _37027_, _37192_);
  and (_37194_, _37193_, _11069_);
  and (_37195_, _37194_, _37191_);
  nor (_37196_, _37044_, _14293_);
  nor (_37197_, _37196_, _37042_);
  and (_37198_, _37197_, _11093_);
  and (_37200_, _37042_, _11090_);
  or (_37201_, _37200_, _37198_);
  and (_37202_, _37201_, _11041_);
  or (_37203_, _37202_, _14297_);
  or (_37204_, _37203_, _37195_);
  nor (_37205_, _37116_, _14299_);
  nor (_37206_, _37205_, _37113_);
  and (_37207_, _37206_, _11121_);
  and (_37208_, _37113_, _11118_);
  or (_37209_, _37208_, _37207_);
  or (_37211_, _37209_, _06541_);
  nor (_37212_, _10521_, _37009_);
  nor (_37213_, _10523_, \oc8051_golden_model_1.ACC [7]);
  nor (_37214_, _37213_, _14305_);
  nor (_37215_, _37214_, _37212_);
  and (_37216_, _37215_, _11149_);
  and (_37217_, _37212_, _11146_);
  or (_37218_, _37217_, _37216_);
  or (_37219_, _37218_, _11127_);
  and (_37220_, _37219_, _11157_);
  and (_37222_, _37220_, _37211_);
  and (_37223_, _37222_, _37204_);
  or (_37224_, _11193_, _10494_);
  nor (_37225_, _14315_, _11192_);
  nor (_37226_, _37225_, _11157_);
  and (_37227_, _37226_, _37224_);
  or (_37228_, _37227_, _11200_);
  or (_37229_, _37228_, _37223_);
  and (_37230_, _37229_, _37018_);
  or (_37231_, _37230_, _11199_);
  or (_37233_, _37017_, _18067_);
  and (_37234_, _37233_, _13012_);
  and (_37235_, _37234_, _37231_);
  or (_37236_, _11277_, _08573_);
  and (_37237_, _37236_, _14331_);
  or (_37238_, _37237_, _37235_);
  or (_37239_, _37238_, _37013_);
  or (_37240_, _37063_, _06926_);
  and (_37241_, _37240_, _05928_);
  and (_37242_, _37241_, _37239_);
  and (_37244_, _37088_, _05927_);
  or (_37245_, _37244_, _06278_);
  or (_37246_, _37245_, _37242_);
  and (_37247_, _14926_, _07935_);
  or (_37248_, _37029_, _06279_);
  or (_37249_, _37248_, _37247_);
  and (_37250_, _37249_, _01347_);
  and (_37251_, _37250_, _37246_);
  or (_37252_, _37251_, _37008_);
  and (_43340_, _37252_, _42618_);
  nor (_37254_, _01347_, _07615_);
  nor (_37255_, _07935_, _07615_);
  nor (_37256_, _14045_, _07594_);
  or (_37257_, _37256_, _37255_);
  or (_37258_, _37257_, _07215_);
  and (_37259_, _14953_, _07935_);
  or (_37260_, _37259_, _37255_);
  or (_37261_, _37260_, _07151_);
  and (_37262_, _07935_, \oc8051_golden_model_1.ACC [3]);
  or (_37263_, _37262_, _37255_);
  and (_37265_, _37263_, _07141_);
  nor (_37266_, _07141_, _07615_);
  or (_37267_, _37266_, _06341_);
  or (_37268_, _37267_, _37265_);
  and (_37269_, _37268_, _06273_);
  and (_37270_, _37269_, _37261_);
  nor (_37271_, _08630_, _07615_);
  and (_37272_, _14950_, _08630_);
  or (_37273_, _37272_, _37271_);
  and (_37274_, _37273_, _06272_);
  or (_37276_, _37274_, _06461_);
  or (_37277_, _37276_, _37270_);
  or (_37278_, _37257_, _07166_);
  and (_37279_, _37278_, _37277_);
  or (_37280_, _37279_, _06464_);
  or (_37281_, _37263_, _06465_);
  and (_37282_, _37281_, _06269_);
  and (_37283_, _37282_, _37280_);
  and (_37284_, _14948_, _08630_);
  or (_37285_, _37284_, _37271_);
  and (_37287_, _37285_, _06268_);
  or (_37288_, _37287_, _06261_);
  or (_37289_, _37288_, _37283_);
  or (_37290_, _37271_, _14979_);
  and (_37291_, _37290_, _37273_);
  or (_37292_, _37291_, _06262_);
  and (_37293_, _37292_, _06258_);
  and (_37294_, _37293_, _37289_);
  or (_37295_, _37271_, _14992_);
  and (_37296_, _37295_, _06257_);
  and (_37298_, _37296_, _37273_);
  or (_37299_, _37298_, _10080_);
  or (_37300_, _37299_, _37294_);
  and (_37301_, _37300_, _37258_);
  or (_37302_, _37301_, _07460_);
  and (_37303_, _09449_, _07935_);
  or (_37304_, _37255_, _07208_);
  or (_37305_, _37304_, _37303_);
  and (_37306_, _37305_, _05982_);
  and (_37307_, _37306_, _37302_);
  and (_37309_, _15048_, _07935_);
  or (_37310_, _37309_, _37255_);
  and (_37311_, _37310_, _10094_);
  or (_37312_, _37311_, _06218_);
  or (_37313_, _37312_, _37307_);
  and (_37314_, _07935_, _08930_);
  or (_37315_, _37314_, _37255_);
  or (_37316_, _37315_, _06219_);
  and (_37317_, _37316_, _37313_);
  or (_37318_, _37317_, _06369_);
  and (_37320_, _14943_, _07935_);
  or (_37321_, _37320_, _37255_);
  or (_37322_, _37321_, _07237_);
  and (_37323_, _37322_, _07240_);
  and (_37324_, _37323_, _37318_);
  and (_37325_, _12577_, _07935_);
  or (_37326_, _37325_, _37255_);
  and (_37327_, _37326_, _06536_);
  or (_37328_, _37327_, _37324_);
  and (_37329_, _37328_, _07242_);
  or (_37331_, _37255_, _08292_);
  and (_37332_, _37315_, _06375_);
  and (_37333_, _37332_, _37331_);
  or (_37334_, _37333_, _37329_);
  and (_37335_, _37334_, _07234_);
  and (_37336_, _37263_, _06545_);
  and (_37337_, _37336_, _37331_);
  or (_37338_, _37337_, _06366_);
  or (_37339_, _37338_, _37335_);
  and (_37340_, _14940_, _07935_);
  or (_37342_, _37255_, _09056_);
  or (_37343_, _37342_, _37340_);
  and (_37344_, _37343_, _09061_);
  and (_37345_, _37344_, _37339_);
  nor (_37346_, _11256_, _14045_);
  or (_37347_, _37346_, _37255_);
  and (_37348_, _37347_, _06528_);
  or (_37349_, _37348_, _06568_);
  or (_37350_, _37349_, _37345_);
  or (_37351_, _37260_, _06926_);
  and (_37353_, _37351_, _05928_);
  and (_37354_, _37353_, _37350_);
  and (_37355_, _37285_, _05927_);
  or (_37356_, _37355_, _06278_);
  or (_37357_, _37356_, _37354_);
  and (_37358_, _15128_, _07935_);
  or (_37359_, _37255_, _06279_);
  or (_37360_, _37359_, _37358_);
  and (_37361_, _37360_, _01347_);
  and (_37362_, _37361_, _37357_);
  or (_37364_, _37362_, _37254_);
  and (_43341_, _37364_, _42618_);
  and (_37365_, _01351_, \oc8051_golden_model_1.PSW [4]);
  and (_37366_, _14045_, \oc8051_golden_model_1.PSW [4]);
  nor (_37367_, _08541_, _14045_);
  or (_37368_, _37367_, _37366_);
  or (_37369_, _37368_, _07215_);
  and (_37370_, _37074_, \oc8051_golden_model_1.PSW [4]);
  and (_37371_, _15176_, _08630_);
  or (_37372_, _37371_, _37370_);
  and (_37374_, _37372_, _06268_);
  and (_37375_, _15162_, _07935_);
  or (_37376_, _37375_, _37366_);
  or (_37377_, _37376_, _07151_);
  and (_37378_, _07935_, \oc8051_golden_model_1.ACC [4]);
  or (_37379_, _37378_, _37366_);
  and (_37380_, _37379_, _07141_);
  and (_37381_, _07142_, \oc8051_golden_model_1.PSW [4]);
  or (_37382_, _37381_, _06341_);
  or (_37383_, _37382_, _37380_);
  and (_37385_, _37383_, _06273_);
  and (_37386_, _37385_, _37377_);
  and (_37387_, _15166_, _08630_);
  or (_37388_, _37387_, _37370_);
  and (_37389_, _37388_, _06272_);
  or (_37390_, _37389_, _06461_);
  or (_37391_, _37390_, _37386_);
  or (_37392_, _37368_, _07166_);
  and (_37393_, _37392_, _37391_);
  or (_37394_, _37393_, _06464_);
  or (_37396_, _37379_, _06465_);
  and (_37397_, _37396_, _06269_);
  and (_37398_, _37397_, _37394_);
  or (_37399_, _37398_, _37374_);
  and (_37400_, _37399_, _06262_);
  or (_37401_, _37370_, _15183_);
  and (_37402_, _37401_, _06261_);
  and (_37403_, _37402_, _37388_);
  or (_37404_, _37403_, _37400_);
  and (_37405_, _37404_, _06258_);
  and (_37407_, _15200_, _08630_);
  or (_37408_, _37407_, _37370_);
  and (_37409_, _37408_, _06257_);
  or (_37410_, _37409_, _10080_);
  or (_37411_, _37410_, _37405_);
  and (_37412_, _37411_, _37369_);
  or (_37413_, _37412_, _07460_);
  and (_37414_, _09448_, _07935_);
  or (_37415_, _37366_, _07208_);
  or (_37416_, _37415_, _37414_);
  and (_37418_, _37416_, _05982_);
  and (_37419_, _37418_, _37413_);
  and (_37420_, _15254_, _07935_);
  or (_37421_, _37420_, _37366_);
  and (_37422_, _37421_, _10094_);
  or (_37423_, _37422_, _06218_);
  or (_37424_, _37423_, _37419_);
  and (_37425_, _08959_, _07935_);
  or (_37426_, _37425_, _37366_);
  or (_37427_, _37426_, _06219_);
  and (_37429_, _37427_, _37424_);
  or (_37430_, _37429_, _06369_);
  and (_37431_, _15269_, _07935_);
  or (_37432_, _37431_, _37366_);
  or (_37433_, _37432_, _07237_);
  and (_37434_, _37433_, _07240_);
  and (_37435_, _37434_, _37430_);
  and (_37436_, _11254_, _07935_);
  or (_37437_, _37436_, _37366_);
  and (_37438_, _37437_, _06536_);
  or (_37440_, _37438_, _37435_);
  and (_37441_, _37440_, _07242_);
  or (_37442_, _37366_, _08544_);
  and (_37443_, _37426_, _06375_);
  and (_37444_, _37443_, _37442_);
  or (_37445_, _37444_, _37441_);
  and (_37446_, _37445_, _07234_);
  and (_37447_, _37379_, _06545_);
  and (_37448_, _37447_, _37442_);
  or (_37449_, _37448_, _06366_);
  or (_37451_, _37449_, _37446_);
  and (_37452_, _15266_, _07935_);
  or (_37453_, _37366_, _09056_);
  or (_37454_, _37453_, _37452_);
  and (_37455_, _37454_, _09061_);
  and (_37456_, _37455_, _37451_);
  nor (_37457_, _11253_, _14045_);
  or (_37458_, _37457_, _37366_);
  and (_37459_, _37458_, _06528_);
  or (_37460_, _37459_, _06568_);
  or (_37462_, _37460_, _37456_);
  or (_37463_, _37376_, _06926_);
  and (_37464_, _37463_, _05928_);
  and (_37465_, _37464_, _37462_);
  and (_37466_, _37372_, _05927_);
  or (_37467_, _37466_, _06278_);
  or (_37468_, _37467_, _37465_);
  and (_37469_, _15329_, _07935_);
  or (_37470_, _37366_, _06279_);
  or (_37471_, _37470_, _37469_);
  and (_37473_, _37471_, _01347_);
  and (_37474_, _37473_, _37468_);
  or (_37475_, _37474_, _37365_);
  and (_43342_, _37475_, _42618_);
  and (_37476_, _01351_, \oc8051_golden_model_1.PSW [5]);
  and (_37477_, _14045_, \oc8051_golden_model_1.PSW [5]);
  and (_37478_, _15358_, _07935_);
  or (_37479_, _37478_, _37477_);
  or (_37480_, _37479_, _07151_);
  and (_37481_, _07935_, \oc8051_golden_model_1.ACC [5]);
  or (_37483_, _37481_, _37477_);
  and (_37484_, _37483_, _07141_);
  and (_37485_, _07142_, \oc8051_golden_model_1.PSW [5]);
  or (_37486_, _37485_, _06341_);
  or (_37487_, _37486_, _37484_);
  and (_37488_, _37487_, _06273_);
  and (_37489_, _37488_, _37480_);
  and (_37490_, _37074_, \oc8051_golden_model_1.PSW [5]);
  and (_37491_, _15372_, _08630_);
  or (_37492_, _37491_, _37490_);
  and (_37494_, _37492_, _06272_);
  or (_37495_, _37494_, _06461_);
  or (_37496_, _37495_, _37489_);
  nor (_37497_, _08244_, _14045_);
  or (_37498_, _37497_, _37477_);
  or (_37499_, _37498_, _07166_);
  and (_37500_, _37499_, _37496_);
  or (_37501_, _37500_, _06464_);
  or (_37502_, _37483_, _06465_);
  and (_37503_, _37502_, _06269_);
  and (_37505_, _37503_, _37501_);
  and (_37506_, _15355_, _08630_);
  or (_37507_, _37506_, _37490_);
  and (_37508_, _37507_, _06268_);
  or (_37509_, _37508_, _06261_);
  or (_37510_, _37509_, _37505_);
  or (_37511_, _37490_, _15387_);
  and (_37512_, _37511_, _37492_);
  or (_37513_, _37512_, _06262_);
  and (_37514_, _37513_, _06258_);
  and (_37516_, _37514_, _37510_);
  or (_37517_, _37490_, _15403_);
  and (_37518_, _37517_, _06257_);
  and (_37519_, _37518_, _37492_);
  or (_37520_, _37519_, _10080_);
  or (_37521_, _37520_, _37516_);
  or (_37522_, _37498_, _07215_);
  and (_37523_, _37522_, _07208_);
  and (_37524_, _37523_, _37521_);
  and (_37525_, _09447_, _07935_);
  or (_37527_, _37525_, _37477_);
  and (_37528_, _37527_, _07460_);
  or (_37529_, _37528_, _10094_);
  or (_37530_, _37529_, _37524_);
  and (_37531_, _15459_, _07935_);
  or (_37532_, _37477_, _05982_);
  or (_37533_, _37532_, _37531_);
  and (_37534_, _37533_, _06219_);
  and (_37535_, _37534_, _37530_);
  and (_37536_, _08946_, _07935_);
  or (_37538_, _37536_, _37477_);
  and (_37539_, _37538_, _06218_);
  or (_37540_, _37539_, _06369_);
  or (_37541_, _37540_, _37535_);
  and (_37542_, _15353_, _07935_);
  or (_37543_, _37542_, _37477_);
  or (_37544_, _37543_, _07237_);
  and (_37545_, _37544_, _07240_);
  and (_37546_, _37545_, _37541_);
  and (_37547_, _11250_, _07935_);
  or (_37549_, _37547_, _37477_);
  and (_37550_, _37549_, _06536_);
  or (_37551_, _37550_, _37546_);
  and (_37552_, _37551_, _07242_);
  or (_37553_, _37477_, _08247_);
  and (_37554_, _37538_, _06375_);
  and (_37555_, _37554_, _37553_);
  or (_37556_, _37555_, _37552_);
  and (_37557_, _37556_, _07234_);
  and (_37558_, _37483_, _06545_);
  and (_37560_, _37558_, _37553_);
  or (_37561_, _37560_, _06366_);
  or (_37562_, _37561_, _37557_);
  and (_37563_, _15350_, _07935_);
  or (_37564_, _37477_, _09056_);
  or (_37565_, _37564_, _37563_);
  and (_37566_, _37565_, _09061_);
  and (_37567_, _37566_, _37562_);
  nor (_37568_, _11249_, _14045_);
  or (_37569_, _37568_, _37477_);
  and (_37571_, _37569_, _06528_);
  or (_37572_, _37571_, _06568_);
  or (_37573_, _37572_, _37567_);
  or (_37574_, _37479_, _06926_);
  and (_37575_, _37574_, _05928_);
  and (_37576_, _37575_, _37573_);
  and (_37577_, _37507_, _05927_);
  or (_37578_, _37577_, _06278_);
  or (_37579_, _37578_, _37576_);
  and (_37580_, _15532_, _07935_);
  or (_37582_, _37477_, _06279_);
  or (_37583_, _37582_, _37580_);
  and (_37584_, _37583_, _01347_);
  and (_37585_, _37584_, _37579_);
  or (_37586_, _37585_, _37476_);
  and (_43344_, _37586_, _42618_);
  nor (_37587_, _01347_, _18157_);
  or (_37588_, _11140_, _10519_);
  and (_37589_, _37588_, _11097_);
  or (_37590_, _11069_, _10592_);
  or (_37592_, _37590_, _11084_);
  not (_37593_, _11033_);
  or (_37594_, _11056_, _10661_);
  or (_37595_, _37594_, _37593_);
  nor (_37596_, _07935_, _18157_);
  nor (_37597_, _08142_, _14045_);
  or (_37598_, _37597_, _37596_);
  or (_37599_, _37598_, _07215_);
  nor (_37600_, _08630_, _18157_);
  and (_37601_, _15570_, _08630_);
  or (_37603_, _37601_, _37600_);
  or (_37604_, _37600_, _15585_);
  and (_37605_, _37604_, _37603_);
  or (_37606_, _37605_, _06262_);
  and (_37607_, _15554_, _07935_);
  or (_37608_, _37607_, _37596_);
  or (_37609_, _37608_, _07151_);
  and (_37610_, _07935_, \oc8051_golden_model_1.ACC [6]);
  or (_37611_, _37610_, _37596_);
  and (_37612_, _37611_, _07141_);
  nor (_37614_, _07141_, _18157_);
  or (_37615_, _37614_, _06341_);
  or (_37616_, _37615_, _37612_);
  and (_37617_, _37616_, _06273_);
  and (_37618_, _37617_, _37609_);
  and (_37619_, _37603_, _06272_);
  or (_37620_, _37619_, _06461_);
  or (_37621_, _37620_, _37618_);
  or (_37622_, _37598_, _07166_);
  and (_37623_, _37622_, _37621_);
  or (_37625_, _37623_, _06464_);
  or (_37626_, _37611_, _06465_);
  and (_37627_, _37626_, _06269_);
  and (_37628_, _37627_, _37625_);
  and (_37629_, _15551_, _08630_);
  or (_37630_, _37629_, _37600_);
  and (_37631_, _37630_, _06268_);
  or (_37632_, _37631_, _06261_);
  or (_37633_, _37632_, _37628_);
  and (_37634_, _37633_, _37606_);
  and (_37636_, _37634_, _10735_);
  or (_37637_, _10661_, _10656_);
  or (_37638_, _37637_, _10717_);
  and (_37639_, _37638_, _26197_);
  or (_37640_, _37639_, _37636_);
  or (_37641_, _10592_, _10588_);
  or (_37642_, _37641_, _10641_);
  and (_37643_, _37642_, _37640_);
  or (_37644_, _37643_, _12644_);
  or (_37645_, _10837_, _06517_);
  or (_37647_, _37645_, _10888_);
  or (_37648_, _10519_, _10517_);
  or (_37649_, _37648_, _10574_);
  and (_37650_, _37649_, _06258_);
  and (_37651_, _37650_, _37647_);
  and (_37652_, _37651_, _37644_);
  and (_37653_, _15602_, _08630_);
  or (_37654_, _37653_, _37600_);
  and (_37655_, _37654_, _06257_);
  or (_37656_, _37655_, _10080_);
  or (_37658_, _37656_, _37652_);
  and (_37659_, _37658_, _37599_);
  or (_37660_, _37659_, _07460_);
  and (_37661_, _09446_, _07935_);
  or (_37662_, _37596_, _07208_);
  or (_37663_, _37662_, _37661_);
  and (_37664_, _37663_, _05982_);
  and (_37665_, _37664_, _37660_);
  and (_37666_, _15657_, _07935_);
  or (_37667_, _37666_, _37596_);
  and (_37669_, _37667_, _10094_);
  or (_37670_, _37669_, _06218_);
  or (_37671_, _37670_, _37665_);
  and (_37672_, _15664_, _07935_);
  or (_37673_, _37672_, _37596_);
  or (_37674_, _37673_, _06219_);
  and (_37675_, _37674_, _37671_);
  or (_37676_, _37675_, _06369_);
  and (_37677_, _15549_, _07935_);
  or (_37678_, _37677_, _37596_);
  or (_37680_, _37678_, _07237_);
  and (_37681_, _37680_, _07240_);
  and (_37682_, _37681_, _37676_);
  and (_37683_, _11247_, _07935_);
  or (_37684_, _37683_, _37596_);
  and (_37685_, _37684_, _06536_);
  or (_37686_, _37685_, _37682_);
  and (_37687_, _37686_, _07242_);
  or (_37688_, _37596_, _08145_);
  and (_37689_, _37673_, _06375_);
  and (_37691_, _37689_, _37688_);
  or (_37692_, _37691_, _37687_);
  and (_37693_, _37692_, _07234_);
  and (_37694_, _37611_, _06545_);
  and (_37695_, _37694_, _37688_);
  or (_37696_, _37695_, _06366_);
  or (_37697_, _37696_, _37693_);
  and (_37698_, _15546_, _07935_);
  or (_37699_, _37698_, _37596_);
  or (_37700_, _37699_, _09056_);
  and (_37702_, _37700_, _37697_);
  or (_37703_, _37702_, _06528_);
  nor (_37704_, _11246_, _14045_);
  or (_37705_, _37704_, _37596_);
  nor (_37706_, _37705_, _09061_);
  nor (_37707_, _37706_, _11034_);
  and (_37708_, _37707_, _37703_);
  and (_37709_, _37594_, _11034_);
  or (_37710_, _37709_, _11033_);
  or (_37711_, _37710_, _37708_);
  and (_37713_, _37711_, _37595_);
  or (_37714_, _37713_, _17504_);
  not (_37715_, _17504_);
  or (_37716_, _37594_, _37715_);
  and (_37717_, _37716_, _17724_);
  and (_37718_, _37717_, _37714_);
  and (_37719_, _37594_, _17723_);
  or (_37720_, _37719_, _11041_);
  or (_37721_, _37720_, _37718_);
  and (_37722_, _37721_, _37592_);
  or (_37724_, _37722_, _06540_);
  or (_37725_, _10837_, _06541_);
  or (_37726_, _37725_, _11112_);
  and (_37727_, _37726_, _11127_);
  and (_37728_, _37727_, _37724_);
  or (_37729_, _37728_, _37589_);
  and (_37730_, _37729_, _11157_);
  and (_37731_, _11186_, _18059_);
  or (_37732_, _37731_, _11201_);
  or (_37733_, _37732_, _37730_);
  or (_37735_, _11230_, _11203_);
  and (_37736_, _37735_, _06285_);
  and (_37737_, _37736_, _37733_);
  and (_37738_, _11270_, _06283_);
  or (_37739_, _37738_, _11243_);
  or (_37740_, _37739_, _37737_);
  or (_37741_, _11313_, _11321_);
  and (_37742_, _37741_, _37740_);
  or (_37743_, _37742_, _06568_);
  or (_37744_, _37608_, _06926_);
  and (_37746_, _37744_, _05928_);
  and (_37747_, _37746_, _37743_);
  and (_37748_, _37630_, _05927_);
  or (_37749_, _37748_, _06278_);
  or (_37750_, _37749_, _37747_);
  and (_37751_, _15734_, _07935_);
  or (_37752_, _37596_, _06279_);
  or (_37753_, _37752_, _37751_);
  and (_37754_, _37753_, _01347_);
  and (_37755_, _37754_, _37750_);
  or (_37757_, _37755_, _37587_);
  and (_43345_, _37757_, _42618_);
  and (_37758_, _05938_, op0_cnst);
  or (_00000_, _37758_, rst);
  and (_37759_, _37758_, _01347_);
  and (_37760_, _25696_, _01960_);
  nor (_37761_, _25696_, _01960_);
  or (_37762_, _37761_, _37760_);
  and (_37763_, _26055_, _01964_);
  nor (_37764_, _26055_, _01964_);
  nand (_37766_, _26747_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  or (_37767_, _26747_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_37768_, _37767_, _37766_);
  nor (_37769_, _27450_, _01979_);
  and (_37770_, _27450_, _01979_);
  or (_37771_, _37770_, _37769_);
  nor (_37772_, _27099_, _01975_);
  nor (_37773_, _26404_, _01968_);
  and (_37774_, _27099_, _01975_);
  or (_37775_, _37774_, _37773_);
  or (_37777_, _37775_, _37772_);
  nor (_37778_, _27805_, _01983_);
  and (_37779_, _28456_, _38291_);
  nor (_37780_, _28456_, _38291_);
  nor (_37781_, _28133_, _38285_);
  and (_37782_, _28133_, _38285_);
  and (_37783_, _29063_, _38281_);
  nor (_37784_, _29063_, _38281_);
  nor (_37785_, _29667_, _38307_);
  or (_37786_, _37785_, _37784_);
  or (_37788_, _37786_, _37783_);
  nor (_37789_, _13073_, _38317_);
  and (_37790_, _13073_, _38317_);
  and (_37791_, _29667_, _38307_);
  and (_37792_, _28759_, _38296_);
  and (_37793_, _25306_, _01956_);
  nor (_37794_, _25306_, _01956_);
  or (_37795_, _37794_, _37793_);
  nor (_37796_, _28759_, _38296_);
  or (_37797_, _37796_, _37795_);
  or (_37799_, _37797_, _37792_);
  and (_37800_, _29366_, _38302_);
  nor (_37801_, _29366_, _38302_);
  or (_37802_, _37801_, _37800_);
  and (_37803_, _29970_, _38312_);
  nor (_37804_, _29970_, _38312_);
  or (_37805_, _37804_, _37803_);
  or (_37806_, _37805_, _37802_);
  or (_37807_, _37806_, _37799_);
  or (_37808_, _37807_, _37791_);
  or (_37810_, _37808_, _37790_);
  or (_37811_, _37810_, _37789_);
  or (_37812_, _37811_, _37788_);
  or (_37813_, _37812_, _37782_);
  or (_37814_, _37813_, _37781_);
  or (_37815_, _37814_, _37780_);
  or (_37816_, _37815_, _37779_);
  or (_37817_, _37816_, _37778_);
  and (_37818_, _26404_, _01968_);
  and (_37819_, _27805_, _01983_);
  or (_37821_, _37819_, _37818_);
  or (_37822_, _37821_, _37817_);
  or (_37823_, _37822_, _37777_);
  or (_37824_, _37823_, _37771_);
  or (_37825_, _37824_, _37768_);
  or (_37826_, _37825_, _37764_);
  or (_37827_, _37826_, _37763_);
  or (_37828_, _37827_, _37762_);
  and (property_invalid_pc, _37828_, _37759_);
  buf (_00543_, _42621_);
  buf (_05076_, _42618_);
  buf (_05127_, _42618_);
  buf (_05179_, _42618_);
  buf (_05230_, _42618_);
  buf (_05282_, _42618_);
  buf (_05334_, _42618_);
  buf (_05385_, _42618_);
  buf (_05437_, _42618_);
  buf (_05488_, _42618_);
  buf (_05540_, _42618_);
  buf (_05591_, _42618_);
  buf (_05644_, _42618_);
  buf (_05697_, _42618_);
  buf (_05750_, _42618_);
  buf (_05803_, _42618_);
  buf (_05856_, _42618_);
  buf (_38745_, _38644_);
  buf (_38747_, _38646_);
  buf (_38760_, _38644_);
  buf (_38761_, _38646_);
  buf (_39074_, _38664_);
  buf (_39075_, _38665_);
  buf (_39076_, _38667_);
  buf (_39077_, _38668_);
  buf (_39078_, _38669_);
  buf (_39079_, _38670_);
  buf (_39080_, _38671_);
  buf (_39081_, _38673_);
  buf (_39082_, _38674_);
  buf (_39084_, _38675_);
  buf (_39085_, _38676_);
  buf (_39086_, _38677_);
  buf (_39087_, _38679_);
  buf (_39088_, _38680_);
  buf (_39140_, _38664_);
  buf (_39141_, _38665_);
  buf (_39142_, _38667_);
  buf (_39143_, _38668_);
  buf (_39144_, _38669_);
  buf (_39145_, _38670_);
  buf (_39146_, _38671_);
  buf (_39147_, _38673_);
  buf (_39148_, _38674_);
  buf (_39150_, _38675_);
  buf (_39151_, _38676_);
  buf (_39152_, _38677_);
  buf (_39153_, _38679_);
  buf (_39154_, _38680_);
  buf (_39685_, _39457_);
  buf (_39845_, _39457_);
  dff (op0_cnst, _00000_);
  dff (\oc8051_gm_cxrom_1.cell0.data [0], _05080_);
  dff (\oc8051_gm_cxrom_1.cell0.data [1], _05083_);
  dff (\oc8051_gm_cxrom_1.cell0.data [2], _05087_);
  dff (\oc8051_gm_cxrom_1.cell0.data [3], _05091_);
  dff (\oc8051_gm_cxrom_1.cell0.data [4], _05095_);
  dff (\oc8051_gm_cxrom_1.cell0.data [5], _05099_);
  dff (\oc8051_gm_cxrom_1.cell0.data [6], _05103_);
  dff (\oc8051_gm_cxrom_1.cell0.data [7], _05073_);
  dff (\oc8051_gm_cxrom_1.cell0.valid , _05076_);
  dff (\oc8051_gm_cxrom_1.cell1.data [0], _05131_);
  dff (\oc8051_gm_cxrom_1.cell1.data [1], _05135_);
  dff (\oc8051_gm_cxrom_1.cell1.data [2], _05139_);
  dff (\oc8051_gm_cxrom_1.cell1.data [3], _05143_);
  dff (\oc8051_gm_cxrom_1.cell1.data [4], _05147_);
  dff (\oc8051_gm_cxrom_1.cell1.data [5], _05151_);
  dff (\oc8051_gm_cxrom_1.cell1.data [6], _05155_);
  dff (\oc8051_gm_cxrom_1.cell1.data [7], _05124_);
  dff (\oc8051_gm_cxrom_1.cell1.valid , _05127_);
  dff (\oc8051_gm_cxrom_1.cell10.data [0], _05595_);
  dff (\oc8051_gm_cxrom_1.cell10.data [1], _05599_);
  dff (\oc8051_gm_cxrom_1.cell10.data [2], _05603_);
  dff (\oc8051_gm_cxrom_1.cell10.data [3], _05607_);
  dff (\oc8051_gm_cxrom_1.cell10.data [4], _05611_);
  dff (\oc8051_gm_cxrom_1.cell10.data [5], _05615_);
  dff (\oc8051_gm_cxrom_1.cell10.data [6], _05619_);
  dff (\oc8051_gm_cxrom_1.cell10.data [7], _05589_);
  dff (\oc8051_gm_cxrom_1.cell10.valid , _05591_);
  dff (\oc8051_gm_cxrom_1.cell11.data [0], _05648_);
  dff (\oc8051_gm_cxrom_1.cell11.data [1], _05652_);
  dff (\oc8051_gm_cxrom_1.cell11.data [2], _05656_);
  dff (\oc8051_gm_cxrom_1.cell11.data [3], _05660_);
  dff (\oc8051_gm_cxrom_1.cell11.data [4], _05664_);
  dff (\oc8051_gm_cxrom_1.cell11.data [5], _05668_);
  dff (\oc8051_gm_cxrom_1.cell11.data [6], _05672_);
  dff (\oc8051_gm_cxrom_1.cell11.data [7], _05641_);
  dff (\oc8051_gm_cxrom_1.cell11.valid , _05644_);
  dff (\oc8051_gm_cxrom_1.cell12.data [0], _05701_);
  dff (\oc8051_gm_cxrom_1.cell12.data [1], _05705_);
  dff (\oc8051_gm_cxrom_1.cell12.data [2], _05709_);
  dff (\oc8051_gm_cxrom_1.cell12.data [3], _05713_);
  dff (\oc8051_gm_cxrom_1.cell12.data [4], _05717_);
  dff (\oc8051_gm_cxrom_1.cell12.data [5], _05721_);
  dff (\oc8051_gm_cxrom_1.cell12.data [6], _05725_);
  dff (\oc8051_gm_cxrom_1.cell12.data [7], _05694_);
  dff (\oc8051_gm_cxrom_1.cell12.valid , _05697_);
  dff (\oc8051_gm_cxrom_1.cell13.data [0], _05754_);
  dff (\oc8051_gm_cxrom_1.cell13.data [1], _05758_);
  dff (\oc8051_gm_cxrom_1.cell13.data [2], _05762_);
  dff (\oc8051_gm_cxrom_1.cell13.data [3], _05766_);
  dff (\oc8051_gm_cxrom_1.cell13.data [4], _05770_);
  dff (\oc8051_gm_cxrom_1.cell13.data [5], _05774_);
  dff (\oc8051_gm_cxrom_1.cell13.data [6], _05778_);
  dff (\oc8051_gm_cxrom_1.cell13.data [7], _05747_);
  dff (\oc8051_gm_cxrom_1.cell13.valid , _05750_);
  dff (\oc8051_gm_cxrom_1.cell14.data [0], _05807_);
  dff (\oc8051_gm_cxrom_1.cell14.data [1], _05811_);
  dff (\oc8051_gm_cxrom_1.cell14.data [2], _05815_);
  dff (\oc8051_gm_cxrom_1.cell14.data [3], _05819_);
  dff (\oc8051_gm_cxrom_1.cell14.data [4], _05823_);
  dff (\oc8051_gm_cxrom_1.cell14.data [5], _05827_);
  dff (\oc8051_gm_cxrom_1.cell14.data [6], _05831_);
  dff (\oc8051_gm_cxrom_1.cell14.data [7], _05800_);
  dff (\oc8051_gm_cxrom_1.cell14.valid , _05803_);
  dff (\oc8051_gm_cxrom_1.cell15.data [0], _05860_);
  dff (\oc8051_gm_cxrom_1.cell15.data [1], _05864_);
  dff (\oc8051_gm_cxrom_1.cell15.data [2], _05868_);
  dff (\oc8051_gm_cxrom_1.cell15.data [3], _05872_);
  dff (\oc8051_gm_cxrom_1.cell15.data [4], _05876_);
  dff (\oc8051_gm_cxrom_1.cell15.data [5], _05880_);
  dff (\oc8051_gm_cxrom_1.cell15.data [6], _05884_);
  dff (\oc8051_gm_cxrom_1.cell15.data [7], _05853_);
  dff (\oc8051_gm_cxrom_1.cell15.valid , _05856_);
  dff (\oc8051_gm_cxrom_1.cell2.data [0], _05183_);
  dff (\oc8051_gm_cxrom_1.cell2.data [1], _05187_);
  dff (\oc8051_gm_cxrom_1.cell2.data [2], _05191_);
  dff (\oc8051_gm_cxrom_1.cell2.data [3], _05194_);
  dff (\oc8051_gm_cxrom_1.cell2.data [4], _05198_);
  dff (\oc8051_gm_cxrom_1.cell2.data [5], _05202_);
  dff (\oc8051_gm_cxrom_1.cell2.data [6], _05206_);
  dff (\oc8051_gm_cxrom_1.cell2.data [7], _05176_);
  dff (\oc8051_gm_cxrom_1.cell2.valid , _05179_);
  dff (\oc8051_gm_cxrom_1.cell3.data [0], _05234_);
  dff (\oc8051_gm_cxrom_1.cell3.data [1], _05238_);
  dff (\oc8051_gm_cxrom_1.cell3.data [2], _05242_);
  dff (\oc8051_gm_cxrom_1.cell3.data [3], _05246_);
  dff (\oc8051_gm_cxrom_1.cell3.data [4], _05250_);
  dff (\oc8051_gm_cxrom_1.cell3.data [5], _05254_);
  dff (\oc8051_gm_cxrom_1.cell3.data [6], _05258_);
  dff (\oc8051_gm_cxrom_1.cell3.data [7], _05227_);
  dff (\oc8051_gm_cxrom_1.cell3.valid , _05230_);
  dff (\oc8051_gm_cxrom_1.cell4.data [0], _05286_);
  dff (\oc8051_gm_cxrom_1.cell4.data [1], _05290_);
  dff (\oc8051_gm_cxrom_1.cell4.data [2], _05294_);
  dff (\oc8051_gm_cxrom_1.cell4.data [3], _05298_);
  dff (\oc8051_gm_cxrom_1.cell4.data [4], _05301_);
  dff (\oc8051_gm_cxrom_1.cell4.data [5], _05305_);
  dff (\oc8051_gm_cxrom_1.cell4.data [6], _05309_);
  dff (\oc8051_gm_cxrom_1.cell4.data [7], _05279_);
  dff (\oc8051_gm_cxrom_1.cell4.valid , _05282_);
  dff (\oc8051_gm_cxrom_1.cell5.data [0], _05337_);
  dff (\oc8051_gm_cxrom_1.cell5.data [1], _05341_);
  dff (\oc8051_gm_cxrom_1.cell5.data [2], _05345_);
  dff (\oc8051_gm_cxrom_1.cell5.data [3], _05349_);
  dff (\oc8051_gm_cxrom_1.cell5.data [4], _05353_);
  dff (\oc8051_gm_cxrom_1.cell5.data [5], _05357_);
  dff (\oc8051_gm_cxrom_1.cell5.data [6], _05361_);
  dff (\oc8051_gm_cxrom_1.cell5.data [7], _05331_);
  dff (\oc8051_gm_cxrom_1.cell5.valid , _05334_);
  dff (\oc8051_gm_cxrom_1.cell6.data [0], _05389_);
  dff (\oc8051_gm_cxrom_1.cell6.data [1], _05393_);
  dff (\oc8051_gm_cxrom_1.cell6.data [2], _05397_);
  dff (\oc8051_gm_cxrom_1.cell6.data [3], _05401_);
  dff (\oc8051_gm_cxrom_1.cell6.data [4], _05405_);
  dff (\oc8051_gm_cxrom_1.cell6.data [5], _05409_);
  dff (\oc8051_gm_cxrom_1.cell6.data [6], _05412_);
  dff (\oc8051_gm_cxrom_1.cell6.data [7], _05382_);
  dff (\oc8051_gm_cxrom_1.cell6.valid , _05385_);
  dff (\oc8051_gm_cxrom_1.cell7.data [0], _05441_);
  dff (\oc8051_gm_cxrom_1.cell7.data [1], _05445_);
  dff (\oc8051_gm_cxrom_1.cell7.data [2], _05448_);
  dff (\oc8051_gm_cxrom_1.cell7.data [3], _05452_);
  dff (\oc8051_gm_cxrom_1.cell7.data [4], _05456_);
  dff (\oc8051_gm_cxrom_1.cell7.data [5], _05460_);
  dff (\oc8051_gm_cxrom_1.cell7.data [6], _05464_);
  dff (\oc8051_gm_cxrom_1.cell7.data [7], _05434_);
  dff (\oc8051_gm_cxrom_1.cell7.valid , _05437_);
  dff (\oc8051_gm_cxrom_1.cell8.data [0], _05492_);
  dff (\oc8051_gm_cxrom_1.cell8.data [1], _05496_);
  dff (\oc8051_gm_cxrom_1.cell8.data [2], _05500_);
  dff (\oc8051_gm_cxrom_1.cell8.data [3], _05504_);
  dff (\oc8051_gm_cxrom_1.cell8.data [4], _05508_);
  dff (\oc8051_gm_cxrom_1.cell8.data [5], _05512_);
  dff (\oc8051_gm_cxrom_1.cell8.data [6], _05516_);
  dff (\oc8051_gm_cxrom_1.cell8.data [7], _05485_);
  dff (\oc8051_gm_cxrom_1.cell8.valid , _05488_);
  dff (\oc8051_gm_cxrom_1.cell9.data [0], _05544_);
  dff (\oc8051_gm_cxrom_1.cell9.data [1], _05548_);
  dff (\oc8051_gm_cxrom_1.cell9.data [2], _05552_);
  dff (\oc8051_gm_cxrom_1.cell9.data [3], _05555_);
  dff (\oc8051_gm_cxrom_1.cell9.data [4], _05559_);
  dff (\oc8051_gm_cxrom_1.cell9.data [5], _05563_);
  dff (\oc8051_gm_cxrom_1.cell9.data [6], _05567_);
  dff (\oc8051_gm_cxrom_1.cell9.data [7], _05537_);
  dff (\oc8051_gm_cxrom_1.cell9.valid , _05540_);
  dff (\oc8051_golden_model_1.IRAM[15] [0], _40795_);
  dff (\oc8051_golden_model_1.IRAM[15] [1], _40796_);
  dff (\oc8051_golden_model_1.IRAM[15] [2], _40797_);
  dff (\oc8051_golden_model_1.IRAM[15] [3], _40799_);
  dff (\oc8051_golden_model_1.IRAM[15] [4], _40800_);
  dff (\oc8051_golden_model_1.IRAM[15] [5], _40801_);
  dff (\oc8051_golden_model_1.IRAM[15] [6], _40802_);
  dff (\oc8051_golden_model_1.IRAM[15] [7], _40572_);
  dff (\oc8051_golden_model_1.IRAM[14] [0], _40783_);
  dff (\oc8051_golden_model_1.IRAM[14] [1], _40784_);
  dff (\oc8051_golden_model_1.IRAM[14] [2], _40785_);
  dff (\oc8051_golden_model_1.IRAM[14] [3], _40787_);
  dff (\oc8051_golden_model_1.IRAM[14] [4], _40788_);
  dff (\oc8051_golden_model_1.IRAM[14] [5], _40789_);
  dff (\oc8051_golden_model_1.IRAM[14] [6], _40790_);
  dff (\oc8051_golden_model_1.IRAM[14] [7], _40791_);
  dff (\oc8051_golden_model_1.IRAM[13] [0], _40771_);
  dff (\oc8051_golden_model_1.IRAM[13] [1], _40772_);
  dff (\oc8051_golden_model_1.IRAM[13] [2], _40773_);
  dff (\oc8051_golden_model_1.IRAM[13] [3], _40774_);
  dff (\oc8051_golden_model_1.IRAM[13] [4], _40776_);
  dff (\oc8051_golden_model_1.IRAM[13] [5], _40777_);
  dff (\oc8051_golden_model_1.IRAM[13] [6], _40778_);
  dff (\oc8051_golden_model_1.IRAM[13] [7], _40779_);
  dff (\oc8051_golden_model_1.IRAM[12] [0], _40759_);
  dff (\oc8051_golden_model_1.IRAM[12] [1], _40760_);
  dff (\oc8051_golden_model_1.IRAM[12] [2], _40761_);
  dff (\oc8051_golden_model_1.IRAM[12] [3], _40762_);
  dff (\oc8051_golden_model_1.IRAM[12] [4], _40764_);
  dff (\oc8051_golden_model_1.IRAM[12] [5], _40765_);
  dff (\oc8051_golden_model_1.IRAM[12] [6], _40766_);
  dff (\oc8051_golden_model_1.IRAM[12] [7], _40767_);
  dff (\oc8051_golden_model_1.IRAM[11] [0], _40746_);
  dff (\oc8051_golden_model_1.IRAM[11] [1], _40748_);
  dff (\oc8051_golden_model_1.IRAM[11] [2], _40749_);
  dff (\oc8051_golden_model_1.IRAM[11] [3], _40750_);
  dff (\oc8051_golden_model_1.IRAM[11] [4], _40751_);
  dff (\oc8051_golden_model_1.IRAM[11] [5], _40752_);
  dff (\oc8051_golden_model_1.IRAM[11] [6], _40754_);
  dff (\oc8051_golden_model_1.IRAM[11] [7], _40755_);
  dff (\oc8051_golden_model_1.IRAM[10] [0], _40734_);
  dff (\oc8051_golden_model_1.IRAM[10] [1], _40736_);
  dff (\oc8051_golden_model_1.IRAM[10] [2], _40737_);
  dff (\oc8051_golden_model_1.IRAM[10] [3], _40738_);
  dff (\oc8051_golden_model_1.IRAM[10] [4], _40739_);
  dff (\oc8051_golden_model_1.IRAM[10] [5], _40740_);
  dff (\oc8051_golden_model_1.IRAM[10] [6], _40742_);
  dff (\oc8051_golden_model_1.IRAM[10] [7], _40743_);
  dff (\oc8051_golden_model_1.IRAM[9] [0], _40723_);
  dff (\oc8051_golden_model_1.IRAM[9] [1], _40724_);
  dff (\oc8051_golden_model_1.IRAM[9] [2], _40726_);
  dff (\oc8051_golden_model_1.IRAM[9] [3], _40727_);
  dff (\oc8051_golden_model_1.IRAM[9] [4], _40728_);
  dff (\oc8051_golden_model_1.IRAM[9] [5], _40729_);
  dff (\oc8051_golden_model_1.IRAM[9] [6], _40730_);
  dff (\oc8051_golden_model_1.IRAM[9] [7], _40732_);
  dff (\oc8051_golden_model_1.IRAM[8] [0], _40711_);
  dff (\oc8051_golden_model_1.IRAM[8] [1], _40712_);
  dff (\oc8051_golden_model_1.IRAM[8] [2], _40714_);
  dff (\oc8051_golden_model_1.IRAM[8] [3], _40715_);
  dff (\oc8051_golden_model_1.IRAM[8] [4], _40716_);
  dff (\oc8051_golden_model_1.IRAM[8] [5], _40717_);
  dff (\oc8051_golden_model_1.IRAM[8] [6], _40718_);
  dff (\oc8051_golden_model_1.IRAM[8] [7], _40720_);
  dff (\oc8051_golden_model_1.IRAM[7] [0], _40698_);
  dff (\oc8051_golden_model_1.IRAM[7] [1], _40700_);
  dff (\oc8051_golden_model_1.IRAM[7] [2], _40701_);
  dff (\oc8051_golden_model_1.IRAM[7] [3], _40702_);
  dff (\oc8051_golden_model_1.IRAM[7] [4], _40703_);
  dff (\oc8051_golden_model_1.IRAM[7] [5], _40704_);
  dff (\oc8051_golden_model_1.IRAM[7] [6], _40706_);
  dff (\oc8051_golden_model_1.IRAM[7] [7], _40707_);
  dff (\oc8051_golden_model_1.IRAM[6] [0], _40685_);
  dff (\oc8051_golden_model_1.IRAM[6] [1], _40688_);
  dff (\oc8051_golden_model_1.IRAM[6] [2], _40689_);
  dff (\oc8051_golden_model_1.IRAM[6] [3], _40690_);
  dff (\oc8051_golden_model_1.IRAM[6] [4], _40691_);
  dff (\oc8051_golden_model_1.IRAM[6] [5], _40692_);
  dff (\oc8051_golden_model_1.IRAM[6] [6], _40694_);
  dff (\oc8051_golden_model_1.IRAM[6] [7], _40695_);
  dff (\oc8051_golden_model_1.IRAM[5] [0], _40673_);
  dff (\oc8051_golden_model_1.IRAM[5] [1], _40674_);
  dff (\oc8051_golden_model_1.IRAM[5] [2], _40677_);
  dff (\oc8051_golden_model_1.IRAM[5] [3], _40678_);
  dff (\oc8051_golden_model_1.IRAM[5] [4], _40679_);
  dff (\oc8051_golden_model_1.IRAM[5] [5], _40680_);
  dff (\oc8051_golden_model_1.IRAM[5] [6], _40681_);
  dff (\oc8051_golden_model_1.IRAM[5] [7], _40683_);
  dff (\oc8051_golden_model_1.IRAM[4] [0], _40662_);
  dff (\oc8051_golden_model_1.IRAM[4] [1], _40663_);
  dff (\oc8051_golden_model_1.IRAM[4] [2], _40665_);
  dff (\oc8051_golden_model_1.IRAM[4] [3], _40666_);
  dff (\oc8051_golden_model_1.IRAM[4] [4], _40667_);
  dff (\oc8051_golden_model_1.IRAM[4] [5], _40668_);
  dff (\oc8051_golden_model_1.IRAM[4] [6], _40669_);
  dff (\oc8051_golden_model_1.IRAM[4] [7], _40671_);
  dff (\oc8051_golden_model_1.IRAM[3] [0], _40649_);
  dff (\oc8051_golden_model_1.IRAM[3] [1], _40651_);
  dff (\oc8051_golden_model_1.IRAM[3] [2], _40652_);
  dff (\oc8051_golden_model_1.IRAM[3] [3], _40653_);
  dff (\oc8051_golden_model_1.IRAM[3] [4], _40654_);
  dff (\oc8051_golden_model_1.IRAM[3] [5], _40655_);
  dff (\oc8051_golden_model_1.IRAM[3] [6], _40657_);
  dff (\oc8051_golden_model_1.IRAM[3] [7], _40658_);
  dff (\oc8051_golden_model_1.IRAM[2] [0], _40637_);
  dff (\oc8051_golden_model_1.IRAM[2] [1], _40638_);
  dff (\oc8051_golden_model_1.IRAM[2] [2], _40640_);
  dff (\oc8051_golden_model_1.IRAM[2] [3], _40641_);
  dff (\oc8051_golden_model_1.IRAM[2] [4], _40642_);
  dff (\oc8051_golden_model_1.IRAM[2] [5], _40643_);
  dff (\oc8051_golden_model_1.IRAM[2] [6], _40644_);
  dff (\oc8051_golden_model_1.IRAM[2] [7], _40646_);
  dff (\oc8051_golden_model_1.IRAM[1] [0], _40623_);
  dff (\oc8051_golden_model_1.IRAM[1] [1], _40626_);
  dff (\oc8051_golden_model_1.IRAM[1] [2], _40627_);
  dff (\oc8051_golden_model_1.IRAM[1] [3], _40628_);
  dff (\oc8051_golden_model_1.IRAM[1] [4], _40629_);
  dff (\oc8051_golden_model_1.IRAM[1] [5], _40630_);
  dff (\oc8051_golden_model_1.IRAM[1] [6], _40632_);
  dff (\oc8051_golden_model_1.IRAM[1] [7], _40633_);
  dff (\oc8051_golden_model_1.B [0], _43153_);
  dff (\oc8051_golden_model_1.B [1], _43154_);
  dff (\oc8051_golden_model_1.B [2], _43155_);
  dff (\oc8051_golden_model_1.B [3], _43156_);
  dff (\oc8051_golden_model_1.B [4], _43157_);
  dff (\oc8051_golden_model_1.B [5], _43159_);
  dff (\oc8051_golden_model_1.B [6], _43160_);
  dff (\oc8051_golden_model_1.B [7], _40573_);
  dff (\oc8051_golden_model_1.ACC [0], _43161_);
  dff (\oc8051_golden_model_1.ACC [1], _43163_);
  dff (\oc8051_golden_model_1.ACC [2], _43164_);
  dff (\oc8051_golden_model_1.ACC [3], _43165_);
  dff (\oc8051_golden_model_1.ACC [4], _43166_);
  dff (\oc8051_golden_model_1.ACC [5], _43167_);
  dff (\oc8051_golden_model_1.ACC [6], _43168_);
  dff (\oc8051_golden_model_1.ACC [7], _40574_);
  dff (\oc8051_golden_model_1.PCON [0], _43170_);
  dff (\oc8051_golden_model_1.PCON [1], _43171_);
  dff (\oc8051_golden_model_1.PCON [2], _43172_);
  dff (\oc8051_golden_model_1.PCON [3], _43173_);
  dff (\oc8051_golden_model_1.PCON [4], _43174_);
  dff (\oc8051_golden_model_1.PCON [5], _43175_);
  dff (\oc8051_golden_model_1.PCON [6], _43176_);
  dff (\oc8051_golden_model_1.PCON [7], _40575_);
  dff (\oc8051_golden_model_1.TMOD [0], _43178_);
  dff (\oc8051_golden_model_1.TMOD [1], _43179_);
  dff (\oc8051_golden_model_1.TMOD [2], _43180_);
  dff (\oc8051_golden_model_1.TMOD [3], _43182_);
  dff (\oc8051_golden_model_1.TMOD [4], _43183_);
  dff (\oc8051_golden_model_1.TMOD [5], _43184_);
  dff (\oc8051_golden_model_1.TMOD [6], _43185_);
  dff (\oc8051_golden_model_1.TMOD [7], _40576_);
  dff (\oc8051_golden_model_1.DPL [0], _43187_);
  dff (\oc8051_golden_model_1.DPL [1], _43188_);
  dff (\oc8051_golden_model_1.DPL [2], _43189_);
  dff (\oc8051_golden_model_1.DPL [3], _43190_);
  dff (\oc8051_golden_model_1.DPL [4], _43191_);
  dff (\oc8051_golden_model_1.DPL [5], _43192_);
  dff (\oc8051_golden_model_1.DPL [6], _43193_);
  dff (\oc8051_golden_model_1.DPL [7], _40577_);
  dff (\oc8051_golden_model_1.DPH [0], _43195_);
  dff (\oc8051_golden_model_1.DPH [1], _43196_);
  dff (\oc8051_golden_model_1.DPH [2], _43197_);
  dff (\oc8051_golden_model_1.DPH [3], _43198_);
  dff (\oc8051_golden_model_1.DPH [4], _43199_);
  dff (\oc8051_golden_model_1.DPH [5], _43200_);
  dff (\oc8051_golden_model_1.DPH [6], _43201_);
  dff (\oc8051_golden_model_1.DPH [7], _40580_);
  dff (\oc8051_golden_model_1.TL1 [0], _43202_);
  dff (\oc8051_golden_model_1.TL1 [1], _43204_);
  dff (\oc8051_golden_model_1.TL1 [2], _43205_);
  dff (\oc8051_golden_model_1.TL1 [3], _43206_);
  dff (\oc8051_golden_model_1.TL1 [4], _43207_);
  dff (\oc8051_golden_model_1.TL1 [5], _43208_);
  dff (\oc8051_golden_model_1.TL1 [6], _43209_);
  dff (\oc8051_golden_model_1.TL1 [7], _40581_);
  dff (\oc8051_golden_model_1.TL0 [0], _43211_);
  dff (\oc8051_golden_model_1.TL0 [1], _43212_);
  dff (\oc8051_golden_model_1.TL0 [2], _43213_);
  dff (\oc8051_golden_model_1.TL0 [3], _43214_);
  dff (\oc8051_golden_model_1.TL0 [4], _43215_);
  dff (\oc8051_golden_model_1.TL0 [5], _43216_);
  dff (\oc8051_golden_model_1.TL0 [6], _43217_);
  dff (\oc8051_golden_model_1.TL0 [7], _40582_);
  dff (\oc8051_golden_model_1.TCON [0], _43219_);
  dff (\oc8051_golden_model_1.TCON [1], _43220_);
  dff (\oc8051_golden_model_1.TCON [2], _43221_);
  dff (\oc8051_golden_model_1.TCON [3], _43223_);
  dff (\oc8051_golden_model_1.TCON [4], _43224_);
  dff (\oc8051_golden_model_1.TCON [5], _43225_);
  dff (\oc8051_golden_model_1.TCON [6], _43226_);
  dff (\oc8051_golden_model_1.TCON [7], _40583_);
  dff (\oc8051_golden_model_1.TH1 [0], _43228_);
  dff (\oc8051_golden_model_1.TH1 [1], _43229_);
  dff (\oc8051_golden_model_1.TH1 [2], _43230_);
  dff (\oc8051_golden_model_1.TH1 [3], _43231_);
  dff (\oc8051_golden_model_1.TH1 [4], _43232_);
  dff (\oc8051_golden_model_1.TH1 [5], _43233_);
  dff (\oc8051_golden_model_1.TH1 [6], _43234_);
  dff (\oc8051_golden_model_1.TH1 [7], _40584_);
  dff (\oc8051_golden_model_1.TH0 [0], _43236_);
  dff (\oc8051_golden_model_1.TH0 [1], _43237_);
  dff (\oc8051_golden_model_1.TH0 [2], _43238_);
  dff (\oc8051_golden_model_1.TH0 [3], _43239_);
  dff (\oc8051_golden_model_1.TH0 [4], _43240_);
  dff (\oc8051_golden_model_1.TH0 [5], _43242_);
  dff (\oc8051_golden_model_1.TH0 [6], _43243_);
  dff (\oc8051_golden_model_1.TH0 [7], _40585_);
  dff (\oc8051_golden_model_1.PC [0], _43245_);
  dff (\oc8051_golden_model_1.PC [1], _43246_);
  dff (\oc8051_golden_model_1.PC [2], _43247_);
  dff (\oc8051_golden_model_1.PC [3], _43249_);
  dff (\oc8051_golden_model_1.PC [4], _43250_);
  dff (\oc8051_golden_model_1.PC [5], _43251_);
  dff (\oc8051_golden_model_1.PC [6], _43252_);
  dff (\oc8051_golden_model_1.PC [7], _43253_);
  dff (\oc8051_golden_model_1.PC [8], _43254_);
  dff (\oc8051_golden_model_1.PC [9], _43255_);
  dff (\oc8051_golden_model_1.PC [10], _43256_);
  dff (\oc8051_golden_model_1.PC [11], _43257_);
  dff (\oc8051_golden_model_1.PC [12], _43258_);
  dff (\oc8051_golden_model_1.PC [13], _43260_);
  dff (\oc8051_golden_model_1.PC [14], _43261_);
  dff (\oc8051_golden_model_1.PC [15], _40586_);
  dff (\oc8051_golden_model_1.P2 [0], _43262_);
  dff (\oc8051_golden_model_1.P2 [1], _43264_);
  dff (\oc8051_golden_model_1.P2 [2], _43265_);
  dff (\oc8051_golden_model_1.P2 [3], _43266_);
  dff (\oc8051_golden_model_1.P2 [4], _43267_);
  dff (\oc8051_golden_model_1.P2 [5], _43268_);
  dff (\oc8051_golden_model_1.P2 [6], _43269_);
  dff (\oc8051_golden_model_1.P2 [7], _40587_);
  dff (\oc8051_golden_model_1.P3 [0], _43271_);
  dff (\oc8051_golden_model_1.P3 [1], _43272_);
  dff (\oc8051_golden_model_1.P3 [2], _43273_);
  dff (\oc8051_golden_model_1.P3 [3], _43274_);
  dff (\oc8051_golden_model_1.P3 [4], _43275_);
  dff (\oc8051_golden_model_1.P3 [5], _43276_);
  dff (\oc8051_golden_model_1.P3 [6], _43277_);
  dff (\oc8051_golden_model_1.P3 [7], _40588_);
  dff (\oc8051_golden_model_1.P0 [0], _43279_);
  dff (\oc8051_golden_model_1.P0 [1], _43280_);
  dff (\oc8051_golden_model_1.P0 [2], _43281_);
  dff (\oc8051_golden_model_1.P0 [3], _43283_);
  dff (\oc8051_golden_model_1.P0 [4], _43284_);
  dff (\oc8051_golden_model_1.P0 [5], _43285_);
  dff (\oc8051_golden_model_1.P0 [6], _43286_);
  dff (\oc8051_golden_model_1.P0 [7], _40589_);
  dff (\oc8051_golden_model_1.P1 [0], _43288_);
  dff (\oc8051_golden_model_1.P1 [1], _43289_);
  dff (\oc8051_golden_model_1.P1 [2], _43290_);
  dff (\oc8051_golden_model_1.P1 [3], _43291_);
  dff (\oc8051_golden_model_1.P1 [4], _43292_);
  dff (\oc8051_golden_model_1.P1 [5], _43293_);
  dff (\oc8051_golden_model_1.P1 [6], _43294_);
  dff (\oc8051_golden_model_1.P1 [7], _40591_);
  dff (\oc8051_golden_model_1.IP [0], _43296_);
  dff (\oc8051_golden_model_1.IP [1], _43297_);
  dff (\oc8051_golden_model_1.IP [2], _43298_);
  dff (\oc8051_golden_model_1.IP [3], _43299_);
  dff (\oc8051_golden_model_1.IP [4], _43300_);
  dff (\oc8051_golden_model_1.IP [5], _43302_);
  dff (\oc8051_golden_model_1.IP [6], _43303_);
  dff (\oc8051_golden_model_1.IP [7], _40592_);
  dff (\oc8051_golden_model_1.IE [0], _43304_);
  dff (\oc8051_golden_model_1.IE [1], _43306_);
  dff (\oc8051_golden_model_1.IE [2], _43307_);
  dff (\oc8051_golden_model_1.IE [3], _43308_);
  dff (\oc8051_golden_model_1.IE [4], _43309_);
  dff (\oc8051_golden_model_1.IE [5], _43310_);
  dff (\oc8051_golden_model_1.IE [6], _43311_);
  dff (\oc8051_golden_model_1.IE [7], _40593_);
  dff (\oc8051_golden_model_1.SCON [0], _43313_);
  dff (\oc8051_golden_model_1.SCON [1], _43314_);
  dff (\oc8051_golden_model_1.SCON [2], _43315_);
  dff (\oc8051_golden_model_1.SCON [3], _43316_);
  dff (\oc8051_golden_model_1.SCON [4], _43317_);
  dff (\oc8051_golden_model_1.SCON [5], _43318_);
  dff (\oc8051_golden_model_1.SCON [6], _43319_);
  dff (\oc8051_golden_model_1.SCON [7], _40594_);
  dff (\oc8051_golden_model_1.SP [0], _43321_);
  dff (\oc8051_golden_model_1.SP [1], _43322_);
  dff (\oc8051_golden_model_1.SP [2], _43323_);
  dff (\oc8051_golden_model_1.SP [3], _43325_);
  dff (\oc8051_golden_model_1.SP [4], _43326_);
  dff (\oc8051_golden_model_1.SP [5], _43327_);
  dff (\oc8051_golden_model_1.SP [6], _43328_);
  dff (\oc8051_golden_model_1.SP [7], _40595_);
  dff (\oc8051_golden_model_1.SBUF [0], _43330_);
  dff (\oc8051_golden_model_1.SBUF [1], _43331_);
  dff (\oc8051_golden_model_1.SBUF [2], _43332_);
  dff (\oc8051_golden_model_1.SBUF [3], _43333_);
  dff (\oc8051_golden_model_1.SBUF [4], _43334_);
  dff (\oc8051_golden_model_1.SBUF [5], _43335_);
  dff (\oc8051_golden_model_1.SBUF [6], _43336_);
  dff (\oc8051_golden_model_1.SBUF [7], _40597_);
  dff (\oc8051_golden_model_1.PSW [0], _43338_);
  dff (\oc8051_golden_model_1.PSW [1], _43339_);
  dff (\oc8051_golden_model_1.PSW [2], _43340_);
  dff (\oc8051_golden_model_1.PSW [3], _43341_);
  dff (\oc8051_golden_model_1.PSW [4], _43342_);
  dff (\oc8051_golden_model_1.PSW [5], _43344_);
  dff (\oc8051_golden_model_1.PSW [6], _43345_);
  dff (\oc8051_golden_model_1.PSW [7], _40598_);
  dff (\oc8051_golden_model_1.IRAM[0] [0], _40612_);
  dff (\oc8051_golden_model_1.IRAM[0] [1], _40613_);
  dff (\oc8051_golden_model_1.IRAM[0] [2], _40614_);
  dff (\oc8051_golden_model_1.IRAM[0] [3], _40615_);
  dff (\oc8051_golden_model_1.IRAM[0] [4], _40616_);
  dff (\oc8051_golden_model_1.IRAM[0] [5], _40618_);
  dff (\oc8051_golden_model_1.IRAM[0] [6], _40619_);
  dff (\oc8051_golden_model_1.IRAM[0] [7], _40620_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _02836_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _02848_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _02870_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _02894_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4], _02916_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5], _00951_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], _02927_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1], _00925_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0], _02940_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1], _02954_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2], _02967_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3], _02981_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4], _02995_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5], _03008_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6], _03022_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7], _00971_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], _02354_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _22124_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0], _02542_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1], _02700_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2], _02882_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3], _03125_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4], _03328_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5], _03527_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6], _03728_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7], _03927_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8], _04023_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9], _04123_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10], _04222_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11], _04321_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12], _04414_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13], _04512_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [14], _04611_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [15], _24283_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [0], _38656_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [1], _38658_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [2], _38659_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [3], _38660_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [4], _38661_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [5], _38662_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [6], _38663_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [7], _38643_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [0], _38664_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [1], _38665_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [2], _38667_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [3], _38668_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [4], _38669_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [5], _38670_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [6], _38671_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [7], _38644_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [0], _38673_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [1], _38674_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [2], _38675_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [3], _38676_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [4], _38677_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [5], _38679_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [6], _38680_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [7], _38646_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _34184_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _34187_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], _09680_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [0], _34189_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [1], _34191_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [2], _09683_);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [0], _34193_);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [1], _09686_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [0], _34195_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [1], _34197_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [2], _34199_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [3], _09689_);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [0], _34201_);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [1], _09692_);
  dff (\oc8051_top_1.oc8051_decoder1.wr , _09695_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], _09754_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], _09756_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], _09659_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [0], _09759_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [1], _09762_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [2], _09662_);
  dff (\oc8051_top_1.oc8051_decoder1.state [0], _09765_);
  dff (\oc8051_top_1.oc8051_decoder1.state [1], _09665_);
  dff (\oc8051_top_1.oc8051_decoder1.op [0], _09768_);
  dff (\oc8051_top_1.oc8051_decoder1.op [1], _09771_);
  dff (\oc8051_top_1.oc8051_decoder1.op [2], _09774_);
  dff (\oc8051_top_1.oc8051_decoder1.op [3], _09777_);
  dff (\oc8051_top_1.oc8051_decoder1.op [4], _09780_);
  dff (\oc8051_top_1.oc8051_decoder1.op [5], _09783_);
  dff (\oc8051_top_1.oc8051_decoder1.op [6], _09786_);
  dff (\oc8051_top_1.oc8051_decoder1.op [7], _09668_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel3 , _09671_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [0], _34182_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [1], _09677_);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [0], _09789_);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [1], _09674_);
  dff (\oc8051_top_1.oc8051_indi_addr1.wr_bit_r , _39457_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [0], _39555_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [1], _39556_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [2], _39557_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [3], _39558_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [4], _39559_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [5], _39560_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [6], _39561_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [7], _39458_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [0], _39562_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [1], _39563_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [2], _39564_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [3], _39566_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [4], _39567_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [5], _39568_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [6], _39569_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [7], _39459_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [0], _39570_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [1], _39571_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [2], _39572_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [3], _39573_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [4], _39574_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [5], _39575_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [6], _39577_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [7], _39460_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [0], _39578_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [1], _39579_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [2], _39580_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [3], _39581_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [4], _39582_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [5], _39583_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [6], _39584_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [7], _39462_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [0], _39585_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [1], _39586_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [2], _39588_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [3], _39589_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [4], _39590_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [5], _39591_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [6], _39592_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [7], _39463_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [0], _39593_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [1], _39594_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [2], _39595_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [3], _39596_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [4], _39597_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [5], _39599_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [6], _39600_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [7], _39464_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [0], _39601_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [1], _39602_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [2], _39603_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [3], _39604_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [4], _39605_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [5], _39606_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [6], _39607_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [7], _39465_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [0], _39608_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [1], _39610_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [2], _39611_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [3], _39612_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [4], _39613_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [5], _39614_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [6], _39615_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [7], _39466_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [0], _39027_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [1], _39028_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [2], _39029_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [3], _39030_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [4], _38743_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [0], _38816_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [1], _38817_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [2], _38818_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [3], _38819_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [4], _38820_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [5], _38822_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [6], _38823_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [7], _38824_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [8], _38825_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [9], _38826_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [10], _38827_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [11], _38828_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [12], _38829_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [13], _38830_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [14], _38831_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [15], _38705_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _38836_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _38837_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _38838_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _38839_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _38840_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _38841_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _38842_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _38843_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _38844_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _38845_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _38847_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _38848_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _38849_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _38850_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _38851_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _38706_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [0], _39031_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [1], _39032_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [2], _39033_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [3], _39034_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [4], _39036_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [5], _39037_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [6], _39038_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [7], _39039_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [8], _39040_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [9], _39041_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [10], _39042_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [11], _39043_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [12], _39044_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [13], _39045_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [14], _39047_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [15], _39048_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [16], _39049_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [17], _39050_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [18], _39051_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [19], _39052_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [20], _39053_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [21], _39054_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [22], _39055_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [23], _39056_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [24], _39058_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [25], _39059_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [26], _39060_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [27], _39061_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [28], _39062_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [29], _39063_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [30], _39064_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [31], _38768_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _38741_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dack_ir , 1'b0);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [0], _39065_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [1], _39067_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [2], _39068_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [3], _39069_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [4], _39070_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [5], _39071_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [6], _39073_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [7], _38744_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [0], _39074_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [1], _39075_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [2], _39076_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [3], _39077_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [4], _39078_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [5], _39079_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [6], _39080_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [7], _38745_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [0], _39081_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [1], _39082_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [2], _39084_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [3], _39085_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [4], _39086_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [5], _39087_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [6], _39088_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [7], _38747_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _38748_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _38749_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], _39089_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _39090_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], _39091_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], _39092_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _39093_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], _39095_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], _39096_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [7], _38750_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [0], _39097_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [1], _39098_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _39099_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [3], _39100_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [4], _39101_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [5], _39102_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [6], _39103_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [7], _39104_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [8], _39106_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [9], _39107_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [10], _39108_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [11], _39109_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [12], _39110_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [13], _39111_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [14], _39112_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [15], _38751_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [0], _39113_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [1], _39114_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [2], _39115_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [3], _39117_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [4], _39118_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [5], _39119_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [6], _39120_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [7], _39121_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [8], _39122_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [9], _39123_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [10], _39124_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [11], _39125_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [12], _39126_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [13], _39128_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [14], _39129_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [15], _38753_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack , _38754_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_t , _38756_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_buff , _38755_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], _39130_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], _39131_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _39132_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], _39133_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _39134_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], _39135_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _39136_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _38758_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [0], _39137_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [1], _39139_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [2], _38759_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [0], _39140_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [1], _39141_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [2], _39142_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [3], _39143_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [4], _39144_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [5], _39145_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [6], _39146_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [7], _38760_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [0], _39147_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [1], _39148_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [2], _39150_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [3], _39151_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [4], _39152_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [5], _39153_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [6], _39154_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [7], _38761_);
  dff (\oc8051_top_1.oc8051_memory_interface1.reti , _38762_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [0], _39155_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [1], _39156_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [2], _39157_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [3], _39158_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [4], _39159_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [5], _39161_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [6], _39162_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [7], _38763_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdone , _38765_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst , _38766_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], _39163_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], _39164_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], _39165_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], _38767_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [0], _39166_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [1], _39167_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [2], _39168_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [3], _39169_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [4], _39170_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [5], _39171_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [6], _39172_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [7], _39173_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [8], _39174_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [9], _39175_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [10], _39176_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [11], _39177_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [12], _39178_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [13], _39179_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [14], _39180_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [15], _39182_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [16], _39183_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [17], _39184_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [18], _39185_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [19], _39186_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [20], _39187_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [21], _39188_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [22], _39189_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [23], _39190_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [24], _39191_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [25], _39193_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [26], _39194_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [27], _39195_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [28], _39196_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [29], _39197_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [30], _39198_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [31], _38769_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [0], _39199_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [1], _39200_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [2], _39201_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [3], _39202_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [4], _39204_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [5], _39205_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [6], _39206_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [7], _38770_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dwe_o , _38771_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dstb_o , _38773_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [0], _39207_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [1], _39208_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [2], _39209_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [3], _39210_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [4], _39211_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [5], _39212_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [6], _39213_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [7], _39215_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [8], _39216_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [9], _39217_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [10], _39218_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [11], _39219_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [12], _39220_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [13], _39221_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [14], _39222_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [15], _38774_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dmem_wait , _38775_);
  dff (\oc8051_top_1.oc8051_memory_interface1.istb_t , _38776_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imem_wait , _38777_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _39223_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _39224_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _39226_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _39227_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [4], _39228_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [5], _39229_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [6], _39230_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [7], _39231_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [8], _39232_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [9], _39233_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [10], _39234_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [11], _39235_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [12], _39237_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [13], _39238_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [14], _39239_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [15], _38778_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_ind , _38779_);
  dff (\oc8051_top_1.oc8051_ram_top1.rd_en_r , _39843_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _39864_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _39865_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _39866_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _39867_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _39868_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _39869_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _39870_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [7], _39844_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_addr_r , _39845_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [0], _39871_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [1], _39872_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [2], _39846_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0], _02798_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1], _02803_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2], _02809_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3], _02814_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4], _02819_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5], _02824_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6], _02829_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7], _02831_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0], _02839_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1], _02842_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2], _02846_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3], _02850_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4], _02853_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5], _02856_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6], _02860_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7], _02862_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0], _02868_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1], _02873_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2], _02876_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3], _02879_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4], _02884_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5], _02887_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6], _02890_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7], _02893_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0], _02929_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1], _02933_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2], _02937_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3], _02941_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4], _02945_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5], _02948_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6], _02952_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7], _02956_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0], _02898_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1], _02902_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2], _02905_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3], _02908_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4], _02911_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5], _02915_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6], _02918_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7], _02921_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0], _03140_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1], _03143_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2], _03146_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3], _03149_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4], _03153_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5], _03156_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6], _03159_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7], _03162_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0], _03112_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1], _03115_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2], _03119_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3], _03122_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4], _03126_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5], _03130_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6], _03133_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7], _03136_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0], _03083_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1], _03087_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2], _03090_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3], _03094_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4], _03097_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5], _03101_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6], _03104_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7], _03107_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0], _03055_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1], _03058_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2], _03062_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3], _03065_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4], _03069_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5], _03072_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6], _03076_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7], _03079_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0], _03026_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1], _03030_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2], _03033_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3], _03037_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4], _03040_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5], _03043_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6], _03046_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7], _03049_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0], _02993_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1], _02998_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2], _03002_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3], _03005_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4], _03010_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5], _03014_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6], _03017_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7], _03020_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0], _02960_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1], _02964_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2], _02969_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3], _02973_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4], _02977_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5], _02982_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6], _02986_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7], _02988_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0], _03248_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1], _03251_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2], _03255_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3], _03258_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4], _03261_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5], _03264_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6], _03268_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7], _02574_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0], _03221_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1], _03225_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2], _03228_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3], _03232_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4], _03235_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5], _03238_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6], _03242_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7], _03244_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0], _03193_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1], _03196_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2], _03200_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3], _03204_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4], _03207_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5], _03211_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6], _03214_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7], _03217_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0], _03166_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1], _03170_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2], _03173_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3], _03176_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4], _03179_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5], _03183_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6], _03186_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7], _03188_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0], _05053_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1], _05055_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2], _05057_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3], _05059_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4], _05061_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5], _05063_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6], _05065_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7], _02564_);
  dff (\oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  dff (\oc8051_top_1.oc8051_rom1.ea_int , 1'b1);
  dff (\oc8051_top_1.oc8051_sfr1.pres_ow , _39679_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [0], _39764_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [1], _39765_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [2], _39766_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [3], _39681_);
  dff (\oc8051_top_1.oc8051_sfr1.bit_out , _39682_);
  dff (\oc8051_top_1.oc8051_sfr1.wait_data , _39683_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [0], _39768_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [1], _39769_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [2], _39770_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [3], _39771_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [4], _39772_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [5], _39773_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [6], _39774_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [7], _39684_);
  dff (\oc8051_top_1.oc8051_sfr1.wr_bit_r , _39685_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], _19757_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], _19769_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], _19780_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3], _19792_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4], _19804_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], _19816_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], _19828_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], _17963_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0], _08867_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1], _08878_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2], _08889_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3], _08900_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4], _08911_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5], _08922_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6], _08933_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7], _06626_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], _13613_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], _13624_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], _13635_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], _13646_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], _13657_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], _13668_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], _13679_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7], _12677_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0], _13690_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1], _13701_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2], _13711_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3], _13722_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4], _13733_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5], _13744_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6], _13755_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7], _12698_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff , _42623_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff , _42621_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff , 1'b0);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie1_buff , _42618_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], _00130_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], _00132_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _00134_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3], _00136_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4], _00138_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], _00139_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _00141_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _42616_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], _00143_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _42615_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc , _42613_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _00145_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _00147_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], _42611_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _00149_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _00150_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], _42609_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], _00152_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [1], _42607_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _00154_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [1], _42605_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , _42570_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , _42568_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , _42566_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , _42564_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0], _00156_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1], _00158_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2], _00160_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], _42561_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0], _00161_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], _00163_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], _00165_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3], _00167_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4], _00169_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5], _00171_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6], _00173_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _42559_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0], _00174_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1], _00176_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2], _00178_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3], _00180_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4], _00182_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5], _00184_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6], _00185_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7], _42556_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0], _40308_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1], _40310_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2], _40312_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3], _40314_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4], _40316_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5], _40318_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6], _40320_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7], _31034_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0], _40322_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1], _40324_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2], _40326_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3], _40327_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4], _40329_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5], _40331_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6], _40333_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7], _31057_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0], _40335_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1], _40337_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2], _40339_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3], _40341_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4], _40343_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5], _40345_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6], _40347_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7], _31079_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0], _40349_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1], _40351_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2], _40353_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3], _40355_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4], _40356_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5], _40358_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6], _40360_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7], _31102_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1], _17339_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], _17350_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3], _17361_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4], _17372_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5], _17383_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6], _17394_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], _15158_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop , _09484_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], _10660_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], _10671_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2], _10682_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3], _10693_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4], _10704_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5], _10715_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6], _10726_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7], _09504_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , _40810_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff , _40813_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0], _41323_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1], _41325_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2], _41327_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3], _41328_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4], _41330_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], _41332_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6], _41334_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7], _40816_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0], _41336_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1], _41338_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2], _41340_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3], _41342_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4], _41344_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5], _41345_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6], _41347_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7], _40819_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , _40822_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _40825_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0], _41349_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1], _41351_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2], _41353_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3], _41355_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4], _41357_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], _41359_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6], _41361_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7], _40828_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0], _41362_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1], _41364_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2], _41366_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3], _41368_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4], _41370_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5], _41372_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6], _41374_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7], _40831_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 , _40834_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _41376_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], _41378_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2], _41379_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3], _41381_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _41383_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], _41385_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6], _41387_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7], _40837_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r , _01626_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _01628_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , _01631_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r , _01634_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0], _02111_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1], _02113_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2], _02115_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3], _02117_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4], _02118_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5], _02120_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6], _02122_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7], _01637_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0], _02124_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1], _02125_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2], _02127_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3], _02129_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4], _02131_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5], _02132_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6], _02134_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7], _01640_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 , _01643_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0], _02136_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1], _02138_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2], _02139_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3], _02141_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4], _02143_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5], _02145_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6], _02146_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7], _01646_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0], _02148_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1], _02150_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2], _02152_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3], _02153_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4], _02155_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5], _02157_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6], _02159_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7], _01649_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set , _01652_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0], _02160_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1], _02162_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2], _02164_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3], _02166_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], _02167_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], _02169_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6], _02171_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], _01655_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0], _01206_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1], _01208_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2], _01210_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _01212_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _01214_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _01216_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _01218_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _01220_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8], _01221_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9], _01223_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], _01225_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _00567_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf , _00543_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , _00545_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , _00548_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive , _00551_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _00554_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r , _00556_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], _01227_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1], _00559_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], _01229_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], _01231_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _01233_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3], _00562_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0], _01235_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1], _01237_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2], _01239_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3], _01241_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4], _01243_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5], _01245_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6], _01247_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7], _00564_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr , _00570_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr , _00572_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd , _00575_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans , _00578_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , _00580_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0], _01249_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1], _01251_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2], _01253_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3], _00583_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0], _01255_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1], _01256_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], _01258_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3], _01260_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4], _01262_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5], _01264_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6], _01266_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7], _01268_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8], _01270_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], _01272_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10], _00586_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0], _01274_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1], _01276_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2], _01278_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3], _01280_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4], _01282_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5], _01284_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6], _01286_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], _00588_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0], _01288_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], _01290_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2], _01291_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3], _01293_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], _01295_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5], _01297_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6], _01299_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], _00591_);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div0 , \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div1 , \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [0], psw[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.p , psw[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [4], \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [5], \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.intr , \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_int , \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell0.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell0.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell0.word [0], word_in[0]);
  buf(\oc8051_gm_cxrom_1.cell0.word [1], word_in[1]);
  buf(\oc8051_gm_cxrom_1.cell0.word [2], word_in[2]);
  buf(\oc8051_gm_cxrom_1.cell0.word [3], word_in[3]);
  buf(\oc8051_gm_cxrom_1.cell0.word [4], word_in[4]);
  buf(\oc8051_gm_cxrom_1.cell0.word [5], word_in[5]);
  buf(\oc8051_gm_cxrom_1.cell0.word [6], word_in[6]);
  buf(\oc8051_gm_cxrom_1.cell0.word [7], word_in[7]);
  buf(\oc8051_gm_cxrom_1.cell1.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell1.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell1.word [0], word_in[8]);
  buf(\oc8051_gm_cxrom_1.cell1.word [1], word_in[9]);
  buf(\oc8051_gm_cxrom_1.cell1.word [2], word_in[10]);
  buf(\oc8051_gm_cxrom_1.cell1.word [3], word_in[11]);
  buf(\oc8051_gm_cxrom_1.cell1.word [4], word_in[12]);
  buf(\oc8051_gm_cxrom_1.cell1.word [5], word_in[13]);
  buf(\oc8051_gm_cxrom_1.cell1.word [6], word_in[14]);
  buf(\oc8051_gm_cxrom_1.cell1.word [7], word_in[15]);
  buf(\oc8051_gm_cxrom_1.cell2.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell2.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell2.word [0], word_in[16]);
  buf(\oc8051_gm_cxrom_1.cell2.word [1], word_in[17]);
  buf(\oc8051_gm_cxrom_1.cell2.word [2], word_in[18]);
  buf(\oc8051_gm_cxrom_1.cell2.word [3], word_in[19]);
  buf(\oc8051_gm_cxrom_1.cell2.word [4], word_in[20]);
  buf(\oc8051_gm_cxrom_1.cell2.word [5], word_in[21]);
  buf(\oc8051_gm_cxrom_1.cell2.word [6], word_in[22]);
  buf(\oc8051_gm_cxrom_1.cell2.word [7], word_in[23]);
  buf(\oc8051_gm_cxrom_1.cell3.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell3.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell3.word [0], word_in[24]);
  buf(\oc8051_gm_cxrom_1.cell3.word [1], word_in[25]);
  buf(\oc8051_gm_cxrom_1.cell3.word [2], word_in[26]);
  buf(\oc8051_gm_cxrom_1.cell3.word [3], word_in[27]);
  buf(\oc8051_gm_cxrom_1.cell3.word [4], word_in[28]);
  buf(\oc8051_gm_cxrom_1.cell3.word [5], word_in[29]);
  buf(\oc8051_gm_cxrom_1.cell3.word [6], word_in[30]);
  buf(\oc8051_gm_cxrom_1.cell3.word [7], word_in[31]);
  buf(\oc8051_gm_cxrom_1.cell4.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell4.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell4.word [0], word_in[32]);
  buf(\oc8051_gm_cxrom_1.cell4.word [1], word_in[33]);
  buf(\oc8051_gm_cxrom_1.cell4.word [2], word_in[34]);
  buf(\oc8051_gm_cxrom_1.cell4.word [3], word_in[35]);
  buf(\oc8051_gm_cxrom_1.cell4.word [4], word_in[36]);
  buf(\oc8051_gm_cxrom_1.cell4.word [5], word_in[37]);
  buf(\oc8051_gm_cxrom_1.cell4.word [6], word_in[38]);
  buf(\oc8051_gm_cxrom_1.cell4.word [7], word_in[39]);
  buf(\oc8051_gm_cxrom_1.cell5.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell5.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell5.word [0], word_in[40]);
  buf(\oc8051_gm_cxrom_1.cell5.word [1], word_in[41]);
  buf(\oc8051_gm_cxrom_1.cell5.word [2], word_in[42]);
  buf(\oc8051_gm_cxrom_1.cell5.word [3], word_in[43]);
  buf(\oc8051_gm_cxrom_1.cell5.word [4], word_in[44]);
  buf(\oc8051_gm_cxrom_1.cell5.word [5], word_in[45]);
  buf(\oc8051_gm_cxrom_1.cell5.word [6], word_in[46]);
  buf(\oc8051_gm_cxrom_1.cell5.word [7], word_in[47]);
  buf(\oc8051_gm_cxrom_1.cell6.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell6.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell6.word [0], word_in[48]);
  buf(\oc8051_gm_cxrom_1.cell6.word [1], word_in[49]);
  buf(\oc8051_gm_cxrom_1.cell6.word [2], word_in[50]);
  buf(\oc8051_gm_cxrom_1.cell6.word [3], word_in[51]);
  buf(\oc8051_gm_cxrom_1.cell6.word [4], word_in[52]);
  buf(\oc8051_gm_cxrom_1.cell6.word [5], word_in[53]);
  buf(\oc8051_gm_cxrom_1.cell6.word [6], word_in[54]);
  buf(\oc8051_gm_cxrom_1.cell6.word [7], word_in[55]);
  buf(\oc8051_gm_cxrom_1.cell7.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell7.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell7.word [0], word_in[56]);
  buf(\oc8051_gm_cxrom_1.cell7.word [1], word_in[57]);
  buf(\oc8051_gm_cxrom_1.cell7.word [2], word_in[58]);
  buf(\oc8051_gm_cxrom_1.cell7.word [3], word_in[59]);
  buf(\oc8051_gm_cxrom_1.cell7.word [4], word_in[60]);
  buf(\oc8051_gm_cxrom_1.cell7.word [5], word_in[61]);
  buf(\oc8051_gm_cxrom_1.cell7.word [6], word_in[62]);
  buf(\oc8051_gm_cxrom_1.cell7.word [7], word_in[63]);
  buf(\oc8051_gm_cxrom_1.cell8.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell8.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell8.word [0], word_in[64]);
  buf(\oc8051_gm_cxrom_1.cell8.word [1], word_in[65]);
  buf(\oc8051_gm_cxrom_1.cell8.word [2], word_in[66]);
  buf(\oc8051_gm_cxrom_1.cell8.word [3], word_in[67]);
  buf(\oc8051_gm_cxrom_1.cell8.word [4], word_in[68]);
  buf(\oc8051_gm_cxrom_1.cell8.word [5], word_in[69]);
  buf(\oc8051_gm_cxrom_1.cell8.word [6], word_in[70]);
  buf(\oc8051_gm_cxrom_1.cell8.word [7], word_in[71]);
  buf(\oc8051_gm_cxrom_1.cell9.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell9.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell9.word [0], word_in[72]);
  buf(\oc8051_gm_cxrom_1.cell9.word [1], word_in[73]);
  buf(\oc8051_gm_cxrom_1.cell9.word [2], word_in[74]);
  buf(\oc8051_gm_cxrom_1.cell9.word [3], word_in[75]);
  buf(\oc8051_gm_cxrom_1.cell9.word [4], word_in[76]);
  buf(\oc8051_gm_cxrom_1.cell9.word [5], word_in[77]);
  buf(\oc8051_gm_cxrom_1.cell9.word [6], word_in[78]);
  buf(\oc8051_gm_cxrom_1.cell9.word [7], word_in[79]);
  buf(\oc8051_gm_cxrom_1.cell10.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell10.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell10.word [0], word_in[80]);
  buf(\oc8051_gm_cxrom_1.cell10.word [1], word_in[81]);
  buf(\oc8051_gm_cxrom_1.cell10.word [2], word_in[82]);
  buf(\oc8051_gm_cxrom_1.cell10.word [3], word_in[83]);
  buf(\oc8051_gm_cxrom_1.cell10.word [4], word_in[84]);
  buf(\oc8051_gm_cxrom_1.cell10.word [5], word_in[85]);
  buf(\oc8051_gm_cxrom_1.cell10.word [6], word_in[86]);
  buf(\oc8051_gm_cxrom_1.cell10.word [7], word_in[87]);
  buf(\oc8051_gm_cxrom_1.cell11.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell11.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell11.word [0], word_in[88]);
  buf(\oc8051_gm_cxrom_1.cell11.word [1], word_in[89]);
  buf(\oc8051_gm_cxrom_1.cell11.word [2], word_in[90]);
  buf(\oc8051_gm_cxrom_1.cell11.word [3], word_in[91]);
  buf(\oc8051_gm_cxrom_1.cell11.word [4], word_in[92]);
  buf(\oc8051_gm_cxrom_1.cell11.word [5], word_in[93]);
  buf(\oc8051_gm_cxrom_1.cell11.word [6], word_in[94]);
  buf(\oc8051_gm_cxrom_1.cell11.word [7], word_in[95]);
  buf(\oc8051_gm_cxrom_1.cell12.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell12.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell12.word [0], word_in[96]);
  buf(\oc8051_gm_cxrom_1.cell12.word [1], word_in[97]);
  buf(\oc8051_gm_cxrom_1.cell12.word [2], word_in[98]);
  buf(\oc8051_gm_cxrom_1.cell12.word [3], word_in[99]);
  buf(\oc8051_gm_cxrom_1.cell12.word [4], word_in[100]);
  buf(\oc8051_gm_cxrom_1.cell12.word [5], word_in[101]);
  buf(\oc8051_gm_cxrom_1.cell12.word [6], word_in[102]);
  buf(\oc8051_gm_cxrom_1.cell12.word [7], word_in[103]);
  buf(\oc8051_gm_cxrom_1.cell13.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell13.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell13.word [0], word_in[104]);
  buf(\oc8051_gm_cxrom_1.cell13.word [1], word_in[105]);
  buf(\oc8051_gm_cxrom_1.cell13.word [2], word_in[106]);
  buf(\oc8051_gm_cxrom_1.cell13.word [3], word_in[107]);
  buf(\oc8051_gm_cxrom_1.cell13.word [4], word_in[108]);
  buf(\oc8051_gm_cxrom_1.cell13.word [5], word_in[109]);
  buf(\oc8051_gm_cxrom_1.cell13.word [6], word_in[110]);
  buf(\oc8051_gm_cxrom_1.cell13.word [7], word_in[111]);
  buf(\oc8051_gm_cxrom_1.cell14.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell14.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell14.word [0], word_in[112]);
  buf(\oc8051_gm_cxrom_1.cell14.word [1], word_in[113]);
  buf(\oc8051_gm_cxrom_1.cell14.word [2], word_in[114]);
  buf(\oc8051_gm_cxrom_1.cell14.word [3], word_in[115]);
  buf(\oc8051_gm_cxrom_1.cell14.word [4], word_in[116]);
  buf(\oc8051_gm_cxrom_1.cell14.word [5], word_in[117]);
  buf(\oc8051_gm_cxrom_1.cell14.word [6], word_in[118]);
  buf(\oc8051_gm_cxrom_1.cell14.word [7], word_in[119]);
  buf(\oc8051_gm_cxrom_1.cell15.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell15.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell15.word [0], word_in[120]);
  buf(\oc8051_gm_cxrom_1.cell15.word [1], word_in[121]);
  buf(\oc8051_gm_cxrom_1.cell15.word [2], word_in[122]);
  buf(\oc8051_gm_cxrom_1.cell15.word [3], word_in[123]);
  buf(\oc8051_gm_cxrom_1.cell15.word [4], word_in[124]);
  buf(\oc8051_gm_cxrom_1.cell15.word [5], word_in[125]);
  buf(\oc8051_gm_cxrom_1.cell15.word [6], word_in[126]);
  buf(\oc8051_gm_cxrom_1.cell15.word [7], word_in[127]);
  buf(\oc8051_top_1.oc8051_decoder1.clk , clk);
  buf(\oc8051_top_1.oc8051_decoder1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.oc8051_decoder1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.oc8051_comp1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_comp1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_comp1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_comp1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_comp1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_comp1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_comp1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_comp1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_comp1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_alu1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_in , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.rst , rst);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.oc8051_indi_addr1.clk , clk);
  buf(\oc8051_top_1.oc8051_indi_addr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [0], psw[0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.txd , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  buf(\oc8051_top_1.oc8051_sfr1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.p , psw[0]);
  buf(\oc8051_top_1.oc8051_sfr1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.ip [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  buf(\oc8051_top_1.oc8051_rom1.rst , rst);
  buf(\oc8051_top_1.oc8051_rom1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.rst , rst);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  buf(\oc8051_gm_cxrom_1.clk , clk);
  buf(\oc8051_gm_cxrom_1.rst , rst);
  buf(\oc8051_gm_cxrom_1.word_in [0], word_in[0]);
  buf(\oc8051_gm_cxrom_1.word_in [1], word_in[1]);
  buf(\oc8051_gm_cxrom_1.word_in [2], word_in[2]);
  buf(\oc8051_gm_cxrom_1.word_in [3], word_in[3]);
  buf(\oc8051_gm_cxrom_1.word_in [4], word_in[4]);
  buf(\oc8051_gm_cxrom_1.word_in [5], word_in[5]);
  buf(\oc8051_gm_cxrom_1.word_in [6], word_in[6]);
  buf(\oc8051_gm_cxrom_1.word_in [7], word_in[7]);
  buf(\oc8051_gm_cxrom_1.word_in [8], word_in[8]);
  buf(\oc8051_gm_cxrom_1.word_in [9], word_in[9]);
  buf(\oc8051_gm_cxrom_1.word_in [10], word_in[10]);
  buf(\oc8051_gm_cxrom_1.word_in [11], word_in[11]);
  buf(\oc8051_gm_cxrom_1.word_in [12], word_in[12]);
  buf(\oc8051_gm_cxrom_1.word_in [13], word_in[13]);
  buf(\oc8051_gm_cxrom_1.word_in [14], word_in[14]);
  buf(\oc8051_gm_cxrom_1.word_in [15], word_in[15]);
  buf(\oc8051_gm_cxrom_1.word_in [16], word_in[16]);
  buf(\oc8051_gm_cxrom_1.word_in [17], word_in[17]);
  buf(\oc8051_gm_cxrom_1.word_in [18], word_in[18]);
  buf(\oc8051_gm_cxrom_1.word_in [19], word_in[19]);
  buf(\oc8051_gm_cxrom_1.word_in [20], word_in[20]);
  buf(\oc8051_gm_cxrom_1.word_in [21], word_in[21]);
  buf(\oc8051_gm_cxrom_1.word_in [22], word_in[22]);
  buf(\oc8051_gm_cxrom_1.word_in [23], word_in[23]);
  buf(\oc8051_gm_cxrom_1.word_in [24], word_in[24]);
  buf(\oc8051_gm_cxrom_1.word_in [25], word_in[25]);
  buf(\oc8051_gm_cxrom_1.word_in [26], word_in[26]);
  buf(\oc8051_gm_cxrom_1.word_in [27], word_in[27]);
  buf(\oc8051_gm_cxrom_1.word_in [28], word_in[28]);
  buf(\oc8051_gm_cxrom_1.word_in [29], word_in[29]);
  buf(\oc8051_gm_cxrom_1.word_in [30], word_in[30]);
  buf(\oc8051_gm_cxrom_1.word_in [31], word_in[31]);
  buf(\oc8051_gm_cxrom_1.word_in [32], word_in[32]);
  buf(\oc8051_gm_cxrom_1.word_in [33], word_in[33]);
  buf(\oc8051_gm_cxrom_1.word_in [34], word_in[34]);
  buf(\oc8051_gm_cxrom_1.word_in [35], word_in[35]);
  buf(\oc8051_gm_cxrom_1.word_in [36], word_in[36]);
  buf(\oc8051_gm_cxrom_1.word_in [37], word_in[37]);
  buf(\oc8051_gm_cxrom_1.word_in [38], word_in[38]);
  buf(\oc8051_gm_cxrom_1.word_in [39], word_in[39]);
  buf(\oc8051_gm_cxrom_1.word_in [40], word_in[40]);
  buf(\oc8051_gm_cxrom_1.word_in [41], word_in[41]);
  buf(\oc8051_gm_cxrom_1.word_in [42], word_in[42]);
  buf(\oc8051_gm_cxrom_1.word_in [43], word_in[43]);
  buf(\oc8051_gm_cxrom_1.word_in [44], word_in[44]);
  buf(\oc8051_gm_cxrom_1.word_in [45], word_in[45]);
  buf(\oc8051_gm_cxrom_1.word_in [46], word_in[46]);
  buf(\oc8051_gm_cxrom_1.word_in [47], word_in[47]);
  buf(\oc8051_gm_cxrom_1.word_in [48], word_in[48]);
  buf(\oc8051_gm_cxrom_1.word_in [49], word_in[49]);
  buf(\oc8051_gm_cxrom_1.word_in [50], word_in[50]);
  buf(\oc8051_gm_cxrom_1.word_in [51], word_in[51]);
  buf(\oc8051_gm_cxrom_1.word_in [52], word_in[52]);
  buf(\oc8051_gm_cxrom_1.word_in [53], word_in[53]);
  buf(\oc8051_gm_cxrom_1.word_in [54], word_in[54]);
  buf(\oc8051_gm_cxrom_1.word_in [55], word_in[55]);
  buf(\oc8051_gm_cxrom_1.word_in [56], word_in[56]);
  buf(\oc8051_gm_cxrom_1.word_in [57], word_in[57]);
  buf(\oc8051_gm_cxrom_1.word_in [58], word_in[58]);
  buf(\oc8051_gm_cxrom_1.word_in [59], word_in[59]);
  buf(\oc8051_gm_cxrom_1.word_in [60], word_in[60]);
  buf(\oc8051_gm_cxrom_1.word_in [61], word_in[61]);
  buf(\oc8051_gm_cxrom_1.word_in [62], word_in[62]);
  buf(\oc8051_gm_cxrom_1.word_in [63], word_in[63]);
  buf(\oc8051_gm_cxrom_1.word_in [64], word_in[64]);
  buf(\oc8051_gm_cxrom_1.word_in [65], word_in[65]);
  buf(\oc8051_gm_cxrom_1.word_in [66], word_in[66]);
  buf(\oc8051_gm_cxrom_1.word_in [67], word_in[67]);
  buf(\oc8051_gm_cxrom_1.word_in [68], word_in[68]);
  buf(\oc8051_gm_cxrom_1.word_in [69], word_in[69]);
  buf(\oc8051_gm_cxrom_1.word_in [70], word_in[70]);
  buf(\oc8051_gm_cxrom_1.word_in [71], word_in[71]);
  buf(\oc8051_gm_cxrom_1.word_in [72], word_in[72]);
  buf(\oc8051_gm_cxrom_1.word_in [73], word_in[73]);
  buf(\oc8051_gm_cxrom_1.word_in [74], word_in[74]);
  buf(\oc8051_gm_cxrom_1.word_in [75], word_in[75]);
  buf(\oc8051_gm_cxrom_1.word_in [76], word_in[76]);
  buf(\oc8051_gm_cxrom_1.word_in [77], word_in[77]);
  buf(\oc8051_gm_cxrom_1.word_in [78], word_in[78]);
  buf(\oc8051_gm_cxrom_1.word_in [79], word_in[79]);
  buf(\oc8051_gm_cxrom_1.word_in [80], word_in[80]);
  buf(\oc8051_gm_cxrom_1.word_in [81], word_in[81]);
  buf(\oc8051_gm_cxrom_1.word_in [82], word_in[82]);
  buf(\oc8051_gm_cxrom_1.word_in [83], word_in[83]);
  buf(\oc8051_gm_cxrom_1.word_in [84], word_in[84]);
  buf(\oc8051_gm_cxrom_1.word_in [85], word_in[85]);
  buf(\oc8051_gm_cxrom_1.word_in [86], word_in[86]);
  buf(\oc8051_gm_cxrom_1.word_in [87], word_in[87]);
  buf(\oc8051_gm_cxrom_1.word_in [88], word_in[88]);
  buf(\oc8051_gm_cxrom_1.word_in [89], word_in[89]);
  buf(\oc8051_gm_cxrom_1.word_in [90], word_in[90]);
  buf(\oc8051_gm_cxrom_1.word_in [91], word_in[91]);
  buf(\oc8051_gm_cxrom_1.word_in [92], word_in[92]);
  buf(\oc8051_gm_cxrom_1.word_in [93], word_in[93]);
  buf(\oc8051_gm_cxrom_1.word_in [94], word_in[94]);
  buf(\oc8051_gm_cxrom_1.word_in [95], word_in[95]);
  buf(\oc8051_gm_cxrom_1.word_in [96], word_in[96]);
  buf(\oc8051_gm_cxrom_1.word_in [97], word_in[97]);
  buf(\oc8051_gm_cxrom_1.word_in [98], word_in[98]);
  buf(\oc8051_gm_cxrom_1.word_in [99], word_in[99]);
  buf(\oc8051_gm_cxrom_1.word_in [100], word_in[100]);
  buf(\oc8051_gm_cxrom_1.word_in [101], word_in[101]);
  buf(\oc8051_gm_cxrom_1.word_in [102], word_in[102]);
  buf(\oc8051_gm_cxrom_1.word_in [103], word_in[103]);
  buf(\oc8051_gm_cxrom_1.word_in [104], word_in[104]);
  buf(\oc8051_gm_cxrom_1.word_in [105], word_in[105]);
  buf(\oc8051_gm_cxrom_1.word_in [106], word_in[106]);
  buf(\oc8051_gm_cxrom_1.word_in [107], word_in[107]);
  buf(\oc8051_gm_cxrom_1.word_in [108], word_in[108]);
  buf(\oc8051_gm_cxrom_1.word_in [109], word_in[109]);
  buf(\oc8051_gm_cxrom_1.word_in [110], word_in[110]);
  buf(\oc8051_gm_cxrom_1.word_in [111], word_in[111]);
  buf(\oc8051_gm_cxrom_1.word_in [112], word_in[112]);
  buf(\oc8051_gm_cxrom_1.word_in [113], word_in[113]);
  buf(\oc8051_gm_cxrom_1.word_in [114], word_in[114]);
  buf(\oc8051_gm_cxrom_1.word_in [115], word_in[115]);
  buf(\oc8051_gm_cxrom_1.word_in [116], word_in[116]);
  buf(\oc8051_gm_cxrom_1.word_in [117], word_in[117]);
  buf(\oc8051_gm_cxrom_1.word_in [118], word_in[118]);
  buf(\oc8051_gm_cxrom_1.word_in [119], word_in[119]);
  buf(\oc8051_gm_cxrom_1.word_in [120], word_in[120]);
  buf(\oc8051_gm_cxrom_1.word_in [121], word_in[121]);
  buf(\oc8051_gm_cxrom_1.word_in [122], word_in[122]);
  buf(\oc8051_gm_cxrom_1.word_in [123], word_in[123]);
  buf(\oc8051_gm_cxrom_1.word_in [124], word_in[124]);
  buf(\oc8051_gm_cxrom_1.word_in [125], word_in[125]);
  buf(\oc8051_gm_cxrom_1.word_in [126], word_in[126]);
  buf(\oc8051_gm_cxrom_1.word_in [127], word_in[127]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [0], \oc8051_golden_model_1.PC [0]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [1], \oc8051_golden_model_1.PC [1]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [2], \oc8051_golden_model_1.PC [2]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [3], \oc8051_golden_model_1.PC [3]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [4], \oc8051_golden_model_1.PC [4]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [5], \oc8051_golden_model_1.PC [5]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [6], \oc8051_golden_model_1.PC [6]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [7], \oc8051_golden_model_1.PC [7]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [8], \oc8051_golden_model_1.PC [8]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [9], \oc8051_golden_model_1.PC [9]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [10], \oc8051_golden_model_1.PC [10]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [11], \oc8051_golden_model_1.PC [11]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [12], \oc8051_golden_model_1.PC [12]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [13], \oc8051_golden_model_1.PC [13]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [14], \oc8051_golden_model_1.PC [14]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [15], \oc8051_golden_model_1.PC [15]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [0], \oc8051_golden_model_1.PC [0]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [1], \oc8051_golden_model_1.PC [1]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [2], \oc8051_golden_model_1.PC [2]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [3], \oc8051_golden_model_1.PC [3]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [4], \oc8051_golden_model_1.PC [4]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [5], \oc8051_golden_model_1.PC [5]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [6], \oc8051_golden_model_1.PC [6]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [7], \oc8051_golden_model_1.PC [7]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [8], \oc8051_golden_model_1.PC [8]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [9], \oc8051_golden_model_1.PC [9]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [10], \oc8051_golden_model_1.PC [10]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [11], \oc8051_golden_model_1.PC [11]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [12], \oc8051_golden_model_1.PC [12]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [13], \oc8051_golden_model_1.PC [13]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [14], \oc8051_golden_model_1.PC [14]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [15], \oc8051_golden_model_1.PC [15]);
  buf(\oc8051_golden_model_1.clk , clk);
  buf(\oc8051_golden_model_1.rst , rst);
  buf(\oc8051_golden_model_1.RD_IRAM_ADDR [0], word_in[0]);
  buf(\oc8051_golden_model_1.RD_IRAM_ADDR [1], word_in[1]);
  buf(\oc8051_golden_model_1.RD_IRAM_ADDR [2], word_in[2]);
  buf(\oc8051_golden_model_1.RD_IRAM_ADDR [3], word_in[3]);
  buf(\oc8051_golden_model_1.ACC_03 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_03 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_03 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_03 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_03 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_03 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_03 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_03 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_13 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_13 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_13 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_13 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_13 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_13 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_13 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_13 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.ACC_23 [0], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_23 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_23 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_23 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_23 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_23 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_23 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_23 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_33 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.ACC_33 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_33 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_33 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_33 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_33 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_33 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_33 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_c4 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_c4 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_c4 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_c4 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_c4 [4], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_c4 [5], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_c4 [6], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_c4 [7], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_d6 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.ACC_d6 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.ACC_d6 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.ACC_d6 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.ACC_d6 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_d6 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_d6 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_d6 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_d7 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.ACC_d7 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.ACC_d7 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.ACC_d7 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.ACC_d7 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_d7 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_d7 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_d7 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_e4 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.ACC_e4 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.ACC_e4 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.ACC_e4 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.ACC_e4 [4], \oc8051_golden_model_1.n1854 [4]);
  buf(\oc8051_golden_model_1.ACC_e4 [5], \oc8051_golden_model_1.n1854 [5]);
  buf(\oc8051_golden_model_1.ACC_e4 [6], \oc8051_golden_model_1.n1854 [6]);
  buf(\oc8051_golden_model_1.ACC_e4 [7], \oc8051_golden_model_1.n1854 [7]);
  buf(\oc8051_golden_model_1.PC_22 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.PC_22 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.PC_22 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.PC_22 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.PC_22 [4], \oc8051_golden_model_1.n1854 [4]);
  buf(\oc8051_golden_model_1.PC_22 [5], \oc8051_golden_model_1.n1854 [5]);
  buf(\oc8051_golden_model_1.PC_22 [6], \oc8051_golden_model_1.n1854 [6]);
  buf(\oc8051_golden_model_1.PC_22 [7], \oc8051_golden_model_1.n1854 [7]);
  buf(\oc8051_golden_model_1.PC_22 [8], \oc8051_golden_model_1.n1268 [0]);
  buf(\oc8051_golden_model_1.PC_22 [9], \oc8051_golden_model_1.n1268 [1]);
  buf(\oc8051_golden_model_1.PC_22 [10], \oc8051_golden_model_1.n1268 [2]);
  buf(\oc8051_golden_model_1.PC_22 [11], \oc8051_golden_model_1.n1268 [3]);
  buf(\oc8051_golden_model_1.PC_22 [12], \oc8051_golden_model_1.n1268 [4]);
  buf(\oc8051_golden_model_1.PC_22 [13], \oc8051_golden_model_1.n1268 [5]);
  buf(\oc8051_golden_model_1.PC_22 [14], \oc8051_golden_model_1.n1268 [6]);
  buf(\oc8051_golden_model_1.PC_22 [15], \oc8051_golden_model_1.n1268 [8]);
  buf(\oc8051_golden_model_1.PC_32 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.PC_32 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.PC_32 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.PC_32 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.PC_32 [4], \oc8051_golden_model_1.n1854 [4]);
  buf(\oc8051_golden_model_1.PC_32 [5], \oc8051_golden_model_1.n1854 [5]);
  buf(\oc8051_golden_model_1.PC_32 [6], \oc8051_golden_model_1.n1854 [6]);
  buf(\oc8051_golden_model_1.PC_32 [7], \oc8051_golden_model_1.n1854 [7]);
  buf(\oc8051_golden_model_1.PC_32 [8], \oc8051_golden_model_1.n1268 [0]);
  buf(\oc8051_golden_model_1.PC_32 [9], \oc8051_golden_model_1.n1268 [1]);
  buf(\oc8051_golden_model_1.PC_32 [10], \oc8051_golden_model_1.n1268 [2]);
  buf(\oc8051_golden_model_1.PC_32 [11], \oc8051_golden_model_1.n1268 [3]);
  buf(\oc8051_golden_model_1.PC_32 [12], \oc8051_golden_model_1.n1268 [4]);
  buf(\oc8051_golden_model_1.PC_32 [13], \oc8051_golden_model_1.n1268 [5]);
  buf(\oc8051_golden_model_1.PC_32 [14], \oc8051_golden_model_1.n1268 [6]);
  buf(\oc8051_golden_model_1.PC_32 [15], \oc8051_golden_model_1.n1268 [8]);
  buf(\oc8051_golden_model_1.PSW_13 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_13 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_13 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_13 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_13 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_13 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_13 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_13 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.PSW_24 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_24 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_24 [2], \oc8051_golden_model_1.n1207 [2]);
  buf(\oc8051_golden_model_1.PSW_24 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_24 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_24 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_24 [6], \oc8051_golden_model_1.n1207 [6]);
  buf(\oc8051_golden_model_1.PSW_24 [7], \oc8051_golden_model_1.n1207 [7]);
  buf(\oc8051_golden_model_1.PSW_25 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_25 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_25 [2], \oc8051_golden_model_1.n1227 [2]);
  buf(\oc8051_golden_model_1.PSW_25 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_25 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_25 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_25 [6], \oc8051_golden_model_1.n1227 [6]);
  buf(\oc8051_golden_model_1.PSW_25 [7], \oc8051_golden_model_1.n1227 [7]);
  buf(\oc8051_golden_model_1.PSW_26 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_26 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_26 [2], \oc8051_golden_model_1.n1246 [2]);
  buf(\oc8051_golden_model_1.PSW_26 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_26 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_26 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_26 [6], \oc8051_golden_model_1.n1258 [6]);
  buf(\oc8051_golden_model_1.PSW_26 [7], \oc8051_golden_model_1.n1246 [7]);
  buf(\oc8051_golden_model_1.PSW_27 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_27 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_27 [2], \oc8051_golden_model_1.n1258 [2]);
  buf(\oc8051_golden_model_1.PSW_27 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_27 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_27 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_27 [6], \oc8051_golden_model_1.n1258 [6]);
  buf(\oc8051_golden_model_1.PSW_27 [7], \oc8051_golden_model_1.n1258 [7]);
  buf(\oc8051_golden_model_1.PSW_28 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_28 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_28 [2], \oc8051_golden_model_1.n1280 [2]);
  buf(\oc8051_golden_model_1.PSW_28 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_28 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_28 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_28 [6], \oc8051_golden_model_1.n1292 [6]);
  buf(\oc8051_golden_model_1.PSW_28 [7], \oc8051_golden_model_1.n1280 [7]);
  buf(\oc8051_golden_model_1.PSW_29 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_29 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_29 [2], \oc8051_golden_model_1.n1280 [2]);
  buf(\oc8051_golden_model_1.PSW_29 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_29 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_29 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_29 [6], \oc8051_golden_model_1.n1292 [6]);
  buf(\oc8051_golden_model_1.PSW_29 [7], \oc8051_golden_model_1.n1280 [7]);
  buf(\oc8051_golden_model_1.PSW_2a [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_2a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2a [2], \oc8051_golden_model_1.n1280 [2]);
  buf(\oc8051_golden_model_1.PSW_2a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2a [6], \oc8051_golden_model_1.n1291 [6]);
  buf(\oc8051_golden_model_1.PSW_2a [7], \oc8051_golden_model_1.n1280 [7]);
  buf(\oc8051_golden_model_1.PSW_2b [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_2b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2b [2], \oc8051_golden_model_1.n1292 [2]);
  buf(\oc8051_golden_model_1.PSW_2b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2b [6], \oc8051_golden_model_1.n1291 [6]);
  buf(\oc8051_golden_model_1.PSW_2b [7], \oc8051_golden_model_1.n1292 [7]);
  buf(\oc8051_golden_model_1.PSW_2c [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_2c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2c [2], \oc8051_golden_model_1.n1292 [2]);
  buf(\oc8051_golden_model_1.PSW_2c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2c [6], \oc8051_golden_model_1.n1291 [6]);
  buf(\oc8051_golden_model_1.PSW_2c [7], \oc8051_golden_model_1.n1292 [7]);
  buf(\oc8051_golden_model_1.PSW_2d [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_2d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2d [2], \oc8051_golden_model_1.n1280 [2]);
  buf(\oc8051_golden_model_1.PSW_2d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2d [6], \oc8051_golden_model_1.n1292 [6]);
  buf(\oc8051_golden_model_1.PSW_2d [7], \oc8051_golden_model_1.n1280 [7]);
  buf(\oc8051_golden_model_1.PSW_2e [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_2e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2e [2], \oc8051_golden_model_1.n1292 [2]);
  buf(\oc8051_golden_model_1.PSW_2e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2e [6], \oc8051_golden_model_1.n1292 [6]);
  buf(\oc8051_golden_model_1.PSW_2e [7], \oc8051_golden_model_1.n1292 [7]);
  buf(\oc8051_golden_model_1.PSW_2f [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_2f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2f [2], \oc8051_golden_model_1.n1292 [2]);
  buf(\oc8051_golden_model_1.PSW_2f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2f [6], \oc8051_golden_model_1.n1292 [6]);
  buf(\oc8051_golden_model_1.PSW_2f [7], \oc8051_golden_model_1.n1292 [7]);
  buf(\oc8051_golden_model_1.PSW_33 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_33 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_33 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_33 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_33 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_33 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_33 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_33 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.PSW_34 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_34 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_34 [2], \oc8051_golden_model_1.n1318 [2]);
  buf(\oc8051_golden_model_1.PSW_34 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_34 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_34 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_34 [6], \oc8051_golden_model_1.n1318 [6]);
  buf(\oc8051_golden_model_1.PSW_34 [7], \oc8051_golden_model_1.n1318 [7]);
  buf(\oc8051_golden_model_1.PSW_35 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_35 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_35 [2], \oc8051_golden_model_1.n1334 [2]);
  buf(\oc8051_golden_model_1.PSW_35 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_35 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_35 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_35 [6], \oc8051_golden_model_1.n1334 [6]);
  buf(\oc8051_golden_model_1.PSW_35 [7], \oc8051_golden_model_1.n1334 [7]);
  buf(\oc8051_golden_model_1.PSW_36 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_36 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_36 [2], \oc8051_golden_model_1.n1350 [2]);
  buf(\oc8051_golden_model_1.PSW_36 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_36 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_36 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_36 [6], \oc8051_golden_model_1.n1350 [6]);
  buf(\oc8051_golden_model_1.PSW_36 [7], \oc8051_golden_model_1.n1350 [7]);
  buf(\oc8051_golden_model_1.PSW_37 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_37 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_37 [2], \oc8051_golden_model_1.n1350 [2]);
  buf(\oc8051_golden_model_1.PSW_37 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_37 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_37 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_37 [6], \oc8051_golden_model_1.n1350 [6]);
  buf(\oc8051_golden_model_1.PSW_37 [7], \oc8051_golden_model_1.n1350 [7]);
  buf(\oc8051_golden_model_1.PSW_38 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_38 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_38 [2], \oc8051_golden_model_1.n1366 [2]);
  buf(\oc8051_golden_model_1.PSW_38 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_38 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_38 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_38 [6], \oc8051_golden_model_1.n1366 [6]);
  buf(\oc8051_golden_model_1.PSW_38 [7], \oc8051_golden_model_1.n1366 [7]);
  buf(\oc8051_golden_model_1.PSW_39 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_39 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_39 [2], \oc8051_golden_model_1.n1366 [2]);
  buf(\oc8051_golden_model_1.PSW_39 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_39 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_39 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_39 [6], \oc8051_golden_model_1.n1366 [6]);
  buf(\oc8051_golden_model_1.PSW_39 [7], \oc8051_golden_model_1.n1366 [7]);
  buf(\oc8051_golden_model_1.PSW_3a [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_3a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3a [2], \oc8051_golden_model_1.n1366 [2]);
  buf(\oc8051_golden_model_1.PSW_3a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3a [6], \oc8051_golden_model_1.n1366 [6]);
  buf(\oc8051_golden_model_1.PSW_3a [7], \oc8051_golden_model_1.n1366 [7]);
  buf(\oc8051_golden_model_1.PSW_3b [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_3b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3b [2], \oc8051_golden_model_1.n1366 [2]);
  buf(\oc8051_golden_model_1.PSW_3b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3b [6], \oc8051_golden_model_1.n1366 [6]);
  buf(\oc8051_golden_model_1.PSW_3b [7], \oc8051_golden_model_1.n1366 [7]);
  buf(\oc8051_golden_model_1.PSW_3c [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_3c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3c [2], \oc8051_golden_model_1.n1366 [2]);
  buf(\oc8051_golden_model_1.PSW_3c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3c [6], \oc8051_golden_model_1.n1366 [6]);
  buf(\oc8051_golden_model_1.PSW_3c [7], \oc8051_golden_model_1.n1366 [7]);
  buf(\oc8051_golden_model_1.PSW_3d [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_3d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3d [2], \oc8051_golden_model_1.n1366 [2]);
  buf(\oc8051_golden_model_1.PSW_3d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3d [6], \oc8051_golden_model_1.n1366 [6]);
  buf(\oc8051_golden_model_1.PSW_3d [7], \oc8051_golden_model_1.n1366 [7]);
  buf(\oc8051_golden_model_1.PSW_3e [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_3e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3e [2], \oc8051_golden_model_1.n1366 [2]);
  buf(\oc8051_golden_model_1.PSW_3e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3e [6], \oc8051_golden_model_1.n1366 [6]);
  buf(\oc8051_golden_model_1.PSW_3e [7], \oc8051_golden_model_1.n1366 [7]);
  buf(\oc8051_golden_model_1.PSW_3f [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_3f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3f [2], \oc8051_golden_model_1.n1366 [2]);
  buf(\oc8051_golden_model_1.PSW_3f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3f [6], \oc8051_golden_model_1.n1366 [6]);
  buf(\oc8051_golden_model_1.PSW_3f [7], \oc8051_golden_model_1.n1366 [7]);
  buf(\oc8051_golden_model_1.PSW_72 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_72 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_72 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_72 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_72 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_72 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_72 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_72 [7], \oc8051_golden_model_1.n1522 [7]);
  buf(\oc8051_golden_model_1.PSW_82 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_82 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_82 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_82 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_82 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_82 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_82 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_82 [7], \oc8051_golden_model_1.n1546 [7]);
  buf(\oc8051_golden_model_1.PSW_84 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_84 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_84 [2], \oc8051_golden_model_1.n1555 [2]);
  buf(\oc8051_golden_model_1.PSW_84 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_84 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_84 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_84 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_84 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_94 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_94 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_94 [2], \oc8051_golden_model_1.n1692 [2]);
  buf(\oc8051_golden_model_1.PSW_94 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_94 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_94 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_94 [6], \oc8051_golden_model_1.n1692 [6]);
  buf(\oc8051_golden_model_1.PSW_94 [7], \oc8051_golden_model_1.n1692 [7]);
  buf(\oc8051_golden_model_1.PSW_95 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_95 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_95 [2], \oc8051_golden_model_1.n1705 [2]);
  buf(\oc8051_golden_model_1.PSW_95 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_95 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_95 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_95 [6], \oc8051_golden_model_1.n1705 [6]);
  buf(\oc8051_golden_model_1.PSW_95 [7], \oc8051_golden_model_1.n1705 [7]);
  buf(\oc8051_golden_model_1.PSW_96 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_96 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_96 [2], \oc8051_golden_model_1.n1718 [2]);
  buf(\oc8051_golden_model_1.PSW_96 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_96 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_96 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_96 [6], \oc8051_golden_model_1.n1718 [6]);
  buf(\oc8051_golden_model_1.PSW_96 [7], \oc8051_golden_model_1.n1718 [7]);
  buf(\oc8051_golden_model_1.PSW_97 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_97 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_97 [2], \oc8051_golden_model_1.n1718 [2]);
  buf(\oc8051_golden_model_1.PSW_97 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_97 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_97 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_97 [6], \oc8051_golden_model_1.n1718 [6]);
  buf(\oc8051_golden_model_1.PSW_97 [7], \oc8051_golden_model_1.n1718 [7]);
  buf(\oc8051_golden_model_1.PSW_98 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_98 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_98 [2], \oc8051_golden_model_1.n1731 [2]);
  buf(\oc8051_golden_model_1.PSW_98 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_98 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_98 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_98 [6], \oc8051_golden_model_1.n1731 [6]);
  buf(\oc8051_golden_model_1.PSW_98 [7], \oc8051_golden_model_1.n1731 [7]);
  buf(\oc8051_golden_model_1.PSW_99 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_99 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_99 [2], \oc8051_golden_model_1.n1731 [2]);
  buf(\oc8051_golden_model_1.PSW_99 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_99 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_99 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_99 [6], \oc8051_golden_model_1.n1731 [6]);
  buf(\oc8051_golden_model_1.PSW_99 [7], \oc8051_golden_model_1.n1731 [7]);
  buf(\oc8051_golden_model_1.PSW_9a [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_9a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9a [2], \oc8051_golden_model_1.n1731 [2]);
  buf(\oc8051_golden_model_1.PSW_9a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9a [6], \oc8051_golden_model_1.n1731 [6]);
  buf(\oc8051_golden_model_1.PSW_9a [7], \oc8051_golden_model_1.n1731 [7]);
  buf(\oc8051_golden_model_1.PSW_9b [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_9b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9b [2], \oc8051_golden_model_1.n1731 [2]);
  buf(\oc8051_golden_model_1.PSW_9b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9b [6], \oc8051_golden_model_1.n1731 [6]);
  buf(\oc8051_golden_model_1.PSW_9b [7], \oc8051_golden_model_1.n1731 [7]);
  buf(\oc8051_golden_model_1.PSW_9c [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_9c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9c [2], \oc8051_golden_model_1.n1731 [2]);
  buf(\oc8051_golden_model_1.PSW_9c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9c [6], \oc8051_golden_model_1.n1731 [6]);
  buf(\oc8051_golden_model_1.PSW_9c [7], \oc8051_golden_model_1.n1731 [7]);
  buf(\oc8051_golden_model_1.PSW_9d [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_9d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9d [2], \oc8051_golden_model_1.n1731 [2]);
  buf(\oc8051_golden_model_1.PSW_9d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9d [6], \oc8051_golden_model_1.n1731 [6]);
  buf(\oc8051_golden_model_1.PSW_9d [7], \oc8051_golden_model_1.n1731 [7]);
  buf(\oc8051_golden_model_1.PSW_9e [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_9e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9e [2], \oc8051_golden_model_1.n1731 [2]);
  buf(\oc8051_golden_model_1.PSW_9e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9e [6], \oc8051_golden_model_1.n1731 [6]);
  buf(\oc8051_golden_model_1.PSW_9e [7], \oc8051_golden_model_1.n1731 [7]);
  buf(\oc8051_golden_model_1.PSW_9f [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_9f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9f [2], \oc8051_golden_model_1.n1731 [2]);
  buf(\oc8051_golden_model_1.PSW_9f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9f [6], \oc8051_golden_model_1.n1731 [6]);
  buf(\oc8051_golden_model_1.PSW_9f [7], \oc8051_golden_model_1.n1731 [7]);
  buf(\oc8051_golden_model_1.PSW_a0 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_a0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a0 [7], \oc8051_golden_model_1.n1734 [7]);
  buf(\oc8051_golden_model_1.PSW_a2 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_a2 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a2 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a2 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a2 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a2 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a2 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a2 [7], \oc8051_golden_model_1.n1735 [7]);
  buf(\oc8051_golden_model_1.PSW_a4 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_a4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a4 [2], \oc8051_golden_model_1.n1746 [2]);
  buf(\oc8051_golden_model_1.PSW_a4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a4 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_b0 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b0 [7], \oc8051_golden_model_1.n1750 [7]);
  buf(\oc8051_golden_model_1.PSW_b3 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b3 [7], \oc8051_golden_model_1.n1766 [7]);
  buf(\oc8051_golden_model_1.PSW_b4 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b4 [7], \oc8051_golden_model_1.n1772 [7]);
  buf(\oc8051_golden_model_1.PSW_b5 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b5 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b5 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b5 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b5 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b5 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b5 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b5 [7], \oc8051_golden_model_1.n1778 [7]);
  buf(\oc8051_golden_model_1.PSW_b6 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b6 [7], \oc8051_golden_model_1.n1784 [7]);
  buf(\oc8051_golden_model_1.PSW_b7 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b7 [7], \oc8051_golden_model_1.n1784 [7]);
  buf(\oc8051_golden_model_1.PSW_b8 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b8 [7], \oc8051_golden_model_1.n1790 [7]);
  buf(\oc8051_golden_model_1.PSW_b9 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b9 [7], \oc8051_golden_model_1.n1790 [7]);
  buf(\oc8051_golden_model_1.PSW_ba [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_ba [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ba [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ba [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ba [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ba [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ba [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ba [7], \oc8051_golden_model_1.n1790 [7]);
  buf(\oc8051_golden_model_1.PSW_bb [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_bb [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bb [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bb [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bb [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bb [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bb [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bb [7], \oc8051_golden_model_1.n1790 [7]);
  buf(\oc8051_golden_model_1.PSW_bc [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_bc [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bc [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bc [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bc [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bc [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bc [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bc [7], \oc8051_golden_model_1.n1790 [7]);
  buf(\oc8051_golden_model_1.PSW_bd [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_bd [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bd [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bd [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bd [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bd [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bd [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bd [7], \oc8051_golden_model_1.n1790 [7]);
  buf(\oc8051_golden_model_1.PSW_be [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_be [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_be [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_be [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_be [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_be [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_be [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_be [7], \oc8051_golden_model_1.n1790 [7]);
  buf(\oc8051_golden_model_1.PSW_bf [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_bf [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bf [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bf [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bf [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bf [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bf [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bf [7], \oc8051_golden_model_1.n1790 [7]);
  buf(\oc8051_golden_model_1.PSW_c3 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_c3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c3 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_d3 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_d3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d3 [7], 1'b1);
  buf(\oc8051_golden_model_1.PSW_d4 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_d4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d4 [7], \oc8051_golden_model_1.n1848 [7]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [0], \oc8051_golden_model_1.n1268 [0]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [1], \oc8051_golden_model_1.n1268 [1]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [2], \oc8051_golden_model_1.n1268 [2]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [3], \oc8051_golden_model_1.n1268 [3]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [4], \oc8051_golden_model_1.n1268 [4]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [5], \oc8051_golden_model_1.n1268 [5]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [6], \oc8051_golden_model_1.n1268 [6]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [7], \oc8051_golden_model_1.n1268 [8]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [4], \oc8051_golden_model_1.n1854 [4]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [5], \oc8051_golden_model_1.n1854 [5]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [6], \oc8051_golden_model_1.n1854 [6]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [7], \oc8051_golden_model_1.n1854 [7]);
  buf(\oc8051_golden_model_1.n0006 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0006 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0007 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0007 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0007 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0011 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0011 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0011 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0019 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0019 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0019 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0023 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0023 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0023 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0023 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0027 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0027 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0027 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0031 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0031 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0031 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0031 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0035 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0035 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0035 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0035 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0039 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0039 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0561 [0], \oc8051_golden_model_1.n1268 [0]);
  buf(\oc8051_golden_model_1.n0561 [1], \oc8051_golden_model_1.n1268 [1]);
  buf(\oc8051_golden_model_1.n0561 [2], \oc8051_golden_model_1.n1268 [2]);
  buf(\oc8051_golden_model_1.n0561 [3], \oc8051_golden_model_1.n1268 [3]);
  buf(\oc8051_golden_model_1.n0561 [4], \oc8051_golden_model_1.n1268 [4]);
  buf(\oc8051_golden_model_1.n0561 [5], \oc8051_golden_model_1.n1268 [5]);
  buf(\oc8051_golden_model_1.n0561 [6], \oc8051_golden_model_1.n1268 [6]);
  buf(\oc8051_golden_model_1.n0561 [7], \oc8051_golden_model_1.n1268 [8]);
  buf(\oc8051_golden_model_1.n0594 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.n0594 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.n0594 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.n0594 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.n0594 [4], \oc8051_golden_model_1.n1854 [4]);
  buf(\oc8051_golden_model_1.n0594 [5], \oc8051_golden_model_1.n1854 [5]);
  buf(\oc8051_golden_model_1.n0594 [6], \oc8051_golden_model_1.n1854 [6]);
  buf(\oc8051_golden_model_1.n0594 [7], \oc8051_golden_model_1.n1854 [7]);
  buf(\oc8051_golden_model_1.n0701 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n0701 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n0701 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n0701 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n0701 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n0701 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n0701 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n0701 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n0701 [8], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [9], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [10], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [11], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [12], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [13], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [14], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [15], 1'b0);
  buf(\oc8051_golden_model_1.n0733 [0], \oc8051_golden_model_1.DPL [0]);
  buf(\oc8051_golden_model_1.n0733 [1], \oc8051_golden_model_1.DPL [1]);
  buf(\oc8051_golden_model_1.n0733 [2], \oc8051_golden_model_1.DPL [2]);
  buf(\oc8051_golden_model_1.n0733 [3], \oc8051_golden_model_1.DPL [3]);
  buf(\oc8051_golden_model_1.n0733 [4], \oc8051_golden_model_1.DPL [4]);
  buf(\oc8051_golden_model_1.n0733 [5], \oc8051_golden_model_1.DPL [5]);
  buf(\oc8051_golden_model_1.n0733 [6], \oc8051_golden_model_1.DPL [6]);
  buf(\oc8051_golden_model_1.n0733 [7], \oc8051_golden_model_1.DPL [7]);
  buf(\oc8051_golden_model_1.n0733 [8], \oc8051_golden_model_1.DPH [0]);
  buf(\oc8051_golden_model_1.n0733 [9], \oc8051_golden_model_1.DPH [1]);
  buf(\oc8051_golden_model_1.n0733 [10], \oc8051_golden_model_1.DPH [2]);
  buf(\oc8051_golden_model_1.n0733 [11], \oc8051_golden_model_1.DPH [3]);
  buf(\oc8051_golden_model_1.n0733 [12], \oc8051_golden_model_1.DPH [4]);
  buf(\oc8051_golden_model_1.n0733 [13], \oc8051_golden_model_1.DPH [5]);
  buf(\oc8051_golden_model_1.n0733 [14], \oc8051_golden_model_1.DPH [6]);
  buf(\oc8051_golden_model_1.n0733 [15], \oc8051_golden_model_1.DPH [7]);
  buf(\oc8051_golden_model_1.n0994 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n0994 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n0994 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n0994 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n0994 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n0994 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n0994 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n0994 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1071 [0], \oc8051_golden_model_1.n1268 [0]);
  buf(\oc8051_golden_model_1.n1071 [1], \oc8051_golden_model_1.n1268 [1]);
  buf(\oc8051_golden_model_1.n1071 [2], \oc8051_golden_model_1.n1268 [2]);
  buf(\oc8051_golden_model_1.n1071 [3], \oc8051_golden_model_1.n1268 [3]);
  buf(\oc8051_golden_model_1.n1073 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1073 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1073 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1073 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1075 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1075 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1075 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1075 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1076 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1076 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1076 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1076 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1077 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1077 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1077 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1077 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1078 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1078 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1078 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1078 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1079 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1079 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1079 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1079 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1080 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1080 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1080 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1080 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1081 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1081 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1081 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1081 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1118 , \oc8051_golden_model_1.n1735 [7]);
  buf(\oc8051_golden_model_1.n1146 , \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1147 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1147 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1147 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1147 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1147 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1147 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1147 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1147 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1147 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1148 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1148 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1148 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1148 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1148 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1148 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1148 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1148 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1148 [8], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1149 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1149 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1149 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1149 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1149 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1149 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1149 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1149 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1150 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1151 , \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1152 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1152 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1152 [2], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1153 , \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1154 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1154 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1155 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1155 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1155 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1155 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1155 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1155 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1155 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1155 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1181 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.n1181 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.n1181 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.n1181 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.n1181 [4], \oc8051_golden_model_1.n1854 [4]);
  buf(\oc8051_golden_model_1.n1181 [5], \oc8051_golden_model_1.n1854 [5]);
  buf(\oc8051_golden_model_1.n1181 [6], \oc8051_golden_model_1.n1854 [6]);
  buf(\oc8051_golden_model_1.n1181 [7], \oc8051_golden_model_1.n1854 [7]);
  buf(\oc8051_golden_model_1.n1181 [8], \oc8051_golden_model_1.n1268 [0]);
  buf(\oc8051_golden_model_1.n1181 [9], \oc8051_golden_model_1.n1268 [1]);
  buf(\oc8051_golden_model_1.n1181 [10], \oc8051_golden_model_1.n1268 [2]);
  buf(\oc8051_golden_model_1.n1181 [11], \oc8051_golden_model_1.n1268 [3]);
  buf(\oc8051_golden_model_1.n1181 [12], \oc8051_golden_model_1.n1268 [4]);
  buf(\oc8051_golden_model_1.n1181 [13], \oc8051_golden_model_1.n1268 [5]);
  buf(\oc8051_golden_model_1.n1181 [14], \oc8051_golden_model_1.n1268 [6]);
  buf(\oc8051_golden_model_1.n1181 [15], \oc8051_golden_model_1.n1268 [8]);
  buf(\oc8051_golden_model_1.n1183 [0], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1183 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1183 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1183 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1183 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1183 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1183 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1183 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1185 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1185 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1185 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1185 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1185 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1185 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1185 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1185 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1185 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1189 [8], \oc8051_golden_model_1.n1207 [7]);
  buf(\oc8051_golden_model_1.n1190 , \oc8051_golden_model_1.n1207 [7]);
  buf(\oc8051_golden_model_1.n1191 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1191 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1191 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1191 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1192 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1192 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1192 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1192 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1192 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1196 [4], \oc8051_golden_model_1.n1207 [6]);
  buf(\oc8051_golden_model_1.n1197 , \oc8051_golden_model_1.n1207 [6]);
  buf(\oc8051_golden_model_1.n1198 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1198 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1198 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1198 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1198 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1198 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1198 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1198 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1198 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1206 , \oc8051_golden_model_1.n1207 [2]);
  buf(\oc8051_golden_model_1.n1207 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1207 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1207 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1207 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1207 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1211 [8], \oc8051_golden_model_1.n1227 [7]);
  buf(\oc8051_golden_model_1.n1212 , \oc8051_golden_model_1.n1227 [7]);
  buf(\oc8051_golden_model_1.n1217 [4], \oc8051_golden_model_1.n1227 [6]);
  buf(\oc8051_golden_model_1.n1218 , \oc8051_golden_model_1.n1227 [6]);
  buf(\oc8051_golden_model_1.n1226 , \oc8051_golden_model_1.n1227 [2]);
  buf(\oc8051_golden_model_1.n1227 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1227 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1227 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1227 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1227 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1229 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.n1229 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.n1229 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.n1229 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.n1229 [4], \oc8051_golden_model_1.n1854 [4]);
  buf(\oc8051_golden_model_1.n1229 [5], \oc8051_golden_model_1.n1854 [5]);
  buf(\oc8051_golden_model_1.n1229 [6], \oc8051_golden_model_1.n1854 [6]);
  buf(\oc8051_golden_model_1.n1229 [7], \oc8051_golden_model_1.n1854 [7]);
  buf(\oc8051_golden_model_1.n1229 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1231 [8], \oc8051_golden_model_1.n1246 [7]);
  buf(\oc8051_golden_model_1.n1232 , \oc8051_golden_model_1.n1246 [7]);
  buf(\oc8051_golden_model_1.n1233 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.n1233 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.n1233 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.n1233 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.n1234 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.n1234 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.n1234 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.n1234 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.n1234 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1236 [4], \oc8051_golden_model_1.n1258 [6]);
  buf(\oc8051_golden_model_1.n1237 , \oc8051_golden_model_1.n1258 [6]);
  buf(\oc8051_golden_model_1.n1238 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.n1238 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.n1238 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.n1238 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.n1238 [4], \oc8051_golden_model_1.n1854 [4]);
  buf(\oc8051_golden_model_1.n1238 [5], \oc8051_golden_model_1.n1854 [5]);
  buf(\oc8051_golden_model_1.n1238 [6], \oc8051_golden_model_1.n1854 [6]);
  buf(\oc8051_golden_model_1.n1238 [7], \oc8051_golden_model_1.n1854 [7]);
  buf(\oc8051_golden_model_1.n1238 [8], \oc8051_golden_model_1.n1854 [7]);
  buf(\oc8051_golden_model_1.n1245 , \oc8051_golden_model_1.n1246 [2]);
  buf(\oc8051_golden_model_1.n1246 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1246 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1246 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1246 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1246 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1246 [6], \oc8051_golden_model_1.n1258 [6]);
  buf(\oc8051_golden_model_1.n1249 [8], \oc8051_golden_model_1.n1258 [7]);
  buf(\oc8051_golden_model_1.n1250 , \oc8051_golden_model_1.n1258 [7]);
  buf(\oc8051_golden_model_1.n1257 , \oc8051_golden_model_1.n1258 [2]);
  buf(\oc8051_golden_model_1.n1258 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1258 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1258 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1258 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1258 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1260 [0], \oc8051_golden_model_1.n1268 [0]);
  buf(\oc8051_golden_model_1.n1260 [1], \oc8051_golden_model_1.n1268 [1]);
  buf(\oc8051_golden_model_1.n1260 [2], \oc8051_golden_model_1.n1268 [2]);
  buf(\oc8051_golden_model_1.n1260 [3], \oc8051_golden_model_1.n1268 [3]);
  buf(\oc8051_golden_model_1.n1260 [4], \oc8051_golden_model_1.n1268 [4]);
  buf(\oc8051_golden_model_1.n1260 [5], \oc8051_golden_model_1.n1268 [5]);
  buf(\oc8051_golden_model_1.n1260 [6], \oc8051_golden_model_1.n1268 [6]);
  buf(\oc8051_golden_model_1.n1260 [7], \oc8051_golden_model_1.n1268 [8]);
  buf(\oc8051_golden_model_1.n1260 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1262 [8], \oc8051_golden_model_1.n1280 [7]);
  buf(\oc8051_golden_model_1.n1263 , \oc8051_golden_model_1.n1280 [7]);
  buf(\oc8051_golden_model_1.n1264 [0], \oc8051_golden_model_1.n1268 [0]);
  buf(\oc8051_golden_model_1.n1264 [1], \oc8051_golden_model_1.n1268 [1]);
  buf(\oc8051_golden_model_1.n1264 [2], \oc8051_golden_model_1.n1268 [2]);
  buf(\oc8051_golden_model_1.n1264 [3], \oc8051_golden_model_1.n1268 [3]);
  buf(\oc8051_golden_model_1.n1264 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1266 [4], \oc8051_golden_model_1.n1292 [6]);
  buf(\oc8051_golden_model_1.n1267 , \oc8051_golden_model_1.n1292 [6]);
  buf(\oc8051_golden_model_1.n1268 [7], \oc8051_golden_model_1.n1268 [8]);
  buf(\oc8051_golden_model_1.n1275 , \oc8051_golden_model_1.n1280 [2]);
  buf(\oc8051_golden_model_1.n1276 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1276 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1276 [2], \oc8051_golden_model_1.n1280 [2]);
  buf(\oc8051_golden_model_1.n1276 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1276 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1276 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1276 [6], \oc8051_golden_model_1.n1292 [6]);
  buf(\oc8051_golden_model_1.n1276 [7], \oc8051_golden_model_1.n1280 [7]);
  buf(\oc8051_golden_model_1.n1278 [4], \oc8051_golden_model_1.n1291 [6]);
  buf(\oc8051_golden_model_1.n1279 , \oc8051_golden_model_1.n1291 [6]);
  buf(\oc8051_golden_model_1.n1280 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1280 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1280 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1280 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1280 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1280 [6], \oc8051_golden_model_1.n1291 [6]);
  buf(\oc8051_golden_model_1.n1282 [8], \oc8051_golden_model_1.n1292 [7]);
  buf(\oc8051_golden_model_1.n1283 , \oc8051_golden_model_1.n1292 [7]);
  buf(\oc8051_golden_model_1.n1290 , \oc8051_golden_model_1.n1292 [2]);
  buf(\oc8051_golden_model_1.n1291 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1291 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1291 [2], \oc8051_golden_model_1.n1292 [2]);
  buf(\oc8051_golden_model_1.n1291 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1291 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1291 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1291 [7], \oc8051_golden_model_1.n1292 [7]);
  buf(\oc8051_golden_model_1.n1292 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1292 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1292 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1292 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1292 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1295 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1295 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1295 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1295 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1295 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1295 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1295 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1295 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1295 [8], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1296 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1296 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1296 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1296 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1296 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1296 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1296 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1296 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1296 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1297 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1297 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1297 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1297 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1297 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1297 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1297 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1297 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1298 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1299 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1299 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1299 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1299 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1299 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1299 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1299 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1299 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1300 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1300 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1300 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1300 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1300 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1300 [5], 1'b0);
  buf(\oc8051_golden_model_1.n1300 [6], 1'b0);
  buf(\oc8051_golden_model_1.n1300 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1303 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1303 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1303 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1303 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1303 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1303 [5], 1'b0);
  buf(\oc8051_golden_model_1.n1303 [6], 1'b0);
  buf(\oc8051_golden_model_1.n1303 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1303 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1305 [8], \oc8051_golden_model_1.n1318 [7]);
  buf(\oc8051_golden_model_1.n1306 , \oc8051_golden_model_1.n1318 [7]);
  buf(\oc8051_golden_model_1.n1307 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1307 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1307 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1307 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1307 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1309 [4], \oc8051_golden_model_1.n1318 [6]);
  buf(\oc8051_golden_model_1.n1310 , \oc8051_golden_model_1.n1318 [6]);
  buf(\oc8051_golden_model_1.n1317 , \oc8051_golden_model_1.n1318 [2]);
  buf(\oc8051_golden_model_1.n1318 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1318 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1318 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1318 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1318 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1322 [8], \oc8051_golden_model_1.n1334 [7]);
  buf(\oc8051_golden_model_1.n1323 , \oc8051_golden_model_1.n1334 [7]);
  buf(\oc8051_golden_model_1.n1325 [4], \oc8051_golden_model_1.n1334 [6]);
  buf(\oc8051_golden_model_1.n1326 , \oc8051_golden_model_1.n1334 [6]);
  buf(\oc8051_golden_model_1.n1333 , \oc8051_golden_model_1.n1334 [2]);
  buf(\oc8051_golden_model_1.n1334 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1334 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1334 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1334 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1334 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1338 [8], \oc8051_golden_model_1.n1350 [7]);
  buf(\oc8051_golden_model_1.n1339 , \oc8051_golden_model_1.n1350 [7]);
  buf(\oc8051_golden_model_1.n1341 [4], \oc8051_golden_model_1.n1350 [6]);
  buf(\oc8051_golden_model_1.n1342 , \oc8051_golden_model_1.n1350 [6]);
  buf(\oc8051_golden_model_1.n1349 , \oc8051_golden_model_1.n1350 [2]);
  buf(\oc8051_golden_model_1.n1350 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1350 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1350 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1350 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1350 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1354 [8], \oc8051_golden_model_1.n1366 [7]);
  buf(\oc8051_golden_model_1.n1355 , \oc8051_golden_model_1.n1366 [7]);
  buf(\oc8051_golden_model_1.n1357 [4], \oc8051_golden_model_1.n1366 [6]);
  buf(\oc8051_golden_model_1.n1358 , \oc8051_golden_model_1.n1366 [6]);
  buf(\oc8051_golden_model_1.n1365 , \oc8051_golden_model_1.n1366 [2]);
  buf(\oc8051_golden_model_1.n1366 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1366 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1366 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1366 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1366 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1520 , \oc8051_golden_model_1.n1522 [7]);
  buf(\oc8051_golden_model_1.n1521 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1521 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1521 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1521 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1521 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1521 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1521 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1522 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1522 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1522 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1522 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1522 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1522 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1522 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1545 , \oc8051_golden_model_1.n1546 [7]);
  buf(\oc8051_golden_model_1.n1546 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1546 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1546 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1546 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1546 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1546 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1546 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1553 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1553 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1553 [2], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1553 [3], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1554 , \oc8051_golden_model_1.n1555 [2]);
  buf(\oc8051_golden_model_1.n1555 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1555 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1555 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1555 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1555 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1555 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1555 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1680 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1680 [1], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1680 [2], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1680 [3], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1680 [4], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1680 [5], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1680 [6], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1680 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1683 , \oc8051_golden_model_1.n1692 [7]);
  buf(\oc8051_golden_model_1.n1685 , \oc8051_golden_model_1.n1692 [6]);
  buf(\oc8051_golden_model_1.n1691 , \oc8051_golden_model_1.n1692 [2]);
  buf(\oc8051_golden_model_1.n1692 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1692 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1692 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1692 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1692 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1696 , \oc8051_golden_model_1.n1705 [7]);
  buf(\oc8051_golden_model_1.n1698 , \oc8051_golden_model_1.n1705 [6]);
  buf(\oc8051_golden_model_1.n1704 , \oc8051_golden_model_1.n1705 [2]);
  buf(\oc8051_golden_model_1.n1705 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1705 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1705 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1705 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1705 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1709 , \oc8051_golden_model_1.n1718 [7]);
  buf(\oc8051_golden_model_1.n1711 , \oc8051_golden_model_1.n1718 [6]);
  buf(\oc8051_golden_model_1.n1717 , \oc8051_golden_model_1.n1718 [2]);
  buf(\oc8051_golden_model_1.n1718 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1718 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1718 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1718 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1718 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1722 , \oc8051_golden_model_1.n1731 [7]);
  buf(\oc8051_golden_model_1.n1724 , \oc8051_golden_model_1.n1731 [6]);
  buf(\oc8051_golden_model_1.n1730 , \oc8051_golden_model_1.n1731 [2]);
  buf(\oc8051_golden_model_1.n1731 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1731 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1731 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1731 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1731 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1733 , \oc8051_golden_model_1.n1734 [7]);
  buf(\oc8051_golden_model_1.n1734 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1734 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1734 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1734 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1734 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1734 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1734 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1735 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1735 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1735 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1735 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1735 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1735 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1735 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1739 [0], \oc8051_golden_model_1.B [0]);
  buf(\oc8051_golden_model_1.n1739 [1], \oc8051_golden_model_1.B [1]);
  buf(\oc8051_golden_model_1.n1739 [2], \oc8051_golden_model_1.B [2]);
  buf(\oc8051_golden_model_1.n1739 [3], \oc8051_golden_model_1.B [3]);
  buf(\oc8051_golden_model_1.n1739 [4], \oc8051_golden_model_1.B [4]);
  buf(\oc8051_golden_model_1.n1739 [5], \oc8051_golden_model_1.B [5]);
  buf(\oc8051_golden_model_1.n1739 [6], \oc8051_golden_model_1.B [6]);
  buf(\oc8051_golden_model_1.n1739 [7], \oc8051_golden_model_1.B [7]);
  buf(\oc8051_golden_model_1.n1739 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1739 [9], 1'b0);
  buf(\oc8051_golden_model_1.n1739 [10], 1'b0);
  buf(\oc8051_golden_model_1.n1739 [11], 1'b0);
  buf(\oc8051_golden_model_1.n1739 [12], 1'b0);
  buf(\oc8051_golden_model_1.n1739 [13], 1'b0);
  buf(\oc8051_golden_model_1.n1739 [14], 1'b0);
  buf(\oc8051_golden_model_1.n1739 [15], 1'b0);
  buf(\oc8051_golden_model_1.n1745 , \oc8051_golden_model_1.n1746 [2]);
  buf(\oc8051_golden_model_1.n1746 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1746 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1746 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1746 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1746 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1746 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1746 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1749 , \oc8051_golden_model_1.n1750 [7]);
  buf(\oc8051_golden_model_1.n1750 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1750 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1750 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1750 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1750 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1750 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1750 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1765 , \oc8051_golden_model_1.n1766 [7]);
  buf(\oc8051_golden_model_1.n1766 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1766 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1766 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1766 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1766 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1766 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1766 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1771 , \oc8051_golden_model_1.n1772 [7]);
  buf(\oc8051_golden_model_1.n1772 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1772 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1772 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1772 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1772 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1772 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1772 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1777 , \oc8051_golden_model_1.n1778 [7]);
  buf(\oc8051_golden_model_1.n1778 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1778 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1778 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1778 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1778 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1778 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1778 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1783 , \oc8051_golden_model_1.n1784 [7]);
  buf(\oc8051_golden_model_1.n1784 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1784 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1784 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1784 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1784 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1784 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1784 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1789 , \oc8051_golden_model_1.n1790 [7]);
  buf(\oc8051_golden_model_1.n1790 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1790 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1790 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1790 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1790 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1790 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1790 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1791 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1791 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1791 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1791 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1791 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1791 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1791 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1791 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1792 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1792 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1792 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1792 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1793 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1793 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1793 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1793 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1793 [4], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1793 [5], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1793 [6], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1793 [7], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1828 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1828 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1828 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1828 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1828 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1828 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1828 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1828 [7], 1'b1);
  buf(\oc8051_golden_model_1.n1847 , \oc8051_golden_model_1.n1848 [7]);
  buf(\oc8051_golden_model_1.n1848 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1848 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1848 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1848 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1848 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1848 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1848 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1852 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1852 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1852 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1852 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1853 [0], \oc8051_golden_model_1.n1854 [4]);
  buf(\oc8051_golden_model_1.n1853 [1], \oc8051_golden_model_1.n1854 [5]);
  buf(\oc8051_golden_model_1.n1853 [2], \oc8051_golden_model_1.n1854 [6]);
  buf(\oc8051_golden_model_1.n1853 [3], \oc8051_golden_model_1.n1854 [7]);
  buf(\oc8051_golden_model_1.n1854 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1854 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1854 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1854 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_top_1.wb_rst_i , rst);
  buf(\oc8051_top_1.wb_clk_i , clk);
  buf(\oc8051_top_1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_top_1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_top_1.pc_log [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_top_1.pc_log [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_top_1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_top_1.pc_log [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_top_1.pc_log [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_top_1.pc_log [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_top_1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_top_1.pc_log [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_top_1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_top_1.pc_log [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_top_1.pc_log [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_top_1.pc_log [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_top_1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_top_1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_top_1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_top_1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_top_1.pc_log_prev [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_top_1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_top_1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_top_1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_top_1.pc_log_prev [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_top_1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_top_1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_top_1.pc_log_prev [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_top_1.pc_log_prev [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_top_1.pc_log_prev [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_top_1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_top_1.pc_log_prev [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_top_1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_top_1.psw [0], psw[0]);
  buf(\oc8051_top_1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.wbd_we_o , \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  buf(\oc8051_top_1.wbd_stb_o , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.wbd_cyc_o , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.wbd_dat_o [0], \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  buf(\oc8051_top_1.wbd_dat_o [1], \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  buf(\oc8051_top_1.wbd_dat_o [2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  buf(\oc8051_top_1.wbd_dat_o [3], \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  buf(\oc8051_top_1.wbd_dat_o [4], \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  buf(\oc8051_top_1.wbd_dat_o [5], \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  buf(\oc8051_top_1.wbd_dat_o [6], \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  buf(\oc8051_top_1.wbd_dat_o [7], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  buf(\oc8051_top_1.wbd_adr_o [0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(\oc8051_top_1.wbd_adr_o [1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(\oc8051_top_1.wbd_adr_o [2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(\oc8051_top_1.wbd_adr_o [3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(\oc8051_top_1.wbd_adr_o [4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(\oc8051_top_1.wbd_adr_o [5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(\oc8051_top_1.wbd_adr_o [6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(\oc8051_top_1.wbd_adr_o [7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(\oc8051_top_1.wbd_adr_o [8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(\oc8051_top_1.wbd_adr_o [9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(\oc8051_top_1.wbd_adr_o [10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(\oc8051_top_1.wbd_adr_o [11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(\oc8051_top_1.wbd_adr_o [12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(\oc8051_top_1.wbd_adr_o [13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(\oc8051_top_1.wbd_adr_o [14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(\oc8051_top_1.wbd_adr_o [15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(\oc8051_top_1.cxrom_data_out [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.cxrom_data_out [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.cxrom_data_out [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.cxrom_data_out [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.cxrom_data_out [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.cxrom_data_out [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.cxrom_data_out [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.cxrom_data_out [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.cxrom_data_out [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.cxrom_data_out [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.cxrom_data_out [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.cxrom_data_out [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.cxrom_data_out [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.cxrom_data_out [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.cxrom_data_out [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.cxrom_data_out [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.cxrom_data_out [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.cxrom_data_out [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.cxrom_data_out [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.cxrom_data_out [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.cxrom_data_out [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.cxrom_data_out [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.cxrom_data_out [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.cxrom_data_out [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.cxrom_data_out [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.cxrom_data_out [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.cxrom_data_out [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.cxrom_data_out [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.cxrom_data_out [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.cxrom_data_out [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.cxrom_data_out [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.cxrom_data_out [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.p0_i [0], p0_in[0]);
  buf(\oc8051_top_1.p0_i [1], p0_in[1]);
  buf(\oc8051_top_1.p0_i [2], p0_in[2]);
  buf(\oc8051_top_1.p0_i [3], p0_in[3]);
  buf(\oc8051_top_1.p0_i [4], p0_in[4]);
  buf(\oc8051_top_1.p0_i [5], p0_in[5]);
  buf(\oc8051_top_1.p0_i [6], p0_in[6]);
  buf(\oc8051_top_1.p0_i [7], p0_in[7]);
  buf(\oc8051_top_1.p0_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.p0_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.p0_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.p0_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.p0_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.p0_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.p0_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.p0_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.p1_i [0], p1_in[0]);
  buf(\oc8051_top_1.p1_i [1], p1_in[1]);
  buf(\oc8051_top_1.p1_i [2], p1_in[2]);
  buf(\oc8051_top_1.p1_i [3], p1_in[3]);
  buf(\oc8051_top_1.p1_i [4], p1_in[4]);
  buf(\oc8051_top_1.p1_i [5], p1_in[5]);
  buf(\oc8051_top_1.p1_i [6], p1_in[6]);
  buf(\oc8051_top_1.p1_i [7], p1_in[7]);
  buf(\oc8051_top_1.p1_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.p1_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.p1_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.p1_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.p1_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.p1_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.p1_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.p1_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.p2_i [0], p2_in[0]);
  buf(\oc8051_top_1.p2_i [1], p2_in[1]);
  buf(\oc8051_top_1.p2_i [2], p2_in[2]);
  buf(\oc8051_top_1.p2_i [3], p2_in[3]);
  buf(\oc8051_top_1.p2_i [4], p2_in[4]);
  buf(\oc8051_top_1.p2_i [5], p2_in[5]);
  buf(\oc8051_top_1.p2_i [6], p2_in[6]);
  buf(\oc8051_top_1.p2_i [7], p2_in[7]);
  buf(\oc8051_top_1.p2_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.p2_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.p2_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.p2_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.p2_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.p2_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.p2_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.p2_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.p3_i [0], p3_in[0]);
  buf(\oc8051_top_1.p3_i [1], p3_in[1]);
  buf(\oc8051_top_1.p3_i [2], p3_in[2]);
  buf(\oc8051_top_1.p3_i [3], p3_in[3]);
  buf(\oc8051_top_1.p3_i [4], p3_in[4]);
  buf(\oc8051_top_1.p3_i [5], p3_in[5]);
  buf(\oc8051_top_1.p3_i [6], p3_in[6]);
  buf(\oc8051_top_1.p3_i [7], p3_in[7]);
  buf(\oc8051_top_1.p3_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.p3_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.p3_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.p3_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.p3_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.p3_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.p3_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.p3_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.rxd_i , rxd_i);
  buf(\oc8051_top_1.txd_o , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  buf(\oc8051_top_1.t0_i , t0_i);
  buf(\oc8051_top_1.t1_i , t1_i);
  buf(\oc8051_top_1.t2_i , t2_i);
  buf(\oc8051_top_1.t2ex_i , t2ex_i);
  buf(\oc8051_top_1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.src_sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.src_sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.sfr_out [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.sfr_out [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.sfr_out [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.sfr_out [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.sfr_out [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.sfr_out [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.sfr_out [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.sfr_out [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.rd_ind , \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  buf(\oc8051_top_1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(rd_iram_addr[0], word_in[0]);
  buf(rd_iram_addr[1], word_in[1]);
  buf(rd_iram_addr[2], word_in[2]);
  buf(rd_iram_addr[3], word_in[3]);
  buf(rd_rom_0_addr[0], \oc8051_golden_model_1.PC [0]);
  buf(rd_rom_0_addr[1], \oc8051_golden_model_1.PC [1]);
  buf(rd_rom_0_addr[2], \oc8051_golden_model_1.PC [2]);
  buf(rd_rom_0_addr[3], \oc8051_golden_model_1.PC [3]);
  buf(rd_rom_0_addr[4], \oc8051_golden_model_1.PC [4]);
  buf(rd_rom_0_addr[5], \oc8051_golden_model_1.PC [5]);
  buf(rd_rom_0_addr[6], \oc8051_golden_model_1.PC [6]);
  buf(rd_rom_0_addr[7], \oc8051_golden_model_1.PC [7]);
  buf(rd_rom_0_addr[8], \oc8051_golden_model_1.PC [8]);
  buf(rd_rom_0_addr[9], \oc8051_golden_model_1.PC [9]);
  buf(rd_rom_0_addr[10], \oc8051_golden_model_1.PC [10]);
  buf(rd_rom_0_addr[11], \oc8051_golden_model_1.PC [11]);
  buf(rd_rom_0_addr[12], \oc8051_golden_model_1.PC [12]);
  buf(rd_rom_0_addr[13], \oc8051_golden_model_1.PC [13]);
  buf(rd_rom_0_addr[14], \oc8051_golden_model_1.PC [14]);
  buf(rd_rom_0_addr[15], \oc8051_golden_model_1.PC [15]);
  buf(ACC_gm[0], \oc8051_golden_model_1.ACC [0]);
  buf(ACC_gm[1], \oc8051_golden_model_1.ACC [1]);
  buf(ACC_gm[2], \oc8051_golden_model_1.ACC [2]);
  buf(ACC_gm[3], \oc8051_golden_model_1.ACC [3]);
  buf(ACC_gm[4], \oc8051_golden_model_1.ACC [4]);
  buf(ACC_gm[5], \oc8051_golden_model_1.ACC [5]);
  buf(ACC_gm[6], \oc8051_golden_model_1.ACC [6]);
  buf(ACC_gm[7], \oc8051_golden_model_1.ACC [7]);
  buf(acc[0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(acc[1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(acc[2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(acc[3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(acc[4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(acc[5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(acc[6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(acc[7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(psw[1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(psw[2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(psw[3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(psw[4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(psw[5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(psw[6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(psw[7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(pc1[0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(pc1[1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(pc1[2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(pc1[3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(pc1[4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(pc1[5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(pc1[6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(pc1[7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(pc1[8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(pc1[9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(pc1[10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(pc1[11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(pc1[12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(pc1[13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(pc1[14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(pc1[15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(pc2[0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(pc2[1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(pc2[2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(pc2[3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(pc2[4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(pc2[5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(pc2[6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(pc2[7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(pc2[8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(pc2[9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(pc2[10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(pc2[11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(pc2[12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(pc2[13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(pc2[14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(pc2[15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(cxrom_data_out[0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(cxrom_data_out[1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(cxrom_data_out[2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(cxrom_data_out[3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(cxrom_data_out[4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(cxrom_data_out[5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(cxrom_data_out[6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(cxrom_data_out[7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(cxrom_data_out[8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(cxrom_data_out[9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(cxrom_data_out[10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(cxrom_data_out[11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(cxrom_data_out[12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(cxrom_data_out[13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(cxrom_data_out[14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(cxrom_data_out[15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(cxrom_data_out[16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(cxrom_data_out[17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(cxrom_data_out[18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(cxrom_data_out[19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(cxrom_data_out[20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(cxrom_data_out[21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(cxrom_data_out[22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(cxrom_data_out[23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(cxrom_data_out[24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(cxrom_data_out[25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(cxrom_data_out[26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(cxrom_data_out[27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(cxrom_data_out[28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(cxrom_data_out[29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(cxrom_data_out[30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(cxrom_data_out[31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(wbd_adr_o[0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(wbd_adr_o[1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(wbd_adr_o[2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(wbd_adr_o[3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(wbd_adr_o[4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(wbd_adr_o[5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(wbd_adr_o[6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(wbd_adr_o[7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(wbd_adr_o[8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(wbd_adr_o[9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(wbd_adr_o[10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(wbd_adr_o[11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(wbd_adr_o[12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(wbd_adr_o[13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(wbd_adr_o[14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(wbd_adr_o[15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(wbd_dat_o[0], \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  buf(wbd_dat_o[1], \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  buf(wbd_dat_o[2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  buf(wbd_dat_o[3], \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  buf(wbd_dat_o[4], \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  buf(wbd_dat_o[5], \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  buf(wbd_dat_o[6], \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  buf(wbd_dat_o[7], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  buf(wbd_cyc_o, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_stb_o, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_we_o, \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  buf(txd_o, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  buf(p3_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(p3_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(p3_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(p3_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(p3_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(p3_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(p3_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(p3_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(p2_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(p2_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(p2_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(p2_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(p2_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(p2_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(p2_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(p2_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(p1_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(p1_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(p1_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(p1_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(p1_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(p1_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(p1_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(p1_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(p0_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(p0_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(p0_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(p0_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(p0_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(p0_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(p0_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(p0_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
endmodule
